i P1_MEMORYFETCH_REG_SCAN_IN
i DATAI_31_
i DATAI_30_
i DATAI_29_
i DATAI_28_
i DATAI_27_
i DATAI_26_
i DATAI_25_
i DATAI_24_
i DATAI_23_
i DATAI_22_
i DATAI_21_
i DATAI_20_
i DATAI_19_
i DATAI_18_
i DATAI_17_
i DATAI_16_
i DATAI_15_
i DATAI_14_
i DATAI_13_
i DATAI_12_
i DATAI_11_
i DATAI_10_
i DATAI_9_
i DATAI_8_
i DATAI_7_
i DATAI_6_
i DATAI_5_
i DATAI_4_
i DATAI_3_
i DATAI_2_
i DATAI_1_
i DATAI_0_
i HOLD
i NA
i BS16
i READY1
i READY2
i P1_READREQUEST_REG_SCAN_IN
i P1_ADS_N_REG_SCAN_IN
i P1_CODEFETCH_REG_SCAN_IN
i P1_M_IO_N_REG_SCAN_IN
i P1_D_C_N_REG_SCAN_IN
i P1_REQUESTPENDING_REG_SCAN_IN
i P1_STATEBS16_REG_SCAN_IN
i P1_MORE_REG_SCAN_IN
i P1_FLUSH_REG_SCAN_IN
i P1_W_R_N_REG_SCAN_IN
i P1_BYTEENABLE_REG_0__SCAN_IN
i P1_BYTEENABLE_REG_1__SCAN_IN
i P1_BYTEENABLE_REG_2__SCAN_IN
i P1_BYTEENABLE_REG_3__SCAN_IN
i P1_REIP_REG_31__SCAN_IN
i P1_REIP_REG_30__SCAN_IN
i P1_REIP_REG_29__SCAN_IN
i P1_REIP_REG_28__SCAN_IN
i P1_REIP_REG_27__SCAN_IN
i P1_REIP_REG_26__SCAN_IN
i P1_REIP_REG_25__SCAN_IN
i P1_REIP_REG_24__SCAN_IN
i P1_REIP_REG_23__SCAN_IN
i P1_REIP_REG_22__SCAN_IN
i P1_REIP_REG_21__SCAN_IN
i P1_REIP_REG_20__SCAN_IN
i P1_REIP_REG_19__SCAN_IN
i P1_REIP_REG_18__SCAN_IN
i P1_REIP_REG_17__SCAN_IN
i P1_REIP_REG_16__SCAN_IN
i P1_REIP_REG_15__SCAN_IN
i P1_REIP_REG_14__SCAN_IN
i P1_REIP_REG_13__SCAN_IN
i P1_REIP_REG_12__SCAN_IN
i P1_REIP_REG_11__SCAN_IN
i P1_REIP_REG_10__SCAN_IN
i P1_REIP_REG_9__SCAN_IN
i P1_REIP_REG_8__SCAN_IN
i P1_REIP_REG_7__SCAN_IN
i P1_REIP_REG_6__SCAN_IN
i P1_REIP_REG_5__SCAN_IN
i P1_REIP_REG_4__SCAN_IN
i P1_REIP_REG_3__SCAN_IN
i P1_REIP_REG_2__SCAN_IN
i P1_REIP_REG_1__SCAN_IN
i P1_REIP_REG_0__SCAN_IN
i P1_EBX_REG_31__SCAN_IN
i P1_EBX_REG_30__SCAN_IN
i P1_EBX_REG_29__SCAN_IN
i P1_EBX_REG_28__SCAN_IN
i P1_EBX_REG_27__SCAN_IN
i P1_EBX_REG_26__SCAN_IN
i P1_EBX_REG_25__SCAN_IN
i P1_EBX_REG_24__SCAN_IN
i P1_EBX_REG_23__SCAN_IN
i P1_EBX_REG_22__SCAN_IN
i P1_EBX_REG_21__SCAN_IN
i P1_EBX_REG_20__SCAN_IN
i P1_EBX_REG_19__SCAN_IN
i P1_EBX_REG_18__SCAN_IN
i P1_EBX_REG_17__SCAN_IN
i P1_EBX_REG_16__SCAN_IN
i P1_EBX_REG_15__SCAN_IN
i P1_EBX_REG_14__SCAN_IN
i P1_EBX_REG_13__SCAN_IN
i P1_EBX_REG_12__SCAN_IN
i P1_EBX_REG_11__SCAN_IN
i P1_EBX_REG_10__SCAN_IN
i P1_EBX_REG_9__SCAN_IN
i P1_EBX_REG_8__SCAN_IN
i P1_EBX_REG_7__SCAN_IN
i P1_EBX_REG_6__SCAN_IN
i P1_EBX_REG_5__SCAN_IN
i P1_EBX_REG_4__SCAN_IN
i P1_EBX_REG_3__SCAN_IN
i P1_EBX_REG_2__SCAN_IN
i P1_EBX_REG_1__SCAN_IN
i P1_EBX_REG_0__SCAN_IN
i P1_EAX_REG_31__SCAN_IN
i P1_EAX_REG_30__SCAN_IN
i P1_EAX_REG_29__SCAN_IN
i P1_EAX_REG_28__SCAN_IN
i P1_EAX_REG_27__SCAN_IN
i P1_EAX_REG_26__SCAN_IN
i P1_EAX_REG_25__SCAN_IN
i P1_EAX_REG_24__SCAN_IN
i P1_EAX_REG_23__SCAN_IN
i P1_EAX_REG_22__SCAN_IN
i P1_EAX_REG_21__SCAN_IN
i P1_EAX_REG_20__SCAN_IN
i P1_EAX_REG_19__SCAN_IN
i P1_EAX_REG_18__SCAN_IN
i P1_EAX_REG_17__SCAN_IN
i P1_EAX_REG_16__SCAN_IN
i P1_EAX_REG_15__SCAN_IN
i P1_EAX_REG_14__SCAN_IN
i P1_EAX_REG_13__SCAN_IN
i P1_EAX_REG_12__SCAN_IN
i P1_EAX_REG_11__SCAN_IN
i P1_EAX_REG_10__SCAN_IN
i P1_EAX_REG_9__SCAN_IN
i P1_EAX_REG_8__SCAN_IN
i P1_EAX_REG_7__SCAN_IN
i P1_EAX_REG_6__SCAN_IN
i P1_EAX_REG_5__SCAN_IN
i P1_EAX_REG_4__SCAN_IN
i P1_EAX_REG_3__SCAN_IN
i P1_EAX_REG_2__SCAN_IN
i P1_EAX_REG_1__SCAN_IN
i P1_EAX_REG_0__SCAN_IN
i P1_DATAO_REG_31__SCAN_IN
i P1_DATAO_REG_30__SCAN_IN
i P1_DATAO_REG_29__SCAN_IN
i P1_DATAO_REG_28__SCAN_IN
i P1_DATAO_REG_27__SCAN_IN
i P1_DATAO_REG_26__SCAN_IN
i P1_DATAO_REG_25__SCAN_IN
i P1_DATAO_REG_24__SCAN_IN
i P1_DATAO_REG_23__SCAN_IN
i P1_DATAO_REG_22__SCAN_IN
i P1_DATAO_REG_21__SCAN_IN
i P1_DATAO_REG_20__SCAN_IN
i P1_DATAO_REG_19__SCAN_IN
i P1_DATAO_REG_18__SCAN_IN
i P1_DATAO_REG_17__SCAN_IN
i P1_DATAO_REG_16__SCAN_IN
i P1_DATAO_REG_15__SCAN_IN
i P1_DATAO_REG_14__SCAN_IN
i P1_DATAO_REG_13__SCAN_IN
i P1_DATAO_REG_12__SCAN_IN
i P1_DATAO_REG_11__SCAN_IN
i P1_DATAO_REG_10__SCAN_IN
i P1_DATAO_REG_9__SCAN_IN
i P1_DATAO_REG_8__SCAN_IN
i P1_DATAO_REG_7__SCAN_IN
i P1_DATAO_REG_6__SCAN_IN
i P1_DATAO_REG_5__SCAN_IN
i P1_DATAO_REG_4__SCAN_IN
i P1_DATAO_REG_3__SCAN_IN
i P1_DATAO_REG_2__SCAN_IN
i P1_DATAO_REG_1__SCAN_IN
i P1_DATAO_REG_0__SCAN_IN
i P1_UWORD_REG_0__SCAN_IN
i P1_UWORD_REG_1__SCAN_IN
i P1_UWORD_REG_2__SCAN_IN
i P1_UWORD_REG_3__SCAN_IN
i P1_UWORD_REG_4__SCAN_IN
i P1_UWORD_REG_5__SCAN_IN
i P1_UWORD_REG_6__SCAN_IN
i P1_UWORD_REG_7__SCAN_IN
i P1_UWORD_REG_8__SCAN_IN
i P1_UWORD_REG_9__SCAN_IN
i P1_UWORD_REG_10__SCAN_IN
i P1_UWORD_REG_11__SCAN_IN
i P1_UWORD_REG_12__SCAN_IN
i P1_UWORD_REG_13__SCAN_IN
i P1_UWORD_REG_14__SCAN_IN
i P1_LWORD_REG_0__SCAN_IN
i P1_LWORD_REG_1__SCAN_IN
i P1_LWORD_REG_2__SCAN_IN
i P1_LWORD_REG_3__SCAN_IN
i P1_LWORD_REG_4__SCAN_IN
i P1_LWORD_REG_5__SCAN_IN
i P1_LWORD_REG_6__SCAN_IN
i P1_LWORD_REG_7__SCAN_IN
i P1_LWORD_REG_8__SCAN_IN
i P1_LWORD_REG_9__SCAN_IN
i P1_LWORD_REG_10__SCAN_IN
i P1_LWORD_REG_11__SCAN_IN
i P1_LWORD_REG_12__SCAN_IN
i P1_LWORD_REG_13__SCAN_IN
i P1_LWORD_REG_14__SCAN_IN
i P1_LWORD_REG_15__SCAN_IN
i P1_PHYADDRPOINTER_REG_31__SCAN_IN
i P1_PHYADDRPOINTER_REG_30__SCAN_IN
i P1_PHYADDRPOINTER_REG_29__SCAN_IN
i P1_PHYADDRPOINTER_REG_28__SCAN_IN
i P1_PHYADDRPOINTER_REG_27__SCAN_IN
i P1_PHYADDRPOINTER_REG_26__SCAN_IN
i P1_PHYADDRPOINTER_REG_25__SCAN_IN
i P1_PHYADDRPOINTER_REG_24__SCAN_IN
i P1_PHYADDRPOINTER_REG_23__SCAN_IN
i P1_PHYADDRPOINTER_REG_22__SCAN_IN
i P1_PHYADDRPOINTER_REG_21__SCAN_IN
i P1_PHYADDRPOINTER_REG_20__SCAN_IN
i P1_PHYADDRPOINTER_REG_19__SCAN_IN
i P1_PHYADDRPOINTER_REG_18__SCAN_IN
i P1_PHYADDRPOINTER_REG_17__SCAN_IN
i P1_PHYADDRPOINTER_REG_16__SCAN_IN
i P1_PHYADDRPOINTER_REG_15__SCAN_IN
i P1_PHYADDRPOINTER_REG_14__SCAN_IN
i P1_PHYADDRPOINTER_REG_13__SCAN_IN
i P1_PHYADDRPOINTER_REG_12__SCAN_IN
i P1_PHYADDRPOINTER_REG_11__SCAN_IN
i P1_PHYADDRPOINTER_REG_10__SCAN_IN
i P1_PHYADDRPOINTER_REG_9__SCAN_IN
i P1_PHYADDRPOINTER_REG_8__SCAN_IN
i P1_PHYADDRPOINTER_REG_7__SCAN_IN
i P1_PHYADDRPOINTER_REG_6__SCAN_IN
i P1_PHYADDRPOINTER_REG_5__SCAN_IN
i P1_PHYADDRPOINTER_REG_4__SCAN_IN
i P1_PHYADDRPOINTER_REG_3__SCAN_IN
i P1_PHYADDRPOINTER_REG_2__SCAN_IN
i P1_PHYADDRPOINTER_REG_1__SCAN_IN
i P1_PHYADDRPOINTER_REG_0__SCAN_IN
i P1_INSTADDRPOINTER_REG_31__SCAN_IN
i P1_INSTADDRPOINTER_REG_30__SCAN_IN
i P1_INSTADDRPOINTER_REG_29__SCAN_IN
i P1_INSTADDRPOINTER_REG_28__SCAN_IN
i P1_INSTADDRPOINTER_REG_27__SCAN_IN
i P1_INSTADDRPOINTER_REG_26__SCAN_IN
i P1_INSTADDRPOINTER_REG_25__SCAN_IN
i P1_INSTADDRPOINTER_REG_24__SCAN_IN
i P1_INSTADDRPOINTER_REG_23__SCAN_IN
i P1_INSTADDRPOINTER_REG_22__SCAN_IN
i P1_INSTADDRPOINTER_REG_21__SCAN_IN
i P1_INSTADDRPOINTER_REG_20__SCAN_IN
i P1_INSTADDRPOINTER_REG_19__SCAN_IN
i P1_INSTADDRPOINTER_REG_18__SCAN_IN
i P1_INSTADDRPOINTER_REG_17__SCAN_IN
i P1_INSTADDRPOINTER_REG_16__SCAN_IN
i P1_INSTADDRPOINTER_REG_15__SCAN_IN
i P1_INSTADDRPOINTER_REG_14__SCAN_IN
i P1_INSTADDRPOINTER_REG_13__SCAN_IN
i P1_INSTADDRPOINTER_REG_12__SCAN_IN
i P1_INSTADDRPOINTER_REG_11__SCAN_IN
i P1_INSTADDRPOINTER_REG_10__SCAN_IN
i P1_INSTADDRPOINTER_REG_9__SCAN_IN
i P1_INSTADDRPOINTER_REG_8__SCAN_IN
i P1_INSTADDRPOINTER_REG_7__SCAN_IN
i P1_INSTADDRPOINTER_REG_6__SCAN_IN
i P1_INSTADDRPOINTER_REG_5__SCAN_IN
i P1_INSTADDRPOINTER_REG_4__SCAN_IN
i P1_INSTADDRPOINTER_REG_3__SCAN_IN
i P1_INSTADDRPOINTER_REG_2__SCAN_IN
i P1_INSTADDRPOINTER_REG_1__SCAN_IN
i P1_INSTADDRPOINTER_REG_0__SCAN_IN
i P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN
i P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN
i P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN
i P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN
i P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN
i P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN
i P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN
i P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN
i P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN
i P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN
i P1_INSTQUEUE_REG_0__0__SCAN_IN
i P1_INSTQUEUE_REG_0__1__SCAN_IN
i P1_INSTQUEUE_REG_0__2__SCAN_IN
i P1_INSTQUEUE_REG_0__3__SCAN_IN
i P1_INSTQUEUE_REG_0__4__SCAN_IN
i P1_INSTQUEUE_REG_0__5__SCAN_IN
i P1_INSTQUEUE_REG_0__6__SCAN_IN
i P1_INSTQUEUE_REG_0__7__SCAN_IN
i P1_INSTQUEUE_REG_1__0__SCAN_IN
i P1_INSTQUEUE_REG_1__1__SCAN_IN
i P1_INSTQUEUE_REG_1__2__SCAN_IN
i P1_INSTQUEUE_REG_1__3__SCAN_IN
i P1_INSTQUEUE_REG_1__4__SCAN_IN
i P1_INSTQUEUE_REG_1__5__SCAN_IN
i P1_INSTQUEUE_REG_1__6__SCAN_IN
i P1_INSTQUEUE_REG_1__7__SCAN_IN
i P1_INSTQUEUE_REG_2__0__SCAN_IN
i P1_INSTQUEUE_REG_2__1__SCAN_IN
i P1_INSTQUEUE_REG_2__2__SCAN_IN
i P1_INSTQUEUE_REG_2__3__SCAN_IN
i P1_INSTQUEUE_REG_2__4__SCAN_IN
i P1_INSTQUEUE_REG_2__5__SCAN_IN
i P1_INSTQUEUE_REG_2__6__SCAN_IN
i P1_INSTQUEUE_REG_2__7__SCAN_IN
i P1_INSTQUEUE_REG_3__0__SCAN_IN
i P1_INSTQUEUE_REG_3__1__SCAN_IN
i P1_INSTQUEUE_REG_3__2__SCAN_IN
i P1_INSTQUEUE_REG_3__3__SCAN_IN
i P1_INSTQUEUE_REG_3__4__SCAN_IN
i P1_INSTQUEUE_REG_3__5__SCAN_IN
i P1_INSTQUEUE_REG_3__6__SCAN_IN
i P1_INSTQUEUE_REG_3__7__SCAN_IN
i P1_INSTQUEUE_REG_4__0__SCAN_IN
i BUF1_REG_0__SCAN_IN
i BUF1_REG_1__SCAN_IN
i BUF1_REG_2__SCAN_IN
i BUF1_REG_3__SCAN_IN
i BUF1_REG_4__SCAN_IN
i BUF1_REG_5__SCAN_IN
i BUF1_REG_6__SCAN_IN
i BUF1_REG_7__SCAN_IN
i BUF1_REG_8__SCAN_IN
i BUF1_REG_9__SCAN_IN
i BUF1_REG_10__SCAN_IN
i BUF1_REG_11__SCAN_IN
i BUF1_REG_12__SCAN_IN
i BUF1_REG_13__SCAN_IN
i BUF1_REG_14__SCAN_IN
i BUF1_REG_15__SCAN_IN
i BUF1_REG_16__SCAN_IN
i BUF1_REG_17__SCAN_IN
i BUF1_REG_18__SCAN_IN
i BUF1_REG_19__SCAN_IN
i BUF1_REG_20__SCAN_IN
i BUF1_REG_21__SCAN_IN
i BUF1_REG_22__SCAN_IN
i BUF1_REG_23__SCAN_IN
i BUF1_REG_24__SCAN_IN
i BUF1_REG_25__SCAN_IN
i BUF1_REG_26__SCAN_IN
i BUF1_REG_27__SCAN_IN
i BUF1_REG_28__SCAN_IN
i BUF1_REG_29__SCAN_IN
i BUF1_REG_30__SCAN_IN
i BUF1_REG_31__SCAN_IN
i BUF2_REG_0__SCAN_IN
i BUF2_REG_1__SCAN_IN
i BUF2_REG_2__SCAN_IN
i BUF2_REG_3__SCAN_IN
i BUF2_REG_4__SCAN_IN
i BUF2_REG_5__SCAN_IN
i BUF2_REG_6__SCAN_IN
i BUF2_REG_7__SCAN_IN
i BUF2_REG_8__SCAN_IN
i BUF2_REG_9__SCAN_IN
i BUF2_REG_10__SCAN_IN
i BUF2_REG_11__SCAN_IN
i BUF2_REG_12__SCAN_IN
i BUF2_REG_13__SCAN_IN
i BUF2_REG_14__SCAN_IN
i BUF2_REG_15__SCAN_IN
i BUF2_REG_16__SCAN_IN
i BUF2_REG_17__SCAN_IN
i BUF2_REG_18__SCAN_IN
i BUF2_REG_19__SCAN_IN
i BUF2_REG_20__SCAN_IN
i BUF2_REG_21__SCAN_IN
i BUF2_REG_22__SCAN_IN
i BUF2_REG_23__SCAN_IN
i BUF2_REG_24__SCAN_IN
i BUF2_REG_25__SCAN_IN
i BUF2_REG_26__SCAN_IN
i BUF2_REG_27__SCAN_IN
i BUF2_REG_28__SCAN_IN
i BUF2_REG_29__SCAN_IN
i BUF2_REG_30__SCAN_IN
i BUF2_REG_31__SCAN_IN
i READY12_REG_SCAN_IN
i READY21_REG_SCAN_IN
i READY22_REG_SCAN_IN
i READY11_REG_SCAN_IN
i P3_BE_N_REG_3__SCAN_IN
i P3_BE_N_REG_2__SCAN_IN
i P3_BE_N_REG_1__SCAN_IN
i P3_BE_N_REG_0__SCAN_IN
i P3_ADDRESS_REG_29__SCAN_IN
i P3_ADDRESS_REG_28__SCAN_IN
i P3_ADDRESS_REG_27__SCAN_IN
i P3_ADDRESS_REG_26__SCAN_IN
i P3_ADDRESS_REG_25__SCAN_IN
i P3_ADDRESS_REG_24__SCAN_IN
i P3_ADDRESS_REG_23__SCAN_IN
i P3_ADDRESS_REG_22__SCAN_IN
i P3_ADDRESS_REG_21__SCAN_IN
i P3_ADDRESS_REG_20__SCAN_IN
i P3_ADDRESS_REG_19__SCAN_IN
i P3_ADDRESS_REG_18__SCAN_IN
i P3_ADDRESS_REG_17__SCAN_IN
i P3_ADDRESS_REG_16__SCAN_IN
i P3_ADDRESS_REG_15__SCAN_IN
i P3_ADDRESS_REG_14__SCAN_IN
i P3_ADDRESS_REG_13__SCAN_IN
i P3_ADDRESS_REG_12__SCAN_IN
i P3_ADDRESS_REG_11__SCAN_IN
i P3_ADDRESS_REG_10__SCAN_IN
i P3_ADDRESS_REG_9__SCAN_IN
i P3_ADDRESS_REG_8__SCAN_IN
i P3_ADDRESS_REG_7__SCAN_IN
i P3_ADDRESS_REG_6__SCAN_IN
i P3_ADDRESS_REG_5__SCAN_IN
i P3_ADDRESS_REG_4__SCAN_IN
i P3_ADDRESS_REG_3__SCAN_IN
i P3_ADDRESS_REG_2__SCAN_IN
i P3_ADDRESS_REG_1__SCAN_IN
i P3_ADDRESS_REG_0__SCAN_IN
i P3_STATE_REG_2__SCAN_IN
i P3_STATE_REG_1__SCAN_IN
i P3_STATE_REG_0__SCAN_IN
i P3_DATAWIDTH_REG_0__SCAN_IN
i P3_DATAWIDTH_REG_1__SCAN_IN
i P3_DATAWIDTH_REG_2__SCAN_IN
i P3_DATAWIDTH_REG_3__SCAN_IN
i P3_DATAWIDTH_REG_4__SCAN_IN
i P3_DATAWIDTH_REG_5__SCAN_IN
i P3_DATAWIDTH_REG_6__SCAN_IN
i P3_DATAWIDTH_REG_7__SCAN_IN
i P3_DATAWIDTH_REG_8__SCAN_IN
i P3_DATAWIDTH_REG_9__SCAN_IN
i P3_DATAWIDTH_REG_10__SCAN_IN
i P3_DATAWIDTH_REG_11__SCAN_IN
i P3_DATAWIDTH_REG_12__SCAN_IN
i P3_DATAWIDTH_REG_13__SCAN_IN
i P3_DATAWIDTH_REG_14__SCAN_IN
i P3_DATAWIDTH_REG_15__SCAN_IN
i P3_DATAWIDTH_REG_16__SCAN_IN
i P3_DATAWIDTH_REG_17__SCAN_IN
i P3_DATAWIDTH_REG_18__SCAN_IN
i P3_DATAWIDTH_REG_19__SCAN_IN
i P3_DATAWIDTH_REG_20__SCAN_IN
i P3_DATAWIDTH_REG_21__SCAN_IN
i P3_DATAWIDTH_REG_22__SCAN_IN
i P3_DATAWIDTH_REG_23__SCAN_IN
i P3_DATAWIDTH_REG_24__SCAN_IN
i P3_DATAWIDTH_REG_25__SCAN_IN
i P3_DATAWIDTH_REG_26__SCAN_IN
i P3_DATAWIDTH_REG_27__SCAN_IN
i P3_DATAWIDTH_REG_28__SCAN_IN
i P3_DATAWIDTH_REG_29__SCAN_IN
i P3_DATAWIDTH_REG_30__SCAN_IN
i P3_DATAWIDTH_REG_31__SCAN_IN
i P3_STATE2_REG_3__SCAN_IN
i P3_STATE2_REG_2__SCAN_IN
i P3_STATE2_REG_1__SCAN_IN
i P3_STATE2_REG_0__SCAN_IN
i P3_INSTQUEUE_REG_15__7__SCAN_IN
i P3_INSTQUEUE_REG_15__6__SCAN_IN
i P3_INSTQUEUE_REG_15__5__SCAN_IN
i P3_INSTQUEUE_REG_15__4__SCAN_IN
i P3_INSTQUEUE_REG_15__3__SCAN_IN
i P3_INSTQUEUE_REG_15__2__SCAN_IN
i P3_INSTQUEUE_REG_15__1__SCAN_IN
i P3_INSTQUEUE_REG_15__0__SCAN_IN
i P3_INSTQUEUE_REG_14__7__SCAN_IN
i P3_INSTQUEUE_REG_14__6__SCAN_IN
i P3_INSTQUEUE_REG_14__5__SCAN_IN
i P3_INSTQUEUE_REG_14__4__SCAN_IN
i P3_INSTQUEUE_REG_14__3__SCAN_IN
i P3_INSTQUEUE_REG_14__2__SCAN_IN
i P3_INSTQUEUE_REG_14__1__SCAN_IN
i P3_INSTQUEUE_REG_14__0__SCAN_IN
i P3_INSTQUEUE_REG_13__7__SCAN_IN
i P3_INSTQUEUE_REG_13__6__SCAN_IN
i P3_INSTQUEUE_REG_13__5__SCAN_IN
i P3_INSTQUEUE_REG_13__4__SCAN_IN
i P3_INSTQUEUE_REG_13__3__SCAN_IN
i P3_INSTQUEUE_REG_13__2__SCAN_IN
i P3_INSTQUEUE_REG_13__1__SCAN_IN
i P3_INSTQUEUE_REG_13__0__SCAN_IN
i P3_INSTQUEUE_REG_12__7__SCAN_IN
i P3_INSTQUEUE_REG_12__6__SCAN_IN
i P3_INSTQUEUE_REG_12__5__SCAN_IN
i P3_INSTQUEUE_REG_12__4__SCAN_IN
i P3_INSTQUEUE_REG_12__3__SCAN_IN
i P3_INSTQUEUE_REG_12__2__SCAN_IN
i P3_INSTQUEUE_REG_12__1__SCAN_IN
i P3_INSTQUEUE_REG_12__0__SCAN_IN
i P3_INSTQUEUE_REG_11__7__SCAN_IN
i P3_INSTQUEUE_REG_11__6__SCAN_IN
i P3_INSTQUEUE_REG_11__5__SCAN_IN
i P3_INSTQUEUE_REG_11__4__SCAN_IN
i P3_INSTQUEUE_REG_11__3__SCAN_IN
i P3_INSTQUEUE_REG_11__2__SCAN_IN
i P3_INSTQUEUE_REG_11__1__SCAN_IN
i P3_INSTQUEUE_REG_11__0__SCAN_IN
i P3_INSTQUEUE_REG_10__7__SCAN_IN
i P3_INSTQUEUE_REG_10__6__SCAN_IN
i P3_INSTQUEUE_REG_10__5__SCAN_IN
i P3_INSTQUEUE_REG_10__4__SCAN_IN
i P3_INSTQUEUE_REG_10__3__SCAN_IN
i P3_INSTQUEUE_REG_10__2__SCAN_IN
i P3_INSTQUEUE_REG_10__1__SCAN_IN
i P3_INSTQUEUE_REG_10__0__SCAN_IN
i P3_INSTQUEUE_REG_9__7__SCAN_IN
i P3_INSTQUEUE_REG_9__6__SCAN_IN
i P3_INSTQUEUE_REG_9__5__SCAN_IN
i P3_INSTQUEUE_REG_9__4__SCAN_IN
i P3_INSTQUEUE_REG_9__3__SCAN_IN
i P3_INSTQUEUE_REG_9__2__SCAN_IN
i P3_INSTQUEUE_REG_9__1__SCAN_IN
i P3_INSTQUEUE_REG_9__0__SCAN_IN
i P3_INSTQUEUE_REG_8__7__SCAN_IN
i P3_INSTQUEUE_REG_8__6__SCAN_IN
i P3_INSTQUEUE_REG_8__5__SCAN_IN
i P3_INSTQUEUE_REG_8__4__SCAN_IN
i P3_INSTQUEUE_REG_8__3__SCAN_IN
i P3_INSTQUEUE_REG_8__2__SCAN_IN
i P3_INSTQUEUE_REG_8__1__SCAN_IN
i P3_INSTQUEUE_REG_8__0__SCAN_IN
i P3_INSTQUEUE_REG_7__7__SCAN_IN
i P3_INSTQUEUE_REG_7__6__SCAN_IN
i P3_INSTQUEUE_REG_7__5__SCAN_IN
i P3_INSTQUEUE_REG_7__4__SCAN_IN
i P3_INSTQUEUE_REG_7__3__SCAN_IN
i P3_INSTQUEUE_REG_7__2__SCAN_IN
i P3_INSTQUEUE_REG_7__1__SCAN_IN
i P3_INSTQUEUE_REG_7__0__SCAN_IN
i P3_INSTQUEUE_REG_6__7__SCAN_IN
i P3_INSTQUEUE_REG_6__6__SCAN_IN
i P3_INSTQUEUE_REG_6__5__SCAN_IN
i P3_INSTQUEUE_REG_6__4__SCAN_IN
i P3_INSTQUEUE_REG_6__3__SCAN_IN
i P3_INSTQUEUE_REG_6__2__SCAN_IN
i P3_INSTQUEUE_REG_6__1__SCAN_IN
i P3_INSTQUEUE_REG_6__0__SCAN_IN
i P3_INSTQUEUE_REG_5__7__SCAN_IN
i P3_INSTQUEUE_REG_5__6__SCAN_IN
i P3_INSTQUEUE_REG_5__5__SCAN_IN
i P3_INSTQUEUE_REG_5__4__SCAN_IN
i P3_INSTQUEUE_REG_5__3__SCAN_IN
i P3_INSTQUEUE_REG_5__2__SCAN_IN
i P3_INSTQUEUE_REG_5__1__SCAN_IN
i P3_INSTQUEUE_REG_5__0__SCAN_IN
i P3_INSTQUEUE_REG_4__7__SCAN_IN
i P3_INSTQUEUE_REG_4__6__SCAN_IN
i P3_INSTQUEUE_REG_4__5__SCAN_IN
i P3_INSTQUEUE_REG_4__4__SCAN_IN
i P3_INSTQUEUE_REG_4__3__SCAN_IN
i P3_INSTQUEUE_REG_4__2__SCAN_IN
i P3_INSTQUEUE_REG_4__1__SCAN_IN
i P3_INSTQUEUE_REG_4__0__SCAN_IN
i P3_INSTQUEUE_REG_3__7__SCAN_IN
i P3_INSTQUEUE_REG_3__6__SCAN_IN
i P3_INSTQUEUE_REG_3__5__SCAN_IN
i P3_INSTQUEUE_REG_3__4__SCAN_IN
i P3_INSTQUEUE_REG_3__3__SCAN_IN
i P3_INSTQUEUE_REG_3__2__SCAN_IN
i P3_INSTQUEUE_REG_3__1__SCAN_IN
i P3_INSTQUEUE_REG_3__0__SCAN_IN
i P3_INSTQUEUE_REG_2__7__SCAN_IN
i P3_INSTQUEUE_REG_2__6__SCAN_IN
i P3_INSTQUEUE_REG_2__5__SCAN_IN
i P3_INSTQUEUE_REG_2__4__SCAN_IN
i P3_INSTQUEUE_REG_2__3__SCAN_IN
i P3_INSTQUEUE_REG_2__2__SCAN_IN
i P3_INSTQUEUE_REG_2__1__SCAN_IN
i P3_INSTQUEUE_REG_2__0__SCAN_IN
i P3_INSTQUEUE_REG_1__7__SCAN_IN
i P3_INSTQUEUE_REG_1__6__SCAN_IN
i P3_INSTQUEUE_REG_1__5__SCAN_IN
i P3_INSTQUEUE_REG_1__4__SCAN_IN
i P3_INSTQUEUE_REG_1__3__SCAN_IN
i P3_INSTQUEUE_REG_1__2__SCAN_IN
i P3_INSTQUEUE_REG_1__1__SCAN_IN
i P3_INSTQUEUE_REG_1__0__SCAN_IN
i P3_INSTQUEUE_REG_0__7__SCAN_IN
i P3_INSTQUEUE_REG_0__6__SCAN_IN
i P3_INSTQUEUE_REG_0__5__SCAN_IN
i P3_INSTQUEUE_REG_0__4__SCAN_IN
i P3_INSTQUEUE_REG_0__3__SCAN_IN
i P3_INSTQUEUE_REG_0__2__SCAN_IN
i P3_INSTQUEUE_REG_0__1__SCAN_IN
i P3_INSTQUEUE_REG_0__0__SCAN_IN
i P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN
i P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN
i P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN
i P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN
i P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN
i P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN
i P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN
i P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN
i P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN
i P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN
i P3_INSTADDRPOINTER_REG_0__SCAN_IN
i P3_INSTADDRPOINTER_REG_1__SCAN_IN
i P3_INSTADDRPOINTER_REG_2__SCAN_IN
i P3_INSTADDRPOINTER_REG_3__SCAN_IN
i P3_INSTADDRPOINTER_REG_4__SCAN_IN
i P3_INSTADDRPOINTER_REG_5__SCAN_IN
i P3_INSTADDRPOINTER_REG_6__SCAN_IN
i P3_INSTADDRPOINTER_REG_7__SCAN_IN
i P3_INSTADDRPOINTER_REG_8__SCAN_IN
i P3_INSTADDRPOINTER_REG_9__SCAN_IN
i P3_INSTADDRPOINTER_REG_10__SCAN_IN
i P3_INSTADDRPOINTER_REG_11__SCAN_IN
i P3_INSTADDRPOINTER_REG_12__SCAN_IN
i P3_INSTADDRPOINTER_REG_13__SCAN_IN
i P3_INSTADDRPOINTER_REG_14__SCAN_IN
i P3_INSTADDRPOINTER_REG_15__SCAN_IN
i P3_INSTADDRPOINTER_REG_16__SCAN_IN
i P3_INSTADDRPOINTER_REG_17__SCAN_IN
i P3_INSTADDRPOINTER_REG_18__SCAN_IN
i P3_INSTADDRPOINTER_REG_19__SCAN_IN
i P3_INSTADDRPOINTER_REG_20__SCAN_IN
i P3_INSTADDRPOINTER_REG_21__SCAN_IN
i P3_INSTADDRPOINTER_REG_22__SCAN_IN
i P3_INSTADDRPOINTER_REG_23__SCAN_IN
i P3_INSTADDRPOINTER_REG_24__SCAN_IN
i P3_INSTADDRPOINTER_REG_25__SCAN_IN
i P3_INSTADDRPOINTER_REG_26__SCAN_IN
i P3_INSTADDRPOINTER_REG_27__SCAN_IN
i P3_INSTADDRPOINTER_REG_28__SCAN_IN
i P3_INSTADDRPOINTER_REG_29__SCAN_IN
i P3_INSTADDRPOINTER_REG_30__SCAN_IN
i P3_INSTADDRPOINTER_REG_31__SCAN_IN
i P3_PHYADDRPOINTER_REG_0__SCAN_IN
i P3_PHYADDRPOINTER_REG_1__SCAN_IN
i P3_PHYADDRPOINTER_REG_2__SCAN_IN
i P3_PHYADDRPOINTER_REG_3__SCAN_IN
i P3_PHYADDRPOINTER_REG_4__SCAN_IN
i P3_PHYADDRPOINTER_REG_5__SCAN_IN
i P3_PHYADDRPOINTER_REG_6__SCAN_IN
i P3_PHYADDRPOINTER_REG_7__SCAN_IN
i P3_PHYADDRPOINTER_REG_8__SCAN_IN
i P3_PHYADDRPOINTER_REG_9__SCAN_IN
i P3_PHYADDRPOINTER_REG_10__SCAN_IN
i P3_PHYADDRPOINTER_REG_11__SCAN_IN
i P3_PHYADDRPOINTER_REG_12__SCAN_IN
i P3_PHYADDRPOINTER_REG_13__SCAN_IN
i P3_PHYADDRPOINTER_REG_14__SCAN_IN
i P3_PHYADDRPOINTER_REG_15__SCAN_IN
i P3_PHYADDRPOINTER_REG_16__SCAN_IN
i P3_PHYADDRPOINTER_REG_17__SCAN_IN
i P3_PHYADDRPOINTER_REG_18__SCAN_IN
i P3_PHYADDRPOINTER_REG_19__SCAN_IN
i P3_PHYADDRPOINTER_REG_20__SCAN_IN
i P3_PHYADDRPOINTER_REG_21__SCAN_IN
i P3_PHYADDRPOINTER_REG_22__SCAN_IN
i P3_PHYADDRPOINTER_REG_23__SCAN_IN
i P3_PHYADDRPOINTER_REG_24__SCAN_IN
i P3_PHYADDRPOINTER_REG_25__SCAN_IN
i P3_PHYADDRPOINTER_REG_26__SCAN_IN
i P3_PHYADDRPOINTER_REG_27__SCAN_IN
i P3_PHYADDRPOINTER_REG_28__SCAN_IN
i P3_PHYADDRPOINTER_REG_29__SCAN_IN
i P3_PHYADDRPOINTER_REG_30__SCAN_IN
i P3_PHYADDRPOINTER_REG_31__SCAN_IN
i P3_LWORD_REG_15__SCAN_IN
i P3_LWORD_REG_14__SCAN_IN
i P3_LWORD_REG_13__SCAN_IN
i P3_LWORD_REG_12__SCAN_IN
i P3_LWORD_REG_11__SCAN_IN
i P3_LWORD_REG_10__SCAN_IN
i P3_LWORD_REG_9__SCAN_IN
i P3_LWORD_REG_8__SCAN_IN
i P3_LWORD_REG_7__SCAN_IN
i P3_LWORD_REG_6__SCAN_IN
i P3_LWORD_REG_5__SCAN_IN
i P3_LWORD_REG_4__SCAN_IN
i P3_LWORD_REG_3__SCAN_IN
i P3_LWORD_REG_2__SCAN_IN
i P3_LWORD_REG_1__SCAN_IN
i P3_LWORD_REG_0__SCAN_IN
i P3_UWORD_REG_14__SCAN_IN
i P3_UWORD_REG_13__SCAN_IN
i P3_UWORD_REG_12__SCAN_IN
i P3_UWORD_REG_11__SCAN_IN
i P3_UWORD_REG_10__SCAN_IN
i P3_UWORD_REG_9__SCAN_IN
i P3_UWORD_REG_8__SCAN_IN
i P3_UWORD_REG_7__SCAN_IN
i P3_UWORD_REG_6__SCAN_IN
i P3_UWORD_REG_5__SCAN_IN
i P3_UWORD_REG_4__SCAN_IN
i P3_UWORD_REG_3__SCAN_IN
i P3_UWORD_REG_2__SCAN_IN
i P3_UWORD_REG_1__SCAN_IN
i P3_UWORD_REG_0__SCAN_IN
i P3_DATAO_REG_0__SCAN_IN
i P3_DATAO_REG_1__SCAN_IN
i P3_DATAO_REG_2__SCAN_IN
i P3_DATAO_REG_3__SCAN_IN
i P3_DATAO_REG_4__SCAN_IN
i P3_DATAO_REG_5__SCAN_IN
i P3_DATAO_REG_6__SCAN_IN
i P3_DATAO_REG_7__SCAN_IN
i P3_DATAO_REG_8__SCAN_IN
i P3_DATAO_REG_9__SCAN_IN
i P3_DATAO_REG_10__SCAN_IN
i P3_DATAO_REG_11__SCAN_IN
i P3_DATAO_REG_12__SCAN_IN
i P3_DATAO_REG_13__SCAN_IN
i P3_DATAO_REG_14__SCAN_IN
i P3_DATAO_REG_15__SCAN_IN
i P3_DATAO_REG_16__SCAN_IN
i P3_DATAO_REG_17__SCAN_IN
i P3_DATAO_REG_18__SCAN_IN
i P3_DATAO_REG_19__SCAN_IN
i P3_DATAO_REG_20__SCAN_IN
i P3_DATAO_REG_21__SCAN_IN
i P3_DATAO_REG_22__SCAN_IN
i P3_DATAO_REG_23__SCAN_IN
i P3_DATAO_REG_24__SCAN_IN
i P3_DATAO_REG_25__SCAN_IN
i P3_DATAO_REG_26__SCAN_IN
i P3_DATAO_REG_27__SCAN_IN
i P3_DATAO_REG_28__SCAN_IN
i P3_DATAO_REG_29__SCAN_IN
i P3_DATAO_REG_30__SCAN_IN
i P3_DATAO_REG_31__SCAN_IN
i P3_EAX_REG_0__SCAN_IN
i P3_EAX_REG_1__SCAN_IN
i P3_EAX_REG_2__SCAN_IN
i P3_EAX_REG_3__SCAN_IN
i P3_EAX_REG_4__SCAN_IN
i P3_EAX_REG_5__SCAN_IN
i P3_EAX_REG_6__SCAN_IN
i P3_EAX_REG_7__SCAN_IN
i P3_EAX_REG_8__SCAN_IN
i P3_EAX_REG_9__SCAN_IN
i P3_EAX_REG_10__SCAN_IN
i P3_EAX_REG_11__SCAN_IN
i P3_EAX_REG_12__SCAN_IN
i P3_EAX_REG_13__SCAN_IN
i P3_EAX_REG_14__SCAN_IN
i P3_EAX_REG_15__SCAN_IN
i P3_EAX_REG_16__SCAN_IN
i P3_EAX_REG_17__SCAN_IN
i P3_EAX_REG_18__SCAN_IN
i P3_EAX_REG_19__SCAN_IN
i P3_EAX_REG_20__SCAN_IN
i P3_EAX_REG_21__SCAN_IN
i P3_EAX_REG_22__SCAN_IN
i P3_EAX_REG_23__SCAN_IN
i P3_EAX_REG_24__SCAN_IN
i P3_EAX_REG_25__SCAN_IN
i P3_EAX_REG_26__SCAN_IN
i P3_EAX_REG_27__SCAN_IN
i P3_EAX_REG_28__SCAN_IN
i P3_EAX_REG_29__SCAN_IN
i P3_EAX_REG_30__SCAN_IN
i P3_EAX_REG_31__SCAN_IN
i P3_EBX_REG_0__SCAN_IN
i P3_EBX_REG_1__SCAN_IN
i P3_EBX_REG_2__SCAN_IN
i P3_EBX_REG_3__SCAN_IN
i P3_EBX_REG_4__SCAN_IN
i P3_EBX_REG_5__SCAN_IN
i P3_EBX_REG_6__SCAN_IN
i P3_EBX_REG_7__SCAN_IN
i P3_EBX_REG_8__SCAN_IN
i P3_EBX_REG_9__SCAN_IN
i P3_EBX_REG_10__SCAN_IN
i P3_EBX_REG_11__SCAN_IN
i P3_EBX_REG_12__SCAN_IN
i P3_EBX_REG_13__SCAN_IN
i P3_EBX_REG_14__SCAN_IN
i P3_EBX_REG_15__SCAN_IN
i P3_EBX_REG_16__SCAN_IN
i P3_EBX_REG_17__SCAN_IN
i P3_EBX_REG_18__SCAN_IN
i P3_EBX_REG_19__SCAN_IN
i P3_EBX_REG_20__SCAN_IN
i P3_EBX_REG_21__SCAN_IN
i P3_EBX_REG_22__SCAN_IN
i P3_EBX_REG_23__SCAN_IN
i P3_EBX_REG_24__SCAN_IN
i P3_EBX_REG_25__SCAN_IN
i P3_EBX_REG_26__SCAN_IN
i P3_EBX_REG_27__SCAN_IN
i P3_EBX_REG_28__SCAN_IN
i P3_EBX_REG_29__SCAN_IN
i P3_EBX_REG_30__SCAN_IN
i P3_EBX_REG_31__SCAN_IN
i P3_REIP_REG_0__SCAN_IN
i P3_REIP_REG_1__SCAN_IN
i P3_REIP_REG_2__SCAN_IN
i P3_REIP_REG_3__SCAN_IN
i P3_REIP_REG_4__SCAN_IN
i P3_REIP_REG_5__SCAN_IN
i P3_REIP_REG_6__SCAN_IN
i P3_REIP_REG_7__SCAN_IN
i P3_REIP_REG_8__SCAN_IN
i P3_REIP_REG_9__SCAN_IN
i P3_REIP_REG_10__SCAN_IN
i P3_REIP_REG_11__SCAN_IN
i P3_REIP_REG_12__SCAN_IN
i P3_REIP_REG_13__SCAN_IN
i P3_REIP_REG_14__SCAN_IN
i P3_REIP_REG_15__SCAN_IN
i P3_REIP_REG_16__SCAN_IN
i P3_REIP_REG_17__SCAN_IN
i P3_REIP_REG_18__SCAN_IN
i P3_REIP_REG_19__SCAN_IN
i P3_REIP_REG_20__SCAN_IN
i P3_REIP_REG_21__SCAN_IN
i P3_REIP_REG_22__SCAN_IN
i P3_REIP_REG_23__SCAN_IN
i P3_REIP_REG_24__SCAN_IN
i P3_REIP_REG_25__SCAN_IN
i P3_REIP_REG_26__SCAN_IN
i P3_REIP_REG_27__SCAN_IN
i P3_REIP_REG_28__SCAN_IN
i P3_REIP_REG_29__SCAN_IN
i P3_REIP_REG_30__SCAN_IN
i P3_REIP_REG_31__SCAN_IN
i P3_BYTEENABLE_REG_3__SCAN_IN
i P3_BYTEENABLE_REG_2__SCAN_IN
i P3_BYTEENABLE_REG_1__SCAN_IN
i P3_BYTEENABLE_REG_0__SCAN_IN
i P3_W_R_N_REG_SCAN_IN
i P3_FLUSH_REG_SCAN_IN
i P3_MORE_REG_SCAN_IN
i P3_STATEBS16_REG_SCAN_IN
i P3_REQUESTPENDING_REG_SCAN_IN
i P3_D_C_N_REG_SCAN_IN
i P3_M_IO_N_REG_SCAN_IN
i P3_CODEFETCH_REG_SCAN_IN
i P3_ADS_N_REG_SCAN_IN
i P3_READREQUEST_REG_SCAN_IN
i P3_MEMORYFETCH_REG_SCAN_IN
i P2_BE_N_REG_3__SCAN_IN
i P2_BE_N_REG_2__SCAN_IN
i P2_BE_N_REG_1__SCAN_IN
i P2_BE_N_REG_0__SCAN_IN
i P2_ADDRESS_REG_29__SCAN_IN
i P2_ADDRESS_REG_28__SCAN_IN
i P2_ADDRESS_REG_27__SCAN_IN
i P2_ADDRESS_REG_26__SCAN_IN
i P2_ADDRESS_REG_25__SCAN_IN
i P2_ADDRESS_REG_24__SCAN_IN
i P2_ADDRESS_REG_23__SCAN_IN
i P2_ADDRESS_REG_22__SCAN_IN
i P2_ADDRESS_REG_21__SCAN_IN
i P2_ADDRESS_REG_20__SCAN_IN
i P2_ADDRESS_REG_19__SCAN_IN
i P2_ADDRESS_REG_18__SCAN_IN
i P2_ADDRESS_REG_17__SCAN_IN
i P2_ADDRESS_REG_16__SCAN_IN
i P2_ADDRESS_REG_15__SCAN_IN
i P2_ADDRESS_REG_14__SCAN_IN
i P2_ADDRESS_REG_13__SCAN_IN
i P2_ADDRESS_REG_12__SCAN_IN
i P2_ADDRESS_REG_11__SCAN_IN
i P2_ADDRESS_REG_10__SCAN_IN
i P2_ADDRESS_REG_9__SCAN_IN
i P2_ADDRESS_REG_8__SCAN_IN
i P2_ADDRESS_REG_7__SCAN_IN
i P2_ADDRESS_REG_6__SCAN_IN
i P2_ADDRESS_REG_5__SCAN_IN
i P2_ADDRESS_REG_4__SCAN_IN
i P2_ADDRESS_REG_3__SCAN_IN
i P2_ADDRESS_REG_2__SCAN_IN
i P2_ADDRESS_REG_1__SCAN_IN
i P2_ADDRESS_REG_0__SCAN_IN
i P2_STATE_REG_2__SCAN_IN
i P2_STATE_REG_1__SCAN_IN
i P2_STATE_REG_0__SCAN_IN
i P2_DATAWIDTH_REG_0__SCAN_IN
i P2_DATAWIDTH_REG_1__SCAN_IN
i P2_DATAWIDTH_REG_2__SCAN_IN
i P2_DATAWIDTH_REG_3__SCAN_IN
i P2_DATAWIDTH_REG_4__SCAN_IN
i P2_DATAWIDTH_REG_5__SCAN_IN
i P2_DATAWIDTH_REG_6__SCAN_IN
i P2_DATAWIDTH_REG_7__SCAN_IN
i P2_DATAWIDTH_REG_8__SCAN_IN
i P2_DATAWIDTH_REG_9__SCAN_IN
i P2_DATAWIDTH_REG_10__SCAN_IN
i P2_DATAWIDTH_REG_11__SCAN_IN
i P2_DATAWIDTH_REG_12__SCAN_IN
i P2_DATAWIDTH_REG_13__SCAN_IN
i P2_DATAWIDTH_REG_14__SCAN_IN
i P2_DATAWIDTH_REG_15__SCAN_IN
i P2_DATAWIDTH_REG_16__SCAN_IN
i P2_DATAWIDTH_REG_17__SCAN_IN
i P2_DATAWIDTH_REG_18__SCAN_IN
i P2_DATAWIDTH_REG_19__SCAN_IN
i P2_DATAWIDTH_REG_20__SCAN_IN
i P2_DATAWIDTH_REG_21__SCAN_IN
i P2_DATAWIDTH_REG_22__SCAN_IN
i P2_DATAWIDTH_REG_23__SCAN_IN
i P2_DATAWIDTH_REG_24__SCAN_IN
i P2_DATAWIDTH_REG_25__SCAN_IN
i P2_DATAWIDTH_REG_26__SCAN_IN
i P2_DATAWIDTH_REG_27__SCAN_IN
i P2_DATAWIDTH_REG_28__SCAN_IN
i P2_DATAWIDTH_REG_29__SCAN_IN
i P2_DATAWIDTH_REG_30__SCAN_IN
i P2_DATAWIDTH_REG_31__SCAN_IN
i P2_STATE2_REG_3__SCAN_IN
i P2_STATE2_REG_2__SCAN_IN
i P2_STATE2_REG_1__SCAN_IN
i P2_STATE2_REG_0__SCAN_IN
i P2_INSTQUEUE_REG_15__7__SCAN_IN
i P2_INSTQUEUE_REG_15__6__SCAN_IN
i P2_INSTQUEUE_REG_15__5__SCAN_IN
i P2_INSTQUEUE_REG_15__4__SCAN_IN
i P2_INSTQUEUE_REG_15__3__SCAN_IN
i P2_INSTQUEUE_REG_15__2__SCAN_IN
i P2_INSTQUEUE_REG_15__1__SCAN_IN
i P2_INSTQUEUE_REG_15__0__SCAN_IN
i P2_INSTQUEUE_REG_14__7__SCAN_IN
i P2_INSTQUEUE_REG_14__6__SCAN_IN
i P2_INSTQUEUE_REG_14__5__SCAN_IN
i P2_INSTQUEUE_REG_14__4__SCAN_IN
i P2_INSTQUEUE_REG_14__3__SCAN_IN
i P2_INSTQUEUE_REG_14__2__SCAN_IN
i P2_INSTQUEUE_REG_14__1__SCAN_IN
i P2_INSTQUEUE_REG_14__0__SCAN_IN
i P2_INSTQUEUE_REG_13__7__SCAN_IN
i P2_INSTQUEUE_REG_13__6__SCAN_IN
i P2_INSTQUEUE_REG_13__5__SCAN_IN
i P2_INSTQUEUE_REG_13__4__SCAN_IN
i P2_INSTQUEUE_REG_13__3__SCAN_IN
i P2_INSTQUEUE_REG_13__2__SCAN_IN
i P2_INSTQUEUE_REG_13__1__SCAN_IN
i P2_INSTQUEUE_REG_13__0__SCAN_IN
i P2_INSTQUEUE_REG_12__7__SCAN_IN
i P2_INSTQUEUE_REG_12__6__SCAN_IN
i P2_INSTQUEUE_REG_12__5__SCAN_IN
i P2_INSTQUEUE_REG_12__4__SCAN_IN
i P2_INSTQUEUE_REG_12__3__SCAN_IN
i P2_INSTQUEUE_REG_12__2__SCAN_IN
i P2_INSTQUEUE_REG_12__1__SCAN_IN
i P2_INSTQUEUE_REG_12__0__SCAN_IN
i P2_INSTQUEUE_REG_11__7__SCAN_IN
i P2_INSTQUEUE_REG_11__6__SCAN_IN
i P2_INSTQUEUE_REG_11__5__SCAN_IN
i P2_INSTQUEUE_REG_11__4__SCAN_IN
i P2_INSTQUEUE_REG_11__3__SCAN_IN
i P2_INSTQUEUE_REG_11__2__SCAN_IN
i P2_INSTQUEUE_REG_11__1__SCAN_IN
i P2_INSTQUEUE_REG_11__0__SCAN_IN
i P2_INSTQUEUE_REG_10__7__SCAN_IN
i P2_INSTQUEUE_REG_10__6__SCAN_IN
i P2_INSTQUEUE_REG_10__5__SCAN_IN
i P2_INSTQUEUE_REG_10__4__SCAN_IN
i P2_INSTQUEUE_REG_10__3__SCAN_IN
i P2_INSTQUEUE_REG_10__2__SCAN_IN
i P2_INSTQUEUE_REG_10__1__SCAN_IN
i P2_INSTQUEUE_REG_10__0__SCAN_IN
i P2_INSTQUEUE_REG_9__7__SCAN_IN
i P2_INSTQUEUE_REG_9__6__SCAN_IN
i P2_INSTQUEUE_REG_9__5__SCAN_IN
i P2_INSTQUEUE_REG_9__4__SCAN_IN
i P2_INSTQUEUE_REG_9__3__SCAN_IN
i P2_INSTQUEUE_REG_9__2__SCAN_IN
i P2_INSTQUEUE_REG_9__1__SCAN_IN
i P2_INSTQUEUE_REG_9__0__SCAN_IN
i P2_INSTQUEUE_REG_8__7__SCAN_IN
i P2_INSTQUEUE_REG_8__6__SCAN_IN
i P2_INSTQUEUE_REG_8__5__SCAN_IN
i P2_INSTQUEUE_REG_8__4__SCAN_IN
i P2_INSTQUEUE_REG_8__3__SCAN_IN
i P2_INSTQUEUE_REG_8__2__SCAN_IN
i P2_INSTQUEUE_REG_8__1__SCAN_IN
i P2_INSTQUEUE_REG_8__0__SCAN_IN
i P2_INSTQUEUE_REG_7__7__SCAN_IN
i P2_INSTQUEUE_REG_7__6__SCAN_IN
i P2_INSTQUEUE_REG_7__5__SCAN_IN
i P2_INSTQUEUE_REG_7__4__SCAN_IN
i P2_INSTQUEUE_REG_7__3__SCAN_IN
i P2_INSTQUEUE_REG_7__2__SCAN_IN
i P2_INSTQUEUE_REG_7__1__SCAN_IN
i P2_INSTQUEUE_REG_7__0__SCAN_IN
i P2_INSTQUEUE_REG_6__7__SCAN_IN
i P2_INSTQUEUE_REG_6__6__SCAN_IN
i P2_INSTQUEUE_REG_6__5__SCAN_IN
i P2_INSTQUEUE_REG_6__4__SCAN_IN
i P2_INSTQUEUE_REG_6__3__SCAN_IN
i P2_INSTQUEUE_REG_6__2__SCAN_IN
i P2_INSTQUEUE_REG_6__1__SCAN_IN
i P2_INSTQUEUE_REG_6__0__SCAN_IN
i P2_INSTQUEUE_REG_5__7__SCAN_IN
i P2_INSTQUEUE_REG_5__6__SCAN_IN
i P2_INSTQUEUE_REG_5__5__SCAN_IN
i P2_INSTQUEUE_REG_5__4__SCAN_IN
i P2_INSTQUEUE_REG_5__3__SCAN_IN
i P2_INSTQUEUE_REG_5__2__SCAN_IN
i P2_INSTQUEUE_REG_5__1__SCAN_IN
i P2_INSTQUEUE_REG_5__0__SCAN_IN
i P2_INSTQUEUE_REG_4__7__SCAN_IN
i P2_INSTQUEUE_REG_4__6__SCAN_IN
i P2_INSTQUEUE_REG_4__5__SCAN_IN
i P2_INSTQUEUE_REG_4__4__SCAN_IN
i P2_INSTQUEUE_REG_4__3__SCAN_IN
i P2_INSTQUEUE_REG_4__2__SCAN_IN
i P2_INSTQUEUE_REG_4__1__SCAN_IN
i P2_INSTQUEUE_REG_4__0__SCAN_IN
i P2_INSTQUEUE_REG_3__7__SCAN_IN
i P2_INSTQUEUE_REG_3__6__SCAN_IN
i P2_INSTQUEUE_REG_3__5__SCAN_IN
i P2_INSTQUEUE_REG_3__4__SCAN_IN
i P2_INSTQUEUE_REG_3__3__SCAN_IN
i P2_INSTQUEUE_REG_3__2__SCAN_IN
i P2_INSTQUEUE_REG_3__1__SCAN_IN
i P2_INSTQUEUE_REG_3__0__SCAN_IN
i P2_INSTQUEUE_REG_2__7__SCAN_IN
i P2_INSTQUEUE_REG_2__6__SCAN_IN
i P2_INSTQUEUE_REG_2__5__SCAN_IN
i P2_INSTQUEUE_REG_2__4__SCAN_IN
i P2_INSTQUEUE_REG_2__3__SCAN_IN
i P2_INSTQUEUE_REG_2__2__SCAN_IN
i P2_INSTQUEUE_REG_2__1__SCAN_IN
i P2_INSTQUEUE_REG_2__0__SCAN_IN
i P2_INSTQUEUE_REG_1__7__SCAN_IN
i P2_INSTQUEUE_REG_1__6__SCAN_IN
i P2_INSTQUEUE_REG_1__5__SCAN_IN
i P2_INSTQUEUE_REG_1__4__SCAN_IN
i P2_INSTQUEUE_REG_1__3__SCAN_IN
i P2_INSTQUEUE_REG_1__2__SCAN_IN
i P2_INSTQUEUE_REG_1__1__SCAN_IN
i P2_INSTQUEUE_REG_1__0__SCAN_IN
i P2_INSTQUEUE_REG_0__7__SCAN_IN
i P2_INSTQUEUE_REG_0__6__SCAN_IN
i P2_INSTQUEUE_REG_0__5__SCAN_IN
i P2_INSTQUEUE_REG_0__4__SCAN_IN
i P2_INSTQUEUE_REG_0__3__SCAN_IN
i P2_INSTQUEUE_REG_0__2__SCAN_IN
i P2_INSTQUEUE_REG_0__1__SCAN_IN
i P2_INSTQUEUE_REG_0__0__SCAN_IN
i P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN
i P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN
i P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN
i P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN
i P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN
i P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN
i P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN
i P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN
i P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN
i P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN
i P2_INSTADDRPOINTER_REG_0__SCAN_IN
i P2_INSTADDRPOINTER_REG_1__SCAN_IN
i P2_INSTADDRPOINTER_REG_2__SCAN_IN
i P2_INSTADDRPOINTER_REG_3__SCAN_IN
i P2_INSTADDRPOINTER_REG_4__SCAN_IN
i P2_INSTADDRPOINTER_REG_5__SCAN_IN
i P2_INSTADDRPOINTER_REG_6__SCAN_IN
i P2_INSTADDRPOINTER_REG_7__SCAN_IN
i P2_INSTADDRPOINTER_REG_8__SCAN_IN
i P2_INSTADDRPOINTER_REG_9__SCAN_IN
i P2_INSTADDRPOINTER_REG_10__SCAN_IN
i P2_INSTADDRPOINTER_REG_11__SCAN_IN
i P2_INSTADDRPOINTER_REG_12__SCAN_IN
i P2_INSTADDRPOINTER_REG_13__SCAN_IN
i P2_INSTADDRPOINTER_REG_14__SCAN_IN
i P2_INSTADDRPOINTER_REG_15__SCAN_IN
i P2_INSTADDRPOINTER_REG_16__SCAN_IN
i P2_INSTADDRPOINTER_REG_17__SCAN_IN
i P2_INSTADDRPOINTER_REG_18__SCAN_IN
i P2_INSTADDRPOINTER_REG_19__SCAN_IN
i P2_INSTADDRPOINTER_REG_20__SCAN_IN
i P2_INSTADDRPOINTER_REG_21__SCAN_IN
i P2_INSTADDRPOINTER_REG_22__SCAN_IN
i P2_INSTADDRPOINTER_REG_23__SCAN_IN
i P2_INSTADDRPOINTER_REG_24__SCAN_IN
i P2_INSTADDRPOINTER_REG_25__SCAN_IN
i P2_INSTADDRPOINTER_REG_26__SCAN_IN
i P2_INSTADDRPOINTER_REG_27__SCAN_IN
i P2_INSTADDRPOINTER_REG_28__SCAN_IN
i P2_INSTADDRPOINTER_REG_29__SCAN_IN
i P2_INSTADDRPOINTER_REG_30__SCAN_IN
i P2_INSTADDRPOINTER_REG_31__SCAN_IN
i P2_PHYADDRPOINTER_REG_0__SCAN_IN
i P2_PHYADDRPOINTER_REG_1__SCAN_IN
i P2_PHYADDRPOINTER_REG_2__SCAN_IN
i P2_PHYADDRPOINTER_REG_3__SCAN_IN
i P2_PHYADDRPOINTER_REG_4__SCAN_IN
i P2_PHYADDRPOINTER_REG_5__SCAN_IN
i P2_PHYADDRPOINTER_REG_6__SCAN_IN
i P2_PHYADDRPOINTER_REG_7__SCAN_IN
i P2_PHYADDRPOINTER_REG_8__SCAN_IN
i P2_PHYADDRPOINTER_REG_9__SCAN_IN
i P2_PHYADDRPOINTER_REG_10__SCAN_IN
i P2_PHYADDRPOINTER_REG_11__SCAN_IN
i P2_PHYADDRPOINTER_REG_12__SCAN_IN
i P2_PHYADDRPOINTER_REG_13__SCAN_IN
i P2_PHYADDRPOINTER_REG_14__SCAN_IN
i P2_PHYADDRPOINTER_REG_15__SCAN_IN
i P2_PHYADDRPOINTER_REG_16__SCAN_IN
i P2_PHYADDRPOINTER_REG_17__SCAN_IN
i P2_PHYADDRPOINTER_REG_18__SCAN_IN
i P2_PHYADDRPOINTER_REG_19__SCAN_IN
i P2_PHYADDRPOINTER_REG_20__SCAN_IN
i P2_PHYADDRPOINTER_REG_21__SCAN_IN
i P2_PHYADDRPOINTER_REG_22__SCAN_IN
i P2_PHYADDRPOINTER_REG_23__SCAN_IN
i P2_PHYADDRPOINTER_REG_24__SCAN_IN
i P2_PHYADDRPOINTER_REG_25__SCAN_IN
i P2_PHYADDRPOINTER_REG_26__SCAN_IN
i P2_PHYADDRPOINTER_REG_27__SCAN_IN
i P2_PHYADDRPOINTER_REG_28__SCAN_IN
i P2_PHYADDRPOINTER_REG_29__SCAN_IN
i P2_PHYADDRPOINTER_REG_30__SCAN_IN
i P2_PHYADDRPOINTER_REG_31__SCAN_IN
i P2_LWORD_REG_15__SCAN_IN
i P2_LWORD_REG_14__SCAN_IN
i P2_LWORD_REG_13__SCAN_IN
i P2_LWORD_REG_12__SCAN_IN
i P2_LWORD_REG_11__SCAN_IN
i P2_LWORD_REG_10__SCAN_IN
i P2_LWORD_REG_9__SCAN_IN
i P2_LWORD_REG_8__SCAN_IN
i P2_LWORD_REG_7__SCAN_IN
i P2_LWORD_REG_6__SCAN_IN
i P2_LWORD_REG_5__SCAN_IN
i P2_LWORD_REG_4__SCAN_IN
i P2_LWORD_REG_3__SCAN_IN
i P2_LWORD_REG_2__SCAN_IN
i P2_LWORD_REG_1__SCAN_IN
i P2_LWORD_REG_0__SCAN_IN
i P2_UWORD_REG_14__SCAN_IN
i P2_UWORD_REG_13__SCAN_IN
i P2_UWORD_REG_12__SCAN_IN
i P2_UWORD_REG_11__SCAN_IN
i P2_UWORD_REG_10__SCAN_IN
i P2_UWORD_REG_9__SCAN_IN
i P2_UWORD_REG_8__SCAN_IN
i P2_UWORD_REG_7__SCAN_IN
i P2_UWORD_REG_6__SCAN_IN
i P2_UWORD_REG_5__SCAN_IN
i P2_UWORD_REG_4__SCAN_IN
i P2_UWORD_REG_3__SCAN_IN
i P2_UWORD_REG_2__SCAN_IN
i P2_UWORD_REG_1__SCAN_IN
i P2_UWORD_REG_0__SCAN_IN
i P2_DATAO_REG_0__SCAN_IN
i P2_DATAO_REG_1__SCAN_IN
i P2_DATAO_REG_2__SCAN_IN
i P2_DATAO_REG_3__SCAN_IN
i P2_DATAO_REG_4__SCAN_IN
i P2_DATAO_REG_5__SCAN_IN
i P2_DATAO_REG_6__SCAN_IN
i P2_DATAO_REG_7__SCAN_IN
i P2_DATAO_REG_8__SCAN_IN
i P2_DATAO_REG_9__SCAN_IN
i P2_DATAO_REG_10__SCAN_IN
i P2_DATAO_REG_11__SCAN_IN
i P2_DATAO_REG_12__SCAN_IN
i P2_DATAO_REG_13__SCAN_IN
i P2_DATAO_REG_14__SCAN_IN
i P2_DATAO_REG_15__SCAN_IN
i P2_DATAO_REG_16__SCAN_IN
i P2_DATAO_REG_17__SCAN_IN
i P2_DATAO_REG_18__SCAN_IN
i P2_DATAO_REG_19__SCAN_IN
i P2_DATAO_REG_20__SCAN_IN
i P2_DATAO_REG_21__SCAN_IN
i P2_DATAO_REG_22__SCAN_IN
i P2_DATAO_REG_23__SCAN_IN
i P2_DATAO_REG_24__SCAN_IN
i P2_DATAO_REG_25__SCAN_IN
i P2_DATAO_REG_26__SCAN_IN
i P2_DATAO_REG_27__SCAN_IN
i P2_DATAO_REG_28__SCAN_IN
i P2_DATAO_REG_29__SCAN_IN
i P2_DATAO_REG_30__SCAN_IN
i P2_DATAO_REG_31__SCAN_IN
i P2_EAX_REG_0__SCAN_IN
i P2_EAX_REG_1__SCAN_IN
i P2_EAX_REG_2__SCAN_IN
i P2_EAX_REG_3__SCAN_IN
i P2_EAX_REG_4__SCAN_IN
i P2_EAX_REG_5__SCAN_IN
i P2_EAX_REG_6__SCAN_IN
i P2_EAX_REG_7__SCAN_IN
i P2_EAX_REG_8__SCAN_IN
i P2_EAX_REG_9__SCAN_IN
i P2_EAX_REG_10__SCAN_IN
i P2_EAX_REG_11__SCAN_IN
i P2_EAX_REG_12__SCAN_IN
i P2_EAX_REG_13__SCAN_IN
i P2_EAX_REG_14__SCAN_IN
i P2_EAX_REG_15__SCAN_IN
i P2_EAX_REG_16__SCAN_IN
i P2_EAX_REG_17__SCAN_IN
i P2_EAX_REG_18__SCAN_IN
i P2_EAX_REG_19__SCAN_IN
i P2_EAX_REG_20__SCAN_IN
i P2_EAX_REG_21__SCAN_IN
i P2_EAX_REG_22__SCAN_IN
i P2_EAX_REG_23__SCAN_IN
i P2_EAX_REG_24__SCAN_IN
i P2_EAX_REG_25__SCAN_IN
i P2_EAX_REG_26__SCAN_IN
i P2_EAX_REG_27__SCAN_IN
i P2_EAX_REG_28__SCAN_IN
i P2_EAX_REG_29__SCAN_IN
i P2_EAX_REG_30__SCAN_IN
i P2_EAX_REG_31__SCAN_IN
i P2_EBX_REG_0__SCAN_IN
i P2_EBX_REG_1__SCAN_IN
i P2_EBX_REG_2__SCAN_IN
i P2_EBX_REG_3__SCAN_IN
i P2_EBX_REG_4__SCAN_IN
i P2_EBX_REG_5__SCAN_IN
i P2_EBX_REG_6__SCAN_IN
i P2_EBX_REG_7__SCAN_IN
i P2_EBX_REG_8__SCAN_IN
i P2_EBX_REG_9__SCAN_IN
i P2_EBX_REG_10__SCAN_IN
i P2_EBX_REG_11__SCAN_IN
i P2_EBX_REG_12__SCAN_IN
i P2_EBX_REG_13__SCAN_IN
i P2_EBX_REG_14__SCAN_IN
i P2_EBX_REG_15__SCAN_IN
i P2_EBX_REG_16__SCAN_IN
i P2_EBX_REG_17__SCAN_IN
i P2_EBX_REG_18__SCAN_IN
i P2_EBX_REG_19__SCAN_IN
i P2_EBX_REG_20__SCAN_IN
i P2_EBX_REG_21__SCAN_IN
i P2_EBX_REG_22__SCAN_IN
i P2_EBX_REG_23__SCAN_IN
i P2_EBX_REG_24__SCAN_IN
i P2_EBX_REG_25__SCAN_IN
i P2_EBX_REG_26__SCAN_IN
i P2_EBX_REG_27__SCAN_IN
i P2_EBX_REG_28__SCAN_IN
i P2_EBX_REG_29__SCAN_IN
i P2_EBX_REG_30__SCAN_IN
i P2_EBX_REG_31__SCAN_IN
i P2_REIP_REG_0__SCAN_IN
i P2_REIP_REG_1__SCAN_IN
i P2_REIP_REG_2__SCAN_IN
i P2_REIP_REG_3__SCAN_IN
i P2_REIP_REG_4__SCAN_IN
i P2_REIP_REG_5__SCAN_IN
i P2_REIP_REG_6__SCAN_IN
i P2_REIP_REG_7__SCAN_IN
i P2_REIP_REG_8__SCAN_IN
i P2_REIP_REG_9__SCAN_IN
i P2_REIP_REG_10__SCAN_IN
i P2_REIP_REG_11__SCAN_IN
i P2_REIP_REG_12__SCAN_IN
i P2_REIP_REG_13__SCAN_IN
i P2_REIP_REG_14__SCAN_IN
i P2_REIP_REG_15__SCAN_IN
i P2_REIP_REG_16__SCAN_IN
i P2_REIP_REG_17__SCAN_IN
i P2_REIP_REG_18__SCAN_IN
i P2_REIP_REG_19__SCAN_IN
i P2_REIP_REG_20__SCAN_IN
i P2_REIP_REG_21__SCAN_IN
i P2_REIP_REG_22__SCAN_IN
i P2_REIP_REG_23__SCAN_IN
i P2_REIP_REG_24__SCAN_IN
i P2_REIP_REG_25__SCAN_IN
i P2_REIP_REG_26__SCAN_IN
i P2_REIP_REG_27__SCAN_IN
i P2_REIP_REG_28__SCAN_IN
i P2_REIP_REG_29__SCAN_IN
i P2_REIP_REG_30__SCAN_IN
i P2_REIP_REG_31__SCAN_IN
i P2_BYTEENABLE_REG_3__SCAN_IN
i P2_BYTEENABLE_REG_2__SCAN_IN
i P2_BYTEENABLE_REG_1__SCAN_IN
i P2_BYTEENABLE_REG_0__SCAN_IN
i P2_W_R_N_REG_SCAN_IN
i P2_FLUSH_REG_SCAN_IN
i P2_MORE_REG_SCAN_IN
i P2_STATEBS16_REG_SCAN_IN
i P2_REQUESTPENDING_REG_SCAN_IN
i P2_D_C_N_REG_SCAN_IN
i P2_M_IO_N_REG_SCAN_IN
i P2_CODEFETCH_REG_SCAN_IN
i P2_ADS_N_REG_SCAN_IN
i P2_READREQUEST_REG_SCAN_IN
i P2_MEMORYFETCH_REG_SCAN_IN
i P1_BE_N_REG_3__SCAN_IN
i P1_BE_N_REG_2__SCAN_IN
i P1_BE_N_REG_1__SCAN_IN
i P1_BE_N_REG_0__SCAN_IN
i P1_ADDRESS_REG_29__SCAN_IN
i P1_ADDRESS_REG_28__SCAN_IN
i P1_ADDRESS_REG_27__SCAN_IN
i P1_ADDRESS_REG_26__SCAN_IN
i P1_ADDRESS_REG_25__SCAN_IN
i P1_ADDRESS_REG_24__SCAN_IN
i P1_ADDRESS_REG_23__SCAN_IN
i P1_ADDRESS_REG_22__SCAN_IN
i P1_ADDRESS_REG_21__SCAN_IN
i P1_ADDRESS_REG_20__SCAN_IN
i P1_ADDRESS_REG_19__SCAN_IN
i P1_ADDRESS_REG_18__SCAN_IN
i P1_ADDRESS_REG_17__SCAN_IN
i P1_ADDRESS_REG_16__SCAN_IN
i P1_ADDRESS_REG_15__SCAN_IN
i P1_ADDRESS_REG_14__SCAN_IN
i P1_ADDRESS_REG_13__SCAN_IN
i P1_ADDRESS_REG_12__SCAN_IN
i P1_ADDRESS_REG_11__SCAN_IN
i P1_ADDRESS_REG_10__SCAN_IN
i P1_ADDRESS_REG_9__SCAN_IN
i P1_ADDRESS_REG_8__SCAN_IN
i P1_ADDRESS_REG_7__SCAN_IN
i P1_ADDRESS_REG_6__SCAN_IN
i P1_ADDRESS_REG_5__SCAN_IN
i P1_ADDRESS_REG_4__SCAN_IN
i P1_ADDRESS_REG_3__SCAN_IN
i P1_ADDRESS_REG_2__SCAN_IN
i P1_ADDRESS_REG_1__SCAN_IN
i P1_ADDRESS_REG_0__SCAN_IN
i P1_STATE_REG_2__SCAN_IN
i P1_STATE_REG_1__SCAN_IN
i P1_STATE_REG_0__SCAN_IN
i P1_DATAWIDTH_REG_0__SCAN_IN
i P1_DATAWIDTH_REG_1__SCAN_IN
i P1_DATAWIDTH_REG_2__SCAN_IN
i P1_DATAWIDTH_REG_3__SCAN_IN
i P1_DATAWIDTH_REG_4__SCAN_IN
i P1_DATAWIDTH_REG_5__SCAN_IN
i P1_DATAWIDTH_REG_6__SCAN_IN
i P1_DATAWIDTH_REG_7__SCAN_IN
i P1_DATAWIDTH_REG_8__SCAN_IN
i P1_DATAWIDTH_REG_9__SCAN_IN
i P1_DATAWIDTH_REG_10__SCAN_IN
i P1_DATAWIDTH_REG_11__SCAN_IN
i P1_DATAWIDTH_REG_12__SCAN_IN
i P1_DATAWIDTH_REG_13__SCAN_IN
i P1_DATAWIDTH_REG_14__SCAN_IN
i P1_DATAWIDTH_REG_15__SCAN_IN
i P1_DATAWIDTH_REG_16__SCAN_IN
i P1_DATAWIDTH_REG_17__SCAN_IN
i P1_DATAWIDTH_REG_18__SCAN_IN
i P1_DATAWIDTH_REG_19__SCAN_IN
i P1_DATAWIDTH_REG_20__SCAN_IN
i P1_DATAWIDTH_REG_21__SCAN_IN
i P1_DATAWIDTH_REG_22__SCAN_IN
i P1_DATAWIDTH_REG_23__SCAN_IN
i P1_DATAWIDTH_REG_24__SCAN_IN
i P1_DATAWIDTH_REG_25__SCAN_IN
i P1_DATAWIDTH_REG_26__SCAN_IN
i P1_DATAWIDTH_REG_27__SCAN_IN
i P1_DATAWIDTH_REG_28__SCAN_IN
i P1_DATAWIDTH_REG_29__SCAN_IN
i P1_DATAWIDTH_REG_30__SCAN_IN
i P1_DATAWIDTH_REG_31__SCAN_IN
i P1_STATE2_REG_3__SCAN_IN
i P1_STATE2_REG_2__SCAN_IN
i P1_STATE2_REG_1__SCAN_IN
i P1_STATE2_REG_0__SCAN_IN
i P1_INSTQUEUE_REG_15__7__SCAN_IN
i P1_INSTQUEUE_REG_15__6__SCAN_IN
i P1_INSTQUEUE_REG_15__5__SCAN_IN
i P1_INSTQUEUE_REG_15__4__SCAN_IN
i P1_INSTQUEUE_REG_15__3__SCAN_IN
i P1_INSTQUEUE_REG_15__2__SCAN_IN
i P1_INSTQUEUE_REG_15__1__SCAN_IN
i P1_INSTQUEUE_REG_15__0__SCAN_IN
i P1_INSTQUEUE_REG_14__7__SCAN_IN
i P1_INSTQUEUE_REG_14__6__SCAN_IN
i P1_INSTQUEUE_REG_14__5__SCAN_IN
i P1_INSTQUEUE_REG_14__4__SCAN_IN
i P1_INSTQUEUE_REG_14__3__SCAN_IN
i P1_INSTQUEUE_REG_14__2__SCAN_IN
i P1_INSTQUEUE_REG_14__1__SCAN_IN
i P1_INSTQUEUE_REG_14__0__SCAN_IN
i P1_INSTQUEUE_REG_13__7__SCAN_IN
i P1_INSTQUEUE_REG_13__6__SCAN_IN
i P1_INSTQUEUE_REG_13__5__SCAN_IN
i P1_INSTQUEUE_REG_13__4__SCAN_IN
i P1_INSTQUEUE_REG_13__3__SCAN_IN
i P1_INSTQUEUE_REG_13__2__SCAN_IN
i P1_INSTQUEUE_REG_13__1__SCAN_IN
i P1_INSTQUEUE_REG_13__0__SCAN_IN
i P1_INSTQUEUE_REG_12__7__SCAN_IN
i P1_INSTQUEUE_REG_12__6__SCAN_IN
i P1_INSTQUEUE_REG_12__5__SCAN_IN
i P1_INSTQUEUE_REG_12__4__SCAN_IN
i P1_INSTQUEUE_REG_12__3__SCAN_IN
i P1_INSTQUEUE_REG_12__2__SCAN_IN
i P1_INSTQUEUE_REG_12__1__SCAN_IN
i P1_INSTQUEUE_REG_12__0__SCAN_IN
i P1_INSTQUEUE_REG_11__7__SCAN_IN
i P1_INSTQUEUE_REG_11__6__SCAN_IN
i P1_INSTQUEUE_REG_11__5__SCAN_IN
i P1_INSTQUEUE_REG_11__4__SCAN_IN
i P1_INSTQUEUE_REG_11__3__SCAN_IN
i P1_INSTQUEUE_REG_11__2__SCAN_IN
i P1_INSTQUEUE_REG_11__1__SCAN_IN
i P1_INSTQUEUE_REG_11__0__SCAN_IN
i P1_INSTQUEUE_REG_10__7__SCAN_IN
i P1_INSTQUEUE_REG_10__6__SCAN_IN
i P1_INSTQUEUE_REG_10__5__SCAN_IN
i P1_INSTQUEUE_REG_10__4__SCAN_IN
i P1_INSTQUEUE_REG_10__3__SCAN_IN
i P1_INSTQUEUE_REG_10__2__SCAN_IN
i P1_INSTQUEUE_REG_10__1__SCAN_IN
i P1_INSTQUEUE_REG_10__0__SCAN_IN
i P1_INSTQUEUE_REG_9__7__SCAN_IN
i P1_INSTQUEUE_REG_9__6__SCAN_IN
i P1_INSTQUEUE_REG_9__5__SCAN_IN
i P1_INSTQUEUE_REG_9__4__SCAN_IN
i P1_INSTQUEUE_REG_9__3__SCAN_IN
i P1_INSTQUEUE_REG_9__2__SCAN_IN
i P1_INSTQUEUE_REG_9__1__SCAN_IN
i P1_INSTQUEUE_REG_9__0__SCAN_IN
i P1_INSTQUEUE_REG_8__7__SCAN_IN
i P1_INSTQUEUE_REG_8__6__SCAN_IN
i P1_INSTQUEUE_REG_8__5__SCAN_IN
i P1_INSTQUEUE_REG_8__4__SCAN_IN
i P1_INSTQUEUE_REG_8__3__SCAN_IN
i P1_INSTQUEUE_REG_8__2__SCAN_IN
i P1_INSTQUEUE_REG_8__1__SCAN_IN
i P1_INSTQUEUE_REG_8__0__SCAN_IN
i P1_INSTQUEUE_REG_7__7__SCAN_IN
i P1_INSTQUEUE_REG_7__6__SCAN_IN
i P1_INSTQUEUE_REG_7__5__SCAN_IN
i P1_INSTQUEUE_REG_7__4__SCAN_IN
i P1_INSTQUEUE_REG_7__3__SCAN_IN
i P1_INSTQUEUE_REG_7__2__SCAN_IN
i P1_INSTQUEUE_REG_7__1__SCAN_IN
i P1_INSTQUEUE_REG_7__0__SCAN_IN
i P1_INSTQUEUE_REG_6__7__SCAN_IN
i P1_INSTQUEUE_REG_6__6__SCAN_IN
i P1_INSTQUEUE_REG_6__5__SCAN_IN
i P1_INSTQUEUE_REG_6__4__SCAN_IN
i P1_INSTQUEUE_REG_6__3__SCAN_IN
i P1_INSTQUEUE_REG_6__2__SCAN_IN
i P1_INSTQUEUE_REG_6__1__SCAN_IN
i P1_INSTQUEUE_REG_6__0__SCAN_IN
i P1_INSTQUEUE_REG_5__7__SCAN_IN
i P1_INSTQUEUE_REG_5__6__SCAN_IN
i P1_INSTQUEUE_REG_5__5__SCAN_IN
i P1_INSTQUEUE_REG_5__4__SCAN_IN
i P1_INSTQUEUE_REG_5__3__SCAN_IN
i P1_INSTQUEUE_REG_5__2__SCAN_IN
i P1_INSTQUEUE_REG_5__1__SCAN_IN
i P1_INSTQUEUE_REG_5__0__SCAN_IN
i P1_INSTQUEUE_REG_4__7__SCAN_IN
i P1_INSTQUEUE_REG_4__6__SCAN_IN
i P1_INSTQUEUE_REG_4__5__SCAN_IN
i P1_INSTQUEUE_REG_4__4__SCAN_IN
i P1_INSTQUEUE_REG_4__3__SCAN_IN
i P1_INSTQUEUE_REG_4__2__SCAN_IN
i P1_INSTQUEUE_REG_4__1__SCAN_IN
o P3_DATAO_REG_31__SCAN_IN
o P3_DATAO_REG_30__SCAN_IN
o P3_DATAO_REG_29__SCAN_IN
o P3_DATAO_REG_28__SCAN_IN
o P3_DATAO_REG_27__SCAN_IN
o P3_DATAO_REG_26__SCAN_IN
o P3_DATAO_REG_25__SCAN_IN
o P3_DATAO_REG_24__SCAN_IN
o P3_DATAO_REG_23__SCAN_IN
o P3_DATAO_REG_22__SCAN_IN
o P3_DATAO_REG_21__SCAN_IN
o P3_DATAO_REG_20__SCAN_IN
o P3_DATAO_REG_19__SCAN_IN
o P3_DATAO_REG_18__SCAN_IN
o P3_DATAO_REG_17__SCAN_IN
o P3_DATAO_REG_16__SCAN_IN
o P3_DATAO_REG_15__SCAN_IN
o P3_DATAO_REG_14__SCAN_IN
o P3_DATAO_REG_13__SCAN_IN
o P3_DATAO_REG_12__SCAN_IN
o P3_DATAO_REG_11__SCAN_IN
o P3_DATAO_REG_10__SCAN_IN
o P3_DATAO_REG_9__SCAN_IN
o P3_DATAO_REG_8__SCAN_IN
o P3_DATAO_REG_7__SCAN_IN
o P3_DATAO_REG_6__SCAN_IN
o P3_DATAO_REG_5__SCAN_IN
o P3_DATAO_REG_4__SCAN_IN
o P3_DATAO_REG_3__SCAN_IN
o P3_DATAO_REG_2__SCAN_IN
o P3_DATAO_REG_1__SCAN_IN
o P3_DATAO_REG_0__SCAN_IN
o P1_ADDRESS_REG_29__SCAN_IN
o P1_ADDRESS_REG_28__SCAN_IN
o P1_ADDRESS_REG_27__SCAN_IN
o P1_ADDRESS_REG_26__SCAN_IN
o P1_ADDRESS_REG_25__SCAN_IN
o P1_ADDRESS_REG_24__SCAN_IN
o P1_ADDRESS_REG_23__SCAN_IN
o P1_ADDRESS_REG_22__SCAN_IN
o P1_ADDRESS_REG_21__SCAN_IN
o P1_ADDRESS_REG_20__SCAN_IN
o P1_ADDRESS_REG_19__SCAN_IN
o P1_ADDRESS_REG_18__SCAN_IN
o P1_ADDRESS_REG_17__SCAN_IN
o P1_ADDRESS_REG_16__SCAN_IN
o P1_ADDRESS_REG_15__SCAN_IN
o P1_ADDRESS_REG_14__SCAN_IN
o P1_ADDRESS_REG_13__SCAN_IN
o P1_ADDRESS_REG_12__SCAN_IN
o P1_ADDRESS_REG_11__SCAN_IN
o P1_ADDRESS_REG_10__SCAN_IN
o P1_ADDRESS_REG_9__SCAN_IN
o P1_ADDRESS_REG_8__SCAN_IN
o P1_ADDRESS_REG_7__SCAN_IN
o P1_ADDRESS_REG_6__SCAN_IN
o P1_ADDRESS_REG_5__SCAN_IN
o P1_ADDRESS_REG_4__SCAN_IN
o P1_ADDRESS_REG_3__SCAN_IN
o P1_ADDRESS_REG_2__SCAN_IN
o P1_ADDRESS_REG_1__SCAN_IN
o P1_ADDRESS_REG_0__SCAN_IN
o U355
o U356
o U357
o U358
o U359
o U360
o U361
o U362
o U363
o U364
o U366
o U367
o U368
o U369
o U370
o U371
o U372
o U373
o U374
o U375
o U347
o U348
o U349
o U350
o U351
o U352
o U353
o U354
o U365
o U376
o P3_W_R_N_REG_SCAN_IN
o P3_D_C_N_REG_SCAN_IN
o P3_M_IO_N_REG_SCAN_IN
o P1_ADS_N_REG_SCAN_IN
o P3_ADS_N_REG_SCAN_IN
o U247
o U246
o U245
o U244
o U243
o U242
o U241
o U240
o U239
o U238
o U237
o U236
o U235
o U234
o U233
o U232
o U231
o U230
o U229
o U228
o U227
o U226
o U225
o U224
o U223
o U222
o U221
o U220
o U219
o U218
o U217
o U216
o U251
o U252
o U253
o U254
o U255
o U256
o U257
o U258
o U259
o U260
o U261
o U262
o U263
o U264
o U265
o U266
o U267
o U268
o U269
o U270
o U271
o U272
o U273
o U274
o U275
o U276
o U277
o U278
o U279
o U280
o U281
o U282
o U212
o U215
o U213
o U214
o P3_U3274
o P3_U3275
o P3_U3276
o P3_U3277
o P3_U3061
o P3_U3060
o P3_U3059
o P3_U3058
o P3_U3057
o P3_U3056
o P3_U3055
o P3_U3054
o P3_U3053
o P3_U3052
o P3_U3051
o P3_U3050
o P3_U3049
o P3_U3048
o P3_U3047
o P3_U3046
o P3_U3045
o P3_U3044
o P3_U3043
o P3_U3042
o P3_U3041
o P3_U3040
o P3_U3039
o P3_U3038
o P3_U3037
o P3_U3036
o P3_U3035
o P3_U3034
o P3_U3033
o P3_U3032
o P3_U3031
o P3_U3030
o P3_U3029
o P3_U3280
o P3_U3281
o P3_U3028
o P3_U3027
o P3_U3026
o P3_U3025
o P3_U3024
o P3_U3023
o P3_U3022
o P3_U3021
o P3_U3020
o P3_U3019
o P3_U3018
o P3_U3017
o P3_U3016
o P3_U3015
o P3_U3014
o P3_U3013
o P3_U3012
o P3_U3011
o P3_U3010
o P3_U3009
o P3_U3008
o P3_U3007
o P3_U3006
o P3_U3005
o P3_U3004
o P3_U3003
o P3_U3002
o P3_U3001
o P3_U3000
o P3_U2999
o P3_U3282
o P3_U2998
o P3_U2997
o P3_U2996
o P3_U2995
o P3_U2994
o P3_U2993
o P3_U2992
o P3_U2991
o P3_U2990
o P3_U2989
o P3_U2988
o P3_U2987
o P3_U2986
o P3_U2985
o P3_U2984
o P3_U2983
o P3_U2982
o P3_U2981
o P3_U2980
o P3_U2979
o P3_U2978
o P3_U2977
o P3_U2976
o P3_U2975
o P3_U2974
o P3_U2973
o P3_U2972
o P3_U2971
o P3_U2970
o P3_U2969
o P3_U2968
o P3_U2967
o P3_U2966
o P3_U2965
o P3_U2964
o P3_U2963
o P3_U2962
o P3_U2961
o P3_U2960
o P3_U2959
o P3_U2958
o P3_U2957
o P3_U2956
o P3_U2955
o P3_U2954
o P3_U2953
o P3_U2952
o P3_U2951
o P3_U2950
o P3_U2949
o P3_U2948
o P3_U2947
o P3_U2946
o P3_U2945
o P3_U2944
o P3_U2943
o P3_U2942
o P3_U2941
o P3_U2940
o P3_U2939
o P3_U2938
o P3_U2937
o P3_U2936
o P3_U2935
o P3_U2934
o P3_U2933
o P3_U2932
o P3_U2931
o P3_U2930
o P3_U2929
o P3_U2928
o P3_U2927
o P3_U2926
o P3_U2925
o P3_U2924
o P3_U2923
o P3_U2922
o P3_U2921
o P3_U2920
o P3_U2919
o P3_U2918
o P3_U2917
o P3_U2916
o P3_U2915
o P3_U2914
o P3_U2913
o P3_U2912
o P3_U2911
o P3_U2910
o P3_U2909
o P3_U2908
o P3_U2907
o P3_U2906
o P3_U2905
o P3_U2904
o P3_U2903
o P3_U2902
o P3_U2901
o P3_U2900
o P3_U2899
o P3_U2898
o P3_U2897
o P3_U2896
o P3_U2895
o P3_U2894
o P3_U2893
o P3_U2892
o P3_U2891
o P3_U2890
o P3_U2889
o P3_U2888
o P3_U2887
o P3_U2886
o P3_U2885
o P3_U2884
o P3_U2883
o P3_U2882
o P3_U2881
o P3_U2880
o P3_U2879
o P3_U2878
o P3_U2877
o P3_U2876
o P3_U2875
o P3_U2874
o P3_U2873
o P3_U2872
o P3_U2871
o P3_U2870
o P3_U2869
o P3_U2868
o P3_U3284
o P3_U3285
o P3_U3288
o P3_U3289
o P3_U3290
o P3_U2867
o P3_U2866
o P3_U2865
o P3_U2864
o P3_U2863
o P3_U2862
o P3_U2861
o P3_U2860
o P3_U2859
o P3_U2858
o P3_U2857
o P3_U2856
o P3_U2855
o P3_U2854
o P3_U2853
o P3_U2852
o P3_U2851
o P3_U2850
o P3_U2849
o P3_U2848
o P3_U2847
o P3_U2846
o P3_U2845
o P3_U2844
o P3_U2843
o P3_U2842
o P3_U2841
o P3_U2840
o P3_U2839
o P3_U2838
o P3_U2837
o P3_U2836
o P3_U2835
o P3_U2834
o P3_U2833
o P3_U2832
o P3_U2831
o P3_U2830
o P3_U2829
o P3_U2828
o P3_U2827
o P3_U2826
o P3_U2825
o P3_U2824
o P3_U2823
o P3_U2822
o P3_U2821
o P3_U2820
o P3_U2819
o P3_U2818
o P3_U2817
o P3_U2816
o P3_U2815
o P3_U2814
o P3_U2813
o P3_U2812
o P3_U2811
o P3_U2810
o P3_U2809
o P3_U2808
o P3_U2807
o P3_U2806
o P3_U2805
o P3_U2804
o P3_U2803
o P3_U2802
o P3_U2801
o P3_U2800
o P3_U2799
o P3_U2798
o P3_U2797
o P3_U2796
o P3_U2795
o P3_U2794
o P3_U2793
o P3_U2792
o P3_U2791
o P3_U2790
o P3_U2789
o P3_U2788
o P3_U2787
o P3_U2786
o P3_U2785
o P3_U2784
o P3_U2783
o P3_U2782
o P3_U2781
o P3_U2780
o P3_U2779
o P3_U2778
o P3_U2777
o P3_U2776
o P3_U2775
o P3_U2774
o P3_U2773
o P3_U2772
o P3_U2771
o P3_U2770
o P3_U2769
o P3_U2768
o P3_U2767
o P3_U2766
o P3_U2765
o P3_U2764
o P3_U2763
o P3_U2762
o P3_U2761
o P3_U2760
o P3_U2759
o P3_U2758
o P3_U2757
o P3_U2756
o P3_U2755
o P3_U2754
o P3_U2753
o P3_U2752
o P3_U2751
o P3_U2750
o P3_U2749
o P3_U2748
o P3_U2747
o P3_U2746
o P3_U2745
o P3_U2744
o P3_U2743
o P3_U2742
o P3_U2741
o P3_U2740
o P3_U2739
o P3_U2738
o P3_U2737
o P3_U2736
o P3_U2735
o P3_U2734
o P3_U2733
o P3_U2732
o P3_U2731
o P3_U2730
o P3_U2729
o P3_U2728
o P3_U2727
o P3_U2726
o P3_U2725
o P3_U2724
o P3_U2723
o P3_U2722
o P3_U2721
o P3_U2720
o P3_U2719
o P3_U2718
o P3_U2717
o P3_U2716
o P3_U2715
o P3_U2714
o P3_U2713
o P3_U2712
o P3_U2711
o P3_U2710
o P3_U2709
o P3_U2708
o P3_U2707
o P3_U2706
o P3_U2705
o P3_U2704
o P3_U2703
o P3_U2702
o P3_U2701
o P3_U2700
o P3_U2699
o P3_U2698
o P3_U2697
o P3_U2696
o P3_U2695
o P3_U2694
o P3_U2693
o P3_U2692
o P3_U2691
o P3_U2690
o P3_U2689
o P3_U2688
o P3_U2687
o P3_U2686
o P3_U2685
o P3_U2684
o P3_U2683
o P3_U2682
o P3_U2681
o P3_U2680
o P3_U2679
o P3_U2678
o P3_U2677
o P3_U2676
o P3_U2675
o P3_U2674
o P3_U2673
o P3_U2672
o P3_U2671
o P3_U2670
o P3_U2669
o P3_U2668
o P3_U2667
o P3_U2666
o P3_U2665
o P3_U2664
o P3_U2663
o P3_U2662
o P3_U2661
o P3_U2660
o P3_U2659
o P3_U2658
o P3_U2657
o P3_U2656
o P3_U2655
o P3_U2654
o P3_U2653
o P3_U2652
o P3_U2651
o P3_U2650
o P3_U2649
o P3_U2648
o P3_U2647
o P3_U2646
o P3_U2645
o P3_U2644
o P3_U2643
o P3_U2642
o P3_U2641
o P3_U2640
o P3_U2639
o P3_U3292
o P3_U2638
o P3_U3293
o P3_U3294
o P3_U2637
o P3_U3295
o P3_U2636
o P3_U3296
o P3_U2635
o P3_U3297
o P3_U2634
o P3_U2633
o P3_U3298
o P3_U3299
o P2_U3585
o P2_U3586
o P2_U3587
o P2_U3588
o P2_U3241
o P2_U3240
o P2_U3239
o P2_U3238
o P2_U3237
o P2_U3236
o P2_U3235
o P2_U3234
o P2_U3233
o P2_U3232
o P2_U3231
o P2_U3230
o P2_U3229
o P2_U3228
o P2_U3227
o P2_U3226
o P2_U3225
o P2_U3224
o P2_U3223
o P2_U3222
o P2_U3221
o P2_U3220
o P2_U3219
o P2_U3218
o P2_U3217
o P2_U3216
o P2_U3215
o P2_U3214
o P2_U3213
o P2_U3212
o P2_U3211
o P2_U3210
o P2_U3209
o P2_U3591
o P2_U3592
o P2_U3208
o P2_U3207
o P2_U3206
o P2_U3205
o P2_U3204
o P2_U3203
o P2_U3202
o P2_U3201
o P2_U3200
o P2_U3199
o P2_U3198
o P2_U3197
o P2_U3196
o P2_U3195
o P2_U3194
o P2_U3193
o P2_U3192
o P2_U3191
o P2_U3190
o P2_U3189
o P2_U3188
o P2_U3187
o P2_U3186
o P2_U3185
o P2_U3184
o P2_U3183
o P2_U3182
o P2_U3181
o P2_U3180
o P2_U3179
o P2_U3593
o P2_U3178
o P2_U3177
o P2_U3176
o P2_U3175
o P2_U3174
o P2_U3173
o P2_U3172
o P2_U3171
o P2_U3170
o P2_U3169
o P2_U3168
o P2_U3167
o P2_U3166
o P2_U3165
o P2_U3164
o P2_U3163
o P2_U3162
o P2_U3161
o P2_U3160
o P2_U3159
o P2_U3158
o P2_U3157
o P2_U3156
o P2_U3155
o P2_U3154
o P2_U3153
o P2_U3152
o P2_U3151
o P2_U3150
o P2_U3149
o P2_U3148
o P2_U3147
o P2_U3146
o P2_U3145
o P2_U3144
o P2_U3143
o P2_U3142
o P2_U3141
o P2_U3140
o P2_U3139
o P2_U3138
o P2_U3137
o P2_U3136
o P2_U3135
o P2_U3134
o P2_U3133
o P2_U3132
o P2_U3131
o P2_U3130
o P2_U3129
o P2_U3128
o P2_U3127
o P2_U3126
o P2_U3125
o P2_U3124
o P2_U3123
o P2_U3122
o P2_U3121
o P2_U3120
o P2_U3119
o P2_U3118
o P2_U3117
o P2_U3116
o P2_U3115
o P2_U3114
o P2_U3113
o P2_U3112
o P2_U3111
o P2_U3110
o P2_U3109
o P2_U3108
o P2_U3107
o P2_U3106
o P2_U3105
o P2_U3104
o P2_U3103
o P2_U3102
o P2_U3101
o P2_U3100
o P2_U3099
o P2_U3098
o P2_U3097
o P2_U3096
o P2_U3095
o P2_U3094
o P2_U3093
o P2_U3092
o P2_U3091
o P2_U3090
o P2_U3089
o P2_U3088
o P2_U3087
o P2_U3086
o P2_U3085
o P2_U3084
o P2_U3083
o P2_U3082
o P2_U3081
o P2_U3080
o P2_U3079
o P2_U3078
o P2_U3077
o P2_U3076
o P2_U3075
o P2_U3074
o P2_U3073
o P2_U3072
o P2_U3071
o P2_U3070
o P2_U3069
o P2_U3068
o P2_U3067
o P2_U3066
o P2_U3065
o P2_U3064
o P2_U3063
o P2_U3062
o P2_U3061
o P2_U3060
o P2_U3059
o P2_U3058
o P2_U3057
o P2_U3056
o P2_U3055
o P2_U3054
o P2_U3053
o P2_U3052
o P2_U3051
o P2_U3050
o P2_U3049
o P2_U3048
o P2_U3595
o P2_U3596
o P2_U3599
o P2_U3600
o P2_U3601
o P2_U3047
o P2_U3602
o P2_U3603
o P2_U3604
o P2_U3605
o P2_U3046
o P2_U3045
o P2_U3044
o P2_U3043
o P2_U3042
o P2_U3041
o P2_U3040
o P2_U3039
o P2_U3038
o P2_U3037
o P2_U3036
o P2_U3035
o P2_U3034
o P2_U3033
o P2_U3032
o P2_U3031
o P2_U3030
o P2_U3029
o P2_U3028
o P2_U3027
o P2_U3026
o P2_U3025
o P2_U3024
o P2_U3023
o P2_U3022
o P2_U3021
o P2_U3020
o P2_U3019
o P2_U3018
o P2_U3017
o P2_U3016
o P2_U3015
o P2_U3014
o P2_U3013
o P2_U3012
o P2_U3011
o P2_U3010
o P2_U3009
o P2_U3008
o P2_U3007
o P2_U3006
o P2_U3005
o P2_U3004
o P2_U3003
o P2_U3002
o P2_U3001
o P2_U3000
o P2_U2999
o P2_U2998
o P2_U2997
o P2_U2996
o P2_U2995
o P2_U2994
o P2_U2993
o P2_U2992
o P2_U2991
o P2_U2990
o P2_U2989
o P2_U2988
o P2_U2987
o P2_U2986
o P2_U2985
o P2_U2984
o P2_U2983
o P2_U2982
o P2_U2981
o P2_U2980
o P2_U2979
o P2_U2978
o P2_U2977
o P2_U2976
o P2_U2975
o P2_U2974
o P2_U2973
o P2_U2972
o P2_U2971
o P2_U2970
o P2_U2969
o P2_U2968
o P2_U2967
o P2_U2966
o P2_U2965
o P2_U2964
o P2_U2963
o P2_U2962
o P2_U2961
o P2_U2960
o P2_U2959
o P2_U2958
o P2_U2957
o P2_U2956
o P2_U2955
o P2_U2954
o P2_U2953
o P2_U2952
o P2_U2951
o P2_U2950
o P2_U2949
o P2_U2948
o P2_U2947
o P2_U2946
o P2_U2945
o P2_U2944
o P2_U2943
o P2_U2942
o P2_U2941
o P2_U2940
o P2_U2939
o P2_U2938
o P2_U2937
o P2_U2936
o P2_U2935
o P2_U2934
o P2_U2933
o P2_U2932
o P2_U2931
o P2_U2930
o P2_U2929
o P2_U2928
o P2_U2927
o P2_U2926
o P2_U2925
o P2_U2924
o P2_U2923
o P2_U2922
o P2_U2921
o P2_U2920
o P2_U2919
o P2_U2918
o P2_U2917
o P2_U2916
o P2_U2915
o P2_U2914
o P2_U2913
o P2_U2912
o P2_U2911
o P2_U2910
o P2_U2909
o P2_U2908
o P2_U2907
o P2_U2906
o P2_U2905
o P2_U2904
o P2_U2903
o P2_U2902
o P2_U2901
o P2_U2900
o P2_U2899
o P2_U2898
o P2_U2897
o P2_U2896
o P2_U2895
o P2_U2894
o P2_U2893
o P2_U2892
o P2_U2891
o P2_U2890
o P2_U2889
o P2_U2888
o P2_U2887
o P2_U2886
o P2_U2885
o P2_U2884
o P2_U2883
o P2_U2882
o P2_U2881
o P2_U2880
o P2_U2879
o P2_U2878
o P2_U2877
o P2_U2876
o P2_U2875
o P2_U2874
o P2_U2873
o P2_U2872
o P2_U2871
o P2_U2870
o P2_U2869
o P2_U2868
o P2_U2867
o P2_U2866
o P2_U2865
o P2_U2864
o P2_U2863
o P2_U2862
o P2_U2861
o P2_U2860
o P2_U2859
o P2_U2858
o P2_U2857
o P2_U2856
o P2_U2855
o P2_U2854
o P2_U2853
o P2_U2852
o P2_U2851
o P2_U2850
o P2_U2849
o P2_U2848
o P2_U2847
o P2_U2846
o P2_U2845
o P2_U2844
o P2_U2843
o P2_U2842
o P2_U2841
o P2_U2840
o P2_U2839
o P2_U2838
o P2_U2837
o P2_U2836
o P2_U2835
o P2_U2834
o P2_U2833
o P2_U2832
o P2_U2831
o P2_U2830
o P2_U2829
o P2_U2828
o P2_U2827
o P2_U2826
o P2_U2825
o P2_U2824
o P2_U2823
o P2_U2822
o P2_U2821
o P2_U2820
o P2_U3608
o P2_U2819
o P2_U3609
o P2_U2818
o P2_U3610
o P2_U2817
o P2_U3611
o P2_U2816
o P2_U2815
o P2_U3612
o P2_U2814
o P1_U3458
o P1_U3459
o P1_U3460
o P1_U3461
o P1_U3226
o P1_U3225
o P1_U3224
o P1_U3223
o P1_U3222
o P1_U3221
o P1_U3220
o P1_U3219
o P1_U3218
o P1_U3217
o P1_U3216
o P1_U3215
o P1_U3214
o P1_U3213
o P1_U3212
o P1_U3211
o P1_U3210
o P1_U3209
o P1_U3208
o P1_U3207
o P1_U3206
o P1_U3205
o P1_U3204
o P1_U3203
o P1_U3202
o P1_U3201
o P1_U3200
o P1_U3199
o P1_U3198
o P1_U3197
o P1_U3196
o P1_U3195
o P1_U3194
o P1_U3464
o P1_U3465
o P1_U3193
o P1_U3192
o P1_U3191
o P1_U3190
o P1_U3189
o P1_U3188
o P1_U3187
o P1_U3186
o P1_U3185
o P1_U3184
o P1_U3183
o P1_U3182
o P1_U3181
o P1_U3180
o P1_U3179
o P1_U3178
o P1_U3177
o P1_U3176
o P1_U3175
o P1_U3174
o P1_U3173
o P1_U3172
o P1_U3171
o P1_U3170
o P1_U3169
o P1_U3168
o P1_U3167
o P1_U3166
o P1_U3165
o P1_U3164
o P1_U3466
o P1_U3163
o P1_U3162
o P1_U3161
o P1_U3160
o P1_U3159
o P1_U3158
o P1_U3157
o P1_U3156
o P1_U3155
o P1_U3154
o P1_U3153
o P1_U3152
o P1_U3151
o P1_U3150
o P1_U3149
o P1_U3148
o P1_U3147
o P1_U3146
o P1_U3145
o P1_U3144
o P1_U3143
o P1_U3142
o P1_U3141
o P1_U3140
o P1_U3139
o P1_U3138
o P1_U3137
o P1_U3136
o P1_U3135
o P1_U3134
o P1_U3133
o P1_U3132
o P1_U3131
o P1_U3130
o P1_U3129
o P1_U3128
o P1_U3127
o P1_U3126
o P1_U3125
o P1_U3124
o P1_U3123
o P1_U3122
o P1_U3121
o P1_U3120
o P1_U3119
o P1_U3118
o P1_U3117
o P1_U3116
o P1_U3115
o P1_U3114
o P1_U3113
o P1_U3112
o P1_U3111
o P1_U3110
o P1_U3109
o P1_U3108
o P1_U3107
o P1_U3106
o P1_U3105
o P1_U3104
o P1_U3103
o P1_U3102
o P1_U3101
o P1_U3100
o P1_U3099
o P1_U3098
o P1_U3097
o P1_U3096
o P1_U3095
o P1_U3094
o P1_U3093
o P1_U3092
o P1_U3091
o P1_U3090
o P1_U3089
o P1_U3088
o P1_U3087
o P1_U3086
o P1_U3085
o P1_U3084
o P1_U3083
o P1_U3082
o P1_U3081
o P1_U3080
o P1_U3079
o P1_U3078
o P1_U3077
o P1_U3076
o P1_U3075
o P1_U3074
o P1_U3073
o P1_U3072
o P1_U3071
o P1_U3070
o P1_U3069
o P1_U3068
o P1_U3067
o P1_U3066
o P1_U3065
o P1_U3064
o P1_U3063
o P1_U3062
o P1_U3061
o P1_U3060
o P1_U3059
o P1_U3058
o P1_U3057
o P1_U3056
o P1_U3055
o P1_U3054
o P1_U3053
o P1_U3052
o P1_U3051
o P1_U3050
o P1_U3049
o P1_U3048
o P1_U3047
o P1_U3046
o P1_U3045
o P1_U3044
o P1_U3043
o P1_U3042
o P1_U3041
o P1_U3040
o P1_U3039
o P1_U3038
o P1_U3037
o P1_U3036
o P1_U3035
o P1_U3034
o P1_U3033
o P1_U3468
o P1_U3469
o P1_U3472
o P1_U3473
o P1_U3474
o P1_U3032
o P1_U3475
o P1_U3476
o P1_U3477
o P1_U3478
o P1_U3031
o P1_U3030
o P1_U3029
o P1_U3028
o P1_U3027
o P1_U3026
o P1_U3025
o P1_U3024
o P1_U3023
o P1_U3022
o P1_U3021
o P1_U3020
o P1_U3019
o P1_U3018
o P1_U3017
o P1_U3016
o P1_U3015
o P1_U3014
o P1_U3013
o P1_U3012
o P1_U3011
o P1_U3010
o P1_U3009
o P1_U3008
o P1_U3007
o P1_U3006
o P1_U3005
o P1_U3004
o P1_U3003
o P1_U3002
o P1_U3001
o P1_U3000
o P1_U2999
o P1_U2998
o P1_U2997
o P1_U2996
o P1_U2995
o P1_U2994
o P1_U2993
o P1_U2992
o P1_U2991
o P1_U2990
o P1_U2989
o P1_U2988
o P1_U2987
o P1_U2986
o P1_U2985
o P1_U2984
o P1_U2983
o P1_U2982
o P1_U2981
o P1_U2980
o P1_U2979
o P1_U2978
o P1_U2977
o P1_U2976
o P1_U2975
o P1_U2974
o P1_U2973
o P1_U2972
o P1_U2971
o P1_U2970
o P1_U2969
o P1_U2968
o P1_U2967
o P1_U2966
o P1_U2965
o P1_U2964
o P1_U2963
o P1_U2962
o P1_U2961
o P1_U2960
o P1_U2959
o P1_U2958
o P1_U2957
o P1_U2956
o P1_U2955
o P1_U2954
o P1_U2953
o P1_U2952
o P1_U2951
o P1_U2950
o P1_U2949
o P1_U2948
o P1_U2947
o P1_U2946
o P1_U2945
o P1_U2944
o P1_U2943
o P1_U2942
o P1_U2941
o P1_U2940
o P1_U2939
o P1_U2938
o P1_U2937
o P1_U2936
o P1_U2935
o P1_U2934
o P1_U2933
o P1_U2932
o P1_U2931
o P1_U2930
o P1_U2929
o P1_U2928
o P1_U2927
o P1_U2926
o P1_U2925
o P1_U2924
o P1_U2923
o P1_U2922
o P1_U2921
o P1_U2920
o P1_U2919
o P1_U2918
o P1_U2917
o P1_U2916
o P1_U2915
o P1_U2914
o P1_U2913
o P1_U2912
o P1_U2911
o P1_U2910
o P1_U2909
o P1_U2908
o P1_U2907
o P1_U2906
o P1_U2905
o P1_U2904
o P1_U2903
o P1_U2902
o P1_U2901
o P1_U2900
o P1_U2899
o P1_U2898
o P1_U2897
o P1_U2896
o P1_U2895
o P1_U2894
o P1_U2893
o P1_U2892
o P1_U2891
o P1_U2890
o P1_U2889
o P1_U2888
o P1_U2887
o P1_U2886
o P1_U2885
o P1_U2884
o P1_U2883
o P1_U2882
o P1_U2881
o P1_U2880
o P1_U2879
o P1_U2878
o P1_U2877
o P1_U2876
o P1_U2875
o P1_U2874
o P1_U2873
o P1_U2872
o P1_U2871
o P1_U2870
o P1_U2869
o P1_U2868
o P1_U2867
o P1_U2866
o P1_U2865
o P1_U2864
o P1_U2863
o P1_U2862
o P1_U2861
o P1_U2860
o P1_U2859
o P1_U2858
o P1_U2857
o P1_U2856
o P1_U2855
o P1_U2854
o P1_U2853
o P1_U2852
o P1_U2851
o P1_U2850
o P1_U2849
o P1_U2848
o P1_U2847
o P1_U2846
o P1_U2845
o P1_U2844
o P1_U2843
o P1_U2842
o P1_U2841
o P1_U2840
o P1_U2839
o P1_U2838
o P1_U2837
o P1_U2836
o P1_U2835
o P1_U2834
o P1_U2833
o P1_U2832
o P1_U2831
o P1_U2830
o P1_U2829
o P1_U2828
o P1_U2827
o P1_U2826
o P1_U2825
o P1_U2824
o P1_U2823
o P1_U2822
o P1_U2821
o P1_U2820
o P1_U2819
o P1_U2818
o P1_U2817
o P1_U2816
o P1_U2815
o P1_U2814
o P1_U2813
o P1_U2812
o P1_U2811
o P1_U2810
o P1_U2809
o P1_U2808
o P1_U3481
o P1_U2807
o P1_U3482
o P1_U3483
o P1_U2806
o P1_U3484
o P1_U2805
o P1_U3485
o P1_U2804
o P1_U3486
o P1_U2803
o P1_U2802
o P1_U3487
o P1_U2801
g1 and U250 U214 ; U207
g2 and U378 U377 P2_W_R_N_REG_SCAN_IN P2_M_IO_N_REG_SCAN_IN ; U208
g3 and READY2 READY22_REG_SCAN_IN ; U209
g4 and READY1 READY11_REG_SCAN_IN ; U210
g5 and READY12_REG_SCAN_IN READY21_REG_SCAN_IN ; U211
g6 nand U208 R170_U6 U214 ; U212
g7 nand U380 U379 U215 P3_M_IO_N_REG_SCAN_IN ; U213
g8 nand U383 U381 R165_U6 P1_W_R_N_REG_SCAN_IN P1_M_IO_N_REG_SCAN_IN ; U214
g9 nand LT_748_U6 U208 ; U215
g10 nand U483 U484 U482 ; U216
g11 nand U480 U481 U479 ; U217
g12 nand U477 U478 U476 ; U218
g13 nand U474 U475 U473 ; U219
g14 nand U471 U472 U470 ; U220
g15 nand U468 U469 U467 ; U221
g16 nand U465 U466 U464 ; U222
g17 nand U462 U463 U461 ; U223
g18 nand U459 U460 U458 ; U224
g19 nand U456 U457 U455 ; U225
g20 nand U453 U454 U452 ; U226
g21 nand U450 U451 U449 ; U227
g22 nand U447 U448 U446 ; U228
g23 nand U444 U445 U443 ; U229
g24 nand U441 U442 U440 ; U230
g25 nand U438 U439 U437 ; U231
g26 nand U435 U436 U434 ; U232
g27 nand U432 U433 U431 ; U233
g28 nand U429 U430 U428 ; U234
g29 nand U426 U427 U425 ; U235
g30 nand U423 U424 U422 ; U236
g31 nand U420 U421 U419 ; U237
g32 nand U417 U418 U416 ; U238
g33 nand U414 U415 U413 ; U239
g34 nand U411 U412 U410 ; U240
g35 nand U408 U409 U407 ; U241
g36 nand U405 U406 U404 ; U242
g37 nand U402 U403 U401 ; U243
g38 nand U399 U400 U398 ; U244
g39 nand U396 U397 U395 ; U245
g40 nand U393 U394 U392 ; U246
g41 nand U390 U391 U389 ; U247
g42 not R165_U6 ; U248
g43 not R170_U6 ; U249
g44 nand U214 U387 ; U250
g45 nand U486 U485 ; U251
g46 nand U488 U487 ; U252
g47 nand U490 U489 ; U253
g48 nand U492 U491 ; U254
g49 nand U494 U493 ; U255
g50 nand U496 U495 ; U256
g51 nand U498 U497 ; U257
g52 nand U500 U499 ; U258
g53 nand U502 U501 ; U259
g54 nand U504 U503 ; U260
g55 nand U506 U505 ; U261
g56 nand U508 U507 ; U262
g57 nand U510 U509 ; U263
g58 nand U512 U511 ; U264
g59 nand U514 U513 ; U265
g60 nand U516 U515 ; U266
g61 nand U518 U517 ; U267
g62 nand U520 U519 ; U268
g63 nand U522 U521 ; U269
g64 nand U524 U523 ; U270
g65 nand U526 U525 ; U271
g66 nand U528 U527 ; U272
g67 nand U530 U529 ; U273
g68 nand U532 U531 ; U274
g69 nand U534 U533 ; U275
g70 nand U536 U535 ; U276
g71 nand U538 U537 ; U277
g72 nand U540 U539 ; U278
g73 nand U542 U541 ; U279
g74 nand U544 U543 ; U280
g75 nand U546 U545 ; U281
g76 nand U548 U547 ; U282
g77 nand U550 U549 ; U283
g78 nand U552 U551 ; U284
g79 nand U554 U553 ; U285
g80 nand U556 U555 ; U286
g81 nand U558 U557 ; U287
g82 nand U560 U559 ; U288
g83 nand U562 U561 ; U289
g84 nand U564 U563 ; U290
g85 nand U566 U565 ; U291
g86 nand U568 U567 ; U292
g87 nand U570 U569 ; U293
g88 nand U572 U571 ; U294
g89 nand U574 U573 ; U295
g90 nand U576 U575 ; U296
g91 nand U578 U577 ; U297
g92 nand U580 U579 ; U298
g93 nand U582 U581 ; U299
g94 nand U584 U583 ; U300
g95 nand U586 U585 ; U301
g96 nand U588 U587 ; U302
g97 nand U590 U589 ; U303
g98 nand U592 U591 ; U304
g99 nand U594 U593 ; U305
g100 nand U596 U595 ; U306
g101 nand U598 U597 ; U307
g102 nand U600 U599 ; U308
g103 nand U602 U601 ; U309
g104 nand U604 U603 ; U310
g105 nand U606 U605 ; U311
g106 nand U608 U607 ; U312
g107 nand U610 U609 ; U313
g108 nand U612 U611 ; U314
g109 nand U614 U613 ; U315
g110 nand U616 U615 ; U316
g111 nand U618 U617 ; U317
g112 nand U620 U619 ; U318
g113 nand U622 U621 ; U319
g114 nand U624 U623 ; U320
g115 nand U626 U625 ; U321
g116 nand U628 U627 ; U322
g117 nand U630 U629 ; U323
g118 nand U632 U631 ; U324
g119 nand U634 U633 ; U325
g120 nand U636 U635 ; U326
g121 nand U638 U637 ; U327
g122 nand U640 U639 ; U328
g123 nand U642 U641 ; U329
g124 nand U644 U643 ; U330
g125 nand U646 U645 ; U331
g126 nand U648 U647 ; U332
g127 nand U650 U649 ; U333
g128 nand U652 U651 ; U334
g129 nand U654 U653 ; U335
g130 nand U656 U655 ; U336
g131 nand U658 U657 ; U337
g132 nand U660 U659 ; U338
g133 nand U662 U661 ; U339
g134 nand U664 U663 ; U340
g135 nand U666 U665 ; U341
g136 nand U668 U667 ; U342
g137 nand U670 U669 ; U343
g138 nand U672 U671 ; U344
g139 nand U674 U673 ; U345
g140 nand U676 U675 ; U346
g141 nand U678 U677 ; U347
g142 nand U680 U679 ; U348
g143 nand U682 U681 ; U349
g144 nand U684 U683 ; U350
g145 nand U686 U685 ; U351
g146 nand U688 U687 ; U352
g147 nand U690 U689 ; U353
g148 nand U692 U691 ; U354
g149 nand U694 U693 ; U355
g150 nand U696 U695 ; U356
g151 nand U698 U697 ; U357
g152 nand U700 U699 ; U358
g153 nand U702 U701 ; U359
g154 nand U704 U703 ; U360
g155 nand U706 U705 ; U361
g156 nand U708 U707 ; U362
g157 nand U710 U709 ; U363
g158 nand U712 U711 ; U364
g159 nand U714 U713 ; U365
g160 nand U716 U715 ; U366
g161 nand U718 U717 ; U367
g162 nand U720 U719 ; U368
g163 nand U722 U721 ; U369
g164 nand U724 U723 ; U370
g165 nand U726 U725 ; U371
g166 nand U728 U727 ; U372
g167 nand U730 U729 ; U373
g168 nand U732 U731 ; U374
g169 nand U734 U733 ; U375
g170 nand U736 U735 ; U376
g171 nor P2_BE_N_REG_2__SCAN_IN P2_BE_N_REG_1__SCAN_IN P2_BE_N_REG_0__SCAN_IN P2_ADS_N_REG_SCAN_IN ; U377
g172 nor P2_BE_N_REG_3__SCAN_IN P2_D_C_N_REG_SCAN_IN ; U378
g173 nor P3_BE_N_REG_1__SCAN_IN P3_BE_N_REG_0__SCAN_IN P3_W_R_N_REG_SCAN_IN P3_D_C_N_REG_SCAN_IN P3_ADS_N_REG_SCAN_IN ; U379
g174 nor P3_BE_N_REG_3__SCAN_IN P3_BE_N_REG_2__SCAN_IN ; U380
g175 nor P1_BE_N_REG_3__SCAN_IN P1_BE_N_REG_1__SCAN_IN P1_BE_N_REG_0__SCAN_IN P1_D_C_N_REG_SCAN_IN P1_ADS_N_REG_SCAN_IN ; U381
g176 nand LT_782_120_U6 LT_782_U6 LT_782_119_U6 ; U382
g177 not P1_BE_N_REG_2__SCAN_IN ; U383
g178 not U382 ; U384
g179 not U214 ; U385
g180 not U215 ; U386
g181 nand R170_U6 U208 ; U387
g182 not U250 ; U388
g183 nand U207 P2_DATAO_REG_0__SCAN_IN ; U389
g184 nand U385 P1_DATAO_REG_0__SCAN_IN ; U390
g185 nand U388 BUF1_REG_0__SCAN_IN ; U391
g186 nand U207 P2_DATAO_REG_1__SCAN_IN ; U392
g187 nand U385 P1_DATAO_REG_1__SCAN_IN ; U393
g188 nand U388 BUF1_REG_1__SCAN_IN ; U394
g189 nand U207 P2_DATAO_REG_2__SCAN_IN ; U395
g190 nand U385 P1_DATAO_REG_2__SCAN_IN ; U396
g191 nand U388 BUF1_REG_2__SCAN_IN ; U397
g192 nand U207 P2_DATAO_REG_3__SCAN_IN ; U398
g193 nand U385 P1_DATAO_REG_3__SCAN_IN ; U399
g194 nand U388 BUF1_REG_3__SCAN_IN ; U400
g195 nand U207 P2_DATAO_REG_4__SCAN_IN ; U401
g196 nand U385 P1_DATAO_REG_4__SCAN_IN ; U402
g197 nand U388 BUF1_REG_4__SCAN_IN ; U403
g198 nand U207 P2_DATAO_REG_5__SCAN_IN ; U404
g199 nand U385 P1_DATAO_REG_5__SCAN_IN ; U405
g200 nand U388 BUF1_REG_5__SCAN_IN ; U406
g201 nand U207 P2_DATAO_REG_6__SCAN_IN ; U407
g202 nand U385 P1_DATAO_REG_6__SCAN_IN ; U408
g203 nand U388 BUF1_REG_6__SCAN_IN ; U409
g204 nand U207 P2_DATAO_REG_7__SCAN_IN ; U410
g205 nand U385 P1_DATAO_REG_7__SCAN_IN ; U411
g206 nand U388 BUF1_REG_7__SCAN_IN ; U412
g207 nand U207 P2_DATAO_REG_8__SCAN_IN ; U413
g208 nand U385 P1_DATAO_REG_8__SCAN_IN ; U414
g209 nand U388 BUF1_REG_8__SCAN_IN ; U415
g210 nand U207 P2_DATAO_REG_9__SCAN_IN ; U416
g211 nand U385 P1_DATAO_REG_9__SCAN_IN ; U417
g212 nand U388 BUF1_REG_9__SCAN_IN ; U418
g213 nand U207 P2_DATAO_REG_10__SCAN_IN ; U419
g214 nand U385 P1_DATAO_REG_10__SCAN_IN ; U420
g215 nand U388 BUF1_REG_10__SCAN_IN ; U421
g216 nand U207 P2_DATAO_REG_11__SCAN_IN ; U422
g217 nand U385 P1_DATAO_REG_11__SCAN_IN ; U423
g218 nand U388 BUF1_REG_11__SCAN_IN ; U424
g219 nand U207 P2_DATAO_REG_12__SCAN_IN ; U425
g220 nand U385 P1_DATAO_REG_12__SCAN_IN ; U426
g221 nand U388 BUF1_REG_12__SCAN_IN ; U427
g222 nand U207 P2_DATAO_REG_13__SCAN_IN ; U428
g223 nand U385 P1_DATAO_REG_13__SCAN_IN ; U429
g224 nand U388 BUF1_REG_13__SCAN_IN ; U430
g225 nand U207 P2_DATAO_REG_14__SCAN_IN ; U431
g226 nand U385 P1_DATAO_REG_14__SCAN_IN ; U432
g227 nand U388 BUF1_REG_14__SCAN_IN ; U433
g228 nand U207 P2_DATAO_REG_15__SCAN_IN ; U434
g229 nand U385 P1_DATAO_REG_15__SCAN_IN ; U435
g230 nand U388 BUF1_REG_15__SCAN_IN ; U436
g231 nand U207 P2_DATAO_REG_16__SCAN_IN ; U437
g232 nand U385 P1_DATAO_REG_16__SCAN_IN ; U438
g233 nand U388 BUF1_REG_16__SCAN_IN ; U439
g234 nand U207 P2_DATAO_REG_17__SCAN_IN ; U440
g235 nand U385 P1_DATAO_REG_17__SCAN_IN ; U441
g236 nand U388 BUF1_REG_17__SCAN_IN ; U442
g237 nand U207 P2_DATAO_REG_18__SCAN_IN ; U443
g238 nand U385 P1_DATAO_REG_18__SCAN_IN ; U444
g239 nand U388 BUF1_REG_18__SCAN_IN ; U445
g240 nand U207 P2_DATAO_REG_19__SCAN_IN ; U446
g241 nand U385 P1_DATAO_REG_19__SCAN_IN ; U447
g242 nand U388 BUF1_REG_19__SCAN_IN ; U448
g243 nand U207 P2_DATAO_REG_20__SCAN_IN ; U449
g244 nand U385 P1_DATAO_REG_20__SCAN_IN ; U450
g245 nand U388 BUF1_REG_20__SCAN_IN ; U451
g246 nand U207 P2_DATAO_REG_21__SCAN_IN ; U452
g247 nand U385 P1_DATAO_REG_21__SCAN_IN ; U453
g248 nand U388 BUF1_REG_21__SCAN_IN ; U454
g249 nand U207 P2_DATAO_REG_22__SCAN_IN ; U455
g250 nand U385 P1_DATAO_REG_22__SCAN_IN ; U456
g251 nand U388 BUF1_REG_22__SCAN_IN ; U457
g252 nand U207 P2_DATAO_REG_23__SCAN_IN ; U458
g253 nand U385 P1_DATAO_REG_23__SCAN_IN ; U459
g254 nand U388 BUF1_REG_23__SCAN_IN ; U460
g255 nand U207 P2_DATAO_REG_24__SCAN_IN ; U461
g256 nand U385 P1_DATAO_REG_24__SCAN_IN ; U462
g257 nand U388 BUF1_REG_24__SCAN_IN ; U463
g258 nand U207 P2_DATAO_REG_25__SCAN_IN ; U464
g259 nand U385 P1_DATAO_REG_25__SCAN_IN ; U465
g260 nand U388 BUF1_REG_25__SCAN_IN ; U466
g261 nand U207 P2_DATAO_REG_26__SCAN_IN ; U467
g262 nand U385 P1_DATAO_REG_26__SCAN_IN ; U468
g263 nand U388 BUF1_REG_26__SCAN_IN ; U469
g264 nand U207 P2_DATAO_REG_27__SCAN_IN ; U470
g265 nand U385 P1_DATAO_REG_27__SCAN_IN ; U471
g266 nand U388 BUF1_REG_27__SCAN_IN ; U472
g267 nand U207 P2_DATAO_REG_28__SCAN_IN ; U473
g268 nand U385 P1_DATAO_REG_28__SCAN_IN ; U474
g269 nand U388 BUF1_REG_28__SCAN_IN ; U475
g270 nand U207 P2_DATAO_REG_29__SCAN_IN ; U476
g271 nand U385 P1_DATAO_REG_29__SCAN_IN ; U477
g272 nand U388 BUF1_REG_29__SCAN_IN ; U478
g273 nand U207 P2_DATAO_REG_30__SCAN_IN ; U479
g274 nand U385 P1_DATAO_REG_30__SCAN_IN ; U480
g275 nand U388 BUF1_REG_30__SCAN_IN ; U481
g276 nand U207 P2_DATAO_REG_31__SCAN_IN ; U482
g277 nand U385 P1_DATAO_REG_31__SCAN_IN ; U483
g278 nand U388 BUF1_REG_31__SCAN_IN ; U484
g279 nand U215 BUF2_REG_0__SCAN_IN ; U485
g280 nand U386 P2_DATAO_REG_0__SCAN_IN ; U486
g281 nand U215 BUF2_REG_1__SCAN_IN ; U487
g282 nand U386 P2_DATAO_REG_1__SCAN_IN ; U488
g283 nand U215 BUF2_REG_2__SCAN_IN ; U489
g284 nand U386 P2_DATAO_REG_2__SCAN_IN ; U490
g285 nand U215 BUF2_REG_3__SCAN_IN ; U491
g286 nand U386 P2_DATAO_REG_3__SCAN_IN ; U492
g287 nand U215 BUF2_REG_4__SCAN_IN ; U493
g288 nand U386 P2_DATAO_REG_4__SCAN_IN ; U494
g289 nand U215 BUF2_REG_5__SCAN_IN ; U495
g290 nand U386 P2_DATAO_REG_5__SCAN_IN ; U496
g291 nand U215 BUF2_REG_6__SCAN_IN ; U497
g292 nand U386 P2_DATAO_REG_6__SCAN_IN ; U498
g293 nand U215 BUF2_REG_7__SCAN_IN ; U499
g294 nand U386 P2_DATAO_REG_7__SCAN_IN ; U500
g295 nand U215 BUF2_REG_8__SCAN_IN ; U501
g296 nand U386 P2_DATAO_REG_8__SCAN_IN ; U502
g297 nand U215 BUF2_REG_9__SCAN_IN ; U503
g298 nand U386 P2_DATAO_REG_9__SCAN_IN ; U504
g299 nand U215 BUF2_REG_10__SCAN_IN ; U505
g300 nand U386 P2_DATAO_REG_10__SCAN_IN ; U506
g301 nand U215 BUF2_REG_11__SCAN_IN ; U507
g302 nand U386 P2_DATAO_REG_11__SCAN_IN ; U508
g303 nand U215 BUF2_REG_12__SCAN_IN ; U509
g304 nand U386 P2_DATAO_REG_12__SCAN_IN ; U510
g305 nand U215 BUF2_REG_13__SCAN_IN ; U511
g306 nand U386 P2_DATAO_REG_13__SCAN_IN ; U512
g307 nand U215 BUF2_REG_14__SCAN_IN ; U513
g308 nand U386 P2_DATAO_REG_14__SCAN_IN ; U514
g309 nand U215 BUF2_REG_15__SCAN_IN ; U515
g310 nand U386 P2_DATAO_REG_15__SCAN_IN ; U516
g311 nand U215 BUF2_REG_16__SCAN_IN ; U517
g312 nand U386 P2_DATAO_REG_16__SCAN_IN ; U518
g313 nand U215 BUF2_REG_17__SCAN_IN ; U519
g314 nand U386 P2_DATAO_REG_17__SCAN_IN ; U520
g315 nand U215 BUF2_REG_18__SCAN_IN ; U521
g316 nand U386 P2_DATAO_REG_18__SCAN_IN ; U522
g317 nand U215 BUF2_REG_19__SCAN_IN ; U523
g318 nand U386 P2_DATAO_REG_19__SCAN_IN ; U524
g319 nand U215 BUF2_REG_20__SCAN_IN ; U525
g320 nand U386 P2_DATAO_REG_20__SCAN_IN ; U526
g321 nand U215 BUF2_REG_21__SCAN_IN ; U527
g322 nand U386 P2_DATAO_REG_21__SCAN_IN ; U528
g323 nand U215 BUF2_REG_22__SCAN_IN ; U529
g324 nand U386 P2_DATAO_REG_22__SCAN_IN ; U530
g325 nand U215 BUF2_REG_23__SCAN_IN ; U531
g326 nand U386 P2_DATAO_REG_23__SCAN_IN ; U532
g327 nand U215 BUF2_REG_24__SCAN_IN ; U533
g328 nand U386 P2_DATAO_REG_24__SCAN_IN ; U534
g329 nand U215 BUF2_REG_25__SCAN_IN ; U535
g330 nand U386 P2_DATAO_REG_25__SCAN_IN ; U536
g331 nand U215 BUF2_REG_26__SCAN_IN ; U537
g332 nand U386 P2_DATAO_REG_26__SCAN_IN ; U538
g333 nand U215 BUF2_REG_27__SCAN_IN ; U539
g334 nand U386 P2_DATAO_REG_27__SCAN_IN ; U540
g335 nand U215 BUF2_REG_28__SCAN_IN ; U541
g336 nand U386 P2_DATAO_REG_28__SCAN_IN ; U542
g337 nand U215 BUF2_REG_29__SCAN_IN ; U543
g338 nand U386 P2_DATAO_REG_29__SCAN_IN ; U544
g339 nand U215 BUF2_REG_30__SCAN_IN ; U545
g340 nand U386 P2_DATAO_REG_30__SCAN_IN ; U546
g341 nand U215 BUF2_REG_31__SCAN_IN ; U547
g342 nand U386 P2_DATAO_REG_31__SCAN_IN ; U548
g343 nand U249 BUF2_REG_9__SCAN_IN ; U549
g344 nand R170_U6 BUF1_REG_9__SCAN_IN ; U550
g345 nand U249 BUF2_REG_8__SCAN_IN ; U551
g346 nand R170_U6 BUF1_REG_8__SCAN_IN ; U552
g347 nand U249 BUF2_REG_7__SCAN_IN ; U553
g348 nand R170_U6 BUF1_REG_7__SCAN_IN ; U554
g349 nand U249 BUF2_REG_6__SCAN_IN ; U555
g350 nand R170_U6 BUF1_REG_6__SCAN_IN ; U556
g351 nand U249 BUF2_REG_5__SCAN_IN ; U557
g352 nand R170_U6 BUF1_REG_5__SCAN_IN ; U558
g353 nand U249 BUF2_REG_4__SCAN_IN ; U559
g354 nand R170_U6 BUF1_REG_4__SCAN_IN ; U560
g355 nand U249 BUF2_REG_3__SCAN_IN ; U561
g356 nand R170_U6 BUF1_REG_3__SCAN_IN ; U562
g357 nand U249 BUF2_REG_31__SCAN_IN ; U563
g358 nand R170_U6 BUF1_REG_31__SCAN_IN ; U564
g359 nand U249 BUF2_REG_30__SCAN_IN ; U565
g360 nand R170_U6 BUF1_REG_30__SCAN_IN ; U566
g361 nand U249 BUF2_REG_2__SCAN_IN ; U567
g362 nand R170_U6 BUF1_REG_2__SCAN_IN ; U568
g363 nand U249 BUF2_REG_29__SCAN_IN ; U569
g364 nand R170_U6 BUF1_REG_29__SCAN_IN ; U570
g365 nand U249 BUF2_REG_28__SCAN_IN ; U571
g366 nand R170_U6 BUF1_REG_28__SCAN_IN ; U572
g367 nand U249 BUF2_REG_27__SCAN_IN ; U573
g368 nand R170_U6 BUF1_REG_27__SCAN_IN ; U574
g369 nand U249 BUF2_REG_26__SCAN_IN ; U575
g370 nand R170_U6 BUF1_REG_26__SCAN_IN ; U576
g371 nand U249 BUF2_REG_25__SCAN_IN ; U577
g372 nand R170_U6 BUF1_REG_25__SCAN_IN ; U578
g373 nand U249 BUF2_REG_24__SCAN_IN ; U579
g374 nand R170_U6 BUF1_REG_24__SCAN_IN ; U580
g375 nand U249 BUF2_REG_23__SCAN_IN ; U581
g376 nand R170_U6 BUF1_REG_23__SCAN_IN ; U582
g377 nand U249 BUF2_REG_22__SCAN_IN ; U583
g378 nand R170_U6 BUF1_REG_22__SCAN_IN ; U584
g379 nand U249 BUF2_REG_21__SCAN_IN ; U585
g380 nand R170_U6 BUF1_REG_21__SCAN_IN ; U586
g381 nand U249 BUF2_REG_20__SCAN_IN ; U587
g382 nand R170_U6 BUF1_REG_20__SCAN_IN ; U588
g383 nand U249 BUF2_REG_1__SCAN_IN ; U589
g384 nand R170_U6 BUF1_REG_1__SCAN_IN ; U590
g385 nand U249 BUF2_REG_19__SCAN_IN ; U591
g386 nand R170_U6 BUF1_REG_19__SCAN_IN ; U592
g387 nand U249 BUF2_REG_18__SCAN_IN ; U593
g388 nand R170_U6 BUF1_REG_18__SCAN_IN ; U594
g389 nand U249 BUF2_REG_17__SCAN_IN ; U595
g390 nand R170_U6 BUF1_REG_17__SCAN_IN ; U596
g391 nand U249 BUF2_REG_16__SCAN_IN ; U597
g392 nand R170_U6 BUF1_REG_16__SCAN_IN ; U598
g393 nand U249 BUF2_REG_15__SCAN_IN ; U599
g394 nand R170_U6 BUF1_REG_15__SCAN_IN ; U600
g395 nand U249 BUF2_REG_14__SCAN_IN ; U601
g396 nand R170_U6 BUF1_REG_14__SCAN_IN ; U602
g397 nand U249 BUF2_REG_13__SCAN_IN ; U603
g398 nand R170_U6 BUF1_REG_13__SCAN_IN ; U604
g399 nand U249 BUF2_REG_12__SCAN_IN ; U605
g400 nand R170_U6 BUF1_REG_12__SCAN_IN ; U606
g401 nand U249 BUF2_REG_11__SCAN_IN ; U607
g402 nand R170_U6 BUF1_REG_11__SCAN_IN ; U608
g403 nand U249 BUF2_REG_10__SCAN_IN ; U609
g404 nand R170_U6 BUF1_REG_10__SCAN_IN ; U610
g405 nand U249 BUF2_REG_0__SCAN_IN ; U611
g406 nand R170_U6 BUF1_REG_0__SCAN_IN ; U612
g407 nand DATAI_9_ U248 ; U613
g408 nand R165_U6 BUF1_REG_9__SCAN_IN ; U614
g409 nand DATAI_8_ U248 ; U615
g410 nand R165_U6 BUF1_REG_8__SCAN_IN ; U616
g411 nand DATAI_7_ U248 ; U617
g412 nand R165_U6 BUF1_REG_7__SCAN_IN ; U618
g413 nand DATAI_6_ U248 ; U619
g414 nand R165_U6 BUF1_REG_6__SCAN_IN ; U620
g415 nand DATAI_5_ U248 ; U621
g416 nand R165_U6 BUF1_REG_5__SCAN_IN ; U622
g417 nand DATAI_4_ U248 ; U623
g418 nand R165_U6 BUF1_REG_4__SCAN_IN ; U624
g419 nand DATAI_3_ U248 ; U625
g420 nand R165_U6 BUF1_REG_3__SCAN_IN ; U626
g421 nand DATAI_31_ U248 ; U627
g422 nand R165_U6 BUF1_REG_31__SCAN_IN ; U628
g423 nand DATAI_30_ U248 ; U629
g424 nand R165_U6 BUF1_REG_30__SCAN_IN ; U630
g425 nand DATAI_2_ U248 ; U631
g426 nand R165_U6 BUF1_REG_2__SCAN_IN ; U632
g427 nand DATAI_29_ U248 ; U633
g428 nand R165_U6 BUF1_REG_29__SCAN_IN ; U634
g429 nand DATAI_28_ U248 ; U635
g430 nand R165_U6 BUF1_REG_28__SCAN_IN ; U636
g431 nand DATAI_27_ U248 ; U637
g432 nand R165_U6 BUF1_REG_27__SCAN_IN ; U638
g433 nand DATAI_26_ U248 ; U639
g434 nand R165_U6 BUF1_REG_26__SCAN_IN ; U640
g435 nand DATAI_25_ U248 ; U641
g436 nand R165_U6 BUF1_REG_25__SCAN_IN ; U642
g437 nand DATAI_24_ U248 ; U643
g438 nand R165_U6 BUF1_REG_24__SCAN_IN ; U644
g439 nand DATAI_23_ U248 ; U645
g440 nand R165_U6 BUF1_REG_23__SCAN_IN ; U646
g441 nand DATAI_22_ U248 ; U647
g442 nand R165_U6 BUF1_REG_22__SCAN_IN ; U648
g443 nand DATAI_21_ U248 ; U649
g444 nand R165_U6 BUF1_REG_21__SCAN_IN ; U650
g445 nand DATAI_20_ U248 ; U651
g446 nand R165_U6 BUF1_REG_20__SCAN_IN ; U652
g447 nand DATAI_1_ U248 ; U653
g448 nand R165_U6 BUF1_REG_1__SCAN_IN ; U654
g449 nand DATAI_19_ U248 ; U655
g450 nand R165_U6 BUF1_REG_19__SCAN_IN ; U656
g451 nand DATAI_18_ U248 ; U657
g452 nand R165_U6 BUF1_REG_18__SCAN_IN ; U658
g453 nand DATAI_17_ U248 ; U659
g454 nand R165_U6 BUF1_REG_17__SCAN_IN ; U660
g455 nand DATAI_16_ U248 ; U661
g456 nand R165_U6 BUF1_REG_16__SCAN_IN ; U662
g457 nand DATAI_15_ U248 ; U663
g458 nand R165_U6 BUF1_REG_15__SCAN_IN ; U664
g459 nand DATAI_14_ U248 ; U665
g460 nand R165_U6 BUF1_REG_14__SCAN_IN ; U666
g461 nand DATAI_13_ U248 ; U667
g462 nand R165_U6 BUF1_REG_13__SCAN_IN ; U668
g463 nand DATAI_12_ U248 ; U669
g464 nand R165_U6 BUF1_REG_12__SCAN_IN ; U670
g465 nand DATAI_11_ U248 ; U671
g466 nand R165_U6 BUF1_REG_11__SCAN_IN ; U672
g467 nand DATAI_10_ U248 ; U673
g468 nand R165_U6 BUF1_REG_10__SCAN_IN ; U674
g469 nand DATAI_0_ U248 ; U675
g470 nand R165_U6 BUF1_REG_0__SCAN_IN ; U676
g471 nand U382 P2_ADDRESS_REG_9__SCAN_IN ; U677
g472 nand U384 P3_ADDRESS_REG_9__SCAN_IN ; U678
g473 nand U382 P2_ADDRESS_REG_8__SCAN_IN ; U679
g474 nand U384 P3_ADDRESS_REG_8__SCAN_IN ; U680
g475 nand U382 P2_ADDRESS_REG_7__SCAN_IN ; U681
g476 nand U384 P3_ADDRESS_REG_7__SCAN_IN ; U682
g477 nand U382 P2_ADDRESS_REG_6__SCAN_IN ; U683
g478 nand U384 P3_ADDRESS_REG_6__SCAN_IN ; U684
g479 nand U382 P2_ADDRESS_REG_5__SCAN_IN ; U685
g480 nand U384 P3_ADDRESS_REG_5__SCAN_IN ; U686
g481 nand U382 P2_ADDRESS_REG_4__SCAN_IN ; U687
g482 nand U384 P3_ADDRESS_REG_4__SCAN_IN ; U688
g483 nand U382 P2_ADDRESS_REG_3__SCAN_IN ; U689
g484 nand U384 P3_ADDRESS_REG_3__SCAN_IN ; U690
g485 nand U382 P2_ADDRESS_REG_2__SCAN_IN ; U691
g486 nand U384 P3_ADDRESS_REG_2__SCAN_IN ; U692
g487 nand U382 P2_ADDRESS_REG_29__SCAN_IN ; U693
g488 nand U384 P3_ADDRESS_REG_29__SCAN_IN ; U694
g489 nand U382 P2_ADDRESS_REG_28__SCAN_IN ; U695
g490 nand U384 P3_ADDRESS_REG_28__SCAN_IN ; U696
g491 nand U382 P2_ADDRESS_REG_27__SCAN_IN ; U697
g492 nand U384 P3_ADDRESS_REG_27__SCAN_IN ; U698
g493 nand U382 P2_ADDRESS_REG_26__SCAN_IN ; U699
g494 nand U384 P3_ADDRESS_REG_26__SCAN_IN ; U700
g495 nand U382 P2_ADDRESS_REG_25__SCAN_IN ; U701
g496 nand U384 P3_ADDRESS_REG_25__SCAN_IN ; U702
g497 nand U382 P2_ADDRESS_REG_24__SCAN_IN ; U703
g498 nand U384 P3_ADDRESS_REG_24__SCAN_IN ; U704
g499 nand U382 P2_ADDRESS_REG_23__SCAN_IN ; U705
g500 nand U384 P3_ADDRESS_REG_23__SCAN_IN ; U706
g501 nand U382 P2_ADDRESS_REG_22__SCAN_IN ; U707
g502 nand U384 P3_ADDRESS_REG_22__SCAN_IN ; U708
g503 nand U382 P2_ADDRESS_REG_21__SCAN_IN ; U709
g504 nand U384 P3_ADDRESS_REG_21__SCAN_IN ; U710
g505 nand U382 P2_ADDRESS_REG_20__SCAN_IN ; U711
g506 nand U384 P3_ADDRESS_REG_20__SCAN_IN ; U712
g507 nand U382 P2_ADDRESS_REG_1__SCAN_IN ; U713
g508 nand U384 P3_ADDRESS_REG_1__SCAN_IN ; U714
g509 nand U382 P2_ADDRESS_REG_19__SCAN_IN ; U715
g510 nand U384 P3_ADDRESS_REG_19__SCAN_IN ; U716
g511 nand U382 P2_ADDRESS_REG_18__SCAN_IN ; U717
g512 nand U384 P3_ADDRESS_REG_18__SCAN_IN ; U718
g513 nand U382 P2_ADDRESS_REG_17__SCAN_IN ; U719
g514 nand U384 P3_ADDRESS_REG_17__SCAN_IN ; U720
g515 nand U382 P2_ADDRESS_REG_16__SCAN_IN ; U721
g516 nand U384 P3_ADDRESS_REG_16__SCAN_IN ; U722
g517 nand U382 P2_ADDRESS_REG_15__SCAN_IN ; U723
g518 nand U384 P3_ADDRESS_REG_15__SCAN_IN ; U724
g519 nand U382 P2_ADDRESS_REG_14__SCAN_IN ; U725
g520 nand U384 P3_ADDRESS_REG_14__SCAN_IN ; U726
g521 nand U382 P2_ADDRESS_REG_13__SCAN_IN ; U727
g522 nand U384 P3_ADDRESS_REG_13__SCAN_IN ; U728
g523 nand U382 P2_ADDRESS_REG_12__SCAN_IN ; U729
g524 nand U384 P3_ADDRESS_REG_12__SCAN_IN ; U730
g525 nand U382 P2_ADDRESS_REG_11__SCAN_IN ; U731
g526 nand U384 P3_ADDRESS_REG_11__SCAN_IN ; U732
g527 nand U382 P2_ADDRESS_REG_10__SCAN_IN ; U733
g528 nand U384 P3_ADDRESS_REG_10__SCAN_IN ; U734
g529 nand U382 P2_ADDRESS_REG_0__SCAN_IN ; U735
g530 nand U384 P3_ADDRESS_REG_0__SCAN_IN ; U736
g531 nor U209 P3_STATEBS16_REG_SCAN_IN ; P3_U2352
g532 and P3_U3354 P3_U2449 ; P3_U2353
g533 and P3_U3688 P3_U4325 ; P3_U2354
g534 and P3_U3689 P3_U4325 ; P3_U2355
g535 and P3_U3355 P3_U2353 ; P3_U2356
g536 and P3_U4323 P3_U2451 ; P3_U2357
g537 and P3_U3690 P3_U4341 ; P3_U2358
g538 and P3_U4324 P3_U2462 ; P3_U2359
g539 and P3_U4296 P3_U2462 ; P3_U2360
g540 and P3_U4297 P3_U2462 ; P3_U2361
g541 and P3_U3691 P3_U4341 ; P3_U2362
g542 and P3_U5442 P3_U5435 ; P3_U2363
g543 and P3_U5392 P3_U3204 ; P3_U2364
g544 and P3_U5341 P3_U3201 ; P3_U2365
g545 and P3_U5290 P3_U3198 ; P3_U2366
g546 and P3_U5239 P3_U5232 ; P3_U2367
g547 and P3_U5189 P3_U3193 ; P3_U2368
g548 and P3_U5137 P3_U3189 ; P3_U2369
g549 and P3_U5085 P3_U3185 ; P3_U2370
g550 and P3_U5036 P3_U5028 ; P3_U2371
g551 and P3_U4985 P3_U3176 ; P3_U2372
g552 and P3_U4933 P3_U3172 ; P3_U2373
g553 and P3_U4881 P3_U3168 ; P3_U2374
g554 and P3_U4829 P3_U4821 ; P3_U2375
g555 and P3_U4778 P3_U3160 ; P3_U2376
g556 and P3_U4726 P3_U3152 ; P3_U2377
g557 and P3_U4674 P3_U3146 ; P3_U2378
g558 and P3_U4322 P3_U4312 ; P3_U2379
g559 and P3_U3260 P3_STATE2_REG_2__SCAN_IN ; P3_U2380
g560 and P3_U4312 P3_STATE2_REG_3__SCAN_IN ; P3_U2381
g561 and P3_U3951 P3_U3249 ; P3_U2382
g562 and P3_U2380 P3_U4296 ; P3_U2383
g563 and P3_U2380 P3_U4297 ; P3_U2384
g564 and P3_U3260 P3_STATE2_REG_1__SCAN_IN ; P3_U2385
g565 and P3_U3249 P3_STATE2_REG_1__SCAN_IN ; P3_U2386
g566 and P3_U3953 P3_U3249 ; P3_U2387
g567 and P3_U3952 P3_U3249 ; P3_U2388
g568 and P3_U4354 P3_U3249 ; P3_U2389
g569 and P3_U4353 P3_STATE2_REG_0__SCAN_IN ; P3_U2390
g570 and P3_U4310 P3_U3218 ; P3_U2391
g571 and P3_U2383 P3_U4293 ; P3_U2392
g572 and P3_U2628 P3_U2361 ; P3_U2393
g573 and P3_U2382 P3_U2628 ; P3_U2394
g574 and P3_U2361 P3_U3241 ; P3_U2395
g575 and P3_U2382 P3_U3241 ; P3_U2396
g576 and P3_U2386 P3_STATEBS16_REG_SCAN_IN ; P3_U2397
g577 and P3_U2386 P3_U2631 ; P3_U2398
g578 and P3_U4309 P3_U4573 ; P3_U2399
g579 and P3_U4310 P3_U4573 ; P3_U2400
g580 and P3_U3260 P3_STATE2_REG_3__SCAN_IN ; P3_U2401
g581 and P3_U3248 P3_U3090 ; P3_U2402
g582 and P3_U2385 P3_U3258 ; P3_U2403
g583 and P3_U2384 P3_U3257 ; P3_U2404
g584 and P3_U7095 P3_U2384 ; P3_U2405
g585 and P3_U4311 P3_U3104 ; P3_U2406
g586 and P3_U4311 P3_U4505 ; P3_U2407
g587 and P3_U4309 P3_U3218 ; P3_U2408
g588 and P3_U3251 P3_STATE2_REG_0__SCAN_IN ; P3_U2409
g589 and P3_U3251 P3_U3121 ; P3_U2410
g590 and P3_U4310 P3_U4608 ; P3_U2411
g591 and P3_U3218 P3_U3107 P3_U4539 ; P3_U2412
g592 and P3_U4312 BUF2_REG_0__SCAN_IN ; P3_U2413
g593 and P3_U4312 BUF2_REG_1__SCAN_IN ; P3_U2414
g594 and P3_U4312 BUF2_REG_2__SCAN_IN ; P3_U2415
g595 and P3_U4312 BUF2_REG_3__SCAN_IN ; P3_U2416
g596 and P3_U4312 BUF2_REG_4__SCAN_IN ; P3_U2417
g597 and P3_U4312 BUF2_REG_5__SCAN_IN ; P3_U2418
g598 and P3_U4312 BUF2_REG_6__SCAN_IN ; P3_U2419
g599 and P3_U4312 BUF2_REG_7__SCAN_IN ; P3_U2420
g600 and P3_U2379 BUF2_REG_24__SCAN_IN ; P3_U2421
g601 and P3_U2379 BUF2_REG_16__SCAN_IN ; P3_U2422
g602 and P3_U2379 BUF2_REG_25__SCAN_IN ; P3_U2423
g603 and P3_U2379 BUF2_REG_17__SCAN_IN ; P3_U2424
g604 and P3_U2379 BUF2_REG_26__SCAN_IN ; P3_U2425
g605 and P3_U2379 BUF2_REG_18__SCAN_IN ; P3_U2426
g606 and P3_U2379 BUF2_REG_27__SCAN_IN ; P3_U2427
g607 and P3_U2379 BUF2_REG_19__SCAN_IN ; P3_U2428
g608 and P3_U2379 BUF2_REG_28__SCAN_IN ; P3_U2429
g609 and P3_U2379 BUF2_REG_20__SCAN_IN ; P3_U2430
g610 and P3_U2379 BUF2_REG_29__SCAN_IN ; P3_U2431
g611 and P3_U2379 BUF2_REG_21__SCAN_IN ; P3_U2432
g612 and P3_U2379 BUF2_REG_30__SCAN_IN ; P3_U2433
g613 and P3_U2379 BUF2_REG_22__SCAN_IN ; P3_U2434
g614 and P3_U2379 BUF2_REG_31__SCAN_IN ; P3_U2435
g615 and P3_U2379 BUF2_REG_23__SCAN_IN ; P3_U2436
g616 and P3_U2381 P3_U3108 ; P3_U2437
g617 and P3_U2381 P3_U3104 ; P3_U2438
g618 and P3_U2381 P3_U3101 ; P3_U2439
g619 and P3_U2381 P3_U3107 ; P3_U2440
g620 and P3_U2381 P3_U3102 ; P3_U2441
g621 and P3_U2381 P3_U3110 ; P3_U2442
g622 and P3_U2381 P3_U3074 ; P3_U2443
g623 and P3_U2391 P3_U3074 ; P3_U2444
g624 and P3_U2381 P3_U3218 ; P3_U2445
g625 and P3_U2391 P3_U3113 ; P3_U2446
g626 and P3_U2409 P3_U3108 ; P3_U2447
g627 and P3_U2391 P3_U4590 ; P3_U2448
g628 and P3_U4344 P3_U4522 ; P3_U2449
g629 and P3_U3660 P3_U4351 ; P3_U2450
g630 and P3_U4608 P3_U3102 P3_U2412 ; P3_U2451
g631 and P3_U2463 P3_U4522 P3_U2412 ; P3_U2452
g632 and P3_STATE2_REG_2__SCAN_IN P3_STATE2_REG_1__SCAN_IN ; P3_U2453
g633 and P3_U2380 P3_U4323 ; P3_U2454
g634 and P3_U2380 P3_U4324 ; P3_U2455
g635 and P3_U4556 P3_U4607 ; P3_U2456
g636 and P3_U3269 P3_U3139 ; P3_U2457
g637 and P3_U4652 P3_U3269 ; P3_U2458
g638 and P3_U7962 P3_U3139 ; P3_U2459
g639 and P3_U7962 P3_U4652 ; P3_U2460
g640 and P3_U4573 P3_U4522 ; P3_U2461
g641 and P3_U2412 P3_U2449 ; P3_U2462
g642 and P3_U4590 P3_U4607 ; P3_U2463
g643 and P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U2464
g644 and P3_U2464 P3_U4332 ; P3_U2465
g645 and P3_U3093 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U2466
g646 and P3_U2464 P3_U2466 ; P3_U2467
g647 and P3_U3094 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U2468
g648 and P3_U2464 P3_U2468 ; P3_U2469
g649 and P3_U2464 P3_U4467 ; P3_U2470
g650 and P3_U4468 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U2471
g651 and P3_U2466 P3_U3097 ; P3_U2472
g652 and P3_U2472 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U2473
g653 and P3_U2468 P3_U3097 ; P3_U2474
g654 and P3_U2474 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U2475
g655 and P3_U4469 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U2476
g656 and P3_U4470 P3_U2466 ; P3_U2477
g657 and P3_U4470 P3_U2468 ; P3_U2478
g658 and P3_U4470 P3_U4467 ; P3_U2479
g659 and P3_U4468 P3_U3100 ; P3_U2480
g660 nor P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U2481
g661 and P3_U2466 P3_U2481 ; P3_U2482
g662 and P3_U2468 P3_U2481 ; P3_U2483
g663 and P3_U4469 P3_U3100 ; P3_U2484
g664 and P3_U4656 P3_U3270 ; P3_U2485
g665 and P3_U3271 P3_U3182 ; P3_U2486
g666 and P3_U3270 P3_U3142 ; P3_U2487
g667 and P3_U4657 P3_U2487 ; P3_U2488
g668 and P3_U3090 P3_U4315 ; P3_U2489
g669 and P3_U3156 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U2490
g670 and P3_U4644 P3_U2487 ; P3_U2491
g671 and P3_U3128 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U2492
g672 and P3_U4646 P3_U3128 ; P3_U2493
g673 and P3_U4645 P3_U2487 ; P3_U2494
g674 and P3_U4646 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U2495
g675 and P3_U4643 P3_U3128 ; P3_U2496
g676 and P3_U2496 P3_U2487 ; P3_U2497
g677 and P3_U7968 P3_U3182 ; P3_U2498
g678 and P3_U4658 P3_U4657 ; P3_U2499
g679 and P3_U4658 P3_U4644 ; P3_U2500
g680 nor P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U2501
g681 and P3_U4658 P3_U4645 ; P3_U2502
g682 and P3_U4658 P3_U2496 ; P3_U2503
g683 and P3_U4660 P3_U3271 ; P3_U2504
g684 and P3_U4644 P3_U2485 ; P3_U2505
g685 and P3_U4645 P3_U2485 ; P3_U2506
g686 and P3_U2496 P3_U2485 ; P3_U2507
g687 and P3_U4660 P3_U7968 ; P3_U2508
g688 and P3_U7965 P3_U4656 ; P3_U2509
g689 and P3_U2509 P3_U4657 ; P3_U2510
g690 and P3_U2509 P3_U4644 ; P3_U2511
g691 and P3_U2509 P3_U4645 ; P3_U2512
g692 and P3_U2509 P3_U2496 ; P3_U2513
g693 and P3_U3218 P3_U3216 ; P3_U2514
g694 and P3_U7970 P3_U7969 P3_U5485 ; P3_U2515
g695 and P3_U5493 P3_U5492 ; P3_U2516
g696 and P3_U3246 P3_U5526 ; P3_U2517
g697 and P3_U3668 P3_U5522 ; P3_U2518
g698 and P3_U3228 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U2519
g699 and P3_U5543 P3_U5548 ; P3_U2520
g700 and P3_U2520 P3_U2519 ; P3_U2521
g701 and P3_U3093 P3_U3228 ; P3_U2522
g702 and P3_U2520 P3_U2522 ; P3_U2523
g703 and P3_U5558 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U2524
g704 and P3_U2520 P3_U2524 ; P3_U2525
g705 and P3_U5558 P3_U3093 ; P3_U2526
g706 and P3_U2520 P3_U2526 ; P3_U2527
g707 and P3_U5543 P3_U3225 ; P3_U2528
g708 and P3_U2528 P3_U2519 ; P3_U2529
g709 and P3_U2528 P3_U2522 ; P3_U2530
g710 and P3_U2528 P3_U2524 ; P3_U2531
g711 and P3_U2528 P3_U2526 ; P3_U2532
g712 and P3_U5548 P3_U3265 ; P3_U2533
g713 and P3_U2533 P3_U2519 ; P3_U2534
g714 and P3_U2533 P3_U2522 ; P3_U2535
g715 and P3_U2533 P3_U2524 ; P3_U2536
g716 and P3_U2533 P3_U2526 ; P3_U2537
g717 and P3_U3265 P3_U3225 ; P3_U2538
g718 and P3_U2519 P3_U2538 ; P3_U2539
g719 and P3_U2522 P3_U2538 ; P3_U2540
g720 and P3_U2524 P3_U2538 ; P3_U2541
g721 and P3_U2526 P3_U2538 ; P3_U2542
g722 and P3_U3272 P3_U3266 ; P3_U2543
g723 and P3_U2543 P3_U2468 ; P3_U2544
g724 and P3_U2543 P3_U4467 ; P3_U2545
g725 and P3_U2543 P3_U4332 ; P3_U2546
g726 and P3_U2543 P3_U2466 ; P3_U2547
g727 and P3_U8034 P3_U3266 ; P3_U2548
g728 and P3_U2548 P3_U2468 ; P3_U2549
g729 and P3_U2548 P3_U4467 ; P3_U2550
g730 and P3_U2548 P3_U4332 ; P3_U2551
g731 and P3_U2548 P3_U2466 ; P3_U2552
g732 and P3_U7516 P3_U3272 ; P3_U2553
g733 and P3_U2553 P3_U2468 ; P3_U2554
g734 and P3_U2553 P3_U4467 ; P3_U2555
g735 and P3_U2553 P3_U4332 ; P3_U2556
g736 and P3_U2553 P3_U2466 ; P3_U2557
g737 and P3_U7516 P3_U8034 ; P3_U2558
g738 and P3_U2558 P3_U2468 ; P3_U2559
g739 and P3_U2558 P3_U4467 ; P3_U2560
g740 and P3_U2558 P3_U4332 ; P3_U2561
g741 and P3_U2558 P3_U2466 ; P3_U2562
g742 and P3_U8037 P3_U4291 ; P3_U2563
g743 and P3_U2563 P3_U2522 ; P3_U2564
g744 and P3_U2563 P3_U2519 ; P3_U2565
g745 and P3_U2563 P3_U2526 ; P3_U2566
g746 and P3_U2563 P3_U2524 ; P3_U2567
g747 and P3_U8037 P3_U3267 ; P3_U2568
g748 and P3_U2568 P3_U2522 ; P3_U2569
g749 and P3_U2568 P3_U2519 ; P3_U2570
g750 and P3_U2568 P3_U2526 ; P3_U2571
g751 and P3_U2568 P3_U2524 ; P3_U2572
g752 and P3_U4291 P3_U3273 ; P3_U2573
g753 and P3_U2573 P3_U2522 ; P3_U2574
g754 and P3_U2573 P3_U2519 ; P3_U2575
g755 and P3_U2573 P3_U2526 ; P3_U2576
g756 and P3_U2573 P3_U2524 ; P3_U2577
g757 and P3_U3273 P3_U3267 ; P3_U2578
g758 and P3_U2578 P3_U2522 ; P3_U2579
g759 and P3_U2578 P3_U2519 ; P3_U2580
g760 and P3_U2578 P3_U2526 ; P3_U2581
g761 and P3_U2578 P3_U2524 ; P3_U2582
g762 and P3_U7775 P3_U4468 ; P3_U2583
g763 and P3_U7775 P3_U2472 ; P3_U2584
g764 and P3_U7775 P3_U2474 ; P3_U2585
g765 and P3_U7775 P3_U4469 ; P3_U2586
g766 and P3_U7775 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U2587
g767 and P3_U2587 P3_U4332 ; P3_U2588
g768 and P3_U2587 P3_U2466 ; P3_U2589
g769 and P3_U2587 P3_U2468 ; P3_U2590
g770 and P3_U2587 P3_U4467 ; P3_U2591
g771 and P3_U4468 P3_U3268 ; P3_U2592
g772 and P3_U2472 P3_U3268 ; P3_U2593
g773 and P3_U2474 P3_U3268 ; P3_U2594
g774 and P3_U4469 P3_U3268 ; P3_U2595
g775 and P3_U3268 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U2596
g776 and P3_U2596 P3_U4332 ; P3_U2597
g777 and P3_U2596 P3_U2466 ; P3_U2598
g778 and P3_U2596 P3_U2468 ; P3_U2599
g779 and P3_U2596 P3_U4467 ; P3_U2600
g780 and P3_U2392 P3_U2352 ; P3_U2601
g781 and P3_U2404 P3_EBX_REG_31__SCAN_IN ; P3_U2602
g782 and P3_U7360 P3_U7358 P3_U7359 P3_U4133 ; P3_U2603
g783 and P3_U7947 P3_U7946 ; P3_U2604
g784 nand P3_U4215 P3_U4214 P3_U4213 P3_U4212 ; P3_U2605
g785 nand P3_U4211 P3_U4210 P3_U4209 P3_U4208 ; P3_U2606
g786 nand P3_U4207 P3_U4206 P3_U4205 P3_U4204 ; P3_U2607
g787 nand P3_U4203 P3_U4202 P3_U4201 P3_U4200 ; P3_U2608
g788 nand P3_U4199 P3_U4198 P3_U4197 P3_U4196 ; P3_U2609
g789 nand P3_U4195 P3_U4194 P3_U4193 P3_U4192 ; P3_U2610
g790 nand P3_U4191 P3_U4190 P3_U4189 P3_U4188 ; P3_U2611
g791 nand P3_U4187 P3_U4186 P3_U4185 P3_U4184 ; P3_U2612
g792 nand P3_U4279 P3_U4278 P3_U4277 P3_U4276 ; P3_U2613
g793 nand P3_U4275 P3_U4274 P3_U4273 P3_U4272 ; P3_U2614
g794 nand P3_U4271 P3_U4270 P3_U4269 P3_U4268 ; P3_U2615
g795 nand P3_U4267 P3_U4266 P3_U4265 P3_U4264 ; P3_U2616
g796 nand P3_U4263 P3_U4262 P3_U4261 P3_U4260 ; P3_U2617
g797 nand P3_U4259 P3_U4258 P3_U4257 P3_U4256 ; P3_U2618
g798 nand P3_U4255 P3_U4254 P3_U4253 P3_U4252 ; P3_U2619
g799 nand P3_U4251 P3_U4250 P3_U4249 P3_U4248 ; P3_U2620
g800 nand P3_U4183 P3_U4182 P3_U4181 P3_U4180 ; P3_U2621
g801 nand P3_U4179 P3_U4178 P3_U4177 P3_U4176 ; P3_U2622
g802 nand P3_U4175 P3_U4174 P3_U4173 P3_U4172 ; P3_U2623
g803 nand P3_U4171 P3_U4170 P3_U4169 P3_U4168 ; P3_U2624
g804 nand P3_U4167 P3_U4166 P3_U4165 P3_U4164 ; P3_U2625
g805 nand P3_U4163 P3_U4162 P3_U4161 P3_U4160 ; P3_U2626
g806 nand P3_U4159 P3_U4158 P3_U4157 P3_U4156 ; P3_U2627
g807 nand P3_U4155 P3_U4154 P3_U4153 P3_U4152 ; P3_U2628
g808 and P3_U3207 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_U2629
g809 not U209 ; P3_U2630
g810 not P3_STATEBS16_REG_SCAN_IN ; P3_U2631
g811 and P3_U3207 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U2632
g812 nand P3_U7937 P3_U7383 ; P3_U2633
g813 nand P3_U7382 P3_U7381 ; P3_U2634
g814 nand P3_U8025 P3_U8024 P3_U4335 ; P3_U2635
g815 nand P3_U8021 P3_U8020 P3_U4335 ; P3_U2636
g816 nand P3_U7370 P3_U7369 ; P3_U2637
g817 nand P3_U8013 P3_U8012 P3_U4327 ; P3_U2638
g818 nand P3_U8003 P3_U8002 P3_U4327 ; P3_U2639
g819 and P3_U7357 P3_U7907 ; P3_U2640
g820 nand P3_U7352 P3_U7351 P3_U4129 P3_U7354 P3_U4130 ; P3_U2641
g821 nand P3_U7344 P3_U7343 P3_U4126 P3_U7346 P3_U4127 ; P3_U2642
g822 nand P3_U7336 P3_U7335 P3_U4123 P3_U7338 P3_U4124 ; P3_U2643
g823 nand P3_U7328 P3_U7327 P3_U4120 P3_U7330 P3_U4121 ; P3_U2644
g824 nand P3_U7320 P3_U7319 P3_U4117 P3_U7322 P3_U4118 ; P3_U2645
g825 nand P3_U7312 P3_U7311 P3_U4114 P3_U7314 P3_U4115 ; P3_U2646
g826 nand P3_U7304 P3_U7303 P3_U4111 P3_U7306 P3_U4112 ; P3_U2647
g827 nand P3_U7296 P3_U7295 P3_U4108 P3_U7298 P3_U4109 ; P3_U2648
g828 nand P3_U7288 P3_U7287 P3_U4105 P3_U7290 P3_U4106 ; P3_U2649
g829 nand P3_U7280 P3_U7279 P3_U4102 P3_U7282 P3_U4103 ; P3_U2650
g830 nand P3_U7272 P3_U7271 P3_U4099 P3_U7274 P3_U4100 ; P3_U2651
g831 nand P3_U7264 P3_U7263 P3_U4096 P3_U7266 P3_U4097 ; P3_U2652
g832 nand P3_U7256 P3_U7255 P3_U4093 P3_U7258 P3_U4094 ; P3_U2653
g833 nand P3_U7248 P3_U7247 P3_U4090 P3_U7250 P3_U4091 ; P3_U2654
g834 nand P3_U7240 P3_U7239 P3_U4087 P3_U7242 P3_U4088 ; P3_U2655
g835 nand P3_U7232 P3_U7231 P3_U4084 P3_U7234 P3_U4085 ; P3_U2656
g836 nand P3_U7224 P3_U7223 P3_U4081 P3_U7226 P3_U4082 ; P3_U2657
g837 nand P3_U7216 P3_U7215 P3_U4078 P3_U7218 P3_U4079 ; P3_U2658
g838 nand P3_U7208 P3_U7207 P3_U4075 P3_U7210 P3_U4076 ; P3_U2659
g839 nand P3_U7200 P3_U7199 P3_U4072 P3_U7202 P3_U4073 ; P3_U2660
g840 nand P3_U7192 P3_U7191 P3_U4069 P3_U7194 P3_U4070 ; P3_U2661
g841 nand P3_U7184 P3_U7183 P3_U4066 P3_U7186 P3_U4067 ; P3_U2662
g842 nand P3_U7176 P3_U7175 P3_U4063 P3_U7178 P3_U4064 ; P3_U2663
g843 nand P3_U7168 P3_U7167 P3_U4060 P3_U7170 P3_U4061 ; P3_U2664
g844 nand P3_U7160 P3_U7159 P3_U4057 P3_U7162 P3_U4058 ; P3_U2665
g845 nand P3_U4056 P3_U4054 ; P3_U2666
g846 nand P3_U4051 P3_U4049 ; P3_U2667
g847 nand P3_U7129 P3_U4043 P3_U7132 P3_U7133 P3_U4045 ; P3_U2668
g848 nand P3_U7119 P3_U4039 P3_U7122 P3_U7123 P3_U4041 ; P3_U2669
g849 nand P3_U7109 P3_U4035 P3_U7112 P3_U7113 P3_U4037 ; P3_U2670
g850 nand P3_U7099 P3_U4031 P3_U7102 P3_U7103 P3_U4033 ; P3_U2671
g851 nand P3_U7092 P3_U7091 ; P3_U2672
g852 nand P3_U7090 P3_U7088 P3_U7089 ; P3_U2673
g853 nand P3_U7087 P3_U7085 P3_U7086 ; P3_U2674
g854 nand P3_U7084 P3_U7082 P3_U7083 ; P3_U2675
g855 nand P3_U7081 P3_U7079 P3_U7080 ; P3_U2676
g856 nand P3_U7078 P3_U7076 P3_U7077 ; P3_U2677
g857 nand P3_U7075 P3_U7073 P3_U7074 ; P3_U2678
g858 nand P3_U7072 P3_U7070 P3_U7071 ; P3_U2679
g859 nand P3_U7069 P3_U7067 P3_U7068 ; P3_U2680
g860 nand P3_U7066 P3_U7064 P3_U7065 ; P3_U2681
g861 nand P3_U7063 P3_U7061 P3_U7062 ; P3_U2682
g862 nand P3_U7060 P3_U7058 P3_U7059 ; P3_U2683
g863 nand P3_U7057 P3_U7055 P3_U7056 ; P3_U2684
g864 nand P3_U7054 P3_U7052 P3_U7053 ; P3_U2685
g865 nand P3_U7051 P3_U7049 P3_U7050 ; P3_U2686
g866 nand P3_U7048 P3_U7046 P3_U7047 ; P3_U2687
g867 nand P3_U7045 P3_U7043 P3_U7044 ; P3_U2688
g868 nand P3_U7042 P3_U7040 P3_U7041 ; P3_U2689
g869 nand P3_U7039 P3_U7037 P3_U7038 ; P3_U2690
g870 nand P3_U7036 P3_U7034 P3_U7035 ; P3_U2691
g871 nand P3_U7033 P3_U7031 P3_U7032 ; P3_U2692
g872 nand P3_U7030 P3_U7028 P3_U7029 ; P3_U2693
g873 nand P3_U7026 P3_U7025 P3_U7027 ; P3_U2694
g874 nand P3_U7023 P3_U7022 P3_U7024 ; P3_U2695
g875 nand P3_U7020 P3_U7019 P3_U7021 ; P3_U2696
g876 nand P3_U7017 P3_U7016 P3_U7018 ; P3_U2697
g877 nand P3_U7014 P3_U7013 P3_U7015 ; P3_U2698
g878 nand P3_U7011 P3_U7010 P3_U7012 ; P3_U2699
g879 nand P3_U7008 P3_U7007 P3_U7009 ; P3_U2700
g880 nand P3_U7005 P3_U7004 P3_U7006 ; P3_U2701
g881 nand P3_U7002 P3_U7001 P3_U7003 ; P3_U2702
g882 nand P3_U6999 P3_U6998 P3_U7000 ; P3_U2703
g883 nand P3_U6995 P3_U6993 P3_U6994 ; P3_U2704
g884 nand P3_U6989 P3_U6988 P3_U6992 P3_U6990 P3_U6991 ; P3_U2705
g885 nand P3_U6984 P3_U6983 P3_U6987 P3_U6985 P3_U6986 ; P3_U2706
g886 nand P3_U6979 P3_U6978 P3_U6982 P3_U6980 P3_U6981 ; P3_U2707
g887 nand P3_U6974 P3_U6973 P3_U4029 P3_U6976 ; P3_U2708
g888 nand P3_U6969 P3_U6968 P3_U4028 P3_U6971 ; P3_U2709
g889 nand P3_U6964 P3_U6963 P3_U4027 P3_U6966 ; P3_U2710
g890 nand P3_U6959 P3_U6958 P3_U4026 P3_U6961 ; P3_U2711
g891 nand P3_U6954 P3_U6953 P3_U4025 P3_U6956 ; P3_U2712
g892 nand P3_U6949 P3_U6948 P3_U4024 P3_U6951 ; P3_U2713
g893 nand P3_U6944 P3_U6943 P3_U4023 P3_U6946 ; P3_U2714
g894 nand P3_U6939 P3_U6938 P3_U4022 P3_U6941 ; P3_U2715
g895 nand P3_U6934 P3_U6933 P3_U4021 P3_U6936 ; P3_U2716
g896 nand P3_U6929 P3_U6928 P3_U4020 P3_U6931 ; P3_U2717
g897 nand P3_U6924 P3_U6923 P3_U4019 P3_U6926 ; P3_U2718
g898 nand P3_U6919 P3_U6918 P3_U4018 P3_U6921 ; P3_U2719
g899 nand P3_U6914 P3_U4017 P3_U6916 ; P3_U2720
g900 nand P3_U6910 P3_U4016 P3_U6912 ; P3_U2721
g901 nand P3_U6906 P3_U4015 P3_U6908 ; P3_U2722
g902 nand P3_U6903 P3_U6902 P3_U4014 ; P3_U2723
g903 nand P3_U6899 P3_U6898 P3_U4013 ; P3_U2724
g904 nand P3_U6895 P3_U6894 P3_U4012 ; P3_U2725
g905 nand P3_U6891 P3_U6890 P3_U4011 ; P3_U2726
g906 nand P3_U6887 P3_U6886 P3_U4010 ; P3_U2727
g907 nand P3_U6883 P3_U6882 P3_U4009 ; P3_U2728
g908 nand P3_U6879 P3_U6878 P3_U4008 ; P3_U2729
g909 nand P3_U6875 P3_U6874 P3_U4007 ; P3_U2730
g910 nand P3_U6871 P3_U6870 P3_U4006 ; P3_U2731
g911 nand P3_U6867 P3_U6866 P3_U4005 ; P3_U2732
g912 nand P3_U6863 P3_U6862 P3_U4004 ; P3_U2733
g913 nand P3_U6859 P3_U6858 P3_U4003 ; P3_U2734
g914 nand P3_U6855 P3_U6854 P3_U4002 ; P3_U2735
g915 and P3_U6759 P3_DATAO_REG_31__SCAN_IN ; P3_U2736
g916 nand P3_U4001 P3_U6850 ; P3_U2737
g917 nand P3_U4000 P3_U6847 ; P3_U2738
g918 nand P3_U3999 P3_U6844 ; P3_U2739
g919 nand P3_U3998 P3_U6841 ; P3_U2740
g920 nand P3_U3997 P3_U6838 ; P3_U2741
g921 nand P3_U3996 P3_U6835 ; P3_U2742
g922 nand P3_U3995 P3_U6832 ; P3_U2743
g923 nand P3_U3994 P3_U6829 ; P3_U2744
g924 nand P3_U3993 P3_U6826 ; P3_U2745
g925 nand P3_U3992 P3_U6823 ; P3_U2746
g926 nand P3_U3991 P3_U6820 ; P3_U2747
g927 nand P3_U3990 P3_U6817 ; P3_U2748
g928 nand P3_U3989 P3_U6814 ; P3_U2749
g929 nand P3_U3988 P3_U6811 ; P3_U2750
g930 nand P3_U3987 P3_U6808 ; P3_U2751
g931 nand P3_U6806 P3_U6805 P3_U6807 ; P3_U2752
g932 nand P3_U6803 P3_U6802 P3_U6804 ; P3_U2753
g933 nand P3_U6800 P3_U6799 P3_U6801 ; P3_U2754
g934 nand P3_U6797 P3_U6796 P3_U6798 ; P3_U2755
g935 nand P3_U6794 P3_U6793 P3_U6795 ; P3_U2756
g936 nand P3_U6791 P3_U6790 P3_U6792 ; P3_U2757
g937 nand P3_U6788 P3_U6787 P3_U6789 ; P3_U2758
g938 nand P3_U6785 P3_U6784 P3_U6786 ; P3_U2759
g939 nand P3_U6782 P3_U6781 P3_U6783 ; P3_U2760
g940 nand P3_U6779 P3_U6778 P3_U6780 ; P3_U2761
g941 nand P3_U6776 P3_U6775 P3_U6777 ; P3_U2762
g942 nand P3_U6773 P3_U6772 P3_U6774 ; P3_U2763
g943 nand P3_U6770 P3_U6769 P3_U6771 ; P3_U2764
g944 nand P3_U6767 P3_U6766 P3_U6768 ; P3_U2765
g945 nand P3_U6764 P3_U6763 P3_U6765 ; P3_U2766
g946 nand P3_U6761 P3_U6760 P3_U6762 ; P3_U2767
g947 nand P3_U6755 P3_U6754 P3_U6756 ; P3_U2768
g948 nand P3_U6752 P3_U6751 P3_U6753 ; P3_U2769
g949 nand P3_U6749 P3_U6748 P3_U6750 ; P3_U2770
g950 nand P3_U6746 P3_U6745 P3_U6747 ; P3_U2771
g951 nand P3_U6743 P3_U6742 P3_U6744 ; P3_U2772
g952 nand P3_U6740 P3_U6739 P3_U6741 ; P3_U2773
g953 nand P3_U6737 P3_U6736 P3_U6738 ; P3_U2774
g954 nand P3_U6734 P3_U6733 P3_U6735 ; P3_U2775
g955 nand P3_U6731 P3_U6730 P3_U6732 ; P3_U2776
g956 nand P3_U6728 P3_U6727 P3_U6729 ; P3_U2777
g957 nand P3_U6725 P3_U6724 P3_U6726 ; P3_U2778
g958 nand P3_U6722 P3_U6721 P3_U6723 ; P3_U2779
g959 nand P3_U6719 P3_U6718 P3_U6720 ; P3_U2780
g960 nand P3_U6716 P3_U6715 P3_U6717 ; P3_U2781
g961 nand P3_U6713 P3_U6712 P3_U6714 ; P3_U2782
g962 nand P3_U6710 P3_U6709 P3_U6711 ; P3_U2783
g963 nand P3_U6707 P3_U6706 P3_U6708 ; P3_U2784
g964 nand P3_U6704 P3_U6703 P3_U6705 ; P3_U2785
g965 nand P3_U6701 P3_U6700 P3_U6702 ; P3_U2786
g966 nand P3_U6698 P3_U6697 P3_U6699 ; P3_U2787
g967 nand P3_U6695 P3_U6694 P3_U6696 ; P3_U2788
g968 nand P3_U6692 P3_U6691 P3_U6693 ; P3_U2789
g969 nand P3_U6689 P3_U6688 P3_U6690 ; P3_U2790
g970 nand P3_U6686 P3_U6685 P3_U6687 ; P3_U2791
g971 nand P3_U6683 P3_U6682 P3_U6684 ; P3_U2792
g972 nand P3_U6680 P3_U6679 P3_U6681 ; P3_U2793
g973 nand P3_U6677 P3_U6676 P3_U6678 ; P3_U2794
g974 nand P3_U6674 P3_U6673 P3_U6675 ; P3_U2795
g975 nand P3_U6671 P3_U6670 P3_U6672 ; P3_U2796
g976 nand P3_U6668 P3_U6667 P3_U6669 ; P3_U2797
g977 nand P3_U6665 P3_U6664 P3_U6666 ; P3_U2798
g978 nand P3_U6656 P3_U6654 P3_U6655 P3_U6653 P3_U3985 ; P3_U2799
g979 nand P3_U6648 P3_U6647 P3_U6646 P3_U6645 P3_U3984 ; P3_U2800
g980 nand P3_U6640 P3_U6639 P3_U6638 P3_U6637 P3_U3983 ; P3_U2801
g981 nand P3_U6632 P3_U6631 P3_U6630 P3_U6629 P3_U3982 ; P3_U2802
g982 nand P3_U6622 P3_U6624 P3_U6621 P3_U6623 P3_U3981 ; P3_U2803
g983 nand P3_U6614 P3_U6616 P3_U6613 P3_U6615 P3_U3980 ; P3_U2804
g984 nand P3_U6606 P3_U6608 P3_U6605 P3_U6607 P3_U3979 ; P3_U2805
g985 nand P3_U6598 P3_U6600 P3_U6597 P3_U6599 P3_U3978 ; P3_U2806
g986 nand P3_U6590 P3_U6589 P3_U6592 P3_U6591 P3_U3977 ; P3_U2807
g987 nand P3_U6582 P3_U6581 P3_U6584 P3_U6583 P3_U3976 ; P3_U2808
g988 nand P3_U6574 P3_U6573 P3_U6575 P3_U3975 P3_U6576 ; P3_U2809
g989 nand P3_U6566 P3_U6565 P3_U6567 P3_U3974 P3_U6568 ; P3_U2810
g990 nand P3_U6558 P3_U6557 P3_U6559 P3_U6560 P3_U3973 ; P3_U2811
g991 nand P3_U6550 P3_U6549 P3_U6551 P3_U6552 P3_U3972 ; P3_U2812
g992 nand P3_U6542 P3_U6541 P3_U6543 P3_U6544 P3_U3971 ; P3_U2813
g993 nand P3_U6534 P3_U6533 P3_U6535 P3_U6536 P3_U3970 ; P3_U2814
g994 nand P3_U6526 P3_U6525 P3_U6528 P3_U6527 P3_U3969 ; P3_U2815
g995 nand P3_U6518 P3_U6517 P3_U6520 P3_U6519 P3_U3968 ; P3_U2816
g996 nand P3_U6510 P3_U6509 P3_U6512 P3_U6511 P3_U3967 ; P3_U2817
g997 nand P3_U6502 P3_U6501 P3_U6504 P3_U6503 P3_U3966 ; P3_U2818
g998 nand P3_U6494 P3_U6493 P3_U6495 P3_U6496 P3_U3965 ; P3_U2819
g999 nand P3_U6486 P3_U6485 P3_U6487 P3_U6488 P3_U3964 ; P3_U2820
g1000 nand P3_U6478 P3_U6477 P3_U6480 P3_U6479 P3_U3963 ; P3_U2821
g1001 nand P3_U6470 P3_U6469 P3_U6472 P3_U6471 P3_U3962 ; P3_U2822
g1002 nand P3_U6462 P3_U6461 P3_U6464 P3_U6463 P3_U3961 ; P3_U2823
g1003 nand P3_U6454 P3_U6453 P3_U6456 P3_U6455 P3_U3960 ; P3_U2824
g1004 nand P3_U6446 P3_U6445 P3_U6448 P3_U6447 P3_U3959 ; P3_U2825
g1005 nand P3_U6438 P3_U6437 P3_U6439 P3_U6440 P3_U3958 ; P3_U2826
g1006 nand P3_U6432 P3_U6431 P3_U6430 P3_U6429 P3_U3957 ; P3_U2827
g1007 nand P3_U6424 P3_U6423 P3_U6422 P3_U6421 P3_U3956 ; P3_U2828
g1008 nand P3_U6416 P3_U6415 P3_U6414 P3_U6413 P3_U3955 ; P3_U2829
g1009 nand P3_U6408 P3_U6407 P3_U6406 P3_U6405 P3_U3954 ; P3_U2830
g1010 and P3_U6396 P3_U7906 ; P3_U2831
g1011 nand P3_U6375 P3_U6373 P3_U6374 ; P3_U2832
g1012 nand P3_U6351 P3_U6349 P3_U6350 ; P3_U2833
g1013 nand P3_U6327 P3_U6325 P3_U6326 ; P3_U2834
g1014 nand P3_U6303 P3_U6301 P3_U6302 ; P3_U2835
g1015 nand P3_U6279 P3_U6277 P3_U6278 ; P3_U2836
g1016 nand P3_U3893 P3_U6254 ; P3_U2837
g1017 nand P3_U3883 P3_U6230 ; P3_U2838
g1018 nand P3_U3873 P3_U6206 ; P3_U2839
g1019 nand P3_U3863 P3_U6182 ; P3_U2840
g1020 nand P3_U3853 P3_U6158 ; P3_U2841
g1021 nand P3_U3845 P3_U6134 ; P3_U2842
g1022 nand P3_U6111 P3_U6109 P3_U6110 ; P3_U2843
g1023 nand P3_U6087 P3_U6085 P3_U6086 ; P3_U2844
g1024 nand P3_U6063 P3_U6061 P3_U6062 ; P3_U2845
g1025 nand P3_U6039 P3_U6037 P3_U6038 ; P3_U2846
g1026 nand P3_U3811 P3_U6014 ; P3_U2847
g1027 nand P3_U3803 P3_U5990 ; P3_U2848
g1028 nand P3_U5967 P3_U5965 P3_U5966 ; P3_U2849
g1029 nand P3_U5943 P3_U5941 P3_U5942 ; P3_U2850
g1030 nand P3_U5919 P3_U5917 P3_U5918 ; P3_U2851
g1031 nand P3_U5895 P3_U5893 P3_U5894 ; P3_U2852
g1032 nand P3_U5871 P3_U5869 P3_U5870 ; P3_U2853
g1033 nand P3_U5847 P3_U5845 P3_U5846 ; P3_U2854
g1034 nand P3_U5823 P3_U5821 P3_U5822 ; P3_U2855
g1035 nand P3_U5799 P3_U5797 P3_U5798 ; P3_U2856
g1036 nand P3_U5775 P3_U5773 P3_U5774 ; P3_U2857
g1037 nand P3_U5751 P3_U5749 P3_U5750 ; P3_U2858
g1038 nand P3_U5727 P3_U5725 P3_U5726 ; P3_U2859
g1039 nand P3_U5703 P3_U5701 P3_U5702 ; P3_U2860
g1040 nand P3_U5679 P3_U5677 P3_U5678 ; P3_U2861
g1041 nand P3_U5654 P3_U5653 P3_U5655 ; P3_U2862
g1042 nand P3_U5616 P3_U5615 ; P3_U2863
g1043 nand P3_U5610 P3_U5609 ; P3_U2864
g1044 nand P3_U5599 P3_U5598 ; P3_U2865
g1045 nand P3_U5591 P3_U5590 ; P3_U2866
g1046 and P3_U5579 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_U2867
g1047 nand P3_U3651 P3_U5482 ; P3_U2868
g1048 nand P3_U3649 P3_U5477 ; P3_U2869
g1049 nand P3_U3647 P3_U5472 ; P3_U2870
g1050 nand P3_U3645 P3_U5467 ; P3_U2871
g1051 nand P3_U3643 P3_U5462 ; P3_U2872
g1052 nand P3_U3641 P3_U5457 ; P3_U2873
g1053 nand P3_U3639 P3_U5452 ; P3_U2874
g1054 nand P3_U3637 P3_U5447 ; P3_U2875
g1055 nand P3_U3633 P3_U5432 ; P3_U2876
g1056 nand P3_U3631 P3_U5427 ; P3_U2877
g1057 nand P3_U3629 P3_U5422 ; P3_U2878
g1058 nand P3_U3627 P3_U5417 ; P3_U2879
g1059 nand P3_U3625 P3_U5412 ; P3_U2880
g1060 nand P3_U3623 P3_U5407 ; P3_U2881
g1061 nand P3_U3621 P3_U5402 ; P3_U2882
g1062 nand P3_U3619 P3_U5397 ; P3_U2883
g1063 nand P3_U3615 P3_U5381 ; P3_U2884
g1064 nand P3_U3613 P3_U5376 ; P3_U2885
g1065 nand P3_U3611 P3_U5371 ; P3_U2886
g1066 nand P3_U3609 P3_U5366 ; P3_U2887
g1067 nand P3_U3607 P3_U5361 ; P3_U2888
g1068 nand P3_U3605 P3_U5356 ; P3_U2889
g1069 nand P3_U3603 P3_U5351 ; P3_U2890
g1070 nand P3_U3601 P3_U5346 ; P3_U2891
g1071 nand P3_U3598 P3_U5330 ; P3_U2892
g1072 nand P3_U3596 P3_U5325 ; P3_U2893
g1073 nand P3_U3594 P3_U5320 ; P3_U2894
g1074 nand P3_U3592 P3_U5315 ; P3_U2895
g1075 nand P3_U3590 P3_U5310 ; P3_U2896
g1076 nand P3_U3588 P3_U5305 ; P3_U2897
g1077 nand P3_U3586 P3_U5300 ; P3_U2898
g1078 nand P3_U3584 P3_U5295 ; P3_U2899
g1079 nand P3_U3580 P3_U5279 ; P3_U2900
g1080 nand P3_U3578 P3_U5274 ; P3_U2901
g1081 nand P3_U3576 P3_U5269 ; P3_U2902
g1082 nand P3_U3574 P3_U5264 ; P3_U2903
g1083 nand P3_U3572 P3_U5259 ; P3_U2904
g1084 nand P3_U3570 P3_U5254 ; P3_U2905
g1085 nand P3_U3568 P3_U5249 ; P3_U2906
g1086 nand P3_U3566 P3_U5244 ; P3_U2907
g1087 nand P3_U5229 P3_U3562 P3_U5228 ; P3_U2908
g1088 nand P3_U5224 P3_U3560 P3_U5223 ; P3_U2909
g1089 nand P3_U5219 P3_U3558 P3_U5218 ; P3_U2910
g1090 nand P3_U5214 P3_U3556 P3_U5213 ; P3_U2911
g1091 nand P3_U5209 P3_U3554 P3_U5208 ; P3_U2912
g1092 nand P3_U5204 P3_U3552 P3_U5203 ; P3_U2913
g1093 nand P3_U5199 P3_U3550 P3_U5198 ; P3_U2914
g1094 nand P3_U5194 P3_U3548 P3_U5193 ; P3_U2915
g1095 nand P3_U5177 P3_U3544 P3_U5176 ; P3_U2916
g1096 nand P3_U5172 P3_U3542 P3_U5171 ; P3_U2917
g1097 nand P3_U5167 P3_U3540 P3_U5166 ; P3_U2918
g1098 nand P3_U5162 P3_U3538 P3_U5161 ; P3_U2919
g1099 nand P3_U5157 P3_U3536 P3_U5156 ; P3_U2920
g1100 nand P3_U5152 P3_U3534 P3_U5151 ; P3_U2921
g1101 nand P3_U5147 P3_U3532 P3_U5146 ; P3_U2922
g1102 nand P3_U5142 P3_U3530 P3_U5141 ; P3_U2923
g1103 nand P3_U5125 P3_U3526 P3_U5124 ; P3_U2924
g1104 nand P3_U5120 P3_U3524 P3_U5119 ; P3_U2925
g1105 nand P3_U5115 P3_U3522 P3_U5114 ; P3_U2926
g1106 nand P3_U5110 P3_U3520 P3_U5109 ; P3_U2927
g1107 nand P3_U5105 P3_U3518 P3_U5104 ; P3_U2928
g1108 nand P3_U5100 P3_U3516 P3_U5099 ; P3_U2929
g1109 nand P3_U5095 P3_U3514 P3_U5094 ; P3_U2930
g1110 nand P3_U5090 P3_U3512 P3_U5089 ; P3_U2931
g1111 nand P3_U5076 P3_U3509 P3_U5075 ; P3_U2932
g1112 nand P3_U5071 P3_U3507 P3_U5070 ; P3_U2933
g1113 nand P3_U5066 P3_U3505 P3_U5065 ; P3_U2934
g1114 nand P3_U5061 P3_U3503 P3_U5060 ; P3_U2935
g1115 nand P3_U5056 P3_U3501 P3_U5055 ; P3_U2936
g1116 nand P3_U5051 P3_U3499 P3_U5050 ; P3_U2937
g1117 nand P3_U5046 P3_U3497 P3_U5045 ; P3_U2938
g1118 nand P3_U5041 P3_U3495 P3_U5040 ; P3_U2939
g1119 nand P3_U5025 P3_U3492 P3_U5024 ; P3_U2940
g1120 nand P3_U5020 P3_U3490 P3_U5019 ; P3_U2941
g1121 nand P3_U5015 P3_U3488 P3_U5014 ; P3_U2942
g1122 nand P3_U5010 P3_U3486 P3_U5009 ; P3_U2943
g1123 nand P3_U5005 P3_U3484 P3_U5004 ; P3_U2944
g1124 nand P3_U5000 P3_U3482 P3_U4999 ; P3_U2945
g1125 nand P3_U4995 P3_U3480 P3_U4994 ; P3_U2946
g1126 nand P3_U4990 P3_U3478 P3_U4989 ; P3_U2947
g1127 nand P3_U4973 P3_U3474 P3_U4972 ; P3_U2948
g1128 nand P3_U4968 P3_U3472 P3_U4967 ; P3_U2949
g1129 nand P3_U4963 P3_U3470 P3_U4962 ; P3_U2950
g1130 nand P3_U4958 P3_U3468 P3_U4957 ; P3_U2951
g1131 nand P3_U4953 P3_U3466 P3_U4952 ; P3_U2952
g1132 nand P3_U4948 P3_U3464 P3_U4947 ; P3_U2953
g1133 nand P3_U4943 P3_U3462 P3_U4942 ; P3_U2954
g1134 nand P3_U4938 P3_U3460 P3_U4937 ; P3_U2955
g1135 nand P3_U4921 P3_U3456 P3_U4920 ; P3_U2956
g1136 nand P3_U4916 P3_U3454 P3_U4915 ; P3_U2957
g1137 nand P3_U4911 P3_U3452 P3_U4910 ; P3_U2958
g1138 nand P3_U4906 P3_U3450 P3_U4905 ; P3_U2959
g1139 nand P3_U4901 P3_U3448 P3_U4900 ; P3_U2960
g1140 nand P3_U4896 P3_U3446 P3_U4895 ; P3_U2961
g1141 nand P3_U4891 P3_U3444 P3_U4890 ; P3_U2962
g1142 nand P3_U4886 P3_U3442 P3_U4885 ; P3_U2963
g1143 nand P3_U4869 P3_U3439 P3_U4868 ; P3_U2964
g1144 nand P3_U4864 P3_U3437 P3_U4863 ; P3_U2965
g1145 nand P3_U4859 P3_U3435 P3_U4858 ; P3_U2966
g1146 nand P3_U4854 P3_U3433 P3_U4853 ; P3_U2967
g1147 nand P3_U4849 P3_U3431 P3_U4848 ; P3_U2968
g1148 nand P3_U4844 P3_U3429 P3_U4843 ; P3_U2969
g1149 nand P3_U4839 P3_U3427 P3_U4838 ; P3_U2970
g1150 nand P3_U4834 P3_U3425 P3_U4833 ; P3_U2971
g1151 nand P3_U4818 P3_U3421 P3_U4817 ; P3_U2972
g1152 nand P3_U4813 P3_U3419 P3_U4812 ; P3_U2973
g1153 nand P3_U4808 P3_U3417 P3_U4807 ; P3_U2974
g1154 nand P3_U4803 P3_U3415 P3_U4802 ; P3_U2975
g1155 nand P3_U4798 P3_U3413 P3_U4797 ; P3_U2976
g1156 nand P3_U4793 P3_U3411 P3_U4792 ; P3_U2977
g1157 nand P3_U4788 P3_U3409 P3_U4787 ; P3_U2978
g1158 nand P3_U4783 P3_U3407 P3_U4782 ; P3_U2979
g1159 nand P3_U4766 P3_U3403 P3_U4765 ; P3_U2980
g1160 nand P3_U4761 P3_U3401 P3_U4760 ; P3_U2981
g1161 nand P3_U4756 P3_U3399 P3_U4755 ; P3_U2982
g1162 nand P3_U4751 P3_U3397 P3_U4750 ; P3_U2983
g1163 nand P3_U4746 P3_U3395 P3_U4745 ; P3_U2984
g1164 nand P3_U4741 P3_U3393 P3_U4740 ; P3_U2985
g1165 nand P3_U4736 P3_U3391 P3_U4735 ; P3_U2986
g1166 nand P3_U4731 P3_U3389 P3_U4730 ; P3_U2987
g1167 nand P3_U4714 P3_U3385 P3_U4713 ; P3_U2988
g1168 nand P3_U4709 P3_U3383 P3_U4708 ; P3_U2989
g1169 nand P3_U4704 P3_U3381 P3_U4703 ; P3_U2990
g1170 nand P3_U4699 P3_U3379 P3_U4698 ; P3_U2991
g1171 nand P3_U4694 P3_U3377 P3_U4693 ; P3_U2992
g1172 nand P3_U4689 P3_U3375 P3_U4688 ; P3_U2993
g1173 nand P3_U4684 P3_U3373 P3_U4683 ; P3_U2994
g1174 nand P3_U4679 P3_U3371 P3_U4678 ; P3_U2995
g1175 nand P3_U7959 P3_U7958 P3_U3367 ; P3_U2996
g1176 nand P3_U4636 P3_U4635 P3_U4634 P3_U4329 ; P3_U2997
g1177 nand P3_U3363 P3_U4632 ; P3_U2998
g1178 and P3_U7937 P3_DATAWIDTH_REG_31__SCAN_IN ; P3_U2999
g1179 and P3_U7937 P3_DATAWIDTH_REG_30__SCAN_IN ; P3_U3000
g1180 and P3_U7937 P3_DATAWIDTH_REG_29__SCAN_IN ; P3_U3001
g1181 and P3_U7937 P3_DATAWIDTH_REG_28__SCAN_IN ; P3_U3002
g1182 and P3_U7937 P3_DATAWIDTH_REG_27__SCAN_IN ; P3_U3003
g1183 and P3_U7937 P3_DATAWIDTH_REG_26__SCAN_IN ; P3_U3004
g1184 and P3_U7937 P3_DATAWIDTH_REG_25__SCAN_IN ; P3_U3005
g1185 and P3_U7937 P3_DATAWIDTH_REG_24__SCAN_IN ; P3_U3006
g1186 and P3_U7937 P3_DATAWIDTH_REG_23__SCAN_IN ; P3_U3007
g1187 and P3_U7937 P3_DATAWIDTH_REG_22__SCAN_IN ; P3_U3008
g1188 and P3_U7937 P3_DATAWIDTH_REG_21__SCAN_IN ; P3_U3009
g1189 and P3_U7937 P3_DATAWIDTH_REG_20__SCAN_IN ; P3_U3010
g1190 and P3_U7937 P3_DATAWIDTH_REG_19__SCAN_IN ; P3_U3011
g1191 and P3_U7937 P3_DATAWIDTH_REG_18__SCAN_IN ; P3_U3012
g1192 and P3_U7937 P3_DATAWIDTH_REG_17__SCAN_IN ; P3_U3013
g1193 and P3_U7937 P3_DATAWIDTH_REG_16__SCAN_IN ; P3_U3014
g1194 and P3_U7937 P3_DATAWIDTH_REG_15__SCAN_IN ; P3_U3015
g1195 and P3_U7937 P3_DATAWIDTH_REG_14__SCAN_IN ; P3_U3016
g1196 and P3_U7937 P3_DATAWIDTH_REG_13__SCAN_IN ; P3_U3017
g1197 and P3_U7937 P3_DATAWIDTH_REG_12__SCAN_IN ; P3_U3018
g1198 and P3_U7937 P3_DATAWIDTH_REG_11__SCAN_IN ; P3_U3019
g1199 and P3_U7937 P3_DATAWIDTH_REG_10__SCAN_IN ; P3_U3020
g1200 and P3_U7937 P3_DATAWIDTH_REG_9__SCAN_IN ; P3_U3021
g1201 and P3_U7937 P3_DATAWIDTH_REG_8__SCAN_IN ; P3_U3022
g1202 and P3_U7937 P3_DATAWIDTH_REG_7__SCAN_IN ; P3_U3023
g1203 and P3_U7937 P3_DATAWIDTH_REG_6__SCAN_IN ; P3_U3024
g1204 and P3_U7937 P3_DATAWIDTH_REG_5__SCAN_IN ; P3_U3025
g1205 and P3_U7937 P3_DATAWIDTH_REG_4__SCAN_IN ; P3_U3026
g1206 and P3_U7937 P3_DATAWIDTH_REG_3__SCAN_IN ; P3_U3027
g1207 and P3_U7937 P3_DATAWIDTH_REG_2__SCAN_IN ; P3_U3028
g1208 nand P3_U7934 P3_U7933 P3_U4463 ; P3_U3029
g1209 nand P3_U7932 P3_U7931 P3_U3311 ; P3_U3030
g1210 nand P3_U3310 P3_U4457 ; P3_U3031
g1211 nand P3_U4443 P3_U4442 P3_U4444 ; P3_U3032
g1212 nand P3_U4440 P3_U4439 P3_U4441 ; P3_U3033
g1213 nand P3_U4437 P3_U4436 P3_U4438 ; P3_U3034
g1214 nand P3_U4434 P3_U4433 P3_U4435 ; P3_U3035
g1215 nand P3_U4431 P3_U4430 P3_U4432 ; P3_U3036
g1216 nand P3_U4428 P3_U4427 P3_U4429 ; P3_U3037
g1217 nand P3_U4425 P3_U4424 P3_U4426 ; P3_U3038
g1218 nand P3_U4422 P3_U4421 P3_U4423 ; P3_U3039
g1219 nand P3_U4419 P3_U4418 P3_U4420 ; P3_U3040
g1220 nand P3_U4416 P3_U4415 P3_U4417 ; P3_U3041
g1221 nand P3_U4413 P3_U4412 P3_U4414 ; P3_U3042
g1222 nand P3_U4410 P3_U4409 P3_U4411 ; P3_U3043
g1223 nand P3_U4407 P3_U4406 P3_U4408 ; P3_U3044
g1224 nand P3_U4404 P3_U4403 P3_U4405 ; P3_U3045
g1225 nand P3_U4401 P3_U4400 P3_U4402 ; P3_U3046
g1226 nand P3_U4398 P3_U4397 P3_U4399 ; P3_U3047
g1227 nand P3_U4395 P3_U4394 P3_U4396 ; P3_U3048
g1228 nand P3_U4392 P3_U4391 P3_U4393 ; P3_U3049
g1229 nand P3_U4389 P3_U4388 P3_U4390 ; P3_U3050
g1230 nand P3_U4386 P3_U4385 P3_U4387 ; P3_U3051
g1231 nand P3_U4383 P3_U4382 P3_U4384 ; P3_U3052
g1232 nand P3_U4380 P3_U4379 P3_U4381 ; P3_U3053
g1233 nand P3_U4377 P3_U4376 P3_U4378 ; P3_U3054
g1234 nand P3_U4374 P3_U4373 P3_U4375 ; P3_U3055
g1235 nand P3_U4371 P3_U4370 P3_U4372 ; P3_U3056
g1236 nand P3_U4368 P3_U4367 P3_U4369 ; P3_U3057
g1237 nand P3_U4365 P3_U4364 P3_U4366 ; P3_U3058
g1238 nand P3_U4362 P3_U4361 P3_U4363 ; P3_U3059
g1239 nand P3_U4359 P3_U4358 P3_U4360 ; P3_U3060
g1240 nand P3_U4356 P3_U4355 P3_U4357 ; P3_U3061
g1241 nand P3_U4247 P3_U4246 P3_U4245 P3_U4244 ; P3_U3062
g1242 nand P3_U4243 P3_U4242 P3_U4241 P3_U4240 ; P3_U3063
g1243 nand P3_U4239 P3_U4238 P3_U4237 P3_U4236 ; P3_U3064
g1244 nand P3_U4235 P3_U4234 P3_U4233 P3_U4232 ; P3_U3065
g1245 nand P3_U4231 P3_U4230 P3_U4229 P3_U4228 ; P3_U3066
g1246 nand P3_U4227 P3_U4226 P3_U4225 P3_U4224 ; P3_U3067
g1247 nand P3_U4223 P3_U4222 P3_U4221 P3_U4220 ; P3_U3068
g1248 nand P3_U4219 P3_U4218 P3_U4217 P3_U4216 ; P3_U3069
g1249 nand P3_U2457 P3_U4642 ; P3_U3070
g1250 nand P3_U2459 P3_U4642 ; P3_U3071
g1251 nand P3_U2458 P3_U4642 ; P3_U3072
g1252 nand P3_U2460 P3_U4642 ; P3_U3073
g1253 nand P3_U3346 P3_U3345 P3_U3347 P3_U3344 P3_U3343 ; P3_U3074
g1254 not P3_REQUESTPENDING_REG_SCAN_IN ; P3_U3075
g1255 not P3_STATE_REG_1__SCAN_IN ; P3_U3076
g1256 nand P3_U3085 P3_STATE_REG_1__SCAN_IN ; P3_U3077
g1257 nand P3_U4308 P3_U3079 ; P3_U3078
g1258 not P3_STATE_REG_2__SCAN_IN ; P3_U3079
g1259 nand P3_U4308 P3_STATE_REG_2__SCAN_IN ; P3_U3080
g1260 not P3_REIP_REG_1__SCAN_IN ; P3_U3081
g1261 nand P3_U3079 P3_STATE_REG_1__SCAN_IN ; P3_U3082
g1262 or P3_STATE_REG_2__SCAN_IN P3_STATE_REG_1__SCAN_IN ; P3_U3083
g1263 not HOLD ; P3_U3084
g1264 not P3_STATE_REG_0__SCAN_IN ; P3_U3085
g1265 nand P3_U3087 P3_STATE_REG_0__SCAN_IN ; P3_U3086
g1266 nand P3_U3084 P3_REQUESTPENDING_REG_SCAN_IN ; P3_U3087
g1267 or HOLD P3_REQUESTPENDING_REG_SCAN_IN ; P3_U3088
g1268 not P3_STATE2_REG_1__SCAN_IN ; P3_U3089
g1269 not P3_STATE2_REG_2__SCAN_IN ; P3_U3090
g1270 or P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U3091
g1271 nand P3_U4467 P3_U3097 ; P3_U3092
g1272 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U3093
g1273 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U3094
g1274 nand P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U3095
g1275 nand P3_U4332 P3_U3097 ; P3_U3096
g1276 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U3097
g1277 nand P3_U3100 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U3098
g1278 nand P3_U4470 P3_U4332 ; P3_U3099
g1279 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U3100
g1280 nand P3_U3341 P3_U3340 P3_U3342 P3_U3339 P3_U3338 ; P3_U3101
g1281 nand P3_U3326 P3_U3325 P3_U3327 P3_U3324 P3_U3323 ; P3_U3102
g1282 nand P3_U3074 P3_U3110 ; P3_U3103
g1283 nand P3_U3321 P3_U3320 P3_U3322 P3_U3319 P3_U3318 ; P3_U3104
g1284 nand P3_U4466 P3_U3085 ; P3_U3105
g1285 nand P3_U4293 P3_U2630 ; P3_U3106
g1286 nand P3_U3331 P3_U3330 P3_U3332 P3_U3329 P3_U3328 ; P3_U3107
g1287 nand P3_U3316 P3_U3315 P3_U3317 P3_U3314 P3_U3313 ; P3_U3108
g1288 nand P3_U2353 P3_U4488 ; P3_U3109
g1289 nand P3_U3351 P3_U3350 P3_U3352 P3_U3349 P3_U3348 ; P3_U3110
g1290 nand P3_U3104 P3_U3108 ; P3_U3111
g1291 nand P3_U4505 P3_U3108 ; P3_U3112
g1292 nand P3_U4607 P3_U3110 ; P3_U3113
g1293 nand P3_U4488 P3_U4505 ; P3_U3114
g1294 nand P3_U2451 P3_U4297 ; P3_U3115
g1295 nand P3_U2452 P3_U4297 ; P3_U3116
g1296 nand P3_U2452 P3_U4296 ; P3_U3117
g1297 nand P3_U4488 P3_U3104 ; P3_U3118
g1298 nand P3_U3356 P3_U2353 ; P3_U3119
g1299 nand P3_U7949 P3_U7948 P3_U3262 P3_U4313 P3_LT_563_U6 ; P3_U3120
g1300 not P3_STATE2_REG_0__SCAN_IN ; P3_U3121
g1301 nand P3_U4629 P3_STATE2_REG_0__SCAN_IN ; P3_U3122
g1302 or P3_STATE2_REG_3__SCAN_IN P3_STATE2_REG_1__SCAN_IN ; P3_U3123
g1303 nand P3_U3089 P3_STATE2_REG_2__SCAN_IN ; P3_U3124
g1304 or P3_STATE2_REG_2__SCAN_IN P3_STATE2_REG_1__SCAN_IN ; P3_U3125
g1305 nand P3_LTE_597_U6 P3_STATE2_REG_3__SCAN_IN ; P3_U3126
g1306 nand P3_U4666 P3_U3121 ; P3_U3127
g1307 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U3128
g1308 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3129
g1309 nand P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U3130
g1310 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U3131
g1311 nand P3_U4648 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U3132
g1312 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U3133
g1313 nand P3_U4649 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U3134
g1314 or P3_STATE2_REG_3__SCAN_IN P3_STATE2_REG_2__SCAN_IN ; P3_U3135
g1315 nand P3_U4295 P3_STATEBS16_REG_SCAN_IN ; P3_U3136
g1316 nand P3_U3153 P3_U4641 ; P3_U3137
g1317 nand P3_U3137 P3_U3128 ; P3_U3138
g1318 nand P3_U3180 P3_U4651 ; P3_U3139
g1319 nand P3_U3141 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U3140
g1320 nand P3_U3150 P3_U3158 ; P3_U3141
g1321 nand P3_U4331 P3_U4655 ; P3_U3142
g1322 nand P3_U3156 P3_U3128 ; P3_U3143
g1323 nand P3_U4647 P3_U2486 ; P3_U3144
g1324 nand P3_U3144 P3_U4667 ; P3_U3145
g1325 nand P3_U3134 P3_U4663 ; P3_U3146
g1326 nand P3_U3386 P3_U2492 ; P3_U3147
g1327 nand P3_U3141 P3_U3128 ; P3_U3148
g1328 nand P3_U2490 P3_U2486 ; P3_U3149
g1329 nand P3_U3137 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U3150
g1330 nand P3_U3149 P3_U4719 ; P3_U3151
g1331 nand P3_U3147 P3_U4717 ; P3_U3152
g1332 nand P3_U3129 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U3153
g1333 nand P3_U3404 P3_U4640 ; P3_U3154
g1334 nand P3_U4643 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U3155
g1335 nand P3_U3148 P3_U3155 ; P3_U3156
g1336 nand P3_U2493 P3_U2486 ; P3_U3157
g1337 nand P3_U4642 P3_U3128 ; P3_U3158
g1338 nand P3_U3157 P3_U4771 ; P3_U3159
g1339 nand P3_U3154 P3_U4769 ; P3_U3160
g1340 nand P3_U3422 P3_U2492 ; P3_U3161
g1341 nand P3_U2495 P3_U2486 ; P3_U3162
g1342 nand P3_U3162 P3_U4822 ; P3_U3163
g1343 nand P3_U3131 P3_U4648 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U3164
g1344 nand P3_U7965 P3_U3142 ; P3_U3165
g1345 nand P3_U2498 P3_U4647 ; P3_U3166
g1346 nand P3_U3166 P3_U4874 ; P3_U3167
g1347 nand P3_U3164 P3_U4872 ; P3_U3168
g1348 nand P3_U3457 P3_U2501 ; P3_U3169
g1349 nand P3_U2498 P3_U2490 ; P3_U3170
g1350 nand P3_U3170 P3_U4926 ; P3_U3171
g1351 nand P3_U3169 P3_U4924 ; P3_U3172
g1352 nand P3_U3475 P3_U4640 ; P3_U3173
g1353 nand P3_U2498 P3_U2493 ; P3_U3174
g1354 nand P3_U3174 P3_U4978 ; P3_U3175
g1355 nand P3_U3173 P3_U4976 ; P3_U3176
g1356 nand P3_U3129 P3_U2501 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U3177
g1357 nand P3_U2498 P3_U2495 ; P3_U3178
g1358 nand P3_U3178 P3_U5029 ; P3_U3179
g1359 nand P3_U4649 P3_U3133 ; P3_U3180
g1360 nand P3_U2485 P3_U4657 ; P3_U3181
g1361 nand P3_U3368 P3_U3181 ; P3_U3182
g1362 nand P3_U2504 P3_U4647 ; P3_U3183
g1363 nand P3_U3183 P3_U3181 ; P3_U3184
g1364 nand P3_U3180 P3_U4331 ; P3_U3185
g1365 nand P3_U3527 P3_U2492 ; P3_U3186
g1366 nand P3_U2504 P3_U2490 ; P3_U3187
g1367 nand P3_U3187 P3_U5130 ; P3_U3188
g1368 nand P3_U3186 P3_U5128 ; P3_U3189
g1369 nand P3_U3545 P3_U4640 ; P3_U3190
g1370 nand P3_U2504 P3_U2493 ; P3_U3191
g1371 nand P3_U3191 P3_U5182 ; P3_U3192
g1372 nand P3_U3190 P3_U5180 ; P3_U3193
g1373 nand P3_U3563 P3_U2492 ; P3_U3194
g1374 nand P3_U2504 P3_U2495 ; P3_U3195
g1375 nand P3_U3581 P3_U4648 ; P3_U3196
g1376 nand P3_U2508 P3_U4647 ; P3_U3197
g1377 nand P3_U3196 P3_U5282 ; P3_U3198
g1378 nand P3_U3133 P3_U2501 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3199
g1379 nand P3_U2508 P3_U2490 ; P3_U3200
g1380 nand P3_U3199 P3_U5333 ; P3_U3201
g1381 nand P3_U3616 P3_U4640 ; P3_U3202
g1382 nand P3_U2508 P3_U2493 ; P3_U3203
g1383 nand P3_U3202 P3_U5384 ; P3_U3204
g1384 nand P3_U3634 P3_U2501 ; P3_U3205
g1385 nand P3_U2508 P3_U2495 ; P3_U3206
g1386 not P3_FLUSH_REG_SCAN_IN ; P3_U3207
g1387 nand P3_U4539 P3_U3102 ; P3_U3208
g1388 nand P3_U2514 P3_U3113 ; P3_U3209
g1389 not P3_GTE_412_U6 ; P3_U3210
g1390 not P3_GTE_485_U6 ; P3_U3211
g1391 not P3_GTE_390_U6 ; P3_U3212
g1392 not P3_GTE_450_U6 ; P3_U3213
g1393 not P3_GTE_504_U6 ; P3_U3214
g1394 not P3_GTE_401_U6 ; P3_U3215
g1395 nand P3_U4590 P3_U3074 ; P3_U3216
g1396 nand P3_U2450 P3_U4323 ; P3_U3217
g1397 nand P3_U3336 P3_U3335 P3_U3337 P3_U3334 P3_U3333 ; P3_U3218
g1398 nand P3_U3662 P3_U2461 ; P3_U3219
g1399 nand P3_U7976 P3_U7975 P3_U3667 ; P3_U3220
g1400 nand P3_U3222 P3_U3119 P3_U5524 ; P3_U3221
g1401 nand P3_U4314 P3_U3218 ; P3_U3222
g1402 nand P3_U5503 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U3223
g1403 nand P3_U5505 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U3224
g1404 nand P3_U3096 P3_U3227 ; P3_U3225
g1405 nand P3_U3674 P3_U2517 ; P3_U3226
g1406 nand P3_U3095 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U3227
g1407 nand P3_U3091 P3_U3095 ; P3_U3228
g1408 nand P3_U4323 P3_U3218 P3_U4350 ; P3_U3229
g1409 nand P3_U2518 P3_U3243 ; P3_U3230
g1410 nand P3_U3115 P3_U5559 ; P3_U3231
g1411 not P3_LT_589_U6 ; P3_U3232
g1412 nand P3_U4330 P3_U3127 P3_U5578 ; P3_U3233
g1413 nand P3_U3135 P3_U3123 ; P3_U3234
g1414 nand P3_U3101 P3_U3104 P3_U4294 ; P3_U3235
g1415 nand P3_U3101 P3_U2630 P3_U4505 ; P3_U3236
g1416 not P3_GTE_370_U6 ; P3_U3237
g1417 not P3_GTE_355_U6 ; P3_U3238
g1418 nand P3_U4295 P3_U3089 ; P3_U3239
g1419 not P3_REIP_REG_0__SCAN_IN ; P3_U3240
g1420 not P3_U2628 ; P3_U3241
g1421 nand P3_U3661 P3_U2450 ; P3_U3242
g1422 nand P3_U2461 P3_U4314 ; P3_U3243
g1423 nand P3_U4352 P3_U4522 ; P3_U3244
g1424 nand P3_U4352 P3_U3102 ; P3_U3245
g1425 nand P3_U3663 P3_U2449 P3_U3664 ; P3_U3246
g1426 nand P3_U3248 P3_STATE2_REG_2__SCAN_IN ; P3_U3247
g1427 nand P3_U4336 P3_U5630 ; P3_U3248
g1428 nand P3_U6403 P3_U6402 ; P3_U3249
g1429 nand P3_U2390 P3_U6663 ; P3_U3250
g1430 nand P3_U6758 P3_U6757 ; P3_U3251
g1431 nand P3_U2390 P3_U6853 ; P3_U3252
g1432 nand P3_U2390 P3_U6997 ; P3_U3253
g1433 nand P3_U5490 P3_U5489 ; P3_U3254
g1434 nand P3_U5487 P3_U5486 ; P3_U3255
g1435 not P3_EBX_REG_31__SCAN_IN ; P3_U3256
g1436 or U209 P3_STATEBS16_REG_SCAN_IN ; P3_U3257
g1437 not P3_ADD_318_U69 ; P3_U3258
g1438 nand P3_ADD_318_U69 P3_U2385 ; P3_U3259
g1439 nand P3_U4030 P3_U4334 ; P3_U3260
g1440 nand P3_U4148 P3_U4144 P3_U4141 P3_U4138 ; P3_U3261
g1441 nand P3_U2462 P3_U3108 P3_U4282 ; P3_U3262
g1442 not P3_CODEFETCH_REG_SCAN_IN ; P3_U3263
g1443 not P3_READREQUEST_REG_SCAN_IN ; P3_U3264
g1444 nand P3_U3099 P3_U3224 ; P3_U3265
g1445 nand P3_U3223 P3_U7515 ; P3_U3266
g1446 nand P3_U4289 P3_U3092 ; P3_U3267
g1447 nand P3_U3098 P3_U7774 ; P3_U3268
g1448 nand P3_U7961 P3_U7960 ; P3_U3269
g1449 nand P3_U7964 P3_U7963 ; P3_U3270
g1450 nand P3_U7967 P3_U7966 ; P3_U3271
g1451 nand P3_U8033 P3_U8032 ; P3_U3272
g1452 nand P3_U8036 P3_U8035 ; P3_U3273
g1453 nand P3_U7921 P3_U7920 ; P3_U3274
g1454 nand P3_U7923 P3_U7922 ; P3_U3275
g1455 nand P3_U7925 P3_U7924 ; P3_U3276
g1456 nand P3_U7927 P3_U7926 ; P3_U3277
g1457 nand P3_U7936 P3_U7935 ; P3_U3278
g1458 and P3_U3083 P3_U4286 ; P3_U3279
g1459 nand P3_U7939 P3_U7938 ; P3_U3280
g1460 nand P3_U7941 P3_U7940 ; P3_U3281
g1461 nand P3_U7955 P3_U7954 ; P3_U3282
g1462 and P3_U3652 P3_U2356 ; P3_U3283
g1463 nand P3_U7972 P3_U7971 ; P3_U3284
g1464 nand P3_U7980 P3_U7979 ; P3_U3285
g1465 nand P3_U7987 P3_U7986 ; P3_U3286
g1466 nand P3_U7984 P3_U7983 ; P3_U3287
g1467 nand P3_U7990 P3_U7989 ; P3_U3288
g1468 nand P3_U7992 P3_U7991 ; P3_U3289
g1469 nand P3_U7996 P3_U7995 ; P3_U3290
g1470 nor P3_DATAWIDTH_REG_1__SCAN_IN P3_REIP_REG_1__SCAN_IN ; P3_U3291
g1471 nand P3_U8011 P3_U8010 ; P3_U3292
g1472 nand P3_U8015 P3_U8014 ; P3_U3293
g1473 nand P3_U8017 P3_U8016 ; P3_U3294
g1474 nand P3_U8019 P3_U8018 ; P3_U3295
g1475 nand P3_U8023 P3_U8022 ; P3_U3296
g1476 nand P3_U8027 P3_U8026 ; P3_U3297
g1477 nand P3_U8029 P3_U8028 ; P3_U3298
g1478 nand P3_U8031 P3_U8030 ; P3_U3299
g1479 nand P3_U8039 P3_U8038 ; P3_U3300
g1480 nand P3_U8041 P3_U8040 ; P3_U3301
g1481 nand P3_U8043 P3_U8042 ; P3_U3302
g1482 and P3_ADD_495_U8 P3_U2356 ; P3_U3303
g1483 nand P3_U8045 P3_U8044 ; P3_U3304
g1484 nand P3_U8047 P3_U8046 ; P3_U3305
g1485 nand P3_U8049 P3_U8048 ; P3_U3306
g1486 nand P3_U8051 P3_U8050 ; P3_U3307
g1487 nand P3_U8053 P3_U8052 ; P3_U3308
g1488 and P3_U4447 P3_STATE_REG_0__SCAN_IN ; P3_U3309
g1489 and P3_U4456 P3_U3080 ; P3_U3310
g1490 and P3_U4458 P3_U3078 ; P3_U3311
g1491 and P3_STATE_REG_0__SCAN_IN P3_REQUESTPENDING_REG_SCAN_IN ; P3_U3312
g1492 and P3_U4475 P3_U4474 P3_U4473 P3_U4472 ; P3_U3313
g1493 and P3_U4479 P3_U4478 P3_U4477 P3_U4476 ; P3_U3314
g1494 and P3_U4481 P3_U4480 ; P3_U3315
g1495 and P3_U4483 P3_U4482 ; P3_U3316
g1496 and P3_U4487 P3_U4486 P3_U4485 P3_U4484 ; P3_U3317
g1497 and P3_U4492 P3_U4491 P3_U4490 P3_U4489 ; P3_U3318
g1498 and P3_U4496 P3_U4495 P3_U4494 P3_U4493 ; P3_U3319
g1499 and P3_U4498 P3_U4497 ; P3_U3320
g1500 and P3_U4500 P3_U4499 ; P3_U3321
g1501 and P3_U4504 P3_U4503 P3_U4502 P3_U4501 ; P3_U3322
g1502 and P3_U4509 P3_U4508 P3_U4507 P3_U4506 ; P3_U3323
g1503 and P3_U4513 P3_U4512 P3_U4511 P3_U4510 ; P3_U3324
g1504 and P3_U4515 P3_U4514 ; P3_U3325
g1505 and P3_U4517 P3_U4516 ; P3_U3326
g1506 and P3_U4521 P3_U4520 P3_U4519 P3_U4518 ; P3_U3327
g1507 and P3_U4543 P3_U4542 P3_U4541 P3_U4540 ; P3_U3328
g1508 and P3_U4547 P3_U4546 P3_U4545 P3_U4544 ; P3_U3329
g1509 and P3_U4549 P3_U4548 ; P3_U3330
g1510 and P3_U4551 P3_U4550 ; P3_U3331
g1511 and P3_U4555 P3_U4554 P3_U4553 P3_U4552 ; P3_U3332
g1512 and P3_U4560 P3_U4559 P3_U4558 P3_U4557 ; P3_U3333
g1513 and P3_U4564 P3_U4563 P3_U4562 P3_U4561 ; P3_U3334
g1514 and P3_U4566 P3_U4565 ; P3_U3335
g1515 and P3_U4568 P3_U4567 ; P3_U3336
g1516 and P3_U4572 P3_U4571 P3_U4570 P3_U4569 ; P3_U3337
g1517 and P3_U4526 P3_U4525 P3_U4524 P3_U4523 ; P3_U3338
g1518 and P3_U4530 P3_U4529 P3_U4528 P3_U4527 ; P3_U3339
g1519 and P3_U4532 P3_U4531 ; P3_U3340
g1520 and P3_U4534 P3_U4533 ; P3_U3341
g1521 and P3_U4538 P3_U4537 P3_U4536 P3_U4535 ; P3_U3342
g1522 and P3_U4594 P3_U4593 P3_U4592 P3_U4591 ; P3_U3343
g1523 and P3_U4598 P3_U4597 P3_U4596 P3_U4595 ; P3_U3344
g1524 and P3_U4600 P3_U4599 ; P3_U3345
g1525 and P3_U4602 P3_U4601 ; P3_U3346
g1526 and P3_U4606 P3_U4605 P3_U4604 P3_U4603 ; P3_U3347
g1527 and P3_U4577 P3_U4576 P3_U4575 P3_U4574 ; P3_U3348
g1528 and P3_U4581 P3_U4580 P3_U4579 P3_U4578 ; P3_U3349
g1529 and P3_U4583 P3_U4582 ; P3_U3350
g1530 and P3_U4585 P3_U4584 ; P3_U3351
g1531 and P3_U4589 P3_U4588 P3_U4587 P3_U4586 ; P3_U3352
g1532 and P3_U2352 P3_U4293 ; P3_U3353
g1533 and P3_U4556 P3_U3218 ; P3_U3354
g1534 and P3_U4323 P3_U3101 ; P3_U3355
g1535 and P3_U4324 P3_U3101 ; P3_U3356
g1536 and P3_U4612 P3_U4611 P3_U4610 P3_U4609 ; P3_U3357
g1537 and P3_U4616 P3_U4615 P3_U4614 P3_U4613 ; P3_U3358
g1538 and P3_U4539 P3_U2630 ; P3_U3359
g1539 and P3_U3107 P3_U3108 P3_U3218 ; P3_U3360
g1540 and P3_U3235 P3_U3236 P3_U4621 ; P3_U3361
g1541 and P3_U4626 P3_U3089 ; P3_U3362
g1542 and P3_U4631 P3_U3124 ; P3_U3363
g1543 and P3_U4340 P3_U2630 ; P3_U3364
g1544 and P3_STATE2_REG_3__SCAN_IN P3_STATE2_REG_0__SCAN_IN ; P3_U3365
g1545 and P3_U4338 P3_U4328 ; P3_U3366
g1546 and P3_U3366 P3_U4639 ; P3_U3367
g1547 and P3_U3165 P3_U4659 ; P3_U3368
g1548 and P3_U4671 P3_U4312 ; P3_U3369
g1549 and P3_U4676 P3_U4675 ; P3_U3370
g1550 and P3_U3370 P3_U4677 ; P3_U3371
g1551 and P3_U4681 P3_U4680 ; P3_U3372
g1552 and P3_U3372 P3_U4682 ; P3_U3373
g1553 and P3_U4686 P3_U4685 ; P3_U3374
g1554 and P3_U3374 P3_U4687 ; P3_U3375
g1555 and P3_U4691 P3_U4690 ; P3_U3376
g1556 and P3_U3376 P3_U4692 ; P3_U3377
g1557 and P3_U4696 P3_U4695 ; P3_U3378
g1558 and P3_U3378 P3_U4697 ; P3_U3379
g1559 and P3_U4701 P3_U4700 ; P3_U3380
g1560 and P3_U3380 P3_U4702 ; P3_U3381
g1561 and P3_U4706 P3_U4705 ; P3_U3382
g1562 and P3_U3382 P3_U4707 ; P3_U3383
g1563 and P3_U4711 P3_U4710 ; P3_U3384
g1564 and P3_U3384 P3_U4712 ; P3_U3385
g1565 and P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3386
g1566 and P3_U4723 P3_U4312 ; P3_U3387
g1567 and P3_U4728 P3_U4727 ; P3_U3388
g1568 and P3_U3388 P3_U4729 ; P3_U3389
g1569 and P3_U4733 P3_U4732 ; P3_U3390
g1570 and P3_U3390 P3_U4734 ; P3_U3391
g1571 and P3_U4738 P3_U4737 ; P3_U3392
g1572 and P3_U3392 P3_U4739 ; P3_U3393
g1573 and P3_U4743 P3_U4742 ; P3_U3394
g1574 and P3_U3394 P3_U4744 ; P3_U3395
g1575 and P3_U4748 P3_U4747 ; P3_U3396
g1576 and P3_U3396 P3_U4749 ; P3_U3397
g1577 and P3_U4753 P3_U4752 ; P3_U3398
g1578 and P3_U3398 P3_U4754 ; P3_U3399
g1579 and P3_U4758 P3_U4757 ; P3_U3400
g1580 and P3_U3400 P3_U4759 ; P3_U3401
g1581 and P3_U4763 P3_U4762 ; P3_U3402
g1582 and P3_U3402 P3_U4764 ; P3_U3403
g1583 and P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U3404
g1584 and P3_U4775 P3_U4312 ; P3_U3405
g1585 and P3_U4780 P3_U4779 ; P3_U3406
g1586 and P3_U3406 P3_U4781 ; P3_U3407
g1587 and P3_U4785 P3_U4784 ; P3_U3408
g1588 and P3_U3408 P3_U4786 ; P3_U3409
g1589 and P3_U4790 P3_U4789 ; P3_U3410
g1590 and P3_U3410 P3_U4791 ; P3_U3411
g1591 and P3_U4795 P3_U4794 ; P3_U3412
g1592 and P3_U3412 P3_U4796 ; P3_U3413
g1593 and P3_U4800 P3_U4799 ; P3_U3414
g1594 and P3_U3414 P3_U4801 ; P3_U3415
g1595 and P3_U4805 P3_U4804 ; P3_U3416
g1596 and P3_U3416 P3_U4806 ; P3_U3417
g1597 and P3_U4810 P3_U4809 ; P3_U3418
g1598 and P3_U3418 P3_U4811 ; P3_U3419
g1599 and P3_U4815 P3_U4814 ; P3_U3420
g1600 and P3_U3420 P3_U4816 ; P3_U3421
g1601 and P3_U3129 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U3422
g1602 and P3_U4826 P3_U4312 ; P3_U3423
g1603 and P3_U4831 P3_U4830 ; P3_U3424
g1604 and P3_U3424 P3_U4832 ; P3_U3425
g1605 and P3_U4836 P3_U4835 ; P3_U3426
g1606 and P3_U3426 P3_U4837 ; P3_U3427
g1607 and P3_U4841 P3_U4840 ; P3_U3428
g1608 and P3_U3428 P3_U4842 ; P3_U3429
g1609 and P3_U4846 P3_U4845 ; P3_U3430
g1610 and P3_U3430 P3_U4847 ; P3_U3431
g1611 and P3_U4851 P3_U4850 ; P3_U3432
g1612 and P3_U3432 P3_U4852 ; P3_U3433
g1613 and P3_U4856 P3_U4855 ; P3_U3434
g1614 and P3_U3434 P3_U4857 ; P3_U3435
g1615 and P3_U4861 P3_U4860 ; P3_U3436
g1616 and P3_U3436 P3_U4862 ; P3_U3437
g1617 and P3_U4866 P3_U4865 ; P3_U3438
g1618 and P3_U3438 P3_U4867 ; P3_U3439
g1619 and P3_U4878 P3_U4312 ; P3_U3440
g1620 and P3_U4883 P3_U4882 ; P3_U3441
g1621 and P3_U3441 P3_U4884 ; P3_U3442
g1622 and P3_U4888 P3_U4887 ; P3_U3443
g1623 and P3_U3443 P3_U4889 ; P3_U3444
g1624 and P3_U4893 P3_U4892 ; P3_U3445
g1625 and P3_U3445 P3_U4894 ; P3_U3446
g1626 and P3_U4898 P3_U4897 ; P3_U3447
g1627 and P3_U3447 P3_U4899 ; P3_U3448
g1628 and P3_U4903 P3_U4902 ; P3_U3449
g1629 and P3_U3449 P3_U4904 ; P3_U3450
g1630 and P3_U4908 P3_U4907 ; P3_U3451
g1631 and P3_U3451 P3_U4909 ; P3_U3452
g1632 and P3_U4913 P3_U4912 ; P3_U3453
g1633 and P3_U3453 P3_U4914 ; P3_U3454
g1634 and P3_U4918 P3_U4917 ; P3_U3455
g1635 and P3_U3455 P3_U4919 ; P3_U3456
g1636 and P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3457
g1637 and P3_U4930 P3_U4312 ; P3_U3458
g1638 and P3_U4935 P3_U4934 ; P3_U3459
g1639 and P3_U3459 P3_U4936 ; P3_U3460
g1640 and P3_U4940 P3_U4939 ; P3_U3461
g1641 and P3_U3461 P3_U4941 ; P3_U3462
g1642 and P3_U4945 P3_U4944 ; P3_U3463
g1643 and P3_U3463 P3_U4946 ; P3_U3464
g1644 and P3_U4950 P3_U4949 ; P3_U3465
g1645 and P3_U3465 P3_U4951 ; P3_U3466
g1646 and P3_U4955 P3_U4954 ; P3_U3467
g1647 and P3_U3467 P3_U4956 ; P3_U3468
g1648 and P3_U4960 P3_U4959 ; P3_U3469
g1649 and P3_U3469 P3_U4961 ; P3_U3470
g1650 and P3_U4965 P3_U4964 ; P3_U3471
g1651 and P3_U3471 P3_U4966 ; P3_U3472
g1652 and P3_U4970 P3_U4969 ; P3_U3473
g1653 and P3_U3473 P3_U4971 ; P3_U3474
g1654 and P3_U3131 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U3475
g1655 and P3_U4982 P3_U4312 ; P3_U3476
g1656 and P3_U4987 P3_U4986 ; P3_U3477
g1657 and P3_U3477 P3_U4988 ; P3_U3478
g1658 and P3_U4992 P3_U4991 ; P3_U3479
g1659 and P3_U3479 P3_U4993 ; P3_U3480
g1660 and P3_U4997 P3_U4996 ; P3_U3481
g1661 and P3_U3481 P3_U4998 ; P3_U3482
g1662 and P3_U5002 P3_U5001 ; P3_U3483
g1663 and P3_U3483 P3_U5003 ; P3_U3484
g1664 and P3_U5007 P3_U5006 ; P3_U3485
g1665 and P3_U3485 P3_U5008 ; P3_U3486
g1666 and P3_U5012 P3_U5011 ; P3_U3487
g1667 and P3_U3487 P3_U5013 ; P3_U3488
g1668 and P3_U5017 P3_U5016 ; P3_U3489
g1669 and P3_U3489 P3_U5018 ; P3_U3490
g1670 and P3_U5022 P3_U5021 ; P3_U3491
g1671 and P3_U3491 P3_U5023 ; P3_U3492
g1672 and P3_U5033 P3_U4312 ; P3_U3493
g1673 and P3_U5038 P3_U5037 ; P3_U3494
g1674 and P3_U3494 P3_U5039 ; P3_U3495
g1675 and P3_U5043 P3_U5042 ; P3_U3496
g1676 and P3_U3496 P3_U5044 ; P3_U3497
g1677 and P3_U5048 P3_U5047 ; P3_U3498
g1678 and P3_U3498 P3_U5049 ; P3_U3499
g1679 and P3_U5053 P3_U5052 ; P3_U3500
g1680 and P3_U3500 P3_U5054 ; P3_U3501
g1681 and P3_U5058 P3_U5057 ; P3_U3502
g1682 and P3_U3502 P3_U5059 ; P3_U3503
g1683 and P3_U5063 P3_U5062 ; P3_U3504
g1684 and P3_U3504 P3_U5064 ; P3_U3505
g1685 and P3_U5068 P3_U5067 ; P3_U3506
g1686 and P3_U3506 P3_U5069 ; P3_U3507
g1687 and P3_U5073 P3_U5072 ; P3_U3508
g1688 and P3_U3508 P3_U5074 ; P3_U3509
g1689 and P3_U5082 P3_U4312 ; P3_U3510
g1690 and P3_U5087 P3_U5086 ; P3_U3511
g1691 and P3_U3511 P3_U5088 ; P3_U3512
g1692 and P3_U5092 P3_U5091 ; P3_U3513
g1693 and P3_U3513 P3_U5093 ; P3_U3514
g1694 and P3_U5097 P3_U5096 ; P3_U3515
g1695 and P3_U3515 P3_U5098 ; P3_U3516
g1696 and P3_U5102 P3_U5101 ; P3_U3517
g1697 and P3_U3517 P3_U5103 ; P3_U3518
g1698 and P3_U5107 P3_U5106 ; P3_U3519
g1699 and P3_U3519 P3_U5108 ; P3_U3520
g1700 and P3_U5112 P3_U5111 ; P3_U3521
g1701 and P3_U3521 P3_U5113 ; P3_U3522
g1702 and P3_U5117 P3_U5116 ; P3_U3523
g1703 and P3_U3523 P3_U5118 ; P3_U3524
g1704 and P3_U5122 P3_U5121 ; P3_U3525
g1705 and P3_U3525 P3_U5123 ; P3_U3526
g1706 and P3_U3133 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3527
g1707 and P3_U5134 P3_U4312 ; P3_U3528
g1708 and P3_U5139 P3_U5138 ; P3_U3529
g1709 and P3_U3529 P3_U5140 ; P3_U3530
g1710 and P3_U5144 P3_U5143 ; P3_U3531
g1711 and P3_U3531 P3_U5145 ; P3_U3532
g1712 and P3_U5149 P3_U5148 ; P3_U3533
g1713 and P3_U3533 P3_U5150 ; P3_U3534
g1714 and P3_U5154 P3_U5153 ; P3_U3535
g1715 and P3_U3535 P3_U5155 ; P3_U3536
g1716 and P3_U5159 P3_U5158 ; P3_U3537
g1717 and P3_U3537 P3_U5160 ; P3_U3538
g1718 and P3_U5164 P3_U5163 ; P3_U3539
g1719 and P3_U3539 P3_U5165 ; P3_U3540
g1720 and P3_U5169 P3_U5168 ; P3_U3541
g1721 and P3_U3541 P3_U5170 ; P3_U3542
g1722 and P3_U5174 P3_U5173 ; P3_U3543
g1723 and P3_U3543 P3_U5175 ; P3_U3544
g1724 and P3_U3133 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U3545
g1725 and P3_U5186 P3_U4312 ; P3_U3546
g1726 and P3_U5191 P3_U5190 ; P3_U3547
g1727 and P3_U3547 P3_U5192 ; P3_U3548
g1728 and P3_U5196 P3_U5195 ; P3_U3549
g1729 and P3_U3549 P3_U5197 ; P3_U3550
g1730 and P3_U5201 P3_U5200 ; P3_U3551
g1731 and P3_U3551 P3_U5202 ; P3_U3552
g1732 and P3_U5206 P3_U5205 ; P3_U3553
g1733 and P3_U3553 P3_U5207 ; P3_U3554
g1734 and P3_U5211 P3_U5210 ; P3_U3555
g1735 and P3_U3555 P3_U5212 ; P3_U3556
g1736 and P3_U5216 P3_U5215 ; P3_U3557
g1737 and P3_U3557 P3_U5217 ; P3_U3558
g1738 and P3_U5221 P3_U5220 ; P3_U3559
g1739 and P3_U3559 P3_U5222 ; P3_U3560
g1740 and P3_U5226 P3_U5225 ; P3_U3561
g1741 and P3_U3561 P3_U5227 ; P3_U3562
g1742 nor P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3563
g1743 and P3_U5237 P3_U4312 ; P3_U3564
g1744 and P3_U5241 P3_U5240 P3_U5243 ; P3_U3565
g1745 and P3_U3565 P3_U5242 ; P3_U3566
g1746 and P3_U5246 P3_U5245 P3_U5248 ; P3_U3567
g1747 and P3_U3567 P3_U5247 ; P3_U3568
g1748 and P3_U5251 P3_U5250 P3_U5253 ; P3_U3569
g1749 and P3_U3569 P3_U5252 ; P3_U3570
g1750 and P3_U5256 P3_U5255 P3_U5258 ; P3_U3571
g1751 and P3_U3571 P3_U5257 ; P3_U3572
g1752 and P3_U5261 P3_U5260 P3_U5263 ; P3_U3573
g1753 and P3_U3573 P3_U5262 ; P3_U3574
g1754 and P3_U5266 P3_U5265 P3_U5268 ; P3_U3575
g1755 and P3_U3575 P3_U5267 ; P3_U3576
g1756 and P3_U5271 P3_U5270 P3_U5273 ; P3_U3577
g1757 and P3_U3577 P3_U5272 ; P3_U3578
g1758 and P3_U5276 P3_U5275 P3_U5278 ; P3_U3579
g1759 and P3_U3579 P3_U5277 ; P3_U3580
g1760 nor P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U3581
g1761 and P3_U5288 P3_U4312 ; P3_U3582
g1762 and P3_U5292 P3_U5291 P3_U5294 ; P3_U3583
g1763 and P3_U3583 P3_U5293 ; P3_U3584
g1764 and P3_U5297 P3_U5296 P3_U5299 ; P3_U3585
g1765 and P3_U3585 P3_U5298 ; P3_U3586
g1766 and P3_U5302 P3_U5301 P3_U5304 ; P3_U3587
g1767 and P3_U3587 P3_U5303 ; P3_U3588
g1768 and P3_U5307 P3_U5306 P3_U5309 ; P3_U3589
g1769 and P3_U3589 P3_U5308 ; P3_U3590
g1770 and P3_U5312 P3_U5311 P3_U5314 ; P3_U3591
g1771 and P3_U3591 P3_U5313 ; P3_U3592
g1772 and P3_U5317 P3_U5316 P3_U5319 ; P3_U3593
g1773 and P3_U3593 P3_U5318 ; P3_U3594
g1774 and P3_U5322 P3_U5321 P3_U5324 ; P3_U3595
g1775 and P3_U3595 P3_U5323 ; P3_U3596
g1776 and P3_U5327 P3_U5326 P3_U5329 ; P3_U3597
g1777 and P3_U3597 P3_U5328 ; P3_U3598
g1778 and P3_U5339 P3_U4312 ; P3_U3599
g1779 and P3_U5343 P3_U5342 P3_U5345 ; P3_U3600
g1780 and P3_U3600 P3_U5344 ; P3_U3601
g1781 and P3_U5348 P3_U5347 P3_U5350 ; P3_U3602
g1782 and P3_U3602 P3_U5349 ; P3_U3603
g1783 and P3_U5353 P3_U5352 P3_U5355 ; P3_U3604
g1784 and P3_U3604 P3_U5354 ; P3_U3605
g1785 and P3_U5358 P3_U5357 P3_U5360 ; P3_U3606
g1786 and P3_U3606 P3_U5359 ; P3_U3607
g1787 and P3_U5363 P3_U5362 P3_U5365 ; P3_U3608
g1788 and P3_U3608 P3_U5364 ; P3_U3609
g1789 and P3_U5368 P3_U5367 P3_U5370 ; P3_U3610
g1790 and P3_U3610 P3_U5369 ; P3_U3611
g1791 and P3_U5373 P3_U5372 P3_U5375 ; P3_U3612
g1792 and P3_U3612 P3_U5374 ; P3_U3613
g1793 and P3_U5378 P3_U5377 P3_U5380 ; P3_U3614
g1794 and P3_U3614 P3_U5379 ; P3_U3615
g1795 nor P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U3616
g1796 and P3_U5390 P3_U4312 ; P3_U3617
g1797 and P3_U5394 P3_U5393 P3_U5396 ; P3_U3618
g1798 and P3_U3618 P3_U5395 ; P3_U3619
g1799 and P3_U5399 P3_U5398 P3_U5401 ; P3_U3620
g1800 and P3_U3620 P3_U5400 ; P3_U3621
g1801 and P3_U5404 P3_U5403 P3_U5406 ; P3_U3622
g1802 and P3_U3622 P3_U5405 ; P3_U3623
g1803 and P3_U5409 P3_U5408 P3_U5411 ; P3_U3624
g1804 and P3_U3624 P3_U5410 ; P3_U3625
g1805 and P3_U5414 P3_U5413 P3_U5416 ; P3_U3626
g1806 and P3_U3626 P3_U5415 ; P3_U3627
g1807 and P3_U5419 P3_U5418 P3_U5421 ; P3_U3628
g1808 and P3_U3628 P3_U5420 ; P3_U3629
g1809 and P3_U5424 P3_U5423 P3_U5426 ; P3_U3630
g1810 and P3_U3630 P3_U5425 ; P3_U3631
g1811 and P3_U5429 P3_U5428 P3_U5431 ; P3_U3632
g1812 and P3_U3632 P3_U5430 ; P3_U3633
g1813 nor P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U3634
g1814 and P3_U5440 P3_U4312 ; P3_U3635
g1815 and P3_U5444 P3_U5443 P3_U5446 ; P3_U3636
g1816 and P3_U3636 P3_U5445 ; P3_U3637
g1817 and P3_U5449 P3_U5448 P3_U5451 ; P3_U3638
g1818 and P3_U3638 P3_U5450 ; P3_U3639
g1819 and P3_U5454 P3_U5453 P3_U5456 ; P3_U3640
g1820 and P3_U3640 P3_U5455 ; P3_U3641
g1821 and P3_U5459 P3_U5458 P3_U5461 ; P3_U3642
g1822 and P3_U3642 P3_U5460 ; P3_U3643
g1823 and P3_U5464 P3_U5463 P3_U5466 ; P3_U3644
g1824 and P3_U3644 P3_U5465 ; P3_U3645
g1825 and P3_U5469 P3_U5468 P3_U5471 ; P3_U3646
g1826 and P3_U3646 P3_U5470 ; P3_U3647
g1827 and P3_U5474 P3_U5473 P3_U5476 ; P3_U3648
g1828 and P3_U3648 P3_U5475 ; P3_U3649
g1829 and P3_U5479 P3_U5478 P3_U5481 ; P3_U3650
g1830 and P3_U3650 P3_U5480 ; P3_U3651
g1831 and P3_U4340 P3_ADD_495_U8 ; P3_U3652
g1832 and P3_STATE2_REG_0__SCAN_IN P3_FLUSH_REG_SCAN_IN ; P3_U3653
g1833 and P3_U4522 P3_U3104 ; P3_U3654
g1834 and P3_U3107 P3_U3118 ; P3_U3655
g1835 and P3_U5495 P3_U4333 ; P3_U3656
g1836 and P3_U3656 P3_U5494 ; P3_U3657
g1837 and P3_U5498 P3_U4330 ; P3_U3658
g1838 and P3_U5502 P3_U5501 ; P3_U3659
g1839 and P3_U4556 P3_U4539 ; P3_U3660
g1840 and P3_U2461 P3_U4297 ; P3_U3661
g1841 and P3_U4590 P3_U3101 ; P3_U3662
g1842 and P3_U4556 P3_U3101 ; P3_U3663
g1843 and P3_U4573 P3_U4324 ; P3_U3664
g1844 and P3_U5511 P3_U5510 P3_U5508 ; P3_U3665
g1845 and P3_U5519 P3_U4339 P3_U5520 ; P3_U3666
g1846 and P3_U7978 P3_U7977 P3_U5521 P3_U3666 ; P3_U3667
g1847 and P3_U5528 P3_U3242 P3_U2517 ; P3_U3668
g1848 and P3_U4470 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U3669
g1849 and P3_U3093 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U3670
g1850 and P3_U3116 P3_U3117 P3_U3119 ; P3_U3671
g1851 and P3_U3245 P3_U3244 P3_U3671 ; P3_U3672
g1852 and P3_U4505 P3_U2456 ; P3_U3673
g1853 and P3_U5533 P3_U5532 ; P3_U3674
g1854 and P3_U5538 P3_U5536 ; P3_U3675
g1855 and P3_U3677 P3_U5539 P3_U3675 ; P3_U3676
g1856 and P3_U5540 P3_U5541 ; P3_U3677
g1857 and P3_U5552 P3_U5550 ; P3_U3678
g1858 and P3_U3678 P3_U5551 ; P3_U3679
g1859 and P3_U5555 P3_U5554 ; P3_U3680
g1860 and P3_U3682 P3_U5562 ; P3_U3681
g1861 and P3_U5565 P3_U5564 ; P3_U3682
g1862 and P3_U5568 P3_U5567 ; P3_U3683
g1863 and P3_U5576 P3_U5574 ; P3_U3684
g1864 and P3_U5587 P3_U5588 ; P3_U3685
g1865 and P3_U5594 P3_U5592 ; P3_U3686
g1866 and P3_U5625 P3_U4333 P3_U5626 ; P3_U3687
g1867 and P3_U2456 P3_U4296 ; P3_U3688
g1868 and P3_U2456 P3_U4323 ; P3_U3689
g1869 and P3_U4608 P3_U4556 ; P3_U3690
g1870 and P3_U2456 P3_U4590 ; P3_U3691
g1871 and P3_U5636 P3_U5635 ; P3_U3692
g1872 and P3_U5638 P3_U5637 P3_U3694 P3_U5633 P3_U5632 ; P3_U3693
g1873 and P3_U3695 P3_U5641 ; P3_U3694
g1874 and P3_U5639 P3_U5640 ; P3_U3695
g1875 and P3_U5643 P3_U5642 P3_U5644 P3_U5646 P3_U5645 ; P3_U3696
g1876 and P3_U5648 P3_U5649 P3_U5647 P3_U5651 P3_U5650 ; P3_U3697
g1877 and P3_U3697 P3_U3696 ; P3_U3698
g1878 and P3_U5660 P3_U5659 ; P3_U3699
g1879 and P3_U5662 P3_U5661 P3_U3701 P3_U5657 ; P3_U3700
g1880 and P3_U3702 P3_U5665 ; P3_U3701
g1881 and P3_U5663 P3_U5664 ; P3_U3702
g1882 and P3_U5667 P3_U5666 P3_U5668 P3_U5670 P3_U5669 ; P3_U3703
g1883 and P3_U5674 P3_U5671 P3_U5672 P3_U5673 ; P3_U3704
g1884 and P3_U3704 P3_U3703 P3_U5675 ; P3_U3705
g1885 and P3_U3707 P3_U5681 ; P3_U3706
g1886 and P3_U5684 P3_U5683 ; P3_U3707
g1887 and P3_U3709 P3_U5689 ; P3_U3708
g1888 and P3_U5687 P3_U5688 ; P3_U3709
g1889 and P3_U5686 P3_U5685 P3_U3708 ; P3_U3710
g1890 and P3_U5691 P3_U5690 P3_U5692 P3_U5694 P3_U5693 ; P3_U3711
g1891 and P3_U5698 P3_U5695 P3_U5696 P3_U5697 ; P3_U3712
g1892 and P3_U3712 P3_U3711 P3_U5699 ; P3_U3713
g1893 and P3_U5705 P3_U5704 ; P3_U3714
g1894 and P3_U5708 P3_U5707 ; P3_U3715
g1895 and P3_U3717 P3_U5713 ; P3_U3716
g1896 and P3_U5711 P3_U5712 ; P3_U3717
g1897 and P3_U5710 P3_U5709 P3_U3716 ; P3_U3718
g1898 and P3_U5715 P3_U5714 P3_U5716 P3_U5718 P3_U5717 ; P3_U3719
g1899 and P3_U5722 P3_U5719 P3_U5720 P3_U5721 ; P3_U3720
g1900 and P3_U3720 P3_U3719 P3_U5723 ; P3_U3721
g1901 and P3_U3723 P3_U5729 ; P3_U3722
g1902 and P3_U5732 P3_U5731 ; P3_U3723
g1903 and P3_U3725 P3_U5737 ; P3_U3724
g1904 and P3_U5735 P3_U5736 ; P3_U3725
g1905 and P3_U5734 P3_U5733 P3_U3724 ; P3_U3726
g1906 and P3_U5739 P3_U5738 P3_U5740 P3_U5742 P3_U5741 ; P3_U3727
g1907 and P3_U5746 P3_U5743 P3_U5744 P3_U5745 ; P3_U3728
g1908 and P3_U3728 P3_U3727 P3_U5747 ; P3_U3729
g1909 and P3_U3731 P3_U5752 ; P3_U3730
g1910 and P3_U5756 P3_U5755 ; P3_U3731
g1911 and P3_U3733 P3_U5761 ; P3_U3732
g1912 and P3_U5759 P3_U5760 ; P3_U3733
g1913 and P3_U5758 P3_U5757 P3_U3732 ; P3_U3734
g1914 and P3_U5763 P3_U5762 P3_U5764 P3_U5766 P3_U5765 ; P3_U3735
g1915 and P3_U5770 P3_U5767 P3_U5768 P3_U5769 ; P3_U3736
g1916 and P3_U3736 P3_U3735 P3_U5771 ; P3_U3737
g1917 and P3_U3739 P3_U5776 ; P3_U3738
g1918 and P3_U5780 P3_U5779 ; P3_U3739
g1919 and P3_U3741 P3_U5785 ; P3_U3740
g1920 and P3_U5783 P3_U5784 ; P3_U3741
g1921 and P3_U5782 P3_U5781 P3_U3740 ; P3_U3742
g1922 and P3_U5787 P3_U5786 P3_U5788 P3_U5790 P3_U5789 ; P3_U3743
g1923 and P3_U5794 P3_U5791 P3_U5792 P3_U5793 ; P3_U3744
g1924 and P3_U3744 P3_U3743 P3_U5795 ; P3_U3745
g1925 and P3_U3747 P3_U5800 ; P3_U3746
g1926 and P3_U5804 P3_U5803 ; P3_U3747
g1927 and P3_U3749 P3_U5809 ; P3_U3748
g1928 and P3_U5807 P3_U5808 ; P3_U3749
g1929 and P3_U5806 P3_U5805 P3_U3748 ; P3_U3750
g1930 and P3_U5811 P3_U5810 P3_U5812 P3_U5814 P3_U5813 ; P3_U3751
g1931 and P3_U5818 P3_U5815 P3_U5816 P3_U5817 ; P3_U3752
g1932 and P3_U3752 P3_U3751 P3_U5819 ; P3_U3753
g1933 and P3_U3755 P3_U5824 ; P3_U3754
g1934 and P3_U5828 P3_U5827 ; P3_U3755
g1935 and P3_U5833 P3_U5832 P3_U5831 ; P3_U3756
g1936 and P3_U5830 P3_U5829 P3_U3756 ; P3_U3757
g1937 and P3_U5835 P3_U5834 P3_U5836 P3_U5838 P3_U5837 ; P3_U3758
g1938 and P3_U5842 P3_U5841 P3_U5840 P3_U5839 ; P3_U3759
g1939 and P3_U3759 P3_U3758 P3_U5843 ; P3_U3760
g1940 and P3_U3762 P3_U5848 ; P3_U3761
g1941 and P3_U5852 P3_U5851 ; P3_U3762
g1942 and P3_U5857 P3_U5856 ; P3_U3763
g1943 and P3_U5854 P3_U5853 P3_U5855 P3_U3763 ; P3_U3764
g1944 and P3_U5859 P3_U5858 P3_U5860 P3_U5862 P3_U5861 ; P3_U3765
g1945 and P3_U5866 P3_U5865 P3_U5864 P3_U5863 ; P3_U3766
g1946 and P3_U3766 P3_U3765 P3_U5867 ; P3_U3767
g1947 and P3_U3769 P3_U5873 ; P3_U3768
g1948 and P3_U5876 P3_U5875 ; P3_U3769
g1949 and P3_U5881 P3_U5880 ; P3_U3770
g1950 and P3_U5878 P3_U5877 P3_U5879 P3_U3770 ; P3_U3771
g1951 and P3_U5883 P3_U5882 P3_U5884 P3_U5886 P3_U5885 ; P3_U3772
g1952 and P3_U5890 P3_U5889 P3_U5888 P3_U5887 ; P3_U3773
g1953 and P3_U3773 P3_U3772 P3_U5891 ; P3_U3774
g1954 and P3_U3776 P3_U5897 ; P3_U3775
g1955 and P3_U5900 P3_U5899 ; P3_U3776
g1956 and P3_U5905 P3_U5904 ; P3_U3777
g1957 and P3_U5902 P3_U5901 P3_U5903 P3_U3777 ; P3_U3778
g1958 and P3_U5907 P3_U5906 P3_U5908 P3_U5910 P3_U5909 ; P3_U3779
g1959 and P3_U5914 P3_U5913 P3_U5912 P3_U5911 ; P3_U3780
g1960 and P3_U3780 P3_U3779 P3_U5915 ; P3_U3781
g1961 and P3_U3783 P3_U5920 ; P3_U3782
g1962 and P3_U5924 P3_U5923 ; P3_U3783
g1963 and P3_U5929 P3_U5928 ; P3_U3784
g1964 and P3_U5926 P3_U5925 P3_U5927 P3_U3784 ; P3_U3785
g1965 and P3_U5931 P3_U5930 P3_U5932 P3_U5934 P3_U5933 ; P3_U3786
g1966 and P3_U5938 P3_U5937 P3_U5936 P3_U5935 ; P3_U3787
g1967 and P3_U3787 P3_U3786 P3_U5939 ; P3_U3788
g1968 and P3_U3790 P3_U5944 ; P3_U3789
g1969 and P3_U5948 P3_U5947 ; P3_U3790
g1970 and P3_U5953 P3_U5952 ; P3_U3791
g1971 and P3_U5950 P3_U5949 P3_U5951 P3_U3791 ; P3_U3792
g1972 and P3_U5955 P3_U5954 P3_U5956 P3_U5958 P3_U5957 ; P3_U3793
g1973 and P3_U5962 P3_U5961 P3_U5960 P3_U5959 ; P3_U3794
g1974 and P3_U3794 P3_U3793 P3_U5963 ; P3_U3795
g1975 and P3_U5972 P3_U5971 ; P3_U3796
g1976 and P3_U5977 P3_U5976 ; P3_U3797
g1977 and P3_U5974 P3_U5973 P3_U5975 P3_U3797 ; P3_U3798
g1978 and P3_U3796 P3_U5970 P3_U3798 P3_U5969 P3_U5968 ; P3_U3799
g1979 and P3_U5979 P3_U5978 P3_U5980 P3_U5982 P3_U5981 ; P3_U3800
g1980 and P3_U5986 P3_U5985 P3_U5984 P3_U5983 ; P3_U3801
g1981 and P3_U3801 P3_U3800 P3_U5987 ; P3_U3802
g1982 and P3_U5991 P3_U5989 ; P3_U3803
g1983 and P3_U5996 P3_U5995 ; P3_U3804
g1984 and P3_U6001 P3_U6000 ; P3_U3805
g1985 and P3_U5998 P3_U5997 P3_U5999 P3_U3805 ; P3_U3806
g1986 and P3_U3804 P3_U5994 P3_U3806 P3_U5993 P3_U5992 ; P3_U3807
g1987 and P3_U6003 P3_U6002 P3_U6004 P3_U6006 P3_U6005 ; P3_U3808
g1988 and P3_U6010 P3_U6009 P3_U6008 P3_U6007 ; P3_U3809
g1989 and P3_U3809 P3_U3808 P3_U6011 ; P3_U3810
g1990 and P3_U6015 P3_U6013 ; P3_U3811
g1991 and P3_U3813 P3_U6017 ; P3_U3812
g1992 and P3_U6020 P3_U6019 ; P3_U3813
g1993 and P3_U6025 P3_U6024 ; P3_U3814
g1994 and P3_U6022 P3_U6021 P3_U6023 P3_U3814 ; P3_U3815
g1995 and P3_U6027 P3_U6026 P3_U6028 P3_U6030 P3_U6029 ; P3_U3816
g1996 and P3_U6034 P3_U6033 P3_U6032 P3_U6031 ; P3_U3817
g1997 and P3_U3817 P3_U3816 P3_U6035 ; P3_U3818
g1998 and P3_U6044 P3_U6043 ; P3_U3819
g1999 and P3_U6046 P3_U6045 P3_U6047 P3_U3821 P3_U6041 ; P3_U3820
g2000 and P3_U6049 P3_U6048 ; P3_U3821
g2001 and P3_U6051 P3_U6050 P3_U6052 P3_U6054 P3_U6053 ; P3_U3822
g2002 and P3_U6058 P3_U6057 P3_U6056 P3_U6055 ; P3_U3823
g2003 and P3_U3823 P3_U3822 P3_U6059 ; P3_U3824
g2004 and P3_U3826 P3_U6065 ; P3_U3825
g2005 and P3_U6068 P3_U6067 ; P3_U3826
g2006 and P3_U6073 P3_U6072 ; P3_U3827
g2007 and P3_U6070 P3_U6069 P3_U6071 P3_U3827 ; P3_U3828
g2008 and P3_U6075 P3_U6074 P3_U6076 P3_U6078 P3_U6077 ; P3_U3829
g2009 and P3_U6082 P3_U6081 P3_U6080 P3_U6079 ; P3_U3830
g2010 and P3_U3830 P3_U3829 P3_U6083 ; P3_U3831
g2011 and P3_U6092 P3_U6091 ; P3_U3832
g2012 and P3_U6094 P3_U6093 P3_U6095 P3_U3834 P3_U6089 ; P3_U3833
g2013 and P3_U6097 P3_U6096 ; P3_U3834
g2014 and P3_U6099 P3_U6098 P3_U6100 P3_U6102 P3_U6101 ; P3_U3835
g2015 and P3_U6106 P3_U6105 P3_U6104 P3_U6103 ; P3_U3836
g2016 and P3_U3836 P3_U3835 P3_U6107 ; P3_U3837
g2017 and P3_U6116 P3_U6115 ; P3_U3838
g2018 and P3_U6121 P3_U6120 ; P3_U3839
g2019 and P3_U6118 P3_U6117 P3_U6119 P3_U3839 ; P3_U3840
g2020 and P3_U6114 P3_U3838 P3_U3840 P3_U6112 P3_U3844 ; P3_U3841
g2021 and P3_U6123 P3_U6122 P3_U6124 P3_U6126 P3_U6125 ; P3_U3842
g2022 and P3_U6130 P3_U6129 P3_U6128 P3_U6127 ; P3_U3843
g2023 and P3_U3843 P3_U3842 P3_U6131 ; P3_U3844
g2024 and P3_U6135 P3_U6133 ; P3_U3845
g2025 and P3_U6140 P3_U6139 ; P3_U3846
g2026 and P3_U6145 P3_U6144 ; P3_U3847
g2027 and P3_U6142 P3_U6141 P3_U6143 P3_U3847 ; P3_U3848
g2028 and P3_U6138 P3_U3846 P3_U3848 P3_U6136 P3_U3852 ; P3_U3849
g2029 and P3_U6147 P3_U6146 P3_U6148 P3_U6150 P3_U6149 ; P3_U3850
g2030 and P3_U6154 P3_U6153 P3_U6152 P3_U6151 ; P3_U3851
g2031 and P3_U3850 P3_U3851 P3_U6155 ; P3_U3852
g2032 and P3_U6159 P3_U6157 ; P3_U3853
g2033 and P3_U6164 P3_U6163 ; P3_U3854
g2034 and P3_U6169 P3_U6168 ; P3_U3855
g2035 and P3_U6166 P3_U6165 P3_U6167 P3_U3855 ; P3_U3856
g2036 and P3_U6161 P3_U6162 P3_U3854 P3_U3856 P3_U6160 ; P3_U3857
g2037 and P3_U6171 P3_U6170 P3_U6172 ; P3_U3858
g2038 and P3_U6174 P3_U6173 ; P3_U3859
g2039 and P3_U6176 P3_U6175 P3_U6177 ; P3_U3860
g2040 and P3_U6179 P3_U6178 ; P3_U3861
g2041 and P3_U3859 P3_U3858 P3_U3860 P3_U3861 ; P3_U3862
g2042 and P3_U6183 P3_U6181 ; P3_U3863
g2043 and P3_U6188 P3_U6187 ; P3_U3864
g2044 and P3_U6193 P3_U6192 ; P3_U3865
g2045 and P3_U6190 P3_U6189 P3_U6191 P3_U3865 ; P3_U3866
g2046 and P3_U6185 P3_U6186 P3_U3864 P3_U3866 P3_U6184 ; P3_U3867
g2047 and P3_U6195 P3_U6194 P3_U6196 ; P3_U3868
g2048 and P3_U6198 P3_U6197 ; P3_U3869
g2049 and P3_U6200 P3_U6199 P3_U6201 ; P3_U3870
g2050 and P3_U6203 P3_U6202 ; P3_U3871
g2051 and P3_U3869 P3_U3868 P3_U3870 P3_U3871 ; P3_U3872
g2052 and P3_U6207 P3_U6205 ; P3_U3873
g2053 and P3_U6212 P3_U6211 ; P3_U3874
g2054 and P3_U6217 P3_U6216 ; P3_U3875
g2055 and P3_U6214 P3_U6213 P3_U6215 P3_U3875 ; P3_U3876
g2056 and P3_U6209 P3_U6210 P3_U3874 P3_U6208 P3_U3876 ; P3_U3877
g2057 and P3_U6219 P3_U6218 P3_U6220 ; P3_U3878
g2058 and P3_U6222 P3_U6221 ; P3_U3879
g2059 and P3_U6224 P3_U6223 P3_U6225 ; P3_U3880
g2060 and P3_U6227 P3_U6226 ; P3_U3881
g2061 and P3_U3879 P3_U3878 P3_U3881 P3_U3880 ; P3_U3882
g2062 and P3_U6231 P3_U6229 ; P3_U3883
g2063 and P3_U6236 P3_U6235 ; P3_U3884
g2064 and P3_U6241 P3_U6240 ; P3_U3885
g2065 and P3_U6238 P3_U6237 P3_U6239 P3_U3885 ; P3_U3886
g2066 and P3_U6233 P3_U6234 P3_U6232 P3_U3884 P3_U3886 ; P3_U3887
g2067 and P3_U6243 P3_U6242 P3_U6244 ; P3_U3888
g2068 and P3_U6246 P3_U6245 ; P3_U3889
g2069 and P3_U6248 P3_U6247 P3_U6249 ; P3_U3890
g2070 and P3_U6251 P3_U6250 ; P3_U3891
g2071 and P3_U3889 P3_U3888 P3_U3891 P3_U3890 ; P3_U3892
g2072 and P3_U6255 P3_U6253 ; P3_U3893
g2073 and P3_U6257 P3_U6256 ; P3_U3894
g2074 and P3_U6260 P3_U6259 ; P3_U3895
g2075 and P3_U6265 P3_U6264 ; P3_U3896
g2076 and P3_U6262 P3_U6261 P3_U6263 P3_U3896 ; P3_U3897
g2077 and P3_U6267 P3_U6266 P3_U6268 ; P3_U3898
g2078 and P3_U6270 P3_U6269 ; P3_U3899
g2079 and P3_U6272 P3_U6271 P3_U6273 ; P3_U3900
g2080 and P3_U6275 P3_U6274 ; P3_U3901
g2081 and P3_U3899 P3_U3898 P3_U3901 P3_U3900 ; P3_U3902
g2082 and P3_U6281 P3_U6280 ; P3_U3903
g2083 and P3_U6284 P3_U6283 ; P3_U3904
g2084 and P3_U6289 P3_U6288 ; P3_U3905
g2085 and P3_U6286 P3_U6285 P3_U6287 P3_U3905 ; P3_U3906
g2086 and P3_U6291 P3_U6290 P3_U6292 ; P3_U3907
g2087 and P3_U6294 P3_U6293 ; P3_U3908
g2088 and P3_U6296 P3_U6295 P3_U6297 ; P3_U3909
g2089 and P3_U6299 P3_U6298 ; P3_U3910
g2090 and P3_U3908 P3_U3907 P3_U3910 P3_U3909 ; P3_U3911
g2091 and P3_U6305 P3_U6304 ; P3_U3912
g2092 and P3_U6308 P3_U6307 ; P3_U3913
g2093 and P3_U6313 P3_U6312 ; P3_U3914
g2094 and P3_U6310 P3_U6309 P3_U6311 P3_U3914 ; P3_U3915
g2095 and P3_U6315 P3_U6314 P3_U6316 ; P3_U3916
g2096 and P3_U6318 P3_U6317 ; P3_U3917
g2097 and P3_U6320 P3_U6319 P3_U6321 ; P3_U3918
g2098 and P3_U6323 P3_U6322 ; P3_U3919
g2099 and P3_U3917 P3_U3916 P3_U3919 P3_U3918 ; P3_U3920
g2100 and P3_U6329 P3_U6328 ; P3_U3921
g2101 and P3_U6332 P3_U6331 ; P3_U3922
g2102 and P3_U6337 P3_U6336 ; P3_U3923
g2103 and P3_U6334 P3_U6333 P3_U6335 P3_U3923 ; P3_U3924
g2104 and P3_U6339 P3_U6338 P3_U6340 ; P3_U3925
g2105 and P3_U6342 P3_U6341 ; P3_U3926
g2106 and P3_U6344 P3_U6343 P3_U6345 ; P3_U3927
g2107 and P3_U6347 P3_U6346 ; P3_U3928
g2108 and P3_U3926 P3_U3925 P3_U3928 P3_U3927 ; P3_U3929
g2109 and P3_U6353 P3_U6352 ; P3_U3930
g2110 and P3_U6356 P3_U6355 ; P3_U3931
g2111 and P3_U6361 P3_U6360 ; P3_U3932
g2112 and P3_U6358 P3_U6357 P3_U6359 P3_U3932 ; P3_U3933
g2113 and P3_U6363 P3_U6362 P3_U6364 ; P3_U3934
g2114 and P3_U6366 P3_U6365 ; P3_U3935
g2115 and P3_U6368 P3_U6367 P3_U6369 ; P3_U3936
g2116 and P3_U6371 P3_U6370 ; P3_U3937
g2117 and P3_U3935 P3_U3934 P3_U3937 P3_U3936 ; P3_U3938
g2118 and P3_U6398 P3_U3247 ; P3_U3939
g2119 and P3_U6377 P3_U6376 ; P3_U3940
g2120 and P3_U6380 P3_U6379 ; P3_U3941
g2121 and P3_U3941 P3_U6381 ; P3_U3942
g2122 and P3_U6386 P3_U6385 P3_U6384 ; P3_U3943
g2123 and P3_U6383 P3_U6382 P3_U3943 ; P3_U3944
g2124 and P3_U3940 P3_U6378 P3_U3942 P3_U3944 ; P3_U3945
g2125 and P3_U6388 P3_U6387 P3_U6389 ; P3_U3946
g2126 and P3_U6391 P3_U6390 ; P3_U3947
g2127 and P3_U3946 P3_U6392 P3_U3947 ; P3_U3948
g2128 and P3_U6394 P3_U6393 ; P3_U3949
g2129 and P3_U6398 P3_U6397 P3_U6395 P3_U3949 P3_U3948 ; P3_U3950
g2130 and P3_U3104 P3_STATE2_REG_0__SCAN_IN ; P3_U3951
g2131 and P3_U3121 P3_STATE2_REG_2__SCAN_IN ; P3_U3952
g2132 and P3_U4505 P3_STATE2_REG_0__SCAN_IN ; P3_U3953
g2133 and P3_U6412 P3_U6411 P3_U6410 P3_U6409 ; P3_U3954
g2134 and P3_U6420 P3_U6419 P3_U6418 P3_U6417 ; P3_U3955
g2135 and P3_U6426 P3_U6425 P3_U6428 P3_U6427 ; P3_U3956
g2136 and P3_U6434 P3_U6433 P3_U6436 P3_U6435 ; P3_U3957
g2137 and P3_U6442 P3_U6441 P3_U6444 P3_U6443 ; P3_U3958
g2138 and P3_U6450 P3_U6449 P3_U6452 P3_U6451 ; P3_U3959
g2139 and P3_U6458 P3_U6457 P3_U6460 P3_U6459 ; P3_U3960
g2140 and P3_U6466 P3_U6465 P3_U6468 P3_U6467 ; P3_U3961
g2141 and P3_U6474 P3_U6473 P3_U6476 P3_U6475 ; P3_U3962
g2142 and P3_U6482 P3_U6481 P3_U6484 P3_U6483 ; P3_U3963
g2143 and P3_U6490 P3_U6489 P3_U6492 P3_U6491 ; P3_U3964
g2144 and P3_U6498 P3_U6497 P3_U6500 P3_U6499 ; P3_U3965
g2145 and P3_U6508 P3_U6505 P3_U6506 P3_U6507 ; P3_U3966
g2146 and P3_U6516 P3_U6513 P3_U6514 P3_U6515 ; P3_U3967
g2147 and P3_U6524 P3_U6521 P3_U6522 P3_U6523 ; P3_U3968
g2148 and P3_U6532 P3_U6529 P3_U6530 P3_U6531 ; P3_U3969
g2149 and P3_U6540 P3_U6537 P3_U6538 P3_U6539 ; P3_U3970
g2150 and P3_U6548 P3_U6545 P3_U6546 P3_U6547 ; P3_U3971
g2151 and P3_U6556 P3_U6553 P3_U6554 P3_U6555 ; P3_U3972
g2152 and P3_U6564 P3_U6561 P3_U6562 P3_U6563 ; P3_U3973
g2153 and P3_U6572 P3_U6569 P3_U6570 P3_U6571 ; P3_U3974
g2154 and P3_U6580 P3_U6577 P3_U6578 P3_U6579 ; P3_U3975
g2155 and P3_U6588 P3_U6585 P3_U6586 P3_U6587 ; P3_U3976
g2156 and P3_U6596 P3_U6593 P3_U6594 P3_U6595 ; P3_U3977
g2157 and P3_U6604 P3_U6601 P3_U6602 P3_U6603 ; P3_U3978
g2158 and P3_U6612 P3_U6609 P3_U6610 P3_U6611 ; P3_U3979
g2159 and P3_U6620 P3_U6619 P3_U6618 P3_U6617 ; P3_U3980
g2160 and P3_U6628 P3_U6627 P3_U6626 P3_U6625 ; P3_U3981
g2161 and P3_U6636 P3_U6635 P3_U6634 P3_U6633 ; P3_U3982
g2162 and P3_U6644 P3_U6641 P3_U6643 P3_U6642 ; P3_U3983
g2163 and P3_U6652 P3_U6649 P3_U6651 P3_U6650 ; P3_U3984
g2164 and P3_U6660 P3_U6657 P3_U6659 P3_U6658 ; P3_U3985
g2165 and P3_U4293 P3_U2390 ; P3_U3986
g2166 and P3_U6809 P3_U6810 ; P3_U3987
g2167 and P3_U6812 P3_U6813 ; P3_U3988
g2168 and P3_U6815 P3_U6816 ; P3_U3989
g2169 and P3_U6818 P3_U6819 ; P3_U3990
g2170 and P3_U6821 P3_U6822 ; P3_U3991
g2171 and P3_U6824 P3_U6825 ; P3_U3992
g2172 and P3_U6827 P3_U6828 ; P3_U3993
g2173 and P3_U6830 P3_U6831 ; P3_U3994
g2174 and P3_U6833 P3_U6834 ; P3_U3995
g2175 and P3_U6836 P3_U6837 ; P3_U3996
g2176 and P3_U6839 P3_U6840 ; P3_U3997
g2177 and P3_U6842 P3_U6843 ; P3_U3998
g2178 and P3_U6845 P3_U6846 ; P3_U3999
g2179 and P3_U6848 P3_U6849 ; P3_U4000
g2180 and P3_U6851 P3_U6852 ; P3_U4001
g2181 and P3_U6857 P3_U6856 ; P3_U4002
g2182 and P3_U6861 P3_U6860 ; P3_U4003
g2183 and P3_U6865 P3_U6864 ; P3_U4004
g2184 and P3_U6869 P3_U6868 ; P3_U4005
g2185 and P3_U6873 P3_U6872 ; P3_U4006
g2186 and P3_U6877 P3_U6876 ; P3_U4007
g2187 and P3_U6881 P3_U6880 ; P3_U4008
g2188 and P3_U6885 P3_U6884 ; P3_U4009
g2189 and P3_U6889 P3_U6888 ; P3_U4010
g2190 and P3_U6893 P3_U6892 ; P3_U4011
g2191 and P3_U6897 P3_U6896 ; P3_U4012
g2192 and P3_U6901 P3_U6900 ; P3_U4013
g2193 and P3_U6905 P3_U6904 ; P3_U4014
g2194 and P3_U6907 P3_U6909 ; P3_U4015
g2195 and P3_U6911 P3_U6913 ; P3_U4016
g2196 and P3_U6915 P3_U6917 ; P3_U4017
g2197 and P3_U6922 P3_U6920 ; P3_U4018
g2198 and P3_U6927 P3_U6925 ; P3_U4019
g2199 and P3_U6932 P3_U6930 ; P3_U4020
g2200 and P3_U6937 P3_U6935 ; P3_U4021
g2201 and P3_U6942 P3_U6940 ; P3_U4022
g2202 and P3_U6947 P3_U6945 ; P3_U4023
g2203 and P3_U6952 P3_U6950 ; P3_U4024
g2204 and P3_U6957 P3_U6955 ; P3_U4025
g2205 and P3_U6962 P3_U6960 ; P3_U4026
g2206 and P3_U6967 P3_U6965 ; P3_U4027
g2207 and P3_U6972 P3_U6970 ; P3_U4028
g2208 and P3_U6977 P3_U6975 ; P3_U4029
g2209 and P3_U4329 P3_U4328 P3_U4336 ; P3_U4030
g2210 and P3_U7098 P3_U7097 P3_U4032 ; P3_U4031
g2211 and P3_U7101 P3_U7100 ; P3_U4032
g2212 and P3_U4034 P3_U7104 ; P3_U4033
g2213 and P3_U7106 P3_U7105 ; P3_U4034
g2214 and P3_U7108 P3_U7107 P3_U4036 ; P3_U4035
g2215 and P3_U7111 P3_U7110 ; P3_U4036
g2216 and P3_U4038 P3_U7114 ; P3_U4037
g2217 and P3_U7116 P3_U7115 ; P3_U4038
g2218 and P3_U7118 P3_U7117 P3_U4040 ; P3_U4039
g2219 and P3_U7121 P3_U7120 ; P3_U4040
g2220 and P3_U4042 P3_U7124 ; P3_U4041
g2221 and P3_U7126 P3_U7125 ; P3_U4042
g2222 and P3_U7128 P3_U7127 P3_U4044 ; P3_U4043
g2223 and P3_U7131 P3_U7130 ; P3_U4044
g2224 and P3_U4046 P3_U7134 ; P3_U4045
g2225 and P3_U7136 P3_U7135 ; P3_U4046
g2226 and P3_U7137 P3_U4316 P3_U7138 ; P3_U4047
g2227 and P3_U7140 P3_U7141 ; P3_U4048
g2228 and P3_U4050 P3_U7144 ; P3_U4049
g2229 and P3_U7146 P3_U7145 ; P3_U4050
g2230 and P3_U4048 P3_U7139 P3_U4047 P3_U7142 P3_U7143 ; P3_U4051
g2231 and P3_U7147 P3_U4316 P3_U7148 ; P3_U4052
g2232 and P3_U7150 P3_U7151 ; P3_U4053
g2233 and P3_U4055 P3_U7154 ; P3_U4054
g2234 and P3_U7156 P3_U7155 ; P3_U4055
g2235 and P3_U4053 P3_U7149 P3_U4052 P3_U7152 P3_U7153 ; P3_U4056
g2236 and P3_U7157 P3_U4316 P3_U7158 ; P3_U4057
g2237 and P3_U4059 P3_U7161 ; P3_U4058
g2238 and P3_U7164 P3_U7163 ; P3_U4059
g2239 and P3_U7165 P3_U4316 P3_U7166 ; P3_U4060
g2240 and P3_U4062 P3_U7169 ; P3_U4061
g2241 and P3_U7172 P3_U7171 ; P3_U4062
g2242 and P3_U7173 P3_U4316 P3_U7174 ; P3_U4063
g2243 and P3_U4065 P3_U7177 ; P3_U4064
g2244 and P3_U7180 P3_U7179 ; P3_U4065
g2245 and P3_U7181 P3_U4316 P3_U7182 ; P3_U4066
g2246 and P3_U4068 P3_U7185 ; P3_U4067
g2247 and P3_U7188 P3_U7187 ; P3_U4068
g2248 and P3_U7189 P3_U4316 P3_U7190 ; P3_U4069
g2249 and P3_U4071 P3_U7193 ; P3_U4070
g2250 and P3_U7196 P3_U7195 ; P3_U4071
g2251 and P3_U7197 P3_U4316 P3_U7198 ; P3_U4072
g2252 and P3_U4074 P3_U7201 ; P3_U4073
g2253 and P3_U7204 P3_U7203 ; P3_U4074
g2254 and P3_U7205 P3_U4316 P3_U7206 ; P3_U4075
g2255 and P3_U4077 P3_U7209 ; P3_U4076
g2256 and P3_U7212 P3_U7211 ; P3_U4077
g2257 and P3_U7213 P3_U4316 P3_U7214 ; P3_U4078
g2258 and P3_U4080 P3_U7217 ; P3_U4079
g2259 and P3_U7220 P3_U7219 ; P3_U4080
g2260 and P3_U7221 P3_U4316 P3_U7222 ; P3_U4081
g2261 and P3_U4083 P3_U7225 ; P3_U4082
g2262 and P3_U7228 P3_U7227 ; P3_U4083
g2263 and P3_U7229 P3_U4316 P3_U7230 ; P3_U4084
g2264 and P3_U4086 P3_U7233 ; P3_U4085
g2265 and P3_U7236 P3_U7235 ; P3_U4086
g2266 and P3_U7237 P3_U4316 P3_U7238 ; P3_U4087
g2267 and P3_U4089 P3_U7241 ; P3_U4088
g2268 and P3_U7244 P3_U7243 ; P3_U4089
g2269 and P3_U7245 P3_U4316 P3_U7246 ; P3_U4090
g2270 and P3_U4092 P3_U7249 ; P3_U4091
g2271 and P3_U7252 P3_U7251 ; P3_U4092
g2272 and P3_U7253 P3_U4316 P3_U7254 ; P3_U4093
g2273 and P3_U4095 P3_U7257 ; P3_U4094
g2274 and P3_U7260 P3_U7259 ; P3_U4095
g2275 and P3_U7261 P3_U4316 P3_U7262 ; P3_U4096
g2276 and P3_U4098 P3_U7265 ; P3_U4097
g2277 and P3_U7268 P3_U7267 ; P3_U4098
g2278 and P3_U7270 P3_U7269 ; P3_U4099
g2279 and P3_U4101 P3_U7273 ; P3_U4100
g2280 and P3_U7276 P3_U7275 ; P3_U4101
g2281 and P3_U7278 P3_U7277 ; P3_U4102
g2282 and P3_U4104 P3_U7281 ; P3_U4103
g2283 and P3_U7284 P3_U7283 ; P3_U4104
g2284 and P3_U7286 P3_U7285 ; P3_U4105
g2285 and P3_U4107 P3_U7289 ; P3_U4106
g2286 and P3_U7292 P3_U7291 ; P3_U4107
g2287 and P3_U7294 P3_U7293 ; P3_U4108
g2288 and P3_U4110 P3_U7297 ; P3_U4109
g2289 and P3_U7300 P3_U7299 ; P3_U4110
g2290 and P3_U7302 P3_U7301 ; P3_U4111
g2291 and P3_U4113 P3_U7305 ; P3_U4112
g2292 and P3_U7308 P3_U7307 ; P3_U4113
g2293 and P3_U7310 P3_U7309 ; P3_U4114
g2294 and P3_U4116 P3_U7313 ; P3_U4115
g2295 and P3_U7316 P3_U7315 ; P3_U4116
g2296 and P3_U7318 P3_U7317 ; P3_U4117
g2297 and P3_U4119 P3_U7321 ; P3_U4118
g2298 and P3_U7324 P3_U7323 ; P3_U4119
g2299 and P3_U7326 P3_U7325 ; P3_U4120
g2300 and P3_U4122 P3_U7329 ; P3_U4121
g2301 and P3_U7332 P3_U7331 ; P3_U4122
g2302 and P3_U7334 P3_U7333 ; P3_U4123
g2303 and P3_U4125 P3_U7337 ; P3_U4124
g2304 and P3_U7340 P3_U7339 ; P3_U4125
g2305 and P3_U7342 P3_U7341 ; P3_U4126
g2306 and P3_U4128 P3_U7345 ; P3_U4127
g2307 and P3_U7348 P3_U7347 ; P3_U4128
g2308 and P3_U7350 P3_U7349 ; P3_U4129
g2309 and P3_U4131 P3_U7353 ; P3_U4130
g2310 and P3_U7356 P3_U7355 ; P3_U4131
g2311 and P3_U7364 P3_U7365 ; P3_U4132
g2312 and P3_U4132 P3_U7361 ; P3_U4133
g2313 and P3_U7362 P3_U3259 ; P3_U4134
g2314 nor P3_SUB_320_U51 P3_U7363 ; P3_U4135
g2315 nor P3_DATAWIDTH_REG_2__SCAN_IN P3_DATAWIDTH_REG_3__SCAN_IN P3_DATAWIDTH_REG_4__SCAN_IN P3_DATAWIDTH_REG_5__SCAN_IN ; P3_U4136
g2316 nor P3_DATAWIDTH_REG_6__SCAN_IN P3_DATAWIDTH_REG_7__SCAN_IN P3_DATAWIDTH_REG_8__SCAN_IN P3_DATAWIDTH_REG_9__SCAN_IN ; P3_U4137
g2317 and P3_U4137 P3_U4136 ; P3_U4138
g2318 nor P3_DATAWIDTH_REG_10__SCAN_IN P3_DATAWIDTH_REG_11__SCAN_IN P3_DATAWIDTH_REG_12__SCAN_IN P3_DATAWIDTH_REG_13__SCAN_IN ; P3_U4139
g2319 nor P3_DATAWIDTH_REG_14__SCAN_IN P3_DATAWIDTH_REG_15__SCAN_IN P3_DATAWIDTH_REG_16__SCAN_IN P3_DATAWIDTH_REG_17__SCAN_IN ; P3_U4140
g2320 and P3_U4140 P3_U4139 ; P3_U4141
g2321 nor P3_DATAWIDTH_REG_18__SCAN_IN P3_DATAWIDTH_REG_19__SCAN_IN P3_DATAWIDTH_REG_20__SCAN_IN P3_DATAWIDTH_REG_21__SCAN_IN ; P3_U4142
g2322 nor P3_DATAWIDTH_REG_22__SCAN_IN P3_DATAWIDTH_REG_23__SCAN_IN P3_DATAWIDTH_REG_24__SCAN_IN P3_DATAWIDTH_REG_25__SCAN_IN ; P3_U4143
g2323 and P3_U4143 P3_U4142 ; P3_U4144
g2324 nor P3_DATAWIDTH_REG_26__SCAN_IN P3_DATAWIDTH_REG_27__SCAN_IN ; P3_U4145
g2325 nor P3_DATAWIDTH_REG_28__SCAN_IN P3_DATAWIDTH_REG_29__SCAN_IN ; P3_U4146
g2326 nor P3_DATAWIDTH_REG_30__SCAN_IN P3_DATAWIDTH_REG_31__SCAN_IN ; P3_U4147
g2327 and P3_U4147 P3_U7366 P3_U4146 P3_U4145 ; P3_U4148
g2328 nor P3_DATAWIDTH_REG_0__SCAN_IN P3_DATAWIDTH_REG_1__SCAN_IN P3_REIP_REG_0__SCAN_IN ; P3_U4149
g2329 and P3_U7375 P3_U2630 ; P3_U4150
g2330 and P3_U7373 P3_U3135 ; P3_U4151
g2331 and P3_U7390 P3_U7389 P3_U7388 P3_U7387 ; P3_U4152
g2332 and P3_U7394 P3_U7393 P3_U7392 P3_U7391 ; P3_U4153
g2333 and P3_U7398 P3_U7397 P3_U7396 P3_U7395 ; P3_U4154
g2334 and P3_U7402 P3_U7401 P3_U7400 P3_U7399 ; P3_U4155
g2335 and P3_U7406 P3_U7405 P3_U7404 P3_U7403 ; P3_U4156
g2336 and P3_U7410 P3_U7409 P3_U7408 P3_U7407 ; P3_U4157
g2337 and P3_U7414 P3_U7413 P3_U7412 P3_U7411 ; P3_U4158
g2338 and P3_U7418 P3_U7417 P3_U7416 P3_U7415 ; P3_U4159
g2339 and P3_U7422 P3_U7421 P3_U7420 P3_U7419 ; P3_U4160
g2340 and P3_U7426 P3_U7425 P3_U7424 P3_U7423 ; P3_U4161
g2341 and P3_U7430 P3_U7429 P3_U7428 P3_U7427 ; P3_U4162
g2342 and P3_U7434 P3_U7433 P3_U7432 P3_U7431 ; P3_U4163
g2343 and P3_U7438 P3_U7437 P3_U7436 P3_U7435 ; P3_U4164
g2344 and P3_U7442 P3_U7441 P3_U7440 P3_U7439 ; P3_U4165
g2345 and P3_U7446 P3_U7445 P3_U7444 P3_U7443 ; P3_U4166
g2346 and P3_U7450 P3_U7449 P3_U7448 P3_U7447 ; P3_U4167
g2347 and P3_U7454 P3_U7453 P3_U7452 P3_U7451 ; P3_U4168
g2348 and P3_U7458 P3_U7457 P3_U7456 P3_U7455 ; P3_U4169
g2349 and P3_U7462 P3_U7461 P3_U7460 P3_U7459 ; P3_U4170
g2350 and P3_U7466 P3_U7465 P3_U7464 P3_U7463 ; P3_U4171
g2351 and P3_U7470 P3_U7469 P3_U7468 P3_U7467 ; P3_U4172
g2352 and P3_U7474 P3_U7473 P3_U7472 P3_U7471 ; P3_U4173
g2353 and P3_U7478 P3_U7477 P3_U7476 P3_U7475 ; P3_U4174
g2354 and P3_U7482 P3_U7481 P3_U7480 P3_U7479 ; P3_U4175
g2355 and P3_U7486 P3_U7485 P3_U7484 P3_U7483 ; P3_U4176
g2356 and P3_U7490 P3_U7489 P3_U7488 P3_U7487 ; P3_U4177
g2357 and P3_U7494 P3_U7493 P3_U7492 P3_U7491 ; P3_U4178
g2358 and P3_U7498 P3_U7497 P3_U7496 P3_U7495 ; P3_U4179
g2359 and P3_U7502 P3_U7501 P3_U7500 P3_U7499 ; P3_U4180
g2360 and P3_U7506 P3_U7505 P3_U7504 P3_U7503 ; P3_U4181
g2361 and P3_U7510 P3_U7509 P3_U7508 P3_U7507 ; P3_U4182
g2362 and P3_U7514 P3_U7513 P3_U7512 P3_U7511 ; P3_U4183
g2363 and P3_U7520 P3_U7519 P3_U7518 P3_U7517 ; P3_U4184
g2364 and P3_U7524 P3_U7523 P3_U7522 P3_U7521 ; P3_U4185
g2365 and P3_U7528 P3_U7527 P3_U7526 P3_U7525 ; P3_U4186
g2366 and P3_U7532 P3_U7531 P3_U7530 P3_U7529 ; P3_U4187
g2367 and P3_U7536 P3_U7535 P3_U7534 P3_U7533 ; P3_U4188
g2368 and P3_U7540 P3_U7539 P3_U7538 P3_U7537 ; P3_U4189
g2369 and P3_U7544 P3_U7543 P3_U7542 P3_U7541 ; P3_U4190
g2370 and P3_U7548 P3_U7547 P3_U7546 P3_U7545 ; P3_U4191
g2371 and P3_U7552 P3_U7551 P3_U7550 P3_U7549 ; P3_U4192
g2372 and P3_U7556 P3_U7555 P3_U7554 P3_U7553 ; P3_U4193
g2373 and P3_U7560 P3_U7559 P3_U7558 P3_U7557 ; P3_U4194
g2374 and P3_U7564 P3_U7563 P3_U7562 P3_U7561 ; P3_U4195
g2375 and P3_U7568 P3_U7567 P3_U7566 P3_U7565 ; P3_U4196
g2376 and P3_U7572 P3_U7571 P3_U7570 P3_U7569 ; P3_U4197
g2377 and P3_U7576 P3_U7575 P3_U7574 P3_U7573 ; P3_U4198
g2378 and P3_U7580 P3_U7579 P3_U7578 P3_U7577 ; P3_U4199
g2379 and P3_U7584 P3_U7583 P3_U7582 P3_U7581 ; P3_U4200
g2380 and P3_U7588 P3_U7587 P3_U7586 P3_U7585 ; P3_U4201
g2381 and P3_U7592 P3_U7591 P3_U7590 P3_U7589 ; P3_U4202
g2382 and P3_U7596 P3_U7595 P3_U7594 P3_U7593 ; P3_U4203
g2383 and P3_U7600 P3_U7599 P3_U7598 P3_U7597 ; P3_U4204
g2384 and P3_U7604 P3_U7603 P3_U7602 P3_U7601 ; P3_U4205
g2385 and P3_U7608 P3_U7607 P3_U7606 P3_U7605 ; P3_U4206
g2386 and P3_U7612 P3_U7611 P3_U7610 P3_U7609 ; P3_U4207
g2387 and P3_U7616 P3_U7615 P3_U7614 P3_U7613 ; P3_U4208
g2388 and P3_U7620 P3_U7619 P3_U7618 P3_U7617 ; P3_U4209
g2389 and P3_U7624 P3_U7623 P3_U7622 P3_U7621 ; P3_U4210
g2390 and P3_U7628 P3_U7627 P3_U7626 P3_U7625 ; P3_U4211
g2391 and P3_U7632 P3_U7631 P3_U7630 P3_U7629 ; P3_U4212
g2392 and P3_U7636 P3_U7635 P3_U7634 P3_U7633 ; P3_U4213
g2393 and P3_U7640 P3_U7639 P3_U7638 P3_U7637 ; P3_U4214
g2394 and P3_U7644 P3_U7643 P3_U7642 P3_U7641 ; P3_U4215
g2395 and P3_U7649 P3_U7648 P3_U7647 P3_U7646 ; P3_U4216
g2396 and P3_U7653 P3_U7652 P3_U7651 P3_U7650 ; P3_U4217
g2397 and P3_U7657 P3_U7656 P3_U7655 P3_U7654 ; P3_U4218
g2398 and P3_U7661 P3_U7660 P3_U7659 P3_U7658 ; P3_U4219
g2399 and P3_U7665 P3_U7664 P3_U7663 P3_U7662 ; P3_U4220
g2400 and P3_U7669 P3_U7668 P3_U7667 P3_U7666 ; P3_U4221
g2401 and P3_U7673 P3_U7672 P3_U7671 P3_U7670 ; P3_U4222
g2402 and P3_U7677 P3_U7676 P3_U7675 P3_U7674 ; P3_U4223
g2403 and P3_U7681 P3_U7680 P3_U7679 P3_U7678 ; P3_U4224
g2404 and P3_U7685 P3_U7684 P3_U7683 P3_U7682 ; P3_U4225
g2405 and P3_U7689 P3_U7688 P3_U7687 P3_U7686 ; P3_U4226
g2406 and P3_U7693 P3_U7692 P3_U7691 P3_U7690 ; P3_U4227
g2407 and P3_U7697 P3_U7696 P3_U7695 P3_U7694 ; P3_U4228
g2408 and P3_U7701 P3_U7700 P3_U7699 P3_U7698 ; P3_U4229
g2409 and P3_U7705 P3_U7704 P3_U7703 P3_U7702 ; P3_U4230
g2410 and P3_U7709 P3_U7708 P3_U7707 P3_U7706 ; P3_U4231
g2411 and P3_U7713 P3_U7712 P3_U7711 P3_U7710 ; P3_U4232
g2412 and P3_U7717 P3_U7716 P3_U7715 P3_U7714 ; P3_U4233
g2413 and P3_U7721 P3_U7720 P3_U7719 P3_U7718 ; P3_U4234
g2414 and P3_U7725 P3_U7724 P3_U7723 P3_U7722 ; P3_U4235
g2415 and P3_U7729 P3_U7728 P3_U7727 P3_U7726 ; P3_U4236
g2416 and P3_U7733 P3_U7732 P3_U7731 P3_U7730 ; P3_U4237
g2417 and P3_U7737 P3_U7736 P3_U7735 P3_U7734 ; P3_U4238
g2418 and P3_U7741 P3_U7740 P3_U7739 P3_U7738 ; P3_U4239
g2419 and P3_U7745 P3_U7744 P3_U7743 P3_U7742 ; P3_U4240
g2420 and P3_U7749 P3_U7748 P3_U7747 P3_U7746 ; P3_U4241
g2421 and P3_U7753 P3_U7752 P3_U7751 P3_U7750 ; P3_U4242
g2422 and P3_U7757 P3_U7756 P3_U7755 P3_U7754 ; P3_U4243
g2423 and P3_U7761 P3_U7760 P3_U7759 P3_U7758 ; P3_U4244
g2424 and P3_U7765 P3_U7764 P3_U7763 P3_U7762 ; P3_U4245
g2425 and P3_U7769 P3_U7768 P3_U7767 P3_U7766 ; P3_U4246
g2426 and P3_U7773 P3_U7772 P3_U7771 P3_U7770 ; P3_U4247
g2427 and P3_U7779 P3_U7778 P3_U7777 P3_U7776 ; P3_U4248
g2428 and P3_U7783 P3_U7782 P3_U7781 P3_U7780 ; P3_U4249
g2429 and P3_U7787 P3_U7786 P3_U7785 P3_U7784 ; P3_U4250
g2430 and P3_U7791 P3_U7790 P3_U7789 P3_U7788 ; P3_U4251
g2431 and P3_U7795 P3_U7794 P3_U7793 P3_U7792 ; P3_U4252
g2432 and P3_U7799 P3_U7798 P3_U7797 P3_U7796 ; P3_U4253
g2433 and P3_U7803 P3_U7802 P3_U7801 P3_U7800 ; P3_U4254
g2434 and P3_U7807 P3_U7806 P3_U7805 P3_U7804 ; P3_U4255
g2435 and P3_U7811 P3_U7810 P3_U7809 P3_U7808 ; P3_U4256
g2436 and P3_U7815 P3_U7814 P3_U7813 P3_U7812 ; P3_U4257
g2437 and P3_U7819 P3_U7818 P3_U7817 P3_U7816 ; P3_U4258
g2438 and P3_U7823 P3_U7822 P3_U7821 P3_U7820 ; P3_U4259
g2439 and P3_U7827 P3_U7826 P3_U7825 P3_U7824 ; P3_U4260
g2440 and P3_U7831 P3_U7830 P3_U7829 P3_U7828 ; P3_U4261
g2441 and P3_U7835 P3_U7834 P3_U7833 P3_U7832 ; P3_U4262
g2442 and P3_U7839 P3_U7838 P3_U7837 P3_U7836 ; P3_U4263
g2443 and P3_U7843 P3_U7842 P3_U7841 P3_U7840 ; P3_U4264
g2444 and P3_U7847 P3_U7846 P3_U7845 P3_U7844 ; P3_U4265
g2445 and P3_U7851 P3_U7850 P3_U7849 P3_U7848 ; P3_U4266
g2446 and P3_U7855 P3_U7854 P3_U7853 P3_U7852 ; P3_U4267
g2447 and P3_U7859 P3_U7858 P3_U7857 P3_U7856 ; P3_U4268
g2448 and P3_U7863 P3_U7862 P3_U7861 P3_U7860 ; P3_U4269
g2449 and P3_U7867 P3_U7866 P3_U7865 P3_U7864 ; P3_U4270
g2450 and P3_U7871 P3_U7870 P3_U7869 P3_U7868 ; P3_U4271
g2451 and P3_U7875 P3_U7874 P3_U7873 P3_U7872 ; P3_U4272
g2452 and P3_U7879 P3_U7878 P3_U7877 P3_U7876 ; P3_U4273
g2453 and P3_U7883 P3_U7882 P3_U7881 P3_U7880 ; P3_U4274
g2454 and P3_U7887 P3_U7886 P3_U7885 P3_U7884 ; P3_U4275
g2455 and P3_U7891 P3_U7890 P3_U7889 P3_U7888 ; P3_U4276
g2456 and P3_U7895 P3_U7894 P3_U7893 P3_U7892 ; P3_U4277
g2457 and P3_U7899 P3_U7898 P3_U7897 P3_U7896 ; P3_U4278
g2458 and P3_U7903 P3_U7902 P3_U7901 P3_U7900 ; P3_U4279
g2459 and P3_U7943 P3_U7942 ; P3_U4280
g2460 nand P3_U3361 P3_U2604 ; P3_U4281
g2461 and P3_U7951 P3_U7950 ; P3_U4282
g2462 nand P3_U3658 P3_U5497 ; P3_U4283
g2463 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_U4284
g2464 nand P3_U2390 P3_U4281 ; P3_U4285
g2465 not BS16 ; P3_U4286
g2466 nand P3_U4151 P3_U4334 ; P3_U4287
g2467 nand P3_U4334 P3_U3239 ; P3_U4288
g2468 nand P3_U3091 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U4289
g2469 nand P3_U2515 P3_U2516 P3_U3657 ; P3_U4290
g2470 not P3_U3267 ; P3_U4291
g2471 nand HOLD P3_U2630 ; P3_U4292
g2472 not P3_U3105 ; P3_U4293
g2473 not P3_U3106 ; P3_U4294
g2474 not P3_U3135 ; P3_U4295
g2475 not P3_U3112 ; P3_U4296
g2476 not P3_U3111 ; P3_U4297
g2477 not P3_U3242 ; P3_U4298
g2478 not P3_U3243 ; P3_U4299
g2479 not P3_U3244 ; P3_U4300
g2480 not P3_U3245 ; P3_U4301
g2481 not P3_U3119 ; P3_U4302
g2482 not P3_U3117 ; P3_U4303
g2483 not P3_U3116 ; P3_U4304
g2484 not P3_U3115 ; P3_U4305
g2485 not P3_U3246 ; P3_U4306
g2486 not P3_U3261 ; P3_U4307
g2487 not P3_U3077 ; P3_U4308
g2488 not P3_U3253 ; P3_U4309
g2489 not P3_U3252 ; P3_U4310
g2490 not P3_U3250 ; P3_U4311
g2491 not P3_U3127 ; P3_U4312
g2492 not P3_LT_563_1260_U6 ; P3_U4313
g2493 not P3_U3217 ; P3_U4314
g2494 nand P3_U4295 P3_U2631 ; P3_U4315
g2495 nand P3_U4347 P3_U3260 ; P3_U4316
g2496 nand P3_U2383 P3_U3105 ; P3_U4317
g2497 not P3_U3247 ; P3_U4318
g2498 not P3_U3259 ; P3_U4319
g2499 not P3_U3080 ; P3_U4320
g2500 not P3_U3078 ; P3_U4321
g2501 not P3_U3136 ; P3_U4322
g2502 not P3_U3114 ; P3_U4323
g2503 not P3_U3118 ; P3_U4324
g2504 not P3_U3219 ; P3_U4325
g2505 not P3_U3181 ; P3_U4326
g2506 nand P3_U4149 P3_U4307 ; P3_U4327
g2507 nand P3_U3365 P3_U4354 ; P3_U4328
g2508 nand P3_U3121 P3_U3090 P3_U2631 P3_STATE2_REG_1__SCAN_IN ; P3_U4329
g2509 nand P3_U3653 P3_U2453 ; P3_U4330
g2510 nand P3_U2458 P3_U4653 ; P3_U4331
g2511 not P3_U3095 ; P3_U4332
g2512 nand P3_U4350 P3_U3113 ; P3_U4333
g2513 nand P3_U2390 P3_U7093 ; P3_U4334
g2514 nand P3_U4452 P3_U3085 ; P3_U4335
g2515 nand P3_U4347 P3_U3121 ; P3_U4336
g2516 nand P3_U2453 P3_U3232 ; P3_U4337
g2517 nand P3_U3090 U209 P3_STATE2_REG_0__SCAN_IN ; P3_U4338
g2518 nand P3_U3654 P3_U4608 ; P3_U4339
g2519 not P3_U3123 ; P3_U4340
g2520 not P3_U3229 ; P3_U4341
g2521 not P3_U3150 ; P3_U4342
g2522 not P3_U3158 ; P3_U4343
g2523 not P3_U3103 ; P3_U4344
g2524 not P3_U3126 ; P3_U4345
g2525 not P3_U3082 ; P3_U4346
g2526 not P3_U3239 ; P3_U4347
g2527 not P3_U3236 ; P3_U4348
g2528 not P3_U3235 ; P3_U4349
g2529 not P3_U3208 ; P3_U4350
g2530 not P3_U3216 ; P3_U4351
g2531 not P3_U3222 ; P3_U4352
g2532 not P3_U3124 ; P3_U4353
g2533 not P3_U3125 ; P3_U4354
g2534 nand P3_U4321 P3_REIP_REG_31__SCAN_IN ; P3_U4355
g2535 nand P3_U4320 P3_REIP_REG_30__SCAN_IN ; P3_U4356
g2536 nand P3_U3077 P3_ADDRESS_REG_29__SCAN_IN ; P3_U4357
g2537 nand P3_U4321 P3_REIP_REG_30__SCAN_IN ; P3_U4358
g2538 nand P3_U4320 P3_REIP_REG_29__SCAN_IN ; P3_U4359
g2539 nand P3_U3077 P3_ADDRESS_REG_28__SCAN_IN ; P3_U4360
g2540 nand P3_U4321 P3_REIP_REG_29__SCAN_IN ; P3_U4361
g2541 nand P3_U4320 P3_REIP_REG_28__SCAN_IN ; P3_U4362
g2542 nand P3_U3077 P3_ADDRESS_REG_27__SCAN_IN ; P3_U4363
g2543 nand P3_U4321 P3_REIP_REG_28__SCAN_IN ; P3_U4364
g2544 nand P3_U4320 P3_REIP_REG_27__SCAN_IN ; P3_U4365
g2545 nand P3_U3077 P3_ADDRESS_REG_26__SCAN_IN ; P3_U4366
g2546 nand P3_U4321 P3_REIP_REG_27__SCAN_IN ; P3_U4367
g2547 nand P3_U4320 P3_REIP_REG_26__SCAN_IN ; P3_U4368
g2548 nand P3_U3077 P3_ADDRESS_REG_25__SCAN_IN ; P3_U4369
g2549 nand P3_U4321 P3_REIP_REG_26__SCAN_IN ; P3_U4370
g2550 nand P3_U4320 P3_REIP_REG_25__SCAN_IN ; P3_U4371
g2551 nand P3_U3077 P3_ADDRESS_REG_24__SCAN_IN ; P3_U4372
g2552 nand P3_U4321 P3_REIP_REG_25__SCAN_IN ; P3_U4373
g2553 nand P3_U4320 P3_REIP_REG_24__SCAN_IN ; P3_U4374
g2554 nand P3_U3077 P3_ADDRESS_REG_23__SCAN_IN ; P3_U4375
g2555 nand P3_U4321 P3_REIP_REG_24__SCAN_IN ; P3_U4376
g2556 nand P3_U4320 P3_REIP_REG_23__SCAN_IN ; P3_U4377
g2557 nand P3_U3077 P3_ADDRESS_REG_22__SCAN_IN ; P3_U4378
g2558 nand P3_U4321 P3_REIP_REG_23__SCAN_IN ; P3_U4379
g2559 nand P3_U4320 P3_REIP_REG_22__SCAN_IN ; P3_U4380
g2560 nand P3_U3077 P3_ADDRESS_REG_21__SCAN_IN ; P3_U4381
g2561 nand P3_U4321 P3_REIP_REG_22__SCAN_IN ; P3_U4382
g2562 nand P3_U4320 P3_REIP_REG_21__SCAN_IN ; P3_U4383
g2563 nand P3_U3077 P3_ADDRESS_REG_20__SCAN_IN ; P3_U4384
g2564 nand P3_U4321 P3_REIP_REG_21__SCAN_IN ; P3_U4385
g2565 nand P3_U4320 P3_REIP_REG_20__SCAN_IN ; P3_U4386
g2566 nand P3_U3077 P3_ADDRESS_REG_19__SCAN_IN ; P3_U4387
g2567 nand P3_U4321 P3_REIP_REG_20__SCAN_IN ; P3_U4388
g2568 nand P3_U4320 P3_REIP_REG_19__SCAN_IN ; P3_U4389
g2569 nand P3_U3077 P3_ADDRESS_REG_18__SCAN_IN ; P3_U4390
g2570 nand P3_U4321 P3_REIP_REG_19__SCAN_IN ; P3_U4391
g2571 nand P3_U4320 P3_REIP_REG_18__SCAN_IN ; P3_U4392
g2572 nand P3_U3077 P3_ADDRESS_REG_17__SCAN_IN ; P3_U4393
g2573 nand P3_U4321 P3_REIP_REG_18__SCAN_IN ; P3_U4394
g2574 nand P3_U4320 P3_REIP_REG_17__SCAN_IN ; P3_U4395
g2575 nand P3_U3077 P3_ADDRESS_REG_16__SCAN_IN ; P3_U4396
g2576 nand P3_U4321 P3_REIP_REG_17__SCAN_IN ; P3_U4397
g2577 nand P3_U4320 P3_REIP_REG_16__SCAN_IN ; P3_U4398
g2578 nand P3_U3077 P3_ADDRESS_REG_15__SCAN_IN ; P3_U4399
g2579 nand P3_U4321 P3_REIP_REG_16__SCAN_IN ; P3_U4400
g2580 nand P3_U4320 P3_REIP_REG_15__SCAN_IN ; P3_U4401
g2581 nand P3_U3077 P3_ADDRESS_REG_14__SCAN_IN ; P3_U4402
g2582 nand P3_U4321 P3_REIP_REG_15__SCAN_IN ; P3_U4403
g2583 nand P3_U4320 P3_REIP_REG_14__SCAN_IN ; P3_U4404
g2584 nand P3_U3077 P3_ADDRESS_REG_13__SCAN_IN ; P3_U4405
g2585 nand P3_U4321 P3_REIP_REG_14__SCAN_IN ; P3_U4406
g2586 nand P3_U4320 P3_REIP_REG_13__SCAN_IN ; P3_U4407
g2587 nand P3_U3077 P3_ADDRESS_REG_12__SCAN_IN ; P3_U4408
g2588 nand P3_U4321 P3_REIP_REG_13__SCAN_IN ; P3_U4409
g2589 nand P3_U4320 P3_REIP_REG_12__SCAN_IN ; P3_U4410
g2590 nand P3_U3077 P3_ADDRESS_REG_11__SCAN_IN ; P3_U4411
g2591 nand P3_U4321 P3_REIP_REG_12__SCAN_IN ; P3_U4412
g2592 nand P3_U4320 P3_REIP_REG_11__SCAN_IN ; P3_U4413
g2593 nand P3_U3077 P3_ADDRESS_REG_10__SCAN_IN ; P3_U4414
g2594 nand P3_U4321 P3_REIP_REG_11__SCAN_IN ; P3_U4415
g2595 nand P3_U4320 P3_REIP_REG_10__SCAN_IN ; P3_U4416
g2596 nand P3_U3077 P3_ADDRESS_REG_9__SCAN_IN ; P3_U4417
g2597 nand P3_U4321 P3_REIP_REG_10__SCAN_IN ; P3_U4418
g2598 nand P3_U4320 P3_REIP_REG_9__SCAN_IN ; P3_U4419
g2599 nand P3_U3077 P3_ADDRESS_REG_8__SCAN_IN ; P3_U4420
g2600 nand P3_U4321 P3_REIP_REG_9__SCAN_IN ; P3_U4421
g2601 nand P3_U4320 P3_REIP_REG_8__SCAN_IN ; P3_U4422
g2602 nand P3_U3077 P3_ADDRESS_REG_7__SCAN_IN ; P3_U4423
g2603 nand P3_U4321 P3_REIP_REG_8__SCAN_IN ; P3_U4424
g2604 nand P3_U4320 P3_REIP_REG_7__SCAN_IN ; P3_U4425
g2605 nand P3_U3077 P3_ADDRESS_REG_6__SCAN_IN ; P3_U4426
g2606 nand P3_U4321 P3_REIP_REG_7__SCAN_IN ; P3_U4427
g2607 nand P3_U4320 P3_REIP_REG_6__SCAN_IN ; P3_U4428
g2608 nand P3_U3077 P3_ADDRESS_REG_5__SCAN_IN ; P3_U4429
g2609 nand P3_U4321 P3_REIP_REG_6__SCAN_IN ; P3_U4430
g2610 nand P3_U4320 P3_REIP_REG_5__SCAN_IN ; P3_U4431
g2611 nand P3_U3077 P3_ADDRESS_REG_4__SCAN_IN ; P3_U4432
g2612 nand P3_U4321 P3_REIP_REG_5__SCAN_IN ; P3_U4433
g2613 nand P3_U4320 P3_REIP_REG_4__SCAN_IN ; P3_U4434
g2614 nand P3_U3077 P3_ADDRESS_REG_3__SCAN_IN ; P3_U4435
g2615 nand P3_U4321 P3_REIP_REG_4__SCAN_IN ; P3_U4436
g2616 nand P3_U4320 P3_REIP_REG_3__SCAN_IN ; P3_U4437
g2617 nand P3_U3077 P3_ADDRESS_REG_2__SCAN_IN ; P3_U4438
g2618 nand P3_U4321 P3_REIP_REG_3__SCAN_IN ; P3_U4439
g2619 nand P3_U4320 P3_REIP_REG_2__SCAN_IN ; P3_U4440
g2620 nand P3_U3077 P3_ADDRESS_REG_1__SCAN_IN ; P3_U4441
g2621 nand P3_U4321 P3_REIP_REG_2__SCAN_IN ; P3_U4442
g2622 nand P3_U4320 P3_REIP_REG_1__SCAN_IN ; P3_U4443
g2623 nand P3_U3077 P3_ADDRESS_REG_0__SCAN_IN ; P3_U4444
g2624 not P3_U3087 ; P3_U4445
g2625 nand P3_U4445 P3_U2630 ; P3_U4446
g2626 nand NA P3_U4346 ; P3_U4447
g2627 not P3_U3088 ; P3_U4448
g2628 nand P3_U4448 P3_U2630 ; P3_U4449
g2629 or NA P3_STATE_REG_0__SCAN_IN ; P3_U4450
g2630 nand P3_U7912 P3_U4450 P3_U7913 ; P3_U4451
g2631 not P3_U3083 ; P3_U4452
g2632 nand P3_U3088 U209 P3_U4346 ; P3_U4453
g2633 nand HOLD P3_U3075 P3_U4452 ; P3_U4454
g2634 nand P3_U4453 P3_U4454 ; P3_U4455
g2635 nand P3_U3309 P3_U4455 ; P3_U4456
g2636 nand P3_U4451 P3_STATE_REG_2__SCAN_IN ; P3_U4457
g2637 nand P3_U4308 U209 ; P3_U4458
g2638 nand P3_U3312 P3_U7915 ; P3_U4459
g2639 nand P3_U3087 P3_STATE_REG_2__SCAN_IN ; P3_U4460
g2640 nand NA P3_U3085 ; P3_U4461
g2641 nand P3_U4461 P3_U4460 ; P3_U4462
g2642 nand P3_U4462 P3_U3076 ; P3_U4463
g2643 nand P3_U4286 P3_U3083 ; P3_U4464
g2644 nand P3_U3076 P3_STATE_REG_2__SCAN_IN ; P3_U4465
g2645 nand P3_U3082 P3_U4465 ; P3_U4466
g2646 not P3_U3091 ; P3_U4467
g2647 not P3_U3096 ; P3_U4468
g2648 not P3_U3092 ; P3_U4469
g2649 not P3_U3098 ; P3_U4470
g2650 not P3_U3099 ; P3_U4471
g2651 nand P3_U2484 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U4472
g2652 nand P3_U2483 P3_INSTQUEUE_REG_1__0__SCAN_IN ; P3_U4473
g2653 nand P3_U2482 P3_INSTQUEUE_REG_2__0__SCAN_IN ; P3_U4474
g2654 nand P3_U2480 P3_INSTQUEUE_REG_3__0__SCAN_IN ; P3_U4475
g2655 nand P3_U2479 P3_INSTQUEUE_REG_4__0__SCAN_IN ; P3_U4476
g2656 nand P3_U2478 P3_INSTQUEUE_REG_5__0__SCAN_IN ; P3_U4477
g2657 nand P3_U2477 P3_INSTQUEUE_REG_6__0__SCAN_IN ; P3_U4478
g2658 nand P3_U4471 P3_INSTQUEUE_REG_7__0__SCAN_IN ; P3_U4479
g2659 nand P3_U2476 P3_INSTQUEUE_REG_8__0__SCAN_IN ; P3_U4480
g2660 nand P3_U2475 P3_INSTQUEUE_REG_9__0__SCAN_IN ; P3_U4481
g2661 nand P3_U2473 P3_INSTQUEUE_REG_10__0__SCAN_IN ; P3_U4482
g2662 nand P3_U2471 P3_INSTQUEUE_REG_11__0__SCAN_IN ; P3_U4483
g2663 nand P3_U2470 P3_INSTQUEUE_REG_12__0__SCAN_IN ; P3_U4484
g2664 nand P3_U2469 P3_INSTQUEUE_REG_13__0__SCAN_IN ; P3_U4485
g2665 nand P3_U2467 P3_INSTQUEUE_REG_14__0__SCAN_IN ; P3_U4486
g2666 nand P3_U2465 P3_INSTQUEUE_REG_15__0__SCAN_IN ; P3_U4487
g2667 not P3_U3108 ; P3_U4488
g2668 nand P3_U2484 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U4489
g2669 nand P3_U2483 P3_INSTQUEUE_REG_1__1__SCAN_IN ; P3_U4490
g2670 nand P3_U2482 P3_INSTQUEUE_REG_2__1__SCAN_IN ; P3_U4491
g2671 nand P3_U2480 P3_INSTQUEUE_REG_3__1__SCAN_IN ; P3_U4492
g2672 nand P3_U2479 P3_INSTQUEUE_REG_4__1__SCAN_IN ; P3_U4493
g2673 nand P3_U2478 P3_INSTQUEUE_REG_5__1__SCAN_IN ; P3_U4494
g2674 nand P3_U2477 P3_INSTQUEUE_REG_6__1__SCAN_IN ; P3_U4495
g2675 nand P3_U4471 P3_INSTQUEUE_REG_7__1__SCAN_IN ; P3_U4496
g2676 nand P3_U2476 P3_INSTQUEUE_REG_8__1__SCAN_IN ; P3_U4497
g2677 nand P3_U2475 P3_INSTQUEUE_REG_9__1__SCAN_IN ; P3_U4498
g2678 nand P3_U2473 P3_INSTQUEUE_REG_10__1__SCAN_IN ; P3_U4499
g2679 nand P3_U2471 P3_INSTQUEUE_REG_11__1__SCAN_IN ; P3_U4500
g2680 nand P3_U2470 P3_INSTQUEUE_REG_12__1__SCAN_IN ; P3_U4501
g2681 nand P3_U2469 P3_INSTQUEUE_REG_13__1__SCAN_IN ; P3_U4502
g2682 nand P3_U2467 P3_INSTQUEUE_REG_14__1__SCAN_IN ; P3_U4503
g2683 nand P3_U2465 P3_INSTQUEUE_REG_15__1__SCAN_IN ; P3_U4504
g2684 not P3_U3104 ; P3_U4505
g2685 nand P3_U2484 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U4506
g2686 nand P3_U2483 P3_INSTQUEUE_REG_1__4__SCAN_IN ; P3_U4507
g2687 nand P3_U2482 P3_INSTQUEUE_REG_2__4__SCAN_IN ; P3_U4508
g2688 nand P3_U2480 P3_INSTQUEUE_REG_3__4__SCAN_IN ; P3_U4509
g2689 nand P3_U2479 P3_INSTQUEUE_REG_4__4__SCAN_IN ; P3_U4510
g2690 nand P3_U2478 P3_INSTQUEUE_REG_5__4__SCAN_IN ; P3_U4511
g2691 nand P3_U2477 P3_INSTQUEUE_REG_6__4__SCAN_IN ; P3_U4512
g2692 nand P3_U4471 P3_INSTQUEUE_REG_7__4__SCAN_IN ; P3_U4513
g2693 nand P3_U2476 P3_INSTQUEUE_REG_8__4__SCAN_IN ; P3_U4514
g2694 nand P3_U2475 P3_INSTQUEUE_REG_9__4__SCAN_IN ; P3_U4515
g2695 nand P3_U2473 P3_INSTQUEUE_REG_10__4__SCAN_IN ; P3_U4516
g2696 nand P3_U2471 P3_INSTQUEUE_REG_11__4__SCAN_IN ; P3_U4517
g2697 nand P3_U2470 P3_INSTQUEUE_REG_12__4__SCAN_IN ; P3_U4518
g2698 nand P3_U2469 P3_INSTQUEUE_REG_13__4__SCAN_IN ; P3_U4519
g2699 nand P3_U2467 P3_INSTQUEUE_REG_14__4__SCAN_IN ; P3_U4520
g2700 nand P3_U2465 P3_INSTQUEUE_REG_15__4__SCAN_IN ; P3_U4521
g2701 not P3_U3102 ; P3_U4522
g2702 nand P3_U2484 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U4523
g2703 nand P3_U2483 P3_INSTQUEUE_REG_1__2__SCAN_IN ; P3_U4524
g2704 nand P3_U2482 P3_INSTQUEUE_REG_2__2__SCAN_IN ; P3_U4525
g2705 nand P3_U2480 P3_INSTQUEUE_REG_3__2__SCAN_IN ; P3_U4526
g2706 nand P3_U2479 P3_INSTQUEUE_REG_4__2__SCAN_IN ; P3_U4527
g2707 nand P3_U2478 P3_INSTQUEUE_REG_5__2__SCAN_IN ; P3_U4528
g2708 nand P3_U2477 P3_INSTQUEUE_REG_6__2__SCAN_IN ; P3_U4529
g2709 nand P3_U4471 P3_INSTQUEUE_REG_7__2__SCAN_IN ; P3_U4530
g2710 nand P3_U2476 P3_INSTQUEUE_REG_8__2__SCAN_IN ; P3_U4531
g2711 nand P3_U2475 P3_INSTQUEUE_REG_9__2__SCAN_IN ; P3_U4532
g2712 nand P3_U2473 P3_INSTQUEUE_REG_10__2__SCAN_IN ; P3_U4533
g2713 nand P3_U2471 P3_INSTQUEUE_REG_11__2__SCAN_IN ; P3_U4534
g2714 nand P3_U2470 P3_INSTQUEUE_REG_12__2__SCAN_IN ; P3_U4535
g2715 nand P3_U2469 P3_INSTQUEUE_REG_13__2__SCAN_IN ; P3_U4536
g2716 nand P3_U2467 P3_INSTQUEUE_REG_14__2__SCAN_IN ; P3_U4537
g2717 nand P3_U2465 P3_INSTQUEUE_REG_15__2__SCAN_IN ; P3_U4538
g2718 not P3_U3101 ; P3_U4539
g2719 nand P3_U2484 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U4540
g2720 nand P3_U2483 P3_INSTQUEUE_REG_1__3__SCAN_IN ; P3_U4541
g2721 nand P3_U2482 P3_INSTQUEUE_REG_2__3__SCAN_IN ; P3_U4542
g2722 nand P3_U2480 P3_INSTQUEUE_REG_3__3__SCAN_IN ; P3_U4543
g2723 nand P3_U2479 P3_INSTQUEUE_REG_4__3__SCAN_IN ; P3_U4544
g2724 nand P3_U2478 P3_INSTQUEUE_REG_5__3__SCAN_IN ; P3_U4545
g2725 nand P3_U2477 P3_INSTQUEUE_REG_6__3__SCAN_IN ; P3_U4546
g2726 nand P3_U4471 P3_INSTQUEUE_REG_7__3__SCAN_IN ; P3_U4547
g2727 nand P3_U2476 P3_INSTQUEUE_REG_8__3__SCAN_IN ; P3_U4548
g2728 nand P3_U2475 P3_INSTQUEUE_REG_9__3__SCAN_IN ; P3_U4549
g2729 nand P3_U2473 P3_INSTQUEUE_REG_10__3__SCAN_IN ; P3_U4550
g2730 nand P3_U2471 P3_INSTQUEUE_REG_11__3__SCAN_IN ; P3_U4551
g2731 nand P3_U2470 P3_INSTQUEUE_REG_12__3__SCAN_IN ; P3_U4552
g2732 nand P3_U2469 P3_INSTQUEUE_REG_13__3__SCAN_IN ; P3_U4553
g2733 nand P3_U2467 P3_INSTQUEUE_REG_14__3__SCAN_IN ; P3_U4554
g2734 nand P3_U2465 P3_INSTQUEUE_REG_15__3__SCAN_IN ; P3_U4555
g2735 not P3_U3107 ; P3_U4556
g2736 nand P3_U2484 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U4557
g2737 nand P3_U2483 P3_INSTQUEUE_REG_1__7__SCAN_IN ; P3_U4558
g2738 nand P3_U2482 P3_INSTQUEUE_REG_2__7__SCAN_IN ; P3_U4559
g2739 nand P3_U2480 P3_INSTQUEUE_REG_3__7__SCAN_IN ; P3_U4560
g2740 nand P3_U2479 P3_INSTQUEUE_REG_4__7__SCAN_IN ; P3_U4561
g2741 nand P3_U2478 P3_INSTQUEUE_REG_5__7__SCAN_IN ; P3_U4562
g2742 nand P3_U2477 P3_INSTQUEUE_REG_6__7__SCAN_IN ; P3_U4563
g2743 nand P3_U4471 P3_INSTQUEUE_REG_7__7__SCAN_IN ; P3_U4564
g2744 nand P3_U2476 P3_INSTQUEUE_REG_8__7__SCAN_IN ; P3_U4565
g2745 nand P3_U2475 P3_INSTQUEUE_REG_9__7__SCAN_IN ; P3_U4566
g2746 nand P3_U2473 P3_INSTQUEUE_REG_10__7__SCAN_IN ; P3_U4567
g2747 nand P3_U2471 P3_INSTQUEUE_REG_11__7__SCAN_IN ; P3_U4568
g2748 nand P3_U2470 P3_INSTQUEUE_REG_12__7__SCAN_IN ; P3_U4569
g2749 nand P3_U2469 P3_INSTQUEUE_REG_13__7__SCAN_IN ; P3_U4570
g2750 nand P3_U2467 P3_INSTQUEUE_REG_14__7__SCAN_IN ; P3_U4571
g2751 nand P3_U2465 P3_INSTQUEUE_REG_15__7__SCAN_IN ; P3_U4572
g2752 not P3_U3218 ; P3_U4573
g2753 nand P3_U2484 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U4574
g2754 nand P3_U2483 P3_INSTQUEUE_REG_1__5__SCAN_IN ; P3_U4575
g2755 nand P3_U2482 P3_INSTQUEUE_REG_2__5__SCAN_IN ; P3_U4576
g2756 nand P3_U2480 P3_INSTQUEUE_REG_3__5__SCAN_IN ; P3_U4577
g2757 nand P3_U2479 P3_INSTQUEUE_REG_4__5__SCAN_IN ; P3_U4578
g2758 nand P3_U2478 P3_INSTQUEUE_REG_5__5__SCAN_IN ; P3_U4579
g2759 nand P3_U2477 P3_INSTQUEUE_REG_6__5__SCAN_IN ; P3_U4580
g2760 nand P3_U4471 P3_INSTQUEUE_REG_7__5__SCAN_IN ; P3_U4581
g2761 nand P3_U2476 P3_INSTQUEUE_REG_8__5__SCAN_IN ; P3_U4582
g2762 nand P3_U2475 P3_INSTQUEUE_REG_9__5__SCAN_IN ; P3_U4583
g2763 nand P3_U2473 P3_INSTQUEUE_REG_10__5__SCAN_IN ; P3_U4584
g2764 nand P3_U2471 P3_INSTQUEUE_REG_11__5__SCAN_IN ; P3_U4585
g2765 nand P3_U2470 P3_INSTQUEUE_REG_12__5__SCAN_IN ; P3_U4586
g2766 nand P3_U2469 P3_INSTQUEUE_REG_13__5__SCAN_IN ; P3_U4587
g2767 nand P3_U2467 P3_INSTQUEUE_REG_14__5__SCAN_IN ; P3_U4588
g2768 nand P3_U2465 P3_INSTQUEUE_REG_15__5__SCAN_IN ; P3_U4589
g2769 not P3_U3110 ; P3_U4590
g2770 nand P3_U2484 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U4591
g2771 nand P3_U2483 P3_INSTQUEUE_REG_1__6__SCAN_IN ; P3_U4592
g2772 nand P3_U2482 P3_INSTQUEUE_REG_2__6__SCAN_IN ; P3_U4593
g2773 nand P3_U2480 P3_INSTQUEUE_REG_3__6__SCAN_IN ; P3_U4594
g2774 nand P3_U2479 P3_INSTQUEUE_REG_4__6__SCAN_IN ; P3_U4595
g2775 nand P3_U2478 P3_INSTQUEUE_REG_5__6__SCAN_IN ; P3_U4596
g2776 nand P3_U2477 P3_INSTQUEUE_REG_6__6__SCAN_IN ; P3_U4597
g2777 nand P3_U4471 P3_INSTQUEUE_REG_7__6__SCAN_IN ; P3_U4598
g2778 nand P3_U2476 P3_INSTQUEUE_REG_8__6__SCAN_IN ; P3_U4599
g2779 nand P3_U2475 P3_INSTQUEUE_REG_9__6__SCAN_IN ; P3_U4600
g2780 nand P3_U2473 P3_INSTQUEUE_REG_10__6__SCAN_IN ; P3_U4601
g2781 nand P3_U2471 P3_INSTQUEUE_REG_11__6__SCAN_IN ; P3_U4602
g2782 nand P3_U2470 P3_INSTQUEUE_REG_12__6__SCAN_IN ; P3_U4603
g2783 nand P3_U2469 P3_INSTQUEUE_REG_13__6__SCAN_IN ; P3_U4604
g2784 nand P3_U2467 P3_INSTQUEUE_REG_14__6__SCAN_IN ; P3_U4605
g2785 nand P3_U2465 P3_INSTQUEUE_REG_15__6__SCAN_IN ; P3_U4606
g2786 not P3_U3074 ; P3_U4607
g2787 not P3_U3113 ; P3_U4608
g2788 nand P3_U2361 P3_U3238 ; P3_U4609
g2789 nand P3_U2360 P3_U3237 ; P3_U4610
g2790 nand P3_U2357 P3_U3212 ; P3_U4611
g2791 nand P3_U4305 P3_U3215 ; P3_U4612
g2792 nand P3_U4304 P3_U3210 ; P3_U4613
g2793 nand P3_U4303 P3_U3213 ; P3_U4614
g2794 nand P3_U2356 P3_U3211 ; P3_U4615
g2795 nand P3_U4302 P3_U3214 ; P3_U4616
g2796 nand P3_U3358 P3_U3357 ; P3_U4617
g2797 nand P3_U2463 P3_U4522 P3_U3360 P3_U7945 P3_U7944 ; P3_U4618
g2798 not P3_U3109 ; P3_U4619
g2799 nand P3_U4280 P3_U4619 ; P3_U4620
g2800 nand P3_U3359 P3_U7916 ; P3_U4621
g2801 not P3_U4281 ; P3_U4622
g2802 not P3_U3262 ; P3_U4623
g2803 or P3_FLUSH_REG_SCAN_IN P3_MORE_REG_SCAN_IN ; P3_U4624
g2804 not P3_U3120 ; P3_U4625
g2805 nand P3_U3353 P3_U4303 ; P3_U4626
g2806 nand P3_U3362 P3_U4625 ; P3_U4627
g2807 nand U209 P3_STATE2_REG_1__SCAN_IN ; P3_U4628
g2808 nand P3_U7953 P3_U7952 P3_STATE2_REG_2__SCAN_IN ; P3_U4629
g2809 not P3_U3122 ; P3_U4630
g2810 nand P3_U7957 P3_U7956 P3_STATE2_REG_1__SCAN_IN ; P3_U4631
g2811 nand P3_U3122 P3_STATE2_REG_2__SCAN_IN ; P3_U4632
g2812 nand P3_U4629 P3_U4338 ; P3_U4633
g2813 nand P3_U3364 P3_U4630 ; P3_U4634
g2814 nand P3_U4633 P3_STATE2_REG_1__SCAN_IN ; P3_U4635
g2815 nand P3_U2390 P3_U4629 ; P3_U4636
g2816 nand P3_U4345 P3_U4354 ; P3_U4637
g2817 nand P3_U4629 P3_U4337 ; P3_U4638
g2818 nand P3_U2390 P3_U3120 ; P3_U4639
g2819 not P3_U3153 ; P3_U4640
g2820 nand P3_U3128 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U4641
g2821 not P3_U3137 ; P3_U4642
g2822 not P3_U3141 ; P3_U4643
g2823 not P3_U3148 ; P3_U4644
g2824 not P3_U3155 ; P3_U4645
g2825 not P3_U3156 ; P3_U4646
g2826 not P3_U3143 ; P3_U4647
g2827 not P3_U3130 ; P3_U4648
g2828 not P3_U3132 ; P3_U4649
g2829 not P3_U3180 ; P3_U4650
g2830 nand P3_U3132 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U4651
g2831 not P3_U3139 ; P3_U4652
g2832 not P3_U3138 ; P3_U4653
g2833 nand P3_U4653 P3_U3269 ; P3_U4654
g2834 nand P3_U4654 P3_U3139 ; P3_U4655
g2835 not P3_U3142 ; P3_U4656
g2836 not P3_U3140 ; P3_U4657
g2837 not P3_U3165 ; P3_U4658
g2838 nand P3_U3140 P3_U3142 ; P3_U4659
g2839 not P3_U3182 ; P3_U4660
g2840 not P3_U3144 ; P3_U4661
g2841 not P3_U3134 ; P3_U4662
g2842 nand P3_U2457 P3_U4653 ; P3_U4663
g2843 not P3_U3146 ; P3_U4664
g2844 nand P3_U3090 P3_STATE2_REG_1__SCAN_IN ; P3_U4665
g2845 nand P3_U3124 P3_U4665 P3_U3126 ; P3_U4666
g2846 nand P3_U4657 P3_U2487 ; P3_U4667
g2847 not P3_U3145 ; P3_U4668
g2848 nand P3_U2489 P3_U3145 ; P3_U4669
g2849 nand P3_U4664 P3_U4669 ; P3_U4670
g2850 nand P3_U3134 P3_STATE2_REG_3__SCAN_IN ; P3_U4671
g2851 nand P3_U3369 P3_U4670 ; P3_U4672
g2852 nand P3_U4668 P3_U4322 ; P3_U4673
g2853 nand P3_U2489 P3_U4673 ; P3_U4674
g2854 nand P3_U2445 P3_U4662 ; P3_U4675
g2855 nand P3_U2436 P3_U2488 ; P3_U4676
g2856 nand P3_U2435 P3_U4661 ; P3_U4677
g2857 nand P3_U2378 P3_U2420 ; P3_U4678
g2858 nand P3_U4672 P3_INSTQUEUE_REG_15__7__SCAN_IN ; P3_U4679
g2859 nand P3_U2443 P3_U4662 ; P3_U4680
g2860 nand P3_U2434 P3_U2488 ; P3_U4681
g2861 nand P3_U2433 P3_U4661 ; P3_U4682
g2862 nand P3_U2419 P3_U2378 ; P3_U4683
g2863 nand P3_U4672 P3_INSTQUEUE_REG_15__6__SCAN_IN ; P3_U4684
g2864 nand P3_U2442 P3_U4662 ; P3_U4685
g2865 nand P3_U2432 P3_U2488 ; P3_U4686
g2866 nand P3_U2431 P3_U4661 ; P3_U4687
g2867 nand P3_U2418 P3_U2378 ; P3_U4688
g2868 nand P3_U4672 P3_INSTQUEUE_REG_15__5__SCAN_IN ; P3_U4689
g2869 nand P3_U2441 P3_U4662 ; P3_U4690
g2870 nand P3_U2430 P3_U2488 ; P3_U4691
g2871 nand P3_U2429 P3_U4661 ; P3_U4692
g2872 nand P3_U2417 P3_U2378 ; P3_U4693
g2873 nand P3_U4672 P3_INSTQUEUE_REG_15__4__SCAN_IN ; P3_U4694
g2874 nand P3_U2440 P3_U4662 ; P3_U4695
g2875 nand P3_U2428 P3_U2488 ; P3_U4696
g2876 nand P3_U2427 P3_U4661 ; P3_U4697
g2877 nand P3_U2416 P3_U2378 ; P3_U4698
g2878 nand P3_U4672 P3_INSTQUEUE_REG_15__3__SCAN_IN ; P3_U4699
g2879 nand P3_U2439 P3_U4662 ; P3_U4700
g2880 nand P3_U2426 P3_U2488 ; P3_U4701
g2881 nand P3_U2425 P3_U4661 ; P3_U4702
g2882 nand P3_U2415 P3_U2378 ; P3_U4703
g2883 nand P3_U4672 P3_INSTQUEUE_REG_15__2__SCAN_IN ; P3_U4704
g2884 nand P3_U2438 P3_U4662 ; P3_U4705
g2885 nand P3_U2424 P3_U2488 ; P3_U4706
g2886 nand P3_U2423 P3_U4661 ; P3_U4707
g2887 nand P3_U2414 P3_U2378 ; P3_U4708
g2888 nand P3_U4672 P3_INSTQUEUE_REG_15__1__SCAN_IN ; P3_U4709
g2889 nand P3_U2437 P3_U4662 ; P3_U4710
g2890 nand P3_U2422 P3_U2488 ; P3_U4711
g2891 nand P3_U2421 P3_U4661 ; P3_U4712
g2892 nand P3_U2413 P3_U2378 ; P3_U4713
g2893 nand P3_U4672 P3_INSTQUEUE_REG_15__0__SCAN_IN ; P3_U4714
g2894 not P3_U3149 ; P3_U4715
g2895 not P3_U3147 ; P3_U4716
g2896 nand P3_U4342 P3_U2457 ; P3_U4717
g2897 not P3_U3152 ; P3_U4718
g2898 nand P3_U4644 P3_U2487 ; P3_U4719
g2899 not P3_U3151 ; P3_U4720
g2900 nand P3_U2489 P3_U3151 ; P3_U4721
g2901 nand P3_U4718 P3_U4721 ; P3_U4722
g2902 nand P3_U3147 P3_STATE2_REG_3__SCAN_IN ; P3_U4723
g2903 nand P3_U3387 P3_U4722 ; P3_U4724
g2904 nand P3_U4720 P3_U4322 ; P3_U4725
g2905 nand P3_U2489 P3_U4725 ; P3_U4726
g2906 nand P3_U4716 P3_U2445 ; P3_U4727
g2907 nand P3_U2491 P3_U2436 ; P3_U4728
g2908 nand P3_U4715 P3_U2435 ; P3_U4729
g2909 nand P3_U2377 P3_U2420 ; P3_U4730
g2910 nand P3_U4724 P3_INSTQUEUE_REG_14__7__SCAN_IN ; P3_U4731
g2911 nand P3_U4716 P3_U2443 ; P3_U4732
g2912 nand P3_U2491 P3_U2434 ; P3_U4733
g2913 nand P3_U4715 P3_U2433 ; P3_U4734
g2914 nand P3_U2377 P3_U2419 ; P3_U4735
g2915 nand P3_U4724 P3_INSTQUEUE_REG_14__6__SCAN_IN ; P3_U4736
g2916 nand P3_U4716 P3_U2442 ; P3_U4737
g2917 nand P3_U2491 P3_U2432 ; P3_U4738
g2918 nand P3_U4715 P3_U2431 ; P3_U4739
g2919 nand P3_U2377 P3_U2418 ; P3_U4740
g2920 nand P3_U4724 P3_INSTQUEUE_REG_14__5__SCAN_IN ; P3_U4741
g2921 nand P3_U4716 P3_U2441 ; P3_U4742
g2922 nand P3_U2491 P3_U2430 ; P3_U4743
g2923 nand P3_U4715 P3_U2429 ; P3_U4744
g2924 nand P3_U2377 P3_U2417 ; P3_U4745
g2925 nand P3_U4724 P3_INSTQUEUE_REG_14__4__SCAN_IN ; P3_U4746
g2926 nand P3_U4716 P3_U2440 ; P3_U4747
g2927 nand P3_U2491 P3_U2428 ; P3_U4748
g2928 nand P3_U4715 P3_U2427 ; P3_U4749
g2929 nand P3_U2377 P3_U2416 ; P3_U4750
g2930 nand P3_U4724 P3_INSTQUEUE_REG_14__3__SCAN_IN ; P3_U4751
g2931 nand P3_U4716 P3_U2439 ; P3_U4752
g2932 nand P3_U2491 P3_U2426 ; P3_U4753
g2933 nand P3_U4715 P3_U2425 ; P3_U4754
g2934 nand P3_U2377 P3_U2415 ; P3_U4755
g2935 nand P3_U4724 P3_INSTQUEUE_REG_14__2__SCAN_IN ; P3_U4756
g2936 nand P3_U4716 P3_U2438 ; P3_U4757
g2937 nand P3_U2491 P3_U2424 ; P3_U4758
g2938 nand P3_U4715 P3_U2423 ; P3_U4759
g2939 nand P3_U2377 P3_U2414 ; P3_U4760
g2940 nand P3_U4724 P3_INSTQUEUE_REG_14__1__SCAN_IN ; P3_U4761
g2941 nand P3_U4716 P3_U2437 ; P3_U4762
g2942 nand P3_U2491 P3_U2422 ; P3_U4763
g2943 nand P3_U4715 P3_U2421 ; P3_U4764
g2944 nand P3_U2377 P3_U2413 ; P3_U4765
g2945 nand P3_U4724 P3_INSTQUEUE_REG_14__0__SCAN_IN ; P3_U4766
g2946 not P3_U3157 ; P3_U4767
g2947 not P3_U3154 ; P3_U4768
g2948 nand P3_U4343 P3_U2457 ; P3_U4769
g2949 not P3_U3160 ; P3_U4770
g2950 nand P3_U4645 P3_U2487 ; P3_U4771
g2951 not P3_U3159 ; P3_U4772
g2952 nand P3_U2489 P3_U3159 ; P3_U4773
g2953 nand P3_U4770 P3_U4773 ; P3_U4774
g2954 nand P3_U3154 P3_STATE2_REG_3__SCAN_IN ; P3_U4775
g2955 nand P3_U3405 P3_U4774 ; P3_U4776
g2956 nand P3_U4772 P3_U4322 ; P3_U4777
g2957 nand P3_U2489 P3_U4777 ; P3_U4778
g2958 nand P3_U4768 P3_U2445 ; P3_U4779
g2959 nand P3_U2494 P3_U2436 ; P3_U4780
g2960 nand P3_U4767 P3_U2435 ; P3_U4781
g2961 nand P3_U2376 P3_U2420 ; P3_U4782
g2962 nand P3_U4776 P3_INSTQUEUE_REG_13__7__SCAN_IN ; P3_U4783
g2963 nand P3_U4768 P3_U2443 ; P3_U4784
g2964 nand P3_U2494 P3_U2434 ; P3_U4785
g2965 nand P3_U4767 P3_U2433 ; P3_U4786
g2966 nand P3_U2376 P3_U2419 ; P3_U4787
g2967 nand P3_U4776 P3_INSTQUEUE_REG_13__6__SCAN_IN ; P3_U4788
g2968 nand P3_U4768 P3_U2442 ; P3_U4789
g2969 nand P3_U2494 P3_U2432 ; P3_U4790
g2970 nand P3_U4767 P3_U2431 ; P3_U4791
g2971 nand P3_U2376 P3_U2418 ; P3_U4792
g2972 nand P3_U4776 P3_INSTQUEUE_REG_13__5__SCAN_IN ; P3_U4793
g2973 nand P3_U4768 P3_U2441 ; P3_U4794
g2974 nand P3_U2494 P3_U2430 ; P3_U4795
g2975 nand P3_U4767 P3_U2429 ; P3_U4796
g2976 nand P3_U2376 P3_U2417 ; P3_U4797
g2977 nand P3_U4776 P3_INSTQUEUE_REG_13__4__SCAN_IN ; P3_U4798
g2978 nand P3_U4768 P3_U2440 ; P3_U4799
g2979 nand P3_U2494 P3_U2428 ; P3_U4800
g2980 nand P3_U4767 P3_U2427 ; P3_U4801
g2981 nand P3_U2376 P3_U2416 ; P3_U4802
g2982 nand P3_U4776 P3_INSTQUEUE_REG_13__3__SCAN_IN ; P3_U4803
g2983 nand P3_U4768 P3_U2439 ; P3_U4804
g2984 nand P3_U2494 P3_U2426 ; P3_U4805
g2985 nand P3_U4767 P3_U2425 ; P3_U4806
g2986 nand P3_U2376 P3_U2415 ; P3_U4807
g2987 nand P3_U4776 P3_INSTQUEUE_REG_13__2__SCAN_IN ; P3_U4808
g2988 nand P3_U4768 P3_U2438 ; P3_U4809
g2989 nand P3_U2494 P3_U2424 ; P3_U4810
g2990 nand P3_U4767 P3_U2423 ; P3_U4811
g2991 nand P3_U2376 P3_U2414 ; P3_U4812
g2992 nand P3_U4776 P3_INSTQUEUE_REG_13__1__SCAN_IN ; P3_U4813
g2993 nand P3_U4768 P3_U2437 ; P3_U4814
g2994 nand P3_U2494 P3_U2422 ; P3_U4815
g2995 nand P3_U4767 P3_U2421 ; P3_U4816
g2996 nand P3_U2376 P3_U2413 ; P3_U4817
g2997 nand P3_U4776 P3_INSTQUEUE_REG_13__0__SCAN_IN ; P3_U4818
g2998 not P3_U3162 ; P3_U4819
g2999 not P3_U3161 ; P3_U4820
g3000 not P3_U3070 ; P3_U4821
g3001 nand P3_U2496 P3_U2487 ; P3_U4822
g3002 not P3_U3163 ; P3_U4823
g3003 nand P3_U2489 P3_U3163 ; P3_U4824
g3004 nand P3_U4824 P3_U3070 ; P3_U4825
g3005 nand P3_U3161 P3_STATE2_REG_3__SCAN_IN ; P3_U4826
g3006 nand P3_U3423 P3_U4825 ; P3_U4827
g3007 nand P3_U4823 P3_U4322 ; P3_U4828
g3008 nand P3_U2489 P3_U4828 ; P3_U4829
g3009 nand P3_U4820 P3_U2445 ; P3_U4830
g3010 nand P3_U2497 P3_U2436 ; P3_U4831
g3011 nand P3_U4819 P3_U2435 ; P3_U4832
g3012 nand P3_U2375 P3_U2420 ; P3_U4833
g3013 nand P3_U4827 P3_INSTQUEUE_REG_12__7__SCAN_IN ; P3_U4834
g3014 nand P3_U4820 P3_U2443 ; P3_U4835
g3015 nand P3_U2497 P3_U2434 ; P3_U4836
g3016 nand P3_U4819 P3_U2433 ; P3_U4837
g3017 nand P3_U2375 P3_U2419 ; P3_U4838
g3018 nand P3_U4827 P3_INSTQUEUE_REG_12__6__SCAN_IN ; P3_U4839
g3019 nand P3_U4820 P3_U2442 ; P3_U4840
g3020 nand P3_U2497 P3_U2432 ; P3_U4841
g3021 nand P3_U4819 P3_U2431 ; P3_U4842
g3022 nand P3_U2375 P3_U2418 ; P3_U4843
g3023 nand P3_U4827 P3_INSTQUEUE_REG_12__5__SCAN_IN ; P3_U4844
g3024 nand P3_U4820 P3_U2441 ; P3_U4845
g3025 nand P3_U2497 P3_U2430 ; P3_U4846
g3026 nand P3_U4819 P3_U2429 ; P3_U4847
g3027 nand P3_U2375 P3_U2417 ; P3_U4848
g3028 nand P3_U4827 P3_INSTQUEUE_REG_12__4__SCAN_IN ; P3_U4849
g3029 nand P3_U4820 P3_U2440 ; P3_U4850
g3030 nand P3_U2497 P3_U2428 ; P3_U4851
g3031 nand P3_U4819 P3_U2427 ; P3_U4852
g3032 nand P3_U2375 P3_U2416 ; P3_U4853
g3033 nand P3_U4827 P3_INSTQUEUE_REG_12__3__SCAN_IN ; P3_U4854
g3034 nand P3_U4820 P3_U2439 ; P3_U4855
g3035 nand P3_U2497 P3_U2426 ; P3_U4856
g3036 nand P3_U4819 P3_U2425 ; P3_U4857
g3037 nand P3_U2375 P3_U2415 ; P3_U4858
g3038 nand P3_U4827 P3_INSTQUEUE_REG_12__2__SCAN_IN ; P3_U4859
g3039 nand P3_U4820 P3_U2438 ; P3_U4860
g3040 nand P3_U2497 P3_U2424 ; P3_U4861
g3041 nand P3_U4819 P3_U2423 ; P3_U4862
g3042 nand P3_U2375 P3_U2414 ; P3_U4863
g3043 nand P3_U4827 P3_INSTQUEUE_REG_12__1__SCAN_IN ; P3_U4864
g3044 nand P3_U4820 P3_U2437 ; P3_U4865
g3045 nand P3_U2497 P3_U2422 ; P3_U4866
g3046 nand P3_U4819 P3_U2421 ; P3_U4867
g3047 nand P3_U2375 P3_U2413 ; P3_U4868
g3048 nand P3_U4827 P3_INSTQUEUE_REG_12__0__SCAN_IN ; P3_U4869
g3049 not P3_U3166 ; P3_U4870
g3050 not P3_U3164 ; P3_U4871
g3051 nand P3_U2459 P3_U4653 ; P3_U4872
g3052 not P3_U3168 ; P3_U4873
g3053 nand P3_U4658 P3_U4657 ; P3_U4874
g3054 not P3_U3167 ; P3_U4875
g3055 nand P3_U2489 P3_U3167 ; P3_U4876
g3056 nand P3_U4873 P3_U4876 ; P3_U4877
g3057 nand P3_U3164 P3_STATE2_REG_3__SCAN_IN ; P3_U4878
g3058 nand P3_U3440 P3_U4877 ; P3_U4879
g3059 nand P3_U4875 P3_U4322 ; P3_U4880
g3060 nand P3_U2489 P3_U4880 ; P3_U4881
g3061 nand P3_U4871 P3_U2445 ; P3_U4882
g3062 nand P3_U2499 P3_U2436 ; P3_U4883
g3063 nand P3_U4870 P3_U2435 ; P3_U4884
g3064 nand P3_U2374 P3_U2420 ; P3_U4885
g3065 nand P3_U4879 P3_INSTQUEUE_REG_11__7__SCAN_IN ; P3_U4886
g3066 nand P3_U4871 P3_U2443 ; P3_U4887
g3067 nand P3_U2499 P3_U2434 ; P3_U4888
g3068 nand P3_U4870 P3_U2433 ; P3_U4889
g3069 nand P3_U2374 P3_U2419 ; P3_U4890
g3070 nand P3_U4879 P3_INSTQUEUE_REG_11__6__SCAN_IN ; P3_U4891
g3071 nand P3_U4871 P3_U2442 ; P3_U4892
g3072 nand P3_U2499 P3_U2432 ; P3_U4893
g3073 nand P3_U4870 P3_U2431 ; P3_U4894
g3074 nand P3_U2374 P3_U2418 ; P3_U4895
g3075 nand P3_U4879 P3_INSTQUEUE_REG_11__5__SCAN_IN ; P3_U4896
g3076 nand P3_U4871 P3_U2441 ; P3_U4897
g3077 nand P3_U2499 P3_U2430 ; P3_U4898
g3078 nand P3_U4870 P3_U2429 ; P3_U4899
g3079 nand P3_U2374 P3_U2417 ; P3_U4900
g3080 nand P3_U4879 P3_INSTQUEUE_REG_11__4__SCAN_IN ; P3_U4901
g3081 nand P3_U4871 P3_U2440 ; P3_U4902
g3082 nand P3_U2499 P3_U2428 ; P3_U4903
g3083 nand P3_U4870 P3_U2427 ; P3_U4904
g3084 nand P3_U2374 P3_U2416 ; P3_U4905
g3085 nand P3_U4879 P3_INSTQUEUE_REG_11__3__SCAN_IN ; P3_U4906
g3086 nand P3_U4871 P3_U2439 ; P3_U4907
g3087 nand P3_U2499 P3_U2426 ; P3_U4908
g3088 nand P3_U4870 P3_U2425 ; P3_U4909
g3089 nand P3_U2374 P3_U2415 ; P3_U4910
g3090 nand P3_U4879 P3_INSTQUEUE_REG_11__2__SCAN_IN ; P3_U4911
g3091 nand P3_U4871 P3_U2438 ; P3_U4912
g3092 nand P3_U2499 P3_U2424 ; P3_U4913
g3093 nand P3_U4870 P3_U2423 ; P3_U4914
g3094 nand P3_U2374 P3_U2414 ; P3_U4915
g3095 nand P3_U4879 P3_INSTQUEUE_REG_11__1__SCAN_IN ; P3_U4916
g3096 nand P3_U4871 P3_U2437 ; P3_U4917
g3097 nand P3_U2499 P3_U2422 ; P3_U4918
g3098 nand P3_U4870 P3_U2421 ; P3_U4919
g3099 nand P3_U2374 P3_U2413 ; P3_U4920
g3100 nand P3_U4879 P3_INSTQUEUE_REG_11__0__SCAN_IN ; P3_U4921
g3101 not P3_U3170 ; P3_U4922
g3102 not P3_U3169 ; P3_U4923
g3103 nand P3_U2459 P3_U4342 ; P3_U4924
g3104 not P3_U3172 ; P3_U4925
g3105 nand P3_U4658 P3_U4644 ; P3_U4926
g3106 not P3_U3171 ; P3_U4927
g3107 nand P3_U2489 P3_U3171 ; P3_U4928
g3108 nand P3_U4925 P3_U4928 ; P3_U4929
g3109 nand P3_U3169 P3_STATE2_REG_3__SCAN_IN ; P3_U4930
g3110 nand P3_U3458 P3_U4929 ; P3_U4931
g3111 nand P3_U4927 P3_U4322 ; P3_U4932
g3112 nand P3_U2489 P3_U4932 ; P3_U4933
g3113 nand P3_U4923 P3_U2445 ; P3_U4934
g3114 nand P3_U2500 P3_U2436 ; P3_U4935
g3115 nand P3_U4922 P3_U2435 ; P3_U4936
g3116 nand P3_U2373 P3_U2420 ; P3_U4937
g3117 nand P3_U4931 P3_INSTQUEUE_REG_10__7__SCAN_IN ; P3_U4938
g3118 nand P3_U4923 P3_U2443 ; P3_U4939
g3119 nand P3_U2500 P3_U2434 ; P3_U4940
g3120 nand P3_U4922 P3_U2433 ; P3_U4941
g3121 nand P3_U2373 P3_U2419 ; P3_U4942
g3122 nand P3_U4931 P3_INSTQUEUE_REG_10__6__SCAN_IN ; P3_U4943
g3123 nand P3_U4923 P3_U2442 ; P3_U4944
g3124 nand P3_U2500 P3_U2432 ; P3_U4945
g3125 nand P3_U4922 P3_U2431 ; P3_U4946
g3126 nand P3_U2373 P3_U2418 ; P3_U4947
g3127 nand P3_U4931 P3_INSTQUEUE_REG_10__5__SCAN_IN ; P3_U4948
g3128 nand P3_U4923 P3_U2441 ; P3_U4949
g3129 nand P3_U2500 P3_U2430 ; P3_U4950
g3130 nand P3_U4922 P3_U2429 ; P3_U4951
g3131 nand P3_U2373 P3_U2417 ; P3_U4952
g3132 nand P3_U4931 P3_INSTQUEUE_REG_10__4__SCAN_IN ; P3_U4953
g3133 nand P3_U4923 P3_U2440 ; P3_U4954
g3134 nand P3_U2500 P3_U2428 ; P3_U4955
g3135 nand P3_U4922 P3_U2427 ; P3_U4956
g3136 nand P3_U2373 P3_U2416 ; P3_U4957
g3137 nand P3_U4931 P3_INSTQUEUE_REG_10__3__SCAN_IN ; P3_U4958
g3138 nand P3_U4923 P3_U2439 ; P3_U4959
g3139 nand P3_U2500 P3_U2426 ; P3_U4960
g3140 nand P3_U4922 P3_U2425 ; P3_U4961
g3141 nand P3_U2373 P3_U2415 ; P3_U4962
g3142 nand P3_U4931 P3_INSTQUEUE_REG_10__2__SCAN_IN ; P3_U4963
g3143 nand P3_U4923 P3_U2438 ; P3_U4964
g3144 nand P3_U2500 P3_U2424 ; P3_U4965
g3145 nand P3_U4922 P3_U2423 ; P3_U4966
g3146 nand P3_U2373 P3_U2414 ; P3_U4967
g3147 nand P3_U4931 P3_INSTQUEUE_REG_10__1__SCAN_IN ; P3_U4968
g3148 nand P3_U4923 P3_U2437 ; P3_U4969
g3149 nand P3_U2500 P3_U2422 ; P3_U4970
g3150 nand P3_U4922 P3_U2421 ; P3_U4971
g3151 nand P3_U2373 P3_U2413 ; P3_U4972
g3152 nand P3_U4931 P3_INSTQUEUE_REG_10__0__SCAN_IN ; P3_U4973
g3153 not P3_U3174 ; P3_U4974
g3154 not P3_U3173 ; P3_U4975
g3155 nand P3_U2459 P3_U4343 ; P3_U4976
g3156 not P3_U3176 ; P3_U4977
g3157 nand P3_U4658 P3_U4645 ; P3_U4978
g3158 not P3_U3175 ; P3_U4979
g3159 nand P3_U2489 P3_U3175 ; P3_U4980
g3160 nand P3_U4977 P3_U4980 ; P3_U4981
g3161 nand P3_U3173 P3_STATE2_REG_3__SCAN_IN ; P3_U4982
g3162 nand P3_U3476 P3_U4981 ; P3_U4983
g3163 nand P3_U4979 P3_U4322 ; P3_U4984
g3164 nand P3_U2489 P3_U4984 ; P3_U4985
g3165 nand P3_U4975 P3_U2445 ; P3_U4986
g3166 nand P3_U2502 P3_U2436 ; P3_U4987
g3167 nand P3_U4974 P3_U2435 ; P3_U4988
g3168 nand P3_U2372 P3_U2420 ; P3_U4989
g3169 nand P3_U4983 P3_INSTQUEUE_REG_9__7__SCAN_IN ; P3_U4990
g3170 nand P3_U4975 P3_U2443 ; P3_U4991
g3171 nand P3_U2502 P3_U2434 ; P3_U4992
g3172 nand P3_U4974 P3_U2433 ; P3_U4993
g3173 nand P3_U2372 P3_U2419 ; P3_U4994
g3174 nand P3_U4983 P3_INSTQUEUE_REG_9__6__SCAN_IN ; P3_U4995
g3175 nand P3_U4975 P3_U2442 ; P3_U4996
g3176 nand P3_U2502 P3_U2432 ; P3_U4997
g3177 nand P3_U4974 P3_U2431 ; P3_U4998
g3178 nand P3_U2372 P3_U2418 ; P3_U4999
g3179 nand P3_U4983 P3_INSTQUEUE_REG_9__5__SCAN_IN ; P3_U5000
g3180 nand P3_U4975 P3_U2441 ; P3_U5001
g3181 nand P3_U2502 P3_U2430 ; P3_U5002
g3182 nand P3_U4974 P3_U2429 ; P3_U5003
g3183 nand P3_U2372 P3_U2417 ; P3_U5004
g3184 nand P3_U4983 P3_INSTQUEUE_REG_9__4__SCAN_IN ; P3_U5005
g3185 nand P3_U4975 P3_U2440 ; P3_U5006
g3186 nand P3_U2502 P3_U2428 ; P3_U5007
g3187 nand P3_U4974 P3_U2427 ; P3_U5008
g3188 nand P3_U2372 P3_U2416 ; P3_U5009
g3189 nand P3_U4983 P3_INSTQUEUE_REG_9__3__SCAN_IN ; P3_U5010
g3190 nand P3_U4975 P3_U2439 ; P3_U5011
g3191 nand P3_U2502 P3_U2426 ; P3_U5012
g3192 nand P3_U4974 P3_U2425 ; P3_U5013
g3193 nand P3_U2372 P3_U2415 ; P3_U5014
g3194 nand P3_U4983 P3_INSTQUEUE_REG_9__2__SCAN_IN ; P3_U5015
g3195 nand P3_U4975 P3_U2438 ; P3_U5016
g3196 nand P3_U2502 P3_U2424 ; P3_U5017
g3197 nand P3_U4974 P3_U2423 ; P3_U5018
g3198 nand P3_U2372 P3_U2414 ; P3_U5019
g3199 nand P3_U4983 P3_INSTQUEUE_REG_9__1__SCAN_IN ; P3_U5020
g3200 nand P3_U4975 P3_U2437 ; P3_U5021
g3201 nand P3_U2502 P3_U2422 ; P3_U5022
g3202 nand P3_U4974 P3_U2421 ; P3_U5023
g3203 nand P3_U2372 P3_U2413 ; P3_U5024
g3204 nand P3_U4983 P3_INSTQUEUE_REG_9__0__SCAN_IN ; P3_U5025
g3205 not P3_U3178 ; P3_U5026
g3206 not P3_U3177 ; P3_U5027
g3207 not P3_U3071 ; P3_U5028
g3208 nand P3_U4658 P3_U2496 ; P3_U5029
g3209 not P3_U3179 ; P3_U5030
g3210 nand P3_U2489 P3_U3179 ; P3_U5031
g3211 nand P3_U5031 P3_U3071 ; P3_U5032
g3212 nand P3_U3177 P3_STATE2_REG_3__SCAN_IN ; P3_U5033
g3213 nand P3_U3493 P3_U5032 ; P3_U5034
g3214 nand P3_U5030 P3_U4322 ; P3_U5035
g3215 nand P3_U2489 P3_U5035 ; P3_U5036
g3216 nand P3_U5027 P3_U2445 ; P3_U5037
g3217 nand P3_U2503 P3_U2436 ; P3_U5038
g3218 nand P3_U5026 P3_U2435 ; P3_U5039
g3219 nand P3_U2371 P3_U2420 ; P3_U5040
g3220 nand P3_U5034 P3_INSTQUEUE_REG_8__7__SCAN_IN ; P3_U5041
g3221 nand P3_U5027 P3_U2443 ; P3_U5042
g3222 nand P3_U2503 P3_U2434 ; P3_U5043
g3223 nand P3_U5026 P3_U2433 ; P3_U5044
g3224 nand P3_U2371 P3_U2419 ; P3_U5045
g3225 nand P3_U5034 P3_INSTQUEUE_REG_8__6__SCAN_IN ; P3_U5046
g3226 nand P3_U5027 P3_U2442 ; P3_U5047
g3227 nand P3_U2503 P3_U2432 ; P3_U5048
g3228 nand P3_U5026 P3_U2431 ; P3_U5049
g3229 nand P3_U2371 P3_U2418 ; P3_U5050
g3230 nand P3_U5034 P3_INSTQUEUE_REG_8__5__SCAN_IN ; P3_U5051
g3231 nand P3_U5027 P3_U2441 ; P3_U5052
g3232 nand P3_U2503 P3_U2430 ; P3_U5053
g3233 nand P3_U5026 P3_U2429 ; P3_U5054
g3234 nand P3_U2371 P3_U2417 ; P3_U5055
g3235 nand P3_U5034 P3_INSTQUEUE_REG_8__4__SCAN_IN ; P3_U5056
g3236 nand P3_U5027 P3_U2440 ; P3_U5057
g3237 nand P3_U2503 P3_U2428 ; P3_U5058
g3238 nand P3_U5026 P3_U2427 ; P3_U5059
g3239 nand P3_U2371 P3_U2416 ; P3_U5060
g3240 nand P3_U5034 P3_INSTQUEUE_REG_8__3__SCAN_IN ; P3_U5061
g3241 nand P3_U5027 P3_U2439 ; P3_U5062
g3242 nand P3_U2503 P3_U2426 ; P3_U5063
g3243 nand P3_U5026 P3_U2425 ; P3_U5064
g3244 nand P3_U2371 P3_U2415 ; P3_U5065
g3245 nand P3_U5034 P3_INSTQUEUE_REG_8__2__SCAN_IN ; P3_U5066
g3246 nand P3_U5027 P3_U2438 ; P3_U5067
g3247 nand P3_U2503 P3_U2424 ; P3_U5068
g3248 nand P3_U5026 P3_U2423 ; P3_U5069
g3249 nand P3_U2371 P3_U2414 ; P3_U5070
g3250 nand P3_U5034 P3_INSTQUEUE_REG_8__1__SCAN_IN ; P3_U5071
g3251 nand P3_U5027 P3_U2437 ; P3_U5072
g3252 nand P3_U2503 P3_U2422 ; P3_U5073
g3253 nand P3_U5026 P3_U2421 ; P3_U5074
g3254 nand P3_U2371 P3_U2413 ; P3_U5075
g3255 nand P3_U5034 P3_INSTQUEUE_REG_8__0__SCAN_IN ; P3_U5076
g3256 not P3_U3183 ; P3_U5077
g3257 not P3_U3185 ; P3_U5078
g3258 not P3_U3184 ; P3_U5079
g3259 nand P3_U2489 P3_U3184 ; P3_U5080
g3260 nand P3_U5078 P3_U5080 ; P3_U5081
g3261 nand P3_U3180 P3_STATE2_REG_3__SCAN_IN ; P3_U5082
g3262 nand P3_U3510 P3_U5081 ; P3_U5083
g3263 nand P3_U5079 P3_U4322 ; P3_U5084
g3264 nand P3_U2489 P3_U5084 ; P3_U5085
g3265 nand P3_U4650 P3_U2445 ; P3_U5086
g3266 nand P3_U4326 P3_U2436 ; P3_U5087
g3267 nand P3_U5077 P3_U2435 ; P3_U5088
g3268 nand P3_U2370 P3_U2420 ; P3_U5089
g3269 nand P3_U5083 P3_INSTQUEUE_REG_7__7__SCAN_IN ; P3_U5090
g3270 nand P3_U4650 P3_U2443 ; P3_U5091
g3271 nand P3_U4326 P3_U2434 ; P3_U5092
g3272 nand P3_U5077 P3_U2433 ; P3_U5093
g3273 nand P3_U2370 P3_U2419 ; P3_U5094
g3274 nand P3_U5083 P3_INSTQUEUE_REG_7__6__SCAN_IN ; P3_U5095
g3275 nand P3_U4650 P3_U2442 ; P3_U5096
g3276 nand P3_U4326 P3_U2432 ; P3_U5097
g3277 nand P3_U5077 P3_U2431 ; P3_U5098
g3278 nand P3_U2370 P3_U2418 ; P3_U5099
g3279 nand P3_U5083 P3_INSTQUEUE_REG_7__5__SCAN_IN ; P3_U5100
g3280 nand P3_U4650 P3_U2441 ; P3_U5101
g3281 nand P3_U4326 P3_U2430 ; P3_U5102
g3282 nand P3_U5077 P3_U2429 ; P3_U5103
g3283 nand P3_U2370 P3_U2417 ; P3_U5104
g3284 nand P3_U5083 P3_INSTQUEUE_REG_7__4__SCAN_IN ; P3_U5105
g3285 nand P3_U4650 P3_U2440 ; P3_U5106
g3286 nand P3_U4326 P3_U2428 ; P3_U5107
g3287 nand P3_U5077 P3_U2427 ; P3_U5108
g3288 nand P3_U2370 P3_U2416 ; P3_U5109
g3289 nand P3_U5083 P3_INSTQUEUE_REG_7__3__SCAN_IN ; P3_U5110
g3290 nand P3_U4650 P3_U2439 ; P3_U5111
g3291 nand P3_U4326 P3_U2426 ; P3_U5112
g3292 nand P3_U5077 P3_U2425 ; P3_U5113
g3293 nand P3_U2370 P3_U2415 ; P3_U5114
g3294 nand P3_U5083 P3_INSTQUEUE_REG_7__2__SCAN_IN ; P3_U5115
g3295 nand P3_U4650 P3_U2438 ; P3_U5116
g3296 nand P3_U4326 P3_U2424 ; P3_U5117
g3297 nand P3_U5077 P3_U2423 ; P3_U5118
g3298 nand P3_U2370 P3_U2414 ; P3_U5119
g3299 nand P3_U5083 P3_INSTQUEUE_REG_7__1__SCAN_IN ; P3_U5120
g3300 nand P3_U4650 P3_U2437 ; P3_U5121
g3301 nand P3_U4326 P3_U2422 ; P3_U5122
g3302 nand P3_U5077 P3_U2421 ; P3_U5123
g3303 nand P3_U2370 P3_U2413 ; P3_U5124
g3304 nand P3_U5083 P3_INSTQUEUE_REG_7__0__SCAN_IN ; P3_U5125
g3305 not P3_U3187 ; P3_U5126
g3306 not P3_U3186 ; P3_U5127
g3307 nand P3_U4342 P3_U2458 ; P3_U5128
g3308 not P3_U3189 ; P3_U5129
g3309 nand P3_U4644 P3_U2485 ; P3_U5130
g3310 not P3_U3188 ; P3_U5131
g3311 nand P3_U2489 P3_U3188 ; P3_U5132
g3312 nand P3_U5129 P3_U5132 ; P3_U5133
g3313 nand P3_U3186 P3_STATE2_REG_3__SCAN_IN ; P3_U5134
g3314 nand P3_U3528 P3_U5133 ; P3_U5135
g3315 nand P3_U5131 P3_U4322 ; P3_U5136
g3316 nand P3_U2489 P3_U5136 ; P3_U5137
g3317 nand P3_U5127 P3_U2445 ; P3_U5138
g3318 nand P3_U2505 P3_U2436 ; P3_U5139
g3319 nand P3_U5126 P3_U2435 ; P3_U5140
g3320 nand P3_U2369 P3_U2420 ; P3_U5141
g3321 nand P3_U5135 P3_INSTQUEUE_REG_6__7__SCAN_IN ; P3_U5142
g3322 nand P3_U5127 P3_U2443 ; P3_U5143
g3323 nand P3_U2505 P3_U2434 ; P3_U5144
g3324 nand P3_U5126 P3_U2433 ; P3_U5145
g3325 nand P3_U2369 P3_U2419 ; P3_U5146
g3326 nand P3_U5135 P3_INSTQUEUE_REG_6__6__SCAN_IN ; P3_U5147
g3327 nand P3_U5127 P3_U2442 ; P3_U5148
g3328 nand P3_U2505 P3_U2432 ; P3_U5149
g3329 nand P3_U5126 P3_U2431 ; P3_U5150
g3330 nand P3_U2369 P3_U2418 ; P3_U5151
g3331 nand P3_U5135 P3_INSTQUEUE_REG_6__5__SCAN_IN ; P3_U5152
g3332 nand P3_U5127 P3_U2441 ; P3_U5153
g3333 nand P3_U2505 P3_U2430 ; P3_U5154
g3334 nand P3_U5126 P3_U2429 ; P3_U5155
g3335 nand P3_U2369 P3_U2417 ; P3_U5156
g3336 nand P3_U5135 P3_INSTQUEUE_REG_6__4__SCAN_IN ; P3_U5157
g3337 nand P3_U5127 P3_U2440 ; P3_U5158
g3338 nand P3_U2505 P3_U2428 ; P3_U5159
g3339 nand P3_U5126 P3_U2427 ; P3_U5160
g3340 nand P3_U2369 P3_U2416 ; P3_U5161
g3341 nand P3_U5135 P3_INSTQUEUE_REG_6__3__SCAN_IN ; P3_U5162
g3342 nand P3_U5127 P3_U2439 ; P3_U5163
g3343 nand P3_U2505 P3_U2426 ; P3_U5164
g3344 nand P3_U5126 P3_U2425 ; P3_U5165
g3345 nand P3_U2369 P3_U2415 ; P3_U5166
g3346 nand P3_U5135 P3_INSTQUEUE_REG_6__2__SCAN_IN ; P3_U5167
g3347 nand P3_U5127 P3_U2438 ; P3_U5168
g3348 nand P3_U2505 P3_U2424 ; P3_U5169
g3349 nand P3_U5126 P3_U2423 ; P3_U5170
g3350 nand P3_U2369 P3_U2414 ; P3_U5171
g3351 nand P3_U5135 P3_INSTQUEUE_REG_6__1__SCAN_IN ; P3_U5172
g3352 nand P3_U5127 P3_U2437 ; P3_U5173
g3353 nand P3_U2505 P3_U2422 ; P3_U5174
g3354 nand P3_U5126 P3_U2421 ; P3_U5175
g3355 nand P3_U2369 P3_U2413 ; P3_U5176
g3356 nand P3_U5135 P3_INSTQUEUE_REG_6__0__SCAN_IN ; P3_U5177
g3357 not P3_U3191 ; P3_U5178
g3358 not P3_U3190 ; P3_U5179
g3359 nand P3_U4343 P3_U2458 ; P3_U5180
g3360 not P3_U3193 ; P3_U5181
g3361 nand P3_U4645 P3_U2485 ; P3_U5182
g3362 not P3_U3192 ; P3_U5183
g3363 nand P3_U2489 P3_U3192 ; P3_U5184
g3364 nand P3_U5181 P3_U5184 ; P3_U5185
g3365 nand P3_U3190 P3_STATE2_REG_3__SCAN_IN ; P3_U5186
g3366 nand P3_U3546 P3_U5185 ; P3_U5187
g3367 nand P3_U5183 P3_U4322 ; P3_U5188
g3368 nand P3_U2489 P3_U5188 ; P3_U5189
g3369 nand P3_U5179 P3_U2445 ; P3_U5190
g3370 nand P3_U2506 P3_U2436 ; P3_U5191
g3371 nand P3_U5178 P3_U2435 ; P3_U5192
g3372 nand P3_U2368 P3_U2420 ; P3_U5193
g3373 nand P3_U5187 P3_INSTQUEUE_REG_5__7__SCAN_IN ; P3_U5194
g3374 nand P3_U5179 P3_U2443 ; P3_U5195
g3375 nand P3_U2506 P3_U2434 ; P3_U5196
g3376 nand P3_U5178 P3_U2433 ; P3_U5197
g3377 nand P3_U2368 P3_U2419 ; P3_U5198
g3378 nand P3_U5187 P3_INSTQUEUE_REG_5__6__SCAN_IN ; P3_U5199
g3379 nand P3_U5179 P3_U2442 ; P3_U5200
g3380 nand P3_U2506 P3_U2432 ; P3_U5201
g3381 nand P3_U5178 P3_U2431 ; P3_U5202
g3382 nand P3_U2368 P3_U2418 ; P3_U5203
g3383 nand P3_U5187 P3_INSTQUEUE_REG_5__5__SCAN_IN ; P3_U5204
g3384 nand P3_U5179 P3_U2441 ; P3_U5205
g3385 nand P3_U2506 P3_U2430 ; P3_U5206
g3386 nand P3_U5178 P3_U2429 ; P3_U5207
g3387 nand P3_U2368 P3_U2417 ; P3_U5208
g3388 nand P3_U5187 P3_INSTQUEUE_REG_5__4__SCAN_IN ; P3_U5209
g3389 nand P3_U5179 P3_U2440 ; P3_U5210
g3390 nand P3_U2506 P3_U2428 ; P3_U5211
g3391 nand P3_U5178 P3_U2427 ; P3_U5212
g3392 nand P3_U2368 P3_U2416 ; P3_U5213
g3393 nand P3_U5187 P3_INSTQUEUE_REG_5__3__SCAN_IN ; P3_U5214
g3394 nand P3_U5179 P3_U2439 ; P3_U5215
g3395 nand P3_U2506 P3_U2426 ; P3_U5216
g3396 nand P3_U5178 P3_U2425 ; P3_U5217
g3397 nand P3_U2368 P3_U2415 ; P3_U5218
g3398 nand P3_U5187 P3_INSTQUEUE_REG_5__2__SCAN_IN ; P3_U5219
g3399 nand P3_U5179 P3_U2438 ; P3_U5220
g3400 nand P3_U2506 P3_U2424 ; P3_U5221
g3401 nand P3_U5178 P3_U2423 ; P3_U5222
g3402 nand P3_U2368 P3_U2414 ; P3_U5223
g3403 nand P3_U5187 P3_INSTQUEUE_REG_5__1__SCAN_IN ; P3_U5224
g3404 nand P3_U5179 P3_U2437 ; P3_U5225
g3405 nand P3_U2506 P3_U2422 ; P3_U5226
g3406 nand P3_U5178 P3_U2421 ; P3_U5227
g3407 nand P3_U2368 P3_U2413 ; P3_U5228
g3408 nand P3_U5187 P3_INSTQUEUE_REG_5__0__SCAN_IN ; P3_U5229
g3409 not P3_U3195 ; P3_U5230
g3410 not P3_U3194 ; P3_U5231
g3411 not P3_U3072 ; P3_U5232
g3412 nand P3_U2496 P3_U2485 ; P3_U5233
g3413 nand P3_U3195 P3_U5233 ; P3_U5234
g3414 nand P3_U2489 P3_U5234 ; P3_U5235
g3415 nand P3_U5235 P3_U3072 ; P3_U5236
g3416 nand P3_U3194 P3_STATE2_REG_3__SCAN_IN ; P3_U5237
g3417 nand P3_U3564 P3_U5236 ; P3_U5238
g3418 nand P3_U2489 P3_U3136 ; P3_U5239
g3419 nand P3_U5231 P3_U2445 ; P3_U5240
g3420 nand P3_U2507 P3_U2436 ; P3_U5241
g3421 nand P3_U5230 P3_U2435 ; P3_U5242
g3422 nand P3_U2367 P3_U2420 ; P3_U5243
g3423 nand P3_U5238 P3_INSTQUEUE_REG_4__7__SCAN_IN ; P3_U5244
g3424 nand P3_U5231 P3_U2443 ; P3_U5245
g3425 nand P3_U2507 P3_U2434 ; P3_U5246
g3426 nand P3_U5230 P3_U2433 ; P3_U5247
g3427 nand P3_U2367 P3_U2419 ; P3_U5248
g3428 nand P3_U5238 P3_INSTQUEUE_REG_4__6__SCAN_IN ; P3_U5249
g3429 nand P3_U5231 P3_U2442 ; P3_U5250
g3430 nand P3_U2507 P3_U2432 ; P3_U5251
g3431 nand P3_U5230 P3_U2431 ; P3_U5252
g3432 nand P3_U2367 P3_U2418 ; P3_U5253
g3433 nand P3_U5238 P3_INSTQUEUE_REG_4__5__SCAN_IN ; P3_U5254
g3434 nand P3_U5231 P3_U2441 ; P3_U5255
g3435 nand P3_U2507 P3_U2430 ; P3_U5256
g3436 nand P3_U5230 P3_U2429 ; P3_U5257
g3437 nand P3_U2367 P3_U2417 ; P3_U5258
g3438 nand P3_U5238 P3_INSTQUEUE_REG_4__4__SCAN_IN ; P3_U5259
g3439 nand P3_U5231 P3_U2440 ; P3_U5260
g3440 nand P3_U2507 P3_U2428 ; P3_U5261
g3441 nand P3_U5230 P3_U2427 ; P3_U5262
g3442 nand P3_U2367 P3_U2416 ; P3_U5263
g3443 nand P3_U5238 P3_INSTQUEUE_REG_4__3__SCAN_IN ; P3_U5264
g3444 nand P3_U5231 P3_U2439 ; P3_U5265
g3445 nand P3_U2507 P3_U2426 ; P3_U5266
g3446 nand P3_U5230 P3_U2425 ; P3_U5267
g3447 nand P3_U2367 P3_U2415 ; P3_U5268
g3448 nand P3_U5238 P3_INSTQUEUE_REG_4__2__SCAN_IN ; P3_U5269
g3449 nand P3_U5231 P3_U2438 ; P3_U5270
g3450 nand P3_U2507 P3_U2424 ; P3_U5271
g3451 nand P3_U5230 P3_U2423 ; P3_U5272
g3452 nand P3_U2367 P3_U2414 ; P3_U5273
g3453 nand P3_U5238 P3_INSTQUEUE_REG_4__1__SCAN_IN ; P3_U5274
g3454 nand P3_U5231 P3_U2437 ; P3_U5275
g3455 nand P3_U2507 P3_U2422 ; P3_U5276
g3456 nand P3_U5230 P3_U2421 ; P3_U5277
g3457 nand P3_U2367 P3_U2413 ; P3_U5278
g3458 nand P3_U5238 P3_INSTQUEUE_REG_4__0__SCAN_IN ; P3_U5279
g3459 not P3_U3197 ; P3_U5280
g3460 not P3_U3196 ; P3_U5281
g3461 nand P3_U2460 P3_U4653 ; P3_U5282
g3462 not P3_U3198 ; P3_U5283
g3463 nand P3_U2509 P3_U4657 ; P3_U5284
g3464 nand P3_U3197 P3_U5284 ; P3_U5285
g3465 nand P3_U2489 P3_U5285 ; P3_U5286
g3466 nand P3_U5283 P3_U5286 ; P3_U5287
g3467 nand P3_U3196 P3_STATE2_REG_3__SCAN_IN ; P3_U5288
g3468 nand P3_U3582 P3_U5287 ; P3_U5289
g3469 nand P3_U2489 P3_U3136 ; P3_U5290
g3470 nand P3_U5281 P3_U2445 ; P3_U5291
g3471 nand P3_U2510 P3_U2436 ; P3_U5292
g3472 nand P3_U5280 P3_U2435 ; P3_U5293
g3473 nand P3_U2366 P3_U2420 ; P3_U5294
g3474 nand P3_U5289 P3_INSTQUEUE_REG_3__7__SCAN_IN ; P3_U5295
g3475 nand P3_U5281 P3_U2443 ; P3_U5296
g3476 nand P3_U2510 P3_U2434 ; P3_U5297
g3477 nand P3_U5280 P3_U2433 ; P3_U5298
g3478 nand P3_U2366 P3_U2419 ; P3_U5299
g3479 nand P3_U5289 P3_INSTQUEUE_REG_3__6__SCAN_IN ; P3_U5300
g3480 nand P3_U5281 P3_U2442 ; P3_U5301
g3481 nand P3_U2510 P3_U2432 ; P3_U5302
g3482 nand P3_U5280 P3_U2431 ; P3_U5303
g3483 nand P3_U2366 P3_U2418 ; P3_U5304
g3484 nand P3_U5289 P3_INSTQUEUE_REG_3__5__SCAN_IN ; P3_U5305
g3485 nand P3_U5281 P3_U2441 ; P3_U5306
g3486 nand P3_U2510 P3_U2430 ; P3_U5307
g3487 nand P3_U5280 P3_U2429 ; P3_U5308
g3488 nand P3_U2366 P3_U2417 ; P3_U5309
g3489 nand P3_U5289 P3_INSTQUEUE_REG_3__4__SCAN_IN ; P3_U5310
g3490 nand P3_U5281 P3_U2440 ; P3_U5311
g3491 nand P3_U2510 P3_U2428 ; P3_U5312
g3492 nand P3_U5280 P3_U2427 ; P3_U5313
g3493 nand P3_U2366 P3_U2416 ; P3_U5314
g3494 nand P3_U5289 P3_INSTQUEUE_REG_3__3__SCAN_IN ; P3_U5315
g3495 nand P3_U5281 P3_U2439 ; P3_U5316
g3496 nand P3_U2510 P3_U2426 ; P3_U5317
g3497 nand P3_U5280 P3_U2425 ; P3_U5318
g3498 nand P3_U2366 P3_U2415 ; P3_U5319
g3499 nand P3_U5289 P3_INSTQUEUE_REG_3__2__SCAN_IN ; P3_U5320
g3500 nand P3_U5281 P3_U2438 ; P3_U5321
g3501 nand P3_U2510 P3_U2424 ; P3_U5322
g3502 nand P3_U5280 P3_U2423 ; P3_U5323
g3503 nand P3_U2366 P3_U2414 ; P3_U5324
g3504 nand P3_U5289 P3_INSTQUEUE_REG_3__1__SCAN_IN ; P3_U5325
g3505 nand P3_U5281 P3_U2437 ; P3_U5326
g3506 nand P3_U2510 P3_U2422 ; P3_U5327
g3507 nand P3_U5280 P3_U2421 ; P3_U5328
g3508 nand P3_U2366 P3_U2413 ; P3_U5329
g3509 nand P3_U5289 P3_INSTQUEUE_REG_3__0__SCAN_IN ; P3_U5330
g3510 not P3_U3200 ; P3_U5331
g3511 not P3_U3199 ; P3_U5332
g3512 nand P3_U2460 P3_U4342 ; P3_U5333
g3513 not P3_U3201 ; P3_U5334
g3514 nand P3_U2509 P3_U4644 ; P3_U5335
g3515 nand P3_U3200 P3_U5335 ; P3_U5336
g3516 nand P3_U2489 P3_U5336 ; P3_U5337
g3517 nand P3_U5334 P3_U5337 ; P3_U5338
g3518 nand P3_U3199 P3_STATE2_REG_3__SCAN_IN ; P3_U5339
g3519 nand P3_U3599 P3_U5338 ; P3_U5340
g3520 nand P3_U2489 P3_U3136 ; P3_U5341
g3521 nand P3_U5332 P3_U2445 ; P3_U5342
g3522 nand P3_U2511 P3_U2436 ; P3_U5343
g3523 nand P3_U5331 P3_U2435 ; P3_U5344
g3524 nand P3_U2365 P3_U2420 ; P3_U5345
g3525 nand P3_U5340 P3_INSTQUEUE_REG_2__7__SCAN_IN ; P3_U5346
g3526 nand P3_U5332 P3_U2443 ; P3_U5347
g3527 nand P3_U2511 P3_U2434 ; P3_U5348
g3528 nand P3_U5331 P3_U2433 ; P3_U5349
g3529 nand P3_U2365 P3_U2419 ; P3_U5350
g3530 nand P3_U5340 P3_INSTQUEUE_REG_2__6__SCAN_IN ; P3_U5351
g3531 nand P3_U5332 P3_U2442 ; P3_U5352
g3532 nand P3_U2511 P3_U2432 ; P3_U5353
g3533 nand P3_U5331 P3_U2431 ; P3_U5354
g3534 nand P3_U2365 P3_U2418 ; P3_U5355
g3535 nand P3_U5340 P3_INSTQUEUE_REG_2__5__SCAN_IN ; P3_U5356
g3536 nand P3_U5332 P3_U2441 ; P3_U5357
g3537 nand P3_U2511 P3_U2430 ; P3_U5358
g3538 nand P3_U5331 P3_U2429 ; P3_U5359
g3539 nand P3_U2365 P3_U2417 ; P3_U5360
g3540 nand P3_U5340 P3_INSTQUEUE_REG_2__4__SCAN_IN ; P3_U5361
g3541 nand P3_U5332 P3_U2440 ; P3_U5362
g3542 nand P3_U2511 P3_U2428 ; P3_U5363
g3543 nand P3_U5331 P3_U2427 ; P3_U5364
g3544 nand P3_U2365 P3_U2416 ; P3_U5365
g3545 nand P3_U5340 P3_INSTQUEUE_REG_2__3__SCAN_IN ; P3_U5366
g3546 nand P3_U5332 P3_U2439 ; P3_U5367
g3547 nand P3_U2511 P3_U2426 ; P3_U5368
g3548 nand P3_U5331 P3_U2425 ; P3_U5369
g3549 nand P3_U2365 P3_U2415 ; P3_U5370
g3550 nand P3_U5340 P3_INSTQUEUE_REG_2__2__SCAN_IN ; P3_U5371
g3551 nand P3_U5332 P3_U2438 ; P3_U5372
g3552 nand P3_U2511 P3_U2424 ; P3_U5373
g3553 nand P3_U5331 P3_U2423 ; P3_U5374
g3554 nand P3_U2365 P3_U2414 ; P3_U5375
g3555 nand P3_U5340 P3_INSTQUEUE_REG_2__1__SCAN_IN ; P3_U5376
g3556 nand P3_U5332 P3_U2437 ; P3_U5377
g3557 nand P3_U2511 P3_U2422 ; P3_U5378
g3558 nand P3_U5331 P3_U2421 ; P3_U5379
g3559 nand P3_U2365 P3_U2413 ; P3_U5380
g3560 nand P3_U5340 P3_INSTQUEUE_REG_2__0__SCAN_IN ; P3_U5381
g3561 not P3_U3203 ; P3_U5382
g3562 not P3_U3202 ; P3_U5383
g3563 nand P3_U2460 P3_U4343 ; P3_U5384
g3564 not P3_U3204 ; P3_U5385
g3565 nand P3_U2509 P3_U4645 ; P3_U5386
g3566 nand P3_U3203 P3_U5386 ; P3_U5387
g3567 nand P3_U2489 P3_U5387 ; P3_U5388
g3568 nand P3_U5385 P3_U5388 ; P3_U5389
g3569 nand P3_U3202 P3_STATE2_REG_3__SCAN_IN ; P3_U5390
g3570 nand P3_U3617 P3_U5389 ; P3_U5391
g3571 nand P3_U2489 P3_U3136 ; P3_U5392
g3572 nand P3_U5383 P3_U2445 ; P3_U5393
g3573 nand P3_U2512 P3_U2436 ; P3_U5394
g3574 nand P3_U5382 P3_U2435 ; P3_U5395
g3575 nand P3_U2364 P3_U2420 ; P3_U5396
g3576 nand P3_U5391 P3_INSTQUEUE_REG_1__7__SCAN_IN ; P3_U5397
g3577 nand P3_U5383 P3_U2443 ; P3_U5398
g3578 nand P3_U2512 P3_U2434 ; P3_U5399
g3579 nand P3_U5382 P3_U2433 ; P3_U5400
g3580 nand P3_U2364 P3_U2419 ; P3_U5401
g3581 nand P3_U5391 P3_INSTQUEUE_REG_1__6__SCAN_IN ; P3_U5402
g3582 nand P3_U5383 P3_U2442 ; P3_U5403
g3583 nand P3_U2512 P3_U2432 ; P3_U5404
g3584 nand P3_U5382 P3_U2431 ; P3_U5405
g3585 nand P3_U2364 P3_U2418 ; P3_U5406
g3586 nand P3_U5391 P3_INSTQUEUE_REG_1__5__SCAN_IN ; P3_U5407
g3587 nand P3_U5383 P3_U2441 ; P3_U5408
g3588 nand P3_U2512 P3_U2430 ; P3_U5409
g3589 nand P3_U5382 P3_U2429 ; P3_U5410
g3590 nand P3_U2364 P3_U2417 ; P3_U5411
g3591 nand P3_U5391 P3_INSTQUEUE_REG_1__4__SCAN_IN ; P3_U5412
g3592 nand P3_U5383 P3_U2440 ; P3_U5413
g3593 nand P3_U2512 P3_U2428 ; P3_U5414
g3594 nand P3_U5382 P3_U2427 ; P3_U5415
g3595 nand P3_U2364 P3_U2416 ; P3_U5416
g3596 nand P3_U5391 P3_INSTQUEUE_REG_1__3__SCAN_IN ; P3_U5417
g3597 nand P3_U5383 P3_U2439 ; P3_U5418
g3598 nand P3_U2512 P3_U2426 ; P3_U5419
g3599 nand P3_U5382 P3_U2425 ; P3_U5420
g3600 nand P3_U2364 P3_U2415 ; P3_U5421
g3601 nand P3_U5391 P3_INSTQUEUE_REG_1__2__SCAN_IN ; P3_U5422
g3602 nand P3_U5383 P3_U2438 ; P3_U5423
g3603 nand P3_U2512 P3_U2424 ; P3_U5424
g3604 nand P3_U5382 P3_U2423 ; P3_U5425
g3605 nand P3_U2364 P3_U2414 ; P3_U5426
g3606 nand P3_U5391 P3_INSTQUEUE_REG_1__1__SCAN_IN ; P3_U5427
g3607 nand P3_U5383 P3_U2437 ; P3_U5428
g3608 nand P3_U2512 P3_U2422 ; P3_U5429
g3609 nand P3_U5382 P3_U2421 ; P3_U5430
g3610 nand P3_U2364 P3_U2413 ; P3_U5431
g3611 nand P3_U5391 P3_INSTQUEUE_REG_1__0__SCAN_IN ; P3_U5432
g3612 not P3_U3206 ; P3_U5433
g3613 not P3_U3205 ; P3_U5434
g3614 not P3_U3073 ; P3_U5435
g3615 nand P3_U2509 P3_U2496 ; P3_U5436
g3616 nand P3_U3206 P3_U5436 ; P3_U5437
g3617 nand P3_U2489 P3_U5437 ; P3_U5438
g3618 nand P3_U5438 P3_U3073 ; P3_U5439
g3619 nand P3_U3205 P3_STATE2_REG_3__SCAN_IN ; P3_U5440
g3620 nand P3_U3635 P3_U5439 ; P3_U5441
g3621 nand P3_U2489 P3_U3136 ; P3_U5442
g3622 nand P3_U5434 P3_U2445 ; P3_U5443
g3623 nand P3_U2513 P3_U2436 ; P3_U5444
g3624 nand P3_U5433 P3_U2435 ; P3_U5445
g3625 nand P3_U2363 P3_U2420 ; P3_U5446
g3626 nand P3_U5441 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U5447
g3627 nand P3_U5434 P3_U2443 ; P3_U5448
g3628 nand P3_U2513 P3_U2434 ; P3_U5449
g3629 nand P3_U5433 P3_U2433 ; P3_U5450
g3630 nand P3_U2363 P3_U2419 ; P3_U5451
g3631 nand P3_U5441 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U5452
g3632 nand P3_U5434 P3_U2442 ; P3_U5453
g3633 nand P3_U2513 P3_U2432 ; P3_U5454
g3634 nand P3_U5433 P3_U2431 ; P3_U5455
g3635 nand P3_U2363 P3_U2418 ; P3_U5456
g3636 nand P3_U5441 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U5457
g3637 nand P3_U5434 P3_U2441 ; P3_U5458
g3638 nand P3_U2513 P3_U2430 ; P3_U5459
g3639 nand P3_U5433 P3_U2429 ; P3_U5460
g3640 nand P3_U2363 P3_U2417 ; P3_U5461
g3641 nand P3_U5441 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U5462
g3642 nand P3_U5434 P3_U2440 ; P3_U5463
g3643 nand P3_U2513 P3_U2428 ; P3_U5464
g3644 nand P3_U5433 P3_U2427 ; P3_U5465
g3645 nand P3_U2363 P3_U2416 ; P3_U5466
g3646 nand P3_U5441 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U5467
g3647 nand P3_U5434 P3_U2439 ; P3_U5468
g3648 nand P3_U2513 P3_U2426 ; P3_U5469
g3649 nand P3_U5433 P3_U2425 ; P3_U5470
g3650 nand P3_U2363 P3_U2415 ; P3_U5471
g3651 nand P3_U5441 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U5472
g3652 nand P3_U5434 P3_U2438 ; P3_U5473
g3653 nand P3_U2513 P3_U2424 ; P3_U5474
g3654 nand P3_U5433 P3_U2423 ; P3_U5475
g3655 nand P3_U2363 P3_U2414 ; P3_U5476
g3656 nand P3_U5441 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U5477
g3657 nand P3_U5434 P3_U2437 ; P3_U5478
g3658 nand P3_U2513 P3_U2422 ; P3_U5479
g3659 nand P3_U5433 P3_U2421 ; P3_U5480
g3660 nand P3_U2363 P3_U2413 ; P3_U5481
g3661 nand P3_U5441 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U5482
g3662 nand P3_U7917 P3_U2514 P3_U3655 P3_U4339 ; P3_U5483
g3663 not P3_U3209 ; P3_U5484
g3664 nand P3_U4296 P3_U3209 ; P3_U5485
g3665 nand P3_GTE_450_U6 P3_U4303 ; P3_U5486
g3666 nand P3_GTE_504_U6 P3_U4302 ; P3_U5487
g3667 not P3_U3255 ; P3_U5488
g3668 nand P3_GTE_412_U6 P3_U4304 ; P3_U5489
g3669 nand P3_GTE_485_U6 P3_U2356 ; P3_U5490
g3670 not P3_U3254 ; P3_U5491
g3671 nand P3_U3254 P3_U2630 ; P3_U5492
g3672 nand P3_GTE_390_U6 P3_U2357 ; P3_U5493
g3673 nand P3_U4294 P3_U3255 ; P3_U5494
g3674 nand P3_GTE_401_U6 P3_U4305 ; P3_U5495
g3675 not P3_U4290 ; P3_U5496
g3676 nand P3_U2390 P3_U4290 ; P3_U5497
g3677 nand P3_U3121 P3_STATE2_REG_3__SCAN_IN ; P3_U5498
g3678 not P3_U4283 ; P3_U5499
g3679 nand P3_U3095 P3_U3097 ; P3_U5500
g3680 nand P3_U5500 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U5501
g3681 nand P3_U2481 P3_U3095 ; P3_U5502
g3682 nand P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U5503
g3683 not P3_U3223 ; P3_U5504
g3684 nand P3_U4332 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U5505
g3685 not P3_U3224 ; P3_U5506
g3686 nand P3_U5484 P3_U3107 ; P3_U5507
g3687 nand P3_U4522 P3_U4607 P3_U4488 ; P3_U5508
g3688 nand P3_U4296 P3_U5507 ; P3_U5509
g3689 nand P3_U7974 P3_U7973 P3_U3104 ; P3_U5510
g3690 nand P3_U4323 P3_U4344 ; P3_U5511
g3691 nand P3_U5509 P3_U3665 ; P3_U5512
g3692 nand P3_U4522 P3_U4607 ; P3_U5513
g3693 nand P3_U4607 P3_U3218 ; P3_U5514
g3694 nand P3_U5514 P3_U3216 P3_U4556 ; P3_U5515
g3695 nand P3_U4573 P3_U4505 ; P3_U5516
g3696 nand P3_U4488 P3_U5516 ; P3_U5517
g3697 nand P3_U3103 P3_U3218 P3_U3112 ; P3_U5518
g3698 nand P3_U4607 P3_U3104 P3_U4573 ; P3_U5519
g3699 nand P3_U4324 P3_U3103 ; P3_U5520
g3700 nand P3_U5518 P3_U3102 ; P3_U5521
g3701 not P3_U3220 ; P3_U5522
g3702 nand P3_U3111 P3_U3114 ; P3_U5523
g3703 nand P3_U2452 P3_U3108 ; P3_U5524
g3704 not P3_U3221 ; P3_U5525
g3705 nand P3_U2462 P3_U3104 ; P3_U5526
g3706 nand P3_U3229 P3_U3219 ; P3_U5527
g3707 nand P3_U2456 P3_U5527 ; P3_U5528
g3708 nand P3_U2518 P3_U3217 ; P3_U5529
g3709 nand P3_U5529 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U5530
g3710 nand P3_U5525 P3_U5530 ; P3_U5531
g3711 nand P3_U2461 P3_U5523 P3_U2450 ; P3_U5532
g3712 nand P3_U3673 P3_U7918 ; P3_U5533
g3713 not P3_U3226 ; P3_U5534
g3714 nand P3_U3672 P3_U5522 ; P3_U5535
g3715 nand P3_U3659 P3_U5523 P3_U2451 ; P3_U5536
g3716 nand P3_U3669 P3_U5531 ; P3_U5537
g3717 nand P3_U3670 P3_U3220 ; P3_U5538
g3718 nand P3_U5504 P3_U5535 ; P3_U5539
g3719 nand P3_U5506 P3_U3226 ; P3_U5540
g3720 nand P3_ADD_495_U9 P3_U2356 ; P3_U5541
g3721 nand P3_U5537 P3_U3676 ; P3_U5542
g3722 not P3_U3265 ; P3_U5543
g3723 nand P3_U4345 P3_U3265 ; P3_U5544
g3724 nand P3_U4340 P3_U5542 ; P3_U5545
g3725 nand P3_U5545 P3_U5544 ; P3_U5546
g3726 not P3_U3227 ; P3_U5547
g3727 not P3_U3225 ; P3_U5548
g3728 nand P3_U5534 P3_U5522 ; P3_U5549
g3729 nand P3_U5548 P3_U5523 P3_U2451 ; P3_U5550
g3730 nand P3_U5547 P3_U5549 ; P3_U5551
g3731 nand P3_ADD_495_U10 P3_U2356 ; P3_U5552
g3732 nand P3_U7982 P3_U7981 P3_U3679 ; P3_U5553
g3733 nand P3_U3286 P3_U3287 P3_STATE2_REG_1__SCAN_IN ; P3_U5554
g3734 nand P3_U4345 P3_U3225 ; P3_U5555
g3735 nand P3_U4340 P3_U5553 ; P3_U5556
g3736 nand P3_U3680 P3_U5556 ; P3_U5557
g3737 not P3_U3228 ; P3_U5558
g3738 nand P3_U4341 P3_U4608 ; P3_U5559
g3739 not P3_U3231 ; P3_U5560
g3740 not P3_U3230 ; P3_U5561
g3741 nand P3_U2466 P3_U3230 ; P3_U5562
g3742 nand P3_U5531 P3_U3094 ; P3_U5563
g3743 nand P3_U5558 P3_U3231 ; P3_U5564
g3744 nand P3_ADD_495_U4 P3_U2356 ; P3_U5565
g3745 nand P3_U5563 P3_U3681 ; P3_U5566
g3746 nand P3_U3286 P3_U7985 P3_STATE2_REG_1__SCAN_IN ; P3_U5567
g3747 nand P3_U5558 P3_U4345 ; P3_U5568
g3748 nand P3_U4340 P3_U5566 ; P3_U5569
g3749 nand P3_U3683 P3_U5569 ; P3_U5570
g3750 nand P3_U5560 P3_U5561 ; P3_U5571
g3751 nand P3_U2356 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U5572
g3752 nand P3_U7994 P3_U7993 P3_U5572 ; P3_U5573
g3753 nand P3_U4345 P3_U3093 ; P3_U5574
g3754 nand P3_U4340 P3_U5573 ; P3_U5575
g3755 nand P3_U7988 P3_STATE2_REG_1__SCAN_IN ; P3_U5576
g3756 nand P3_U3684 P3_U5575 ; P3_U5577
g3757 nand P3_U2453 P3_LT_589_U6 P3_STATE2_REG_0__SCAN_IN ; P3_U5578
g3758 not P3_U3233 ; P3_U5579
g3759 nand P3_U3132 P3_STATE2_REG_3__SCAN_IN ; P3_U5580
g3760 nand P3_U3233 P3_U5580 ; P3_U5581
g3761 nand P3_U4315 P3_U3123 ; P3_U5582
g3762 nand P3_U4647 P3_U3271 ; P3_U5583
g3763 nand P3_U3182 P3_U5583 ; P3_U5584
g3764 nand P3_U3183 P3_U5584 ; P3_U5585
g3765 nand P3_U4322 P3_U5585 ; P3_U5586
g3766 nand P3_U5582 P3_U3142 ; P3_U5587
g3767 nand P3_U4650 P3_STATE2_REG_3__SCAN_IN ; P3_U5588
g3768 nand P3_U3685 P3_U5586 ; P3_U5589
g3769 nand P3_U5589 P3_U3233 ; P3_U5590
g3770 nand P3_U5581 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_U5591
g3771 nand P3_U3131 P3_U4648 P3_STATE2_REG_3__SCAN_IN ; P3_U5592
g3772 nand P3_U4322 P3_U7999 ; P3_U5593
g3773 nand P3_U3270 P3_U5582 ; P3_U5594
g3774 nand P3_U3686 P3_U5593 ; P3_U5595
g3775 nand P3_U3130 P3_STATE2_REG_3__SCAN_IN ; P3_U5596
g3776 nand P3_U3233 P3_U5596 ; P3_U5597
g3777 nand P3_U5597 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U5598
g3778 nand P3_U5595 P3_U3233 ; P3_U5599
g3779 nand P3_U4322 P3_U3156 ; P3_U5600
g3780 nand P3_U3129 P3_STATE2_REG_3__SCAN_IN ; P3_U5601
g3781 nand P3_U5601 P3_U5600 ; P3_U5602
g3782 nand P3_U5602 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U5603
g3783 nand P3_U2493 P3_U4322 ; P3_U5604
g3784 nand P3_U5582 P3_U3141 ; P3_U5605
g3785 nand P3_U5605 P3_U5603 P3_U5604 ; P3_U5606
g3786 nand P3_U3128 P3_STATE2_REG_3__SCAN_IN ; P3_U5607
g3787 nand P3_U3233 P3_U5607 ; P3_U5608
g3788 nand P3_U5608 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_U5609
g3789 nand P3_U5606 P3_U3233 ; P3_U5610
g3790 not P3_U3234 ; P3_U5611
g3791 nand P3_U5611 P3_U3233 ; P3_U5612
g3792 nand P3_U3128 P3_STATE2_REG_3__SCAN_IN ; P3_U5613
g3793 nand P3_U4337 P3_U5613 ; P3_U5614
g3794 nand P3_U5614 P3_U3233 ; P3_U5615
g3795 nand P3_U5612 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_U5616
g3796 nand P3_U2463 P3_U4294 P3_GTE_450_U6 ; P3_U5617
g3797 nand P3_GTE_370_U6 P3_U4344 ; P3_U5618
g3798 nand P3_U5618 P3_U5617 ; P3_U5619
g3799 nand P3_U4590 P3_U2630 P3_GTE_412_U6 ; P3_U5620
g3800 nand P3_GTE_355_U6 P3_U3074 ; P3_U5621
g3801 nand P3_U5621 P3_U5620 ; P3_U5622
g3802 nand P3_GTE_390_U6 P3_U4488 ; P3_U5623
g3803 nand P3_U8001 P3_U8000 P3_U5623 ; P3_U5624
g3804 nand P3_U3102 P3_U3108 P3_GTE_401_U6 ; P3_U5625
g3805 nand P3_U4349 P3_GTE_504_U6 ; P3_U5626
g3806 nand P3_U4348 P3_GTE_485_U6 ; P3_U5627
g3807 nand P3_U4539 P3_U5624 ; P3_U5628
g3808 nand P3_U2515 P3_U5627 P3_U3687 P3_U5628 ; P3_U5629
g3809 nand P3_U2390 P3_U5629 ; P3_U5630
g3810 not P3_U3248 ; P3_U5631
g3811 nand P3_ADD_360_1242_U85 P3_U2395 ; P3_U5632
g3812 nand P3_SUB_357_1258_U69 P3_U2393 ; P3_U5633
g3813 nand P3_ADD_558_U5 P3_U3220 ; P3_U5634
g3814 nand P3_U4298 P3_ADD_553_U5 ; P3_U5635
g3815 nand P3_U4299 P3_ADD_547_U5 ; P3_U5636
g3816 nand P3_U4300 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5637
g3817 nand P3_U4301 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5638
g3818 nand P3_U2354 P3_ADD_531_U5 ; P3_U5639
g3819 nand P3_U2355 P3_ADD_526_U5 ; P3_U5640
g3820 nand P3_U4302 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5641
g3821 nand P3_U2356 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5642
g3822 nand P3_U4303 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5643
g3823 nand P3_U4304 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5644
g3824 nand P3_ADD_405_U4 P3_U4305 ; P3_U5645
g3825 nand P3_ADD_394_U4 P3_U2357 ; P3_U5646
g3826 nand P3_U2358 P3_ADD_385_U5 ; P3_U5647
g3827 nand P3_U2359 P3_ADD_380_U5 ; P3_U5648
g3828 nand P3_U4306 P3_ADD_349_U5 ; P3_U5649
g3829 nand P3_U2362 P3_ADD_344_U5 ; P3_U5650
g3830 nand P3_ADD_371_1212_U87 P3_U2360 ; P3_U5651
g3831 nand P3_U3692 P3_U5634 P3_U3693 P3_U3698 ; P3_U5652
g3832 nand P3_U2402 P3_REIP_REG_0__SCAN_IN ; P3_U5653
g3833 nand P3_U4318 P3_U5652 ; P3_U5654
g3834 nand P3_U5631 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U5655
g3835 nand P3_ADD_360_1242_U19 P3_U2395 ; P3_U5656
g3836 nand P3_SUB_357_1258_U21 P3_U2393 ; P3_U5657
g3837 nand P3_ADD_558_U85 P3_U3220 ; P3_U5658
g3838 nand P3_ADD_553_U85 P3_U4298 ; P3_U5659
g3839 nand P3_ADD_547_U85 P3_U4299 ; P3_U5660
g3840 nand P3_ADD_541_U4 P3_U4300 ; P3_U5661
g3841 nand P3_ADD_536_U4 P3_U4301 ; P3_U5662
g3842 nand P3_ADD_531_U85 P3_U2354 ; P3_U5663
g3843 nand P3_ADD_526_U71 P3_U2355 ; P3_U5664
g3844 nand P3_ADD_515_U4 P3_U4302 ; P3_U5665
g3845 nand P3_ADD_494_U4 P3_U2356 ; P3_U5666
g3846 nand P3_ADD_476_U4 P3_U4303 ; P3_U5667
g3847 nand P3_ADD_441_U4 P3_U4304 ; P3_U5668
g3848 nand P3_ADD_405_U81 P3_U4305 ; P3_U5669
g3849 nand P3_ADD_394_U81 P3_U2357 ; P3_U5670
g3850 nand P3_ADD_385_U85 P3_U2358 ; P3_U5671
g3851 nand P3_ADD_380_U85 P3_U2359 ; P3_U5672
g3852 nand P3_ADD_349_U85 P3_U4306 ; P3_U5673
g3853 nand P3_ADD_344_U85 P3_U2362 ; P3_U5674
g3854 nand P3_ADD_371_1212_U20 P3_U2360 ; P3_U5675
g3855 nand P3_U5658 P3_U3699 P3_U5656 P3_U3705 P3_U3700 ; P3_U5676
g3856 nand P3_U2402 P3_REIP_REG_1__SCAN_IN ; P3_U5677
g3857 nand P3_U4318 P3_U5676 ; P3_U5678
g3858 nand P3_U5631 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_U5679
g3859 nand P3_ADD_360_1242_U91 P3_U2395 ; P3_U5680
g3860 nand P3_SUB_357_1258_U78 P3_U2393 ; P3_U5681
g3861 nand P3_ADD_558_U74 P3_U3220 ; P3_U5682
g3862 nand P3_ADD_553_U74 P3_U4298 ; P3_U5683
g3863 nand P3_ADD_547_U74 P3_U4299 ; P3_U5684
g3864 nand P3_ADD_541_U71 P3_U4300 ; P3_U5685
g3865 nand P3_ADD_536_U71 P3_U4301 ; P3_U5686
g3866 nand P3_ADD_531_U74 P3_U2354 ; P3_U5687
g3867 nand P3_ADD_526_U60 P3_U2355 ; P3_U5688
g3868 nand P3_ADD_515_U71 P3_U4302 ; P3_U5689
g3869 nand P3_ADD_494_U71 P3_U2356 ; P3_U5690
g3870 nand P3_ADD_476_U71 P3_U4303 ; P3_U5691
g3871 nand P3_ADD_441_U71 P3_U4304 ; P3_U5692
g3872 nand P3_ADD_405_U5 P3_U4305 ; P3_U5693
g3873 nand P3_ADD_394_U5 P3_U2357 ; P3_U5694
g3874 nand P3_ADD_385_U74 P3_U2358 ; P3_U5695
g3875 nand P3_ADD_380_U74 P3_U2359 ; P3_U5696
g3876 nand P3_ADD_349_U74 P3_U4306 ; P3_U5697
g3877 nand P3_ADD_344_U74 P3_U2362 ; P3_U5698
g3878 nand P3_ADD_371_1212_U93 P3_U2360 ; P3_U5699
g3879 nand P3_U5682 P3_U3710 P3_U5680 P3_U3706 P3_U3713 ; P3_U5700
g3880 nand P3_U2402 P3_REIP_REG_2__SCAN_IN ; P3_U5701
g3881 nand P3_U4318 P3_U5700 ; P3_U5702
g3882 nand P3_U5631 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_U5703
g3883 nand P3_ADD_360_1242_U17 P3_U2395 ; P3_U5704
g3884 nand P3_SUB_357_1258_U76 P3_U2393 ; P3_U5705
g3885 nand P3_ADD_558_U71 P3_U3220 ; P3_U5706
g3886 nand P3_ADD_553_U71 P3_U4298 ; P3_U5707
g3887 nand P3_ADD_547_U71 P3_U4299 ; P3_U5708
g3888 nand P3_ADD_541_U68 P3_U4300 ; P3_U5709
g3889 nand P3_ADD_536_U68 P3_U4301 ; P3_U5710
g3890 nand P3_ADD_531_U71 P3_U2354 ; P3_U5711
g3891 nand P3_ADD_526_U57 P3_U2355 ; P3_U5712
g3892 nand P3_ADD_515_U68 P3_U4302 ; P3_U5713
g3893 nand P3_ADD_494_U68 P3_U2356 ; P3_U5714
g3894 nand P3_ADD_476_U68 P3_U4303 ; P3_U5715
g3895 nand P3_ADD_441_U68 P3_U4304 ; P3_U5716
g3896 nand P3_ADD_405_U93 P3_U4305 ; P3_U5717
g3897 nand P3_ADD_394_U93 P3_U2357 ; P3_U5718
g3898 nand P3_ADD_385_U71 P3_U2358 ; P3_U5719
g3899 nand P3_ADD_380_U71 P3_U2359 ; P3_U5720
g3900 nand P3_ADD_349_U71 P3_U4306 ; P3_U5721
g3901 nand P3_ADD_344_U71 P3_U2362 ; P3_U5722
g3902 nand P3_ADD_371_1212_U18 P3_U2360 ; P3_U5723
g3903 nand P3_U3715 P3_U5706 P3_U3718 P3_U3714 P3_U3721 ; P3_U5724
g3904 nand P3_U2402 P3_REIP_REG_3__SCAN_IN ; P3_U5725
g3905 nand P3_U4318 P3_U5724 ; P3_U5726
g3906 nand P3_U5631 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_U5727
g3907 nand P3_ADD_360_1242_U18 P3_U2395 ; P3_U5728
g3908 nand P3_SUB_357_1258_U75 P3_U2393 ; P3_U5729
g3909 nand P3_ADD_558_U70 P3_U3220 ; P3_U5730
g3910 nand P3_ADD_553_U70 P3_U4298 ; P3_U5731
g3911 nand P3_ADD_547_U70 P3_U4299 ; P3_U5732
g3912 nand P3_ADD_541_U67 P3_U4300 ; P3_U5733
g3913 nand P3_ADD_536_U67 P3_U4301 ; P3_U5734
g3914 nand P3_ADD_531_U70 P3_U2354 ; P3_U5735
g3915 nand P3_ADD_526_U56 P3_U2355 ; P3_U5736
g3916 nand P3_ADD_515_U67 P3_U4302 ; P3_U5737
g3917 nand P3_ADD_494_U67 P3_U2356 ; P3_U5738
g3918 nand P3_ADD_476_U67 P3_U4303 ; P3_U5739
g3919 nand P3_ADD_441_U67 P3_U4304 ; P3_U5740
g3920 nand P3_ADD_405_U68 P3_U4305 ; P3_U5741
g3921 nand P3_ADD_394_U68 P3_U2357 ; P3_U5742
g3922 nand P3_ADD_385_U70 P3_U2358 ; P3_U5743
g3923 nand P3_ADD_380_U70 P3_U2359 ; P3_U5744
g3924 nand P3_ADD_349_U70 P3_U4306 ; P3_U5745
g3925 nand P3_ADD_344_U70 P3_U2362 ; P3_U5746
g3926 nand P3_ADD_371_1212_U91 P3_U2360 ; P3_U5747
g3927 nand P3_U5730 P3_U3726 P3_U5728 P3_U3722 P3_U3729 ; P3_U5748
g3928 nand P3_U2402 P3_REIP_REG_4__SCAN_IN ; P3_U5749
g3929 nand P3_U4318 P3_U5748 ; P3_U5750
g3930 nand P3_U5631 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_U5751
g3931 nand P3_ADD_360_1242_U89 P3_U2395 ; P3_U5752
g3932 nand P3_SUB_357_1258_U74 P3_U2393 ; P3_U5753
g3933 nand P3_ADD_558_U69 P3_U3220 ; P3_U5754
g3934 nand P3_ADD_553_U69 P3_U4298 ; P3_U5755
g3935 nand P3_ADD_547_U69 P3_U4299 ; P3_U5756
g3936 nand P3_ADD_541_U66 P3_U4300 ; P3_U5757
g3937 nand P3_ADD_536_U66 P3_U4301 ; P3_U5758
g3938 nand P3_ADD_531_U69 P3_U2354 ; P3_U5759
g3939 nand P3_ADD_526_U55 P3_U2355 ; P3_U5760
g3940 nand P3_ADD_515_U66 P3_U4302 ; P3_U5761
g3941 nand P3_ADD_494_U66 P3_U2356 ; P3_U5762
g3942 nand P3_ADD_476_U66 P3_U4303 ; P3_U5763
g3943 nand P3_ADD_441_U66 P3_U4304 ; P3_U5764
g3944 nand P3_ADD_405_U67 P3_U4305 ; P3_U5765
g3945 nand P3_ADD_394_U67 P3_U2357 ; P3_U5766
g3946 nand P3_ADD_385_U69 P3_U2358 ; P3_U5767
g3947 nand P3_ADD_380_U69 P3_U2359 ; P3_U5768
g3948 nand P3_ADD_349_U69 P3_U4306 ; P3_U5769
g3949 nand P3_ADD_344_U69 P3_U2362 ; P3_U5770
g3950 nand P3_ADD_371_1212_U19 P3_U2360 ; P3_U5771
g3951 nand P3_U3734 P3_U5754 P3_U5753 P3_U3730 P3_U3737 ; P3_U5772
g3952 nand P3_U2402 P3_REIP_REG_5__SCAN_IN ; P3_U5773
g3953 nand P3_U4318 P3_U5772 ; P3_U5774
g3954 nand P3_U5631 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_U5775
g3955 nand P3_ADD_360_1242_U88 P3_U2395 ; P3_U5776
g3956 nand P3_SUB_357_1258_U73 P3_U2393 ; P3_U5777
g3957 nand P3_ADD_558_U68 P3_U3220 ; P3_U5778
g3958 nand P3_ADD_553_U68 P3_U4298 ; P3_U5779
g3959 nand P3_ADD_547_U68 P3_U4299 ; P3_U5780
g3960 nand P3_ADD_541_U65 P3_U4300 ; P3_U5781
g3961 nand P3_ADD_536_U65 P3_U4301 ; P3_U5782
g3962 nand P3_ADD_531_U68 P3_U2354 ; P3_U5783
g3963 nand P3_ADD_526_U54 P3_U2355 ; P3_U5784
g3964 nand P3_ADD_515_U65 P3_U4302 ; P3_U5785
g3965 nand P3_ADD_494_U65 P3_U2356 ; P3_U5786
g3966 nand P3_ADD_476_U65 P3_U4303 ; P3_U5787
g3967 nand P3_ADD_441_U65 P3_U4304 ; P3_U5788
g3968 nand P3_ADD_405_U66 P3_U4305 ; P3_U5789
g3969 nand P3_ADD_394_U66 P3_U2357 ; P3_U5790
g3970 nand P3_ADD_385_U68 P3_U2358 ; P3_U5791
g3971 nand P3_ADD_380_U68 P3_U2359 ; P3_U5792
g3972 nand P3_ADD_349_U68 P3_U4306 ; P3_U5793
g3973 nand P3_ADD_344_U68 P3_U2362 ; P3_U5794
g3974 nand P3_ADD_371_1212_U90 P3_U2360 ; P3_U5795
g3975 nand P3_U3742 P3_U5778 P3_U5777 P3_U3738 P3_U3745 ; P3_U5796
g3976 nand P3_U2402 P3_REIP_REG_6__SCAN_IN ; P3_U5797
g3977 nand P3_U4318 P3_U5796 ; P3_U5798
g3978 nand P3_U5631 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_U5799
g3979 nand P3_ADD_360_1242_U87 P3_U2395 ; P3_U5800
g3980 nand P3_SUB_357_1258_U72 P3_U2393 ; P3_U5801
g3981 nand P3_ADD_558_U67 P3_U3220 ; P3_U5802
g3982 nand P3_ADD_553_U67 P3_U4298 ; P3_U5803
g3983 nand P3_ADD_547_U67 P3_U4299 ; P3_U5804
g3984 nand P3_ADD_541_U64 P3_U4300 ; P3_U5805
g3985 nand P3_ADD_536_U64 P3_U4301 ; P3_U5806
g3986 nand P3_ADD_531_U67 P3_U2354 ; P3_U5807
g3987 nand P3_ADD_526_U53 P3_U2355 ; P3_U5808
g3988 nand P3_ADD_515_U64 P3_U4302 ; P3_U5809
g3989 nand P3_ADD_494_U64 P3_U2356 ; P3_U5810
g3990 nand P3_ADD_476_U64 P3_U4303 ; P3_U5811
g3991 nand P3_ADD_441_U64 P3_U4304 ; P3_U5812
g3992 nand P3_ADD_405_U65 P3_U4305 ; P3_U5813
g3993 nand P3_ADD_394_U65 P3_U2357 ; P3_U5814
g3994 nand P3_ADD_385_U67 P3_U2358 ; P3_U5815
g3995 nand P3_ADD_380_U67 P3_U2359 ; P3_U5816
g3996 nand P3_ADD_349_U67 P3_U4306 ; P3_U5817
g3997 nand P3_ADD_344_U67 P3_U2362 ; P3_U5818
g3998 nand P3_ADD_371_1212_U89 P3_U2360 ; P3_U5819
g3999 nand P3_U3750 P3_U5802 P3_U5801 P3_U3746 P3_U3753 ; P3_U5820
g4000 nand P3_U2402 P3_REIP_REG_7__SCAN_IN ; P3_U5821
g4001 nand P3_U4318 P3_U5820 ; P3_U5822
g4002 nand P3_U5631 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_U5823
g4003 nand P3_ADD_360_1242_U86 P3_U2395 ; P3_U5824
g4004 nand P3_SUB_357_1258_U71 P3_U2393 ; P3_U5825
g4005 nand P3_ADD_558_U66 P3_U3220 ; P3_U5826
g4006 nand P3_ADD_553_U66 P3_U4298 ; P3_U5827
g4007 nand P3_ADD_547_U66 P3_U4299 ; P3_U5828
g4008 nand P3_ADD_541_U63 P3_U4300 ; P3_U5829
g4009 nand P3_ADD_536_U63 P3_U4301 ; P3_U5830
g4010 nand P3_ADD_531_U66 P3_U2354 ; P3_U5831
g4011 nand P3_ADD_526_U52 P3_U2355 ; P3_U5832
g4012 nand P3_ADD_515_U63 P3_U4302 ; P3_U5833
g4013 nand P3_ADD_494_U63 P3_U2356 ; P3_U5834
g4014 nand P3_ADD_476_U63 P3_U4303 ; P3_U5835
g4015 nand P3_ADD_441_U63 P3_U4304 ; P3_U5836
g4016 nand P3_ADD_405_U64 P3_U4305 ; P3_U5837
g4017 nand P3_ADD_394_U64 P3_U2357 ; P3_U5838
g4018 nand P3_ADD_385_U66 P3_U2358 ; P3_U5839
g4019 nand P3_ADD_380_U66 P3_U2359 ; P3_U5840
g4020 nand P3_ADD_349_U66 P3_U4306 ; P3_U5841
g4021 nand P3_ADD_344_U66 P3_U2362 ; P3_U5842
g4022 nand P3_ADD_371_1212_U88 P3_U2360 ; P3_U5843
g4023 nand P3_U3757 P3_U5826 P3_U5825 P3_U3754 P3_U3760 ; P3_U5844
g4024 nand P3_U2402 P3_REIP_REG_8__SCAN_IN ; P3_U5845
g4025 nand P3_U4318 P3_U5844 ; P3_U5846
g4026 nand P3_U5631 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_U5847
g4027 nand P3_ADD_360_1242_U106 P3_U2395 ; P3_U5848
g4028 nand P3_SUB_357_1258_U70 P3_U2393 ; P3_U5849
g4029 nand P3_ADD_558_U65 P3_U3220 ; P3_U5850
g4030 nand P3_ADD_553_U65 P3_U4298 ; P3_U5851
g4031 nand P3_ADD_547_U65 P3_U4299 ; P3_U5852
g4032 nand P3_ADD_541_U62 P3_U4300 ; P3_U5853
g4033 nand P3_ADD_536_U62 P3_U4301 ; P3_U5854
g4034 nand P3_ADD_531_U65 P3_U2354 ; P3_U5855
g4035 nand P3_ADD_526_U51 P3_U2355 ; P3_U5856
g4036 nand P3_ADD_515_U62 P3_U4302 ; P3_U5857
g4037 nand P3_ADD_494_U62 P3_U2356 ; P3_U5858
g4038 nand P3_ADD_476_U62 P3_U4303 ; P3_U5859
g4039 nand P3_ADD_441_U62 P3_U4304 ; P3_U5860
g4040 nand P3_ADD_405_U63 P3_U4305 ; P3_U5861
g4041 nand P3_ADD_394_U63 P3_U2357 ; P3_U5862
g4042 nand P3_ADD_385_U65 P3_U2358 ; P3_U5863
g4043 nand P3_ADD_380_U65 P3_U2359 ; P3_U5864
g4044 nand P3_ADD_349_U65 P3_U4306 ; P3_U5865
g4045 nand P3_ADD_344_U65 P3_U2362 ; P3_U5866
g4046 nand P3_ADD_371_1212_U109 P3_U2360 ; P3_U5867
g4047 nand P3_U3764 P3_U5850 P3_U5849 P3_U3761 P3_U3767 ; P3_U5868
g4048 nand P3_U2402 P3_REIP_REG_9__SCAN_IN ; P3_U5869
g4049 nand P3_U4318 P3_U5868 ; P3_U5870
g4050 nand P3_U5631 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_U5871
g4051 nand P3_ADD_360_1242_U4 P3_U2395 ; P3_U5872
g4052 nand P3_SUB_357_1258_U93 P3_U2393 ; P3_U5873
g4053 nand P3_ADD_558_U95 P3_U3220 ; P3_U5874
g4054 nand P3_ADD_553_U95 P3_U4298 ; P3_U5875
g4055 nand P3_ADD_547_U95 P3_U4299 ; P3_U5876
g4056 nand P3_ADD_541_U91 P3_U4300 ; P3_U5877
g4057 nand P3_ADD_536_U91 P3_U4301 ; P3_U5878
g4058 nand P3_ADD_531_U95 P3_U2354 ; P3_U5879
g4059 nand P3_ADD_526_U81 P3_U2355 ; P3_U5880
g4060 nand P3_ADD_515_U91 P3_U4302 ; P3_U5881
g4061 nand P3_ADD_494_U91 P3_U2356 ; P3_U5882
g4062 nand P3_ADD_476_U91 P3_U4303 ; P3_U5883
g4063 nand P3_ADD_441_U91 P3_U4304 ; P3_U5884
g4064 nand P3_ADD_405_U91 P3_U4305 ; P3_U5885
g4065 nand P3_ADD_394_U91 P3_U2357 ; P3_U5886
g4066 nand P3_ADD_385_U95 P3_U2358 ; P3_U5887
g4067 nand P3_ADD_380_U95 P3_U2359 ; P3_U5888
g4068 nand P3_ADD_349_U95 P3_U4306 ; P3_U5889
g4069 nand P3_ADD_344_U95 P3_U2362 ; P3_U5890
g4070 nand P3_ADD_371_1212_U5 P3_U2360 ; P3_U5891
g4071 nand P3_U5874 P3_U3771 P3_U5872 P3_U3774 P3_U3768 ; P3_U5892
g4072 nand P3_U2402 P3_REIP_REG_10__SCAN_IN ; P3_U5893
g4073 nand P3_U4318 P3_U5892 ; P3_U5894
g4074 nand P3_U5631 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_U5895
g4075 nand P3_ADD_360_1242_U84 P3_U2395 ; P3_U5896
g4076 nand P3_SUB_357_1258_U92 P3_U2393 ; P3_U5897
g4077 nand P3_ADD_558_U94 P3_U3220 ; P3_U5898
g4078 nand P3_ADD_553_U94 P3_U4298 ; P3_U5899
g4079 nand P3_ADD_547_U94 P3_U4299 ; P3_U5900
g4080 nand P3_ADD_541_U90 P3_U4300 ; P3_U5901
g4081 nand P3_ADD_536_U90 P3_U4301 ; P3_U5902
g4082 nand P3_ADD_531_U94 P3_U2354 ; P3_U5903
g4083 nand P3_ADD_526_U80 P3_U2355 ; P3_U5904
g4084 nand P3_ADD_515_U90 P3_U4302 ; P3_U5905
g4085 nand P3_ADD_494_U90 P3_U2356 ; P3_U5906
g4086 nand P3_ADD_476_U90 P3_U4303 ; P3_U5907
g4087 nand P3_ADD_441_U90 P3_U4304 ; P3_U5908
g4088 nand P3_ADD_405_U90 P3_U4305 ; P3_U5909
g4089 nand P3_ADD_394_U90 P3_U2357 ; P3_U5910
g4090 nand P3_ADD_385_U94 P3_U2358 ; P3_U5911
g4091 nand P3_ADD_380_U94 P3_U2359 ; P3_U5912
g4092 nand P3_ADD_349_U94 P3_U4306 ; P3_U5913
g4093 nand P3_ADD_344_U94 P3_U2362 ; P3_U5914
g4094 nand P3_ADD_371_1212_U86 P3_U2360 ; P3_U5915
g4095 nand P3_U5898 P3_U3778 P3_U5896 P3_U3775 P3_U3781 ; P3_U5916
g4096 nand P3_U2402 P3_REIP_REG_11__SCAN_IN ; P3_U5917
g4097 nand P3_U4318 P3_U5916 ; P3_U5918
g4098 nand P3_U5631 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_U5919
g4099 nand P3_ADD_360_1242_U5 P3_U2395 ; P3_U5920
g4100 nand P3_SUB_357_1258_U91 P3_U2393 ; P3_U5921
g4101 nand P3_ADD_558_U93 P3_U3220 ; P3_U5922
g4102 nand P3_ADD_553_U93 P3_U4298 ; P3_U5923
g4103 nand P3_ADD_547_U93 P3_U4299 ; P3_U5924
g4104 nand P3_ADD_541_U89 P3_U4300 ; P3_U5925
g4105 nand P3_ADD_536_U89 P3_U4301 ; P3_U5926
g4106 nand P3_ADD_531_U93 P3_U2354 ; P3_U5927
g4107 nand P3_ADD_526_U79 P3_U2355 ; P3_U5928
g4108 nand P3_ADD_515_U89 P3_U4302 ; P3_U5929
g4109 nand P3_ADD_494_U89 P3_U2356 ; P3_U5930
g4110 nand P3_ADD_476_U89 P3_U4303 ; P3_U5931
g4111 nand P3_ADD_441_U89 P3_U4304 ; P3_U5932
g4112 nand P3_ADD_405_U89 P3_U4305 ; P3_U5933
g4113 nand P3_ADD_394_U89 P3_U2357 ; P3_U5934
g4114 nand P3_ADD_385_U93 P3_U2358 ; P3_U5935
g4115 nand P3_ADD_380_U93 P3_U2359 ; P3_U5936
g4116 nand P3_ADD_349_U93 P3_U4306 ; P3_U5937
g4117 nand P3_ADD_344_U93 P3_U2362 ; P3_U5938
g4118 nand P3_ADD_371_1212_U6 P3_U2360 ; P3_U5939
g4119 nand P3_U3785 P3_U5922 P3_U5921 P3_U3782 P3_U3788 ; P3_U5940
g4120 nand P3_U2402 P3_REIP_REG_12__SCAN_IN ; P3_U5941
g4121 nand P3_U4318 P3_U5940 ; P3_U5942
g4122 nand P3_U5631 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_U5943
g4123 nand P3_ADD_360_1242_U6 P3_U2395 ; P3_U5944
g4124 nand P3_SUB_357_1258_U15 P3_U2393 ; P3_U5945
g4125 nand P3_ADD_558_U92 P3_U3220 ; P3_U5946
g4126 nand P3_ADD_553_U92 P3_U4298 ; P3_U5947
g4127 nand P3_ADD_547_U92 P3_U4299 ; P3_U5948
g4128 nand P3_ADD_541_U88 P3_U4300 ; P3_U5949
g4129 nand P3_ADD_536_U88 P3_U4301 ; P3_U5950
g4130 nand P3_ADD_531_U92 P3_U2354 ; P3_U5951
g4131 nand P3_ADD_526_U78 P3_U2355 ; P3_U5952
g4132 nand P3_ADD_515_U88 P3_U4302 ; P3_U5953
g4133 nand P3_ADD_494_U88 P3_U2356 ; P3_U5954
g4134 nand P3_ADD_476_U88 P3_U4303 ; P3_U5955
g4135 nand P3_ADD_441_U88 P3_U4304 ; P3_U5956
g4136 nand P3_ADD_405_U88 P3_U4305 ; P3_U5957
g4137 nand P3_ADD_394_U88 P3_U2357 ; P3_U5958
g4138 nand P3_ADD_385_U92 P3_U2358 ; P3_U5959
g4139 nand P3_ADD_380_U92 P3_U2359 ; P3_U5960
g4140 nand P3_ADD_349_U92 P3_U4306 ; P3_U5961
g4141 nand P3_ADD_344_U92 P3_U2362 ; P3_U5962
g4142 nand P3_ADD_371_1212_U7 P3_U2360 ; P3_U5963
g4143 nand P3_U3792 P3_U5946 P3_U5945 P3_U3789 P3_U3795 ; P3_U5964
g4144 nand P3_U2402 P3_REIP_REG_13__SCAN_IN ; P3_U5965
g4145 nand P3_U4318 P3_U5964 ; P3_U5966
g4146 nand P3_U5631 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_U5967
g4147 nand P3_ADD_360_1242_U83 P3_U2395 ; P3_U5968
g4148 nand P3_SUB_357_1258_U90 P3_U2393 ; P3_U5969
g4149 nand P3_ADD_558_U91 P3_U3220 ; P3_U5970
g4150 nand P3_ADD_553_U91 P3_U4298 ; P3_U5971
g4151 nand P3_ADD_547_U91 P3_U4299 ; P3_U5972
g4152 nand P3_ADD_541_U87 P3_U4300 ; P3_U5973
g4153 nand P3_ADD_536_U87 P3_U4301 ; P3_U5974
g4154 nand P3_ADD_531_U91 P3_U2354 ; P3_U5975
g4155 nand P3_ADD_526_U77 P3_U2355 ; P3_U5976
g4156 nand P3_ADD_515_U87 P3_U4302 ; P3_U5977
g4157 nand P3_ADD_494_U87 P3_U2356 ; P3_U5978
g4158 nand P3_ADD_476_U87 P3_U4303 ; P3_U5979
g4159 nand P3_ADD_441_U87 P3_U4304 ; P3_U5980
g4160 nand P3_ADD_405_U87 P3_U4305 ; P3_U5981
g4161 nand P3_ADD_394_U87 P3_U2357 ; P3_U5982
g4162 nand P3_ADD_385_U91 P3_U2358 ; P3_U5983
g4163 nand P3_ADD_380_U91 P3_U2359 ; P3_U5984
g4164 nand P3_ADD_349_U91 P3_U4306 ; P3_U5985
g4165 nand P3_ADD_344_U91 P3_U2362 ; P3_U5986
g4166 nand P3_ADD_371_1212_U85 P3_U2360 ; P3_U5987
g4167 nand P3_U3802 P3_U3799 ; P3_U5988
g4168 nand P3_U2402 P3_REIP_REG_14__SCAN_IN ; P3_U5989
g4169 nand P3_U4318 P3_U5988 ; P3_U5990
g4170 nand P3_U5631 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_U5991
g4171 nand P3_ADD_360_1242_U7 P3_U2395 ; P3_U5992
g4172 nand P3_SUB_357_1258_U89 P3_U2393 ; P3_U5993
g4173 nand P3_ADD_558_U90 P3_U3220 ; P3_U5994
g4174 nand P3_ADD_553_U90 P3_U4298 ; P3_U5995
g4175 nand P3_ADD_547_U90 P3_U4299 ; P3_U5996
g4176 nand P3_ADD_541_U86 P3_U4300 ; P3_U5997
g4177 nand P3_ADD_536_U86 P3_U4301 ; P3_U5998
g4178 nand P3_ADD_531_U90 P3_U2354 ; P3_U5999
g4179 nand P3_ADD_526_U76 P3_U2355 ; P3_U6000
g4180 nand P3_ADD_515_U86 P3_U4302 ; P3_U6001
g4181 nand P3_ADD_494_U86 P3_U2356 ; P3_U6002
g4182 nand P3_ADD_476_U86 P3_U4303 ; P3_U6003
g4183 nand P3_ADD_441_U86 P3_U4304 ; P3_U6004
g4184 nand P3_ADD_405_U86 P3_U4305 ; P3_U6005
g4185 nand P3_ADD_394_U86 P3_U2357 ; P3_U6006
g4186 nand P3_ADD_385_U90 P3_U2358 ; P3_U6007
g4187 nand P3_ADD_380_U90 P3_U2359 ; P3_U6008
g4188 nand P3_ADD_349_U90 P3_U4306 ; P3_U6009
g4189 nand P3_ADD_344_U90 P3_U2362 ; P3_U6010
g4190 nand P3_ADD_371_1212_U8 P3_U2360 ; P3_U6011
g4191 nand P3_U3810 P3_U3807 ; P3_U6012
g4192 nand P3_U2402 P3_REIP_REG_15__SCAN_IN ; P3_U6013
g4193 nand P3_U4318 P3_U6012 ; P3_U6014
g4194 nand P3_U5631 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_U6015
g4195 nand P3_ADD_360_1242_U82 P3_U2395 ; P3_U6016
g4196 nand P3_SUB_357_1258_U88 P3_U2393 ; P3_U6017
g4197 nand P3_ADD_558_U89 P3_U3220 ; P3_U6018
g4198 nand P3_ADD_553_U89 P3_U4298 ; P3_U6019
g4199 nand P3_ADD_547_U89 P3_U4299 ; P3_U6020
g4200 nand P3_ADD_541_U85 P3_U4300 ; P3_U6021
g4201 nand P3_ADD_536_U85 P3_U4301 ; P3_U6022
g4202 nand P3_ADD_531_U89 P3_U2354 ; P3_U6023
g4203 nand P3_ADD_526_U75 P3_U2355 ; P3_U6024
g4204 nand P3_ADD_515_U85 P3_U4302 ; P3_U6025
g4205 nand P3_ADD_494_U85 P3_U2356 ; P3_U6026
g4206 nand P3_ADD_476_U85 P3_U4303 ; P3_U6027
g4207 nand P3_ADD_441_U85 P3_U4304 ; P3_U6028
g4208 nand P3_ADD_405_U85 P3_U4305 ; P3_U6029
g4209 nand P3_ADD_394_U85 P3_U2357 ; P3_U6030
g4210 nand P3_ADD_385_U89 P3_U2358 ; P3_U6031
g4211 nand P3_ADD_380_U89 P3_U2359 ; P3_U6032
g4212 nand P3_ADD_349_U89 P3_U4306 ; P3_U6033
g4213 nand P3_ADD_344_U89 P3_U2362 ; P3_U6034
g4214 nand P3_ADD_371_1212_U84 P3_U2360 ; P3_U6035
g4215 nand P3_U6018 P3_U3815 P3_U6016 P3_U3812 P3_U3818 ; P3_U6036
g4216 nand P3_U2402 P3_REIP_REG_16__SCAN_IN ; P3_U6037
g4217 nand P3_U4318 P3_U6036 ; P3_U6038
g4218 nand P3_U5631 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_U6039
g4219 nand P3_ADD_360_1242_U8 P3_U2395 ; P3_U6040
g4220 nand P3_SUB_357_1258_U16 P3_U2393 ; P3_U6041
g4221 nand P3_ADD_558_U88 P3_U3220 ; P3_U6042
g4222 nand P3_ADD_553_U88 P3_U4298 ; P3_U6043
g4223 nand P3_ADD_547_U88 P3_U4299 ; P3_U6044
g4224 nand P3_ADD_541_U84 P3_U4300 ; P3_U6045
g4225 nand P3_ADD_536_U84 P3_U4301 ; P3_U6046
g4226 nand P3_ADD_531_U88 P3_U2354 ; P3_U6047
g4227 nand P3_ADD_526_U74 P3_U2355 ; P3_U6048
g4228 nand P3_ADD_515_U84 P3_U4302 ; P3_U6049
g4229 nand P3_ADD_494_U84 P3_U2356 ; P3_U6050
g4230 nand P3_ADD_476_U84 P3_U4303 ; P3_U6051
g4231 nand P3_ADD_441_U84 P3_U4304 ; P3_U6052
g4232 nand P3_ADD_405_U84 P3_U4305 ; P3_U6053
g4233 nand P3_ADD_394_U84 P3_U2357 ; P3_U6054
g4234 nand P3_ADD_385_U88 P3_U2358 ; P3_U6055
g4235 nand P3_ADD_380_U88 P3_U2359 ; P3_U6056
g4236 nand P3_ADD_349_U88 P3_U4306 ; P3_U6057
g4237 nand P3_ADD_344_U88 P3_U2362 ; P3_U6058
g4238 nand P3_ADD_371_1212_U9 P3_U2360 ; P3_U6059
g4239 nand P3_U6042 P3_U3819 P3_U6040 P3_U3824 P3_U3820 ; P3_U6060
g4240 nand P3_U2402 P3_REIP_REG_17__SCAN_IN ; P3_U6061
g4241 nand P3_U4318 P3_U6060 ; P3_U6062
g4242 nand P3_U5631 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_U6063
g4243 nand P3_ADD_360_1242_U81 P3_U2395 ; P3_U6064
g4244 nand P3_SUB_357_1258_U87 P3_U2393 ; P3_U6065
g4245 nand P3_ADD_558_U87 P3_U3220 ; P3_U6066
g4246 nand P3_ADD_553_U87 P3_U4298 ; P3_U6067
g4247 nand P3_ADD_547_U87 P3_U4299 ; P3_U6068
g4248 nand P3_ADD_541_U83 P3_U4300 ; P3_U6069
g4249 nand P3_ADD_536_U83 P3_U4301 ; P3_U6070
g4250 nand P3_ADD_531_U87 P3_U2354 ; P3_U6071
g4251 nand P3_ADD_526_U73 P3_U2355 ; P3_U6072
g4252 nand P3_ADD_515_U83 P3_U4302 ; P3_U6073
g4253 nand P3_ADD_494_U83 P3_U2356 ; P3_U6074
g4254 nand P3_ADD_476_U83 P3_U4303 ; P3_U6075
g4255 nand P3_ADD_441_U83 P3_U4304 ; P3_U6076
g4256 nand P3_ADD_405_U83 P3_U4305 ; P3_U6077
g4257 nand P3_ADD_394_U83 P3_U2357 ; P3_U6078
g4258 nand P3_ADD_385_U87 P3_U2358 ; P3_U6079
g4259 nand P3_ADD_380_U87 P3_U2359 ; P3_U6080
g4260 nand P3_ADD_349_U87 P3_U4306 ; P3_U6081
g4261 nand P3_ADD_344_U87 P3_U2362 ; P3_U6082
g4262 nand P3_ADD_371_1212_U83 P3_U2360 ; P3_U6083
g4263 nand P3_U6066 P3_U3828 P3_U6064 P3_U3825 P3_U3831 ; P3_U6084
g4264 nand P3_U2402 P3_REIP_REG_18__SCAN_IN ; P3_U6085
g4265 nand P3_U4318 P3_U6084 ; P3_U6086
g4266 nand P3_U5631 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_U6087
g4267 nand P3_ADD_360_1242_U9 P3_U2395 ; P3_U6088
g4268 nand P3_SUB_357_1258_U86 P3_U2393 ; P3_U6089
g4269 nand P3_ADD_558_U86 P3_U3220 ; P3_U6090
g4270 nand P3_ADD_553_U86 P3_U4298 ; P3_U6091
g4271 nand P3_ADD_547_U86 P3_U4299 ; P3_U6092
g4272 nand P3_ADD_541_U82 P3_U4300 ; P3_U6093
g4273 nand P3_ADD_536_U82 P3_U4301 ; P3_U6094
g4274 nand P3_ADD_531_U86 P3_U2354 ; P3_U6095
g4275 nand P3_ADD_526_U72 P3_U2355 ; P3_U6096
g4276 nand P3_ADD_515_U82 P3_U4302 ; P3_U6097
g4277 nand P3_ADD_494_U82 P3_U2356 ; P3_U6098
g4278 nand P3_ADD_476_U82 P3_U4303 ; P3_U6099
g4279 nand P3_ADD_441_U82 P3_U4304 ; P3_U6100
g4280 nand P3_ADD_405_U82 P3_U4305 ; P3_U6101
g4281 nand P3_ADD_394_U82 P3_U2357 ; P3_U6102
g4282 nand P3_ADD_385_U86 P3_U2358 ; P3_U6103
g4283 nand P3_ADD_380_U86 P3_U2359 ; P3_U6104
g4284 nand P3_ADD_349_U86 P3_U4306 ; P3_U6105
g4285 nand P3_ADD_344_U86 P3_U2362 ; P3_U6106
g4286 nand P3_ADD_371_1212_U10 P3_U2360 ; P3_U6107
g4287 nand P3_U6090 P3_U3832 P3_U6088 P3_U3837 P3_U3833 ; P3_U6108
g4288 nand P3_U2402 P3_REIP_REG_19__SCAN_IN ; P3_U6109
g4289 nand P3_U4318 P3_U6108 ; P3_U6110
g4290 nand P3_U5631 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_U6111
g4291 nand P3_ADD_360_1242_U10 P3_U2395 ; P3_U6112
g4292 nand P3_SUB_357_1258_U17 P3_U2393 ; P3_U6113
g4293 nand P3_ADD_558_U84 P3_U3220 ; P3_U6114
g4294 nand P3_ADD_553_U84 P3_U4298 ; P3_U6115
g4295 nand P3_ADD_547_U84 P3_U4299 ; P3_U6116
g4296 nand P3_ADD_541_U81 P3_U4300 ; P3_U6117
g4297 nand P3_ADD_536_U81 P3_U4301 ; P3_U6118
g4298 nand P3_ADD_531_U84 P3_U2354 ; P3_U6119
g4299 nand P3_ADD_526_U70 P3_U2355 ; P3_U6120
g4300 nand P3_ADD_515_U81 P3_U4302 ; P3_U6121
g4301 nand P3_ADD_494_U81 P3_U2356 ; P3_U6122
g4302 nand P3_ADD_476_U81 P3_U4303 ; P3_U6123
g4303 nand P3_ADD_441_U81 P3_U4304 ; P3_U6124
g4304 nand P3_ADD_405_U80 P3_U4305 ; P3_U6125
g4305 nand P3_ADD_394_U80 P3_U2357 ; P3_U6126
g4306 nand P3_ADD_385_U84 P3_U2358 ; P3_U6127
g4307 nand P3_ADD_380_U84 P3_U2359 ; P3_U6128
g4308 nand P3_ADD_349_U84 P3_U4306 ; P3_U6129
g4309 nand P3_ADD_344_U84 P3_U2362 ; P3_U6130
g4310 nand P3_ADD_371_1212_U11 P3_U2360 ; P3_U6131
g4311 nand P3_U6113 P3_U3841 ; P3_U6132
g4312 nand P3_U2402 P3_REIP_REG_20__SCAN_IN ; P3_U6133
g4313 nand P3_U4318 P3_U6132 ; P3_U6134
g4314 nand P3_U5631 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_U6135
g4315 nand P3_ADD_360_1242_U11 P3_U2395 ; P3_U6136
g4316 nand P3_SUB_357_1258_U85 P3_U2393 ; P3_U6137
g4317 nand P3_ADD_558_U83 P3_U3220 ; P3_U6138
g4318 nand P3_ADD_553_U83 P3_U4298 ; P3_U6139
g4319 nand P3_ADD_547_U83 P3_U4299 ; P3_U6140
g4320 nand P3_ADD_541_U80 P3_U4300 ; P3_U6141
g4321 nand P3_ADD_536_U80 P3_U4301 ; P3_U6142
g4322 nand P3_ADD_531_U83 P3_U2354 ; P3_U6143
g4323 nand P3_ADD_526_U69 P3_U2355 ; P3_U6144
g4324 nand P3_ADD_515_U80 P3_U4302 ; P3_U6145
g4325 nand P3_ADD_494_U80 P3_U2356 ; P3_U6146
g4326 nand P3_ADD_476_U80 P3_U4303 ; P3_U6147
g4327 nand P3_ADD_441_U80 P3_U4304 ; P3_U6148
g4328 nand P3_ADD_405_U79 P3_U4305 ; P3_U6149
g4329 nand P3_ADD_394_U79 P3_U2357 ; P3_U6150
g4330 nand P3_ADD_385_U83 P3_U2358 ; P3_U6151
g4331 nand P3_ADD_380_U83 P3_U2359 ; P3_U6152
g4332 nand P3_ADD_349_U83 P3_U4306 ; P3_U6153
g4333 nand P3_ADD_344_U83 P3_U2362 ; P3_U6154
g4334 nand P3_ADD_371_1212_U12 P3_U2360 ; P3_U6155
g4335 nand P3_U6137 P3_U3849 ; P3_U6156
g4336 nand P3_U2402 P3_REIP_REG_21__SCAN_IN ; P3_U6157
g4337 nand P3_U4318 P3_U6156 ; P3_U6158
g4338 nand P3_U5631 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_U6159
g4339 nand P3_ADD_360_1242_U80 P3_U2395 ; P3_U6160
g4340 nand P3_SUB_357_1258_U84 P3_U2393 ; P3_U6161
g4341 nand P3_ADD_558_U82 P3_U3220 ; P3_U6162
g4342 nand P3_ADD_553_U82 P3_U4298 ; P3_U6163
g4343 nand P3_ADD_547_U82 P3_U4299 ; P3_U6164
g4344 nand P3_ADD_541_U79 P3_U4300 ; P3_U6165
g4345 nand P3_ADD_536_U79 P3_U4301 ; P3_U6166
g4346 nand P3_ADD_531_U82 P3_U2354 ; P3_U6167
g4347 nand P3_ADD_526_U68 P3_U2355 ; P3_U6168
g4348 nand P3_ADD_515_U79 P3_U4302 ; P3_U6169
g4349 nand P3_ADD_494_U79 P3_U2356 ; P3_U6170
g4350 nand P3_ADD_476_U79 P3_U4303 ; P3_U6171
g4351 nand P3_ADD_441_U79 P3_U4304 ; P3_U6172
g4352 nand P3_ADD_405_U78 P3_U4305 ; P3_U6173
g4353 nand P3_ADD_394_U78 P3_U2357 ; P3_U6174
g4354 nand P3_ADD_385_U82 P3_U2358 ; P3_U6175
g4355 nand P3_ADD_380_U82 P3_U2359 ; P3_U6176
g4356 nand P3_ADD_349_U82 P3_U4306 ; P3_U6177
g4357 nand P3_ADD_344_U82 P3_U2362 ; P3_U6178
g4358 nand P3_ADD_371_1212_U82 P3_U2360 ; P3_U6179
g4359 nand P3_U3862 P3_U3857 ; P3_U6180
g4360 nand P3_U2402 P3_REIP_REG_22__SCAN_IN ; P3_U6181
g4361 nand P3_U4318 P3_U6180 ; P3_U6182
g4362 nand P3_U5631 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_U6183
g4363 nand P3_ADD_360_1242_U12 P3_U2395 ; P3_U6184
g4364 nand P3_SUB_357_1258_U83 P3_U2393 ; P3_U6185
g4365 nand P3_ADD_558_U81 P3_U3220 ; P3_U6186
g4366 nand P3_ADD_553_U81 P3_U4298 ; P3_U6187
g4367 nand P3_ADD_547_U81 P3_U4299 ; P3_U6188
g4368 nand P3_ADD_541_U78 P3_U4300 ; P3_U6189
g4369 nand P3_ADD_536_U78 P3_U4301 ; P3_U6190
g4370 nand P3_ADD_531_U81 P3_U2354 ; P3_U6191
g4371 nand P3_ADD_526_U67 P3_U2355 ; P3_U6192
g4372 nand P3_ADD_515_U78 P3_U4302 ; P3_U6193
g4373 nand P3_ADD_494_U78 P3_U2356 ; P3_U6194
g4374 nand P3_ADD_476_U78 P3_U4303 ; P3_U6195
g4375 nand P3_ADD_441_U78 P3_U4304 ; P3_U6196
g4376 nand P3_ADD_405_U77 P3_U4305 ; P3_U6197
g4377 nand P3_ADD_394_U77 P3_U2357 ; P3_U6198
g4378 nand P3_ADD_385_U81 P3_U2358 ; P3_U6199
g4379 nand P3_ADD_380_U81 P3_U2359 ; P3_U6200
g4380 nand P3_ADD_349_U81 P3_U4306 ; P3_U6201
g4381 nand P3_ADD_344_U81 P3_U2362 ; P3_U6202
g4382 nand P3_ADD_371_1212_U13 P3_U2360 ; P3_U6203
g4383 nand P3_U3872 P3_U3867 ; P3_U6204
g4384 nand P3_U2402 P3_REIP_REG_23__SCAN_IN ; P3_U6205
g4385 nand P3_U4318 P3_U6204 ; P3_U6206
g4386 nand P3_U5631 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_U6207
g4387 nand P3_ADD_360_1242_U79 P3_U2395 ; P3_U6208
g4388 nand P3_SUB_357_1258_U82 P3_U2393 ; P3_U6209
g4389 nand P3_ADD_558_U80 P3_U3220 ; P3_U6210
g4390 nand P3_ADD_553_U80 P3_U4298 ; P3_U6211
g4391 nand P3_ADD_547_U80 P3_U4299 ; P3_U6212
g4392 nand P3_ADD_541_U77 P3_U4300 ; P3_U6213
g4393 nand P3_ADD_536_U77 P3_U4301 ; P3_U6214
g4394 nand P3_ADD_531_U80 P3_U2354 ; P3_U6215
g4395 nand P3_ADD_526_U66 P3_U2355 ; P3_U6216
g4396 nand P3_ADD_515_U77 P3_U4302 ; P3_U6217
g4397 nand P3_ADD_494_U77 P3_U2356 ; P3_U6218
g4398 nand P3_ADD_476_U77 P3_U4303 ; P3_U6219
g4399 nand P3_ADD_441_U77 P3_U4304 ; P3_U6220
g4400 nand P3_ADD_405_U76 P3_U4305 ; P3_U6221
g4401 nand P3_ADD_394_U76 P3_U2357 ; P3_U6222
g4402 nand P3_ADD_385_U80 P3_U2358 ; P3_U6223
g4403 nand P3_ADD_380_U80 P3_U2359 ; P3_U6224
g4404 nand P3_ADD_349_U80 P3_U4306 ; P3_U6225
g4405 nand P3_ADD_344_U80 P3_U2362 ; P3_U6226
g4406 nand P3_ADD_371_1212_U81 P3_U2360 ; P3_U6227
g4407 nand P3_U3882 P3_U3877 ; P3_U6228
g4408 nand P3_U2402 P3_REIP_REG_24__SCAN_IN ; P3_U6229
g4409 nand P3_U4318 P3_U6228 ; P3_U6230
g4410 nand P3_U5631 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_U6231
g4411 nand P3_ADD_360_1242_U13 P3_U2395 ; P3_U6232
g4412 nand P3_SUB_357_1258_U81 P3_U2393 ; P3_U6233
g4413 nand P3_ADD_558_U79 P3_U3220 ; P3_U6234
g4414 nand P3_ADD_553_U79 P3_U4298 ; P3_U6235
g4415 nand P3_ADD_547_U79 P3_U4299 ; P3_U6236
g4416 nand P3_ADD_541_U76 P3_U4300 ; P3_U6237
g4417 nand P3_ADD_536_U76 P3_U4301 ; P3_U6238
g4418 nand P3_ADD_531_U79 P3_U2354 ; P3_U6239
g4419 nand P3_ADD_526_U65 P3_U2355 ; P3_U6240
g4420 nand P3_ADD_515_U76 P3_U4302 ; P3_U6241
g4421 nand P3_ADD_494_U76 P3_U2356 ; P3_U6242
g4422 nand P3_ADD_476_U76 P3_U4303 ; P3_U6243
g4423 nand P3_ADD_441_U76 P3_U4304 ; P3_U6244
g4424 nand P3_ADD_405_U75 P3_U4305 ; P3_U6245
g4425 nand P3_ADD_394_U75 P3_U2357 ; P3_U6246
g4426 nand P3_ADD_385_U79 P3_U2358 ; P3_U6247
g4427 nand P3_ADD_380_U79 P3_U2359 ; P3_U6248
g4428 nand P3_ADD_349_U79 P3_U4306 ; P3_U6249
g4429 nand P3_ADD_344_U79 P3_U2362 ; P3_U6250
g4430 nand P3_ADD_371_1212_U14 P3_U2360 ; P3_U6251
g4431 nand P3_U3892 P3_U3887 ; P3_U6252
g4432 nand P3_U2402 P3_REIP_REG_25__SCAN_IN ; P3_U6253
g4433 nand P3_U4318 P3_U6252 ; P3_U6254
g4434 nand P3_U5631 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_U6255
g4435 nand P3_ADD_360_1242_U14 P3_U2395 ; P3_U6256
g4436 nand P3_SUB_357_1258_U18 P3_U2393 ; P3_U6257
g4437 nand P3_ADD_558_U78 P3_U3220 ; P3_U6258
g4438 nand P3_ADD_553_U78 P3_U4298 ; P3_U6259
g4439 nand P3_ADD_547_U78 P3_U4299 ; P3_U6260
g4440 nand P3_ADD_541_U75 P3_U4300 ; P3_U6261
g4441 nand P3_ADD_536_U75 P3_U4301 ; P3_U6262
g4442 nand P3_ADD_531_U78 P3_U2354 ; P3_U6263
g4443 nand P3_ADD_526_U64 P3_U2355 ; P3_U6264
g4444 nand P3_ADD_515_U75 P3_U4302 ; P3_U6265
g4445 nand P3_ADD_494_U75 P3_U2356 ; P3_U6266
g4446 nand P3_ADD_476_U75 P3_U4303 ; P3_U6267
g4447 nand P3_ADD_441_U75 P3_U4304 ; P3_U6268
g4448 nand P3_ADD_405_U74 P3_U4305 ; P3_U6269
g4449 nand P3_ADD_394_U74 P3_U2357 ; P3_U6270
g4450 nand P3_ADD_385_U78 P3_U2358 ; P3_U6271
g4451 nand P3_ADD_380_U78 P3_U2359 ; P3_U6272
g4452 nand P3_ADD_349_U78 P3_U4306 ; P3_U6273
g4453 nand P3_ADD_344_U78 P3_U2362 ; P3_U6274
g4454 nand P3_ADD_371_1212_U15 P3_U2360 ; P3_U6275
g4455 nand P3_U3894 P3_U6258 P3_U3895 P3_U3897 P3_U3902 ; P3_U6276
g4456 nand P3_U2402 P3_REIP_REG_26__SCAN_IN ; P3_U6277
g4457 nand P3_U4318 P3_U6276 ; P3_U6278
g4458 nand P3_U5631 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_U6279
g4459 nand P3_ADD_360_1242_U78 P3_U2395 ; P3_U6280
g4460 nand P3_SUB_357_1258_U80 P3_U2393 ; P3_U6281
g4461 nand P3_ADD_558_U77 P3_U3220 ; P3_U6282
g4462 nand P3_ADD_553_U77 P3_U4298 ; P3_U6283
g4463 nand P3_ADD_547_U77 P3_U4299 ; P3_U6284
g4464 nand P3_ADD_541_U74 P3_U4300 ; P3_U6285
g4465 nand P3_ADD_536_U74 P3_U4301 ; P3_U6286
g4466 nand P3_ADD_531_U77 P3_U2354 ; P3_U6287
g4467 nand P3_ADD_526_U63 P3_U2355 ; P3_U6288
g4468 nand P3_ADD_515_U74 P3_U4302 ; P3_U6289
g4469 nand P3_ADD_494_U74 P3_U2356 ; P3_U6290
g4470 nand P3_ADD_476_U74 P3_U4303 ; P3_U6291
g4471 nand P3_ADD_441_U74 P3_U4304 ; P3_U6292
g4472 nand P3_ADD_405_U73 P3_U4305 ; P3_U6293
g4473 nand P3_ADD_394_U73 P3_U2357 ; P3_U6294
g4474 nand P3_ADD_385_U77 P3_U2358 ; P3_U6295
g4475 nand P3_ADD_380_U77 P3_U2359 ; P3_U6296
g4476 nand P3_ADD_349_U77 P3_U4306 ; P3_U6297
g4477 nand P3_ADD_344_U77 P3_U2362 ; P3_U6298
g4478 nand P3_ADD_371_1212_U80 P3_U2360 ; P3_U6299
g4479 nand P3_U3903 P3_U6282 P3_U3904 P3_U3906 P3_U3911 ; P3_U6300
g4480 nand P3_U2402 P3_REIP_REG_27__SCAN_IN ; P3_U6301
g4481 nand P3_U4318 P3_U6300 ; P3_U6302
g4482 nand P3_U5631 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_U6303
g4483 nand P3_ADD_360_1242_U15 P3_U2395 ; P3_U6304
g4484 nand P3_SUB_357_1258_U19 P3_U2393 ; P3_U6305
g4485 nand P3_ADD_558_U76 P3_U3220 ; P3_U6306
g4486 nand P3_ADD_553_U76 P3_U4298 ; P3_U6307
g4487 nand P3_ADD_547_U76 P3_U4299 ; P3_U6308
g4488 nand P3_ADD_541_U73 P3_U4300 ; P3_U6309
g4489 nand P3_ADD_536_U73 P3_U4301 ; P3_U6310
g4490 nand P3_ADD_531_U76 P3_U2354 ; P3_U6311
g4491 nand P3_ADD_526_U62 P3_U2355 ; P3_U6312
g4492 nand P3_ADD_515_U73 P3_U4302 ; P3_U6313
g4493 nand P3_ADD_494_U73 P3_U2356 ; P3_U6314
g4494 nand P3_ADD_476_U73 P3_U4303 ; P3_U6315
g4495 nand P3_ADD_441_U73 P3_U4304 ; P3_U6316
g4496 nand P3_ADD_405_U72 P3_U4305 ; P3_U6317
g4497 nand P3_ADD_394_U72 P3_U2357 ; P3_U6318
g4498 nand P3_ADD_385_U76 P3_U2358 ; P3_U6319
g4499 nand P3_ADD_380_U76 P3_U2359 ; P3_U6320
g4500 nand P3_ADD_349_U76 P3_U4306 ; P3_U6321
g4501 nand P3_ADD_344_U76 P3_U2362 ; P3_U6322
g4502 nand P3_ADD_371_1212_U16 P3_U2360 ; P3_U6323
g4503 nand P3_U3912 P3_U6306 P3_U3913 P3_U3915 P3_U3920 ; P3_U6324
g4504 nand P3_U2402 P3_REIP_REG_28__SCAN_IN ; P3_U6325
g4505 nand P3_U4318 P3_U6324 ; P3_U6326
g4506 nand P3_U5631 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_U6327
g4507 nand P3_ADD_360_1242_U16 P3_U2395 ; P3_U6328
g4508 nand P3_SUB_357_1258_U79 P3_U2393 ; P3_U6329
g4509 nand P3_ADD_558_U75 P3_U3220 ; P3_U6330
g4510 nand P3_ADD_553_U75 P3_U4298 ; P3_U6331
g4511 nand P3_ADD_547_U75 P3_U4299 ; P3_U6332
g4512 nand P3_ADD_541_U72 P3_U4300 ; P3_U6333
g4513 nand P3_ADD_536_U72 P3_U4301 ; P3_U6334
g4514 nand P3_ADD_531_U75 P3_U2354 ; P3_U6335
g4515 nand P3_ADD_526_U61 P3_U2355 ; P3_U6336
g4516 nand P3_ADD_515_U72 P3_U4302 ; P3_U6337
g4517 nand P3_ADD_494_U72 P3_U2356 ; P3_U6338
g4518 nand P3_ADD_476_U72 P3_U4303 ; P3_U6339
g4519 nand P3_ADD_441_U72 P3_U4304 ; P3_U6340
g4520 nand P3_ADD_405_U71 P3_U4305 ; P3_U6341
g4521 nand P3_ADD_394_U71 P3_U2357 ; P3_U6342
g4522 nand P3_ADD_385_U75 P3_U2358 ; P3_U6343
g4523 nand P3_ADD_380_U75 P3_U2359 ; P3_U6344
g4524 nand P3_ADD_349_U75 P3_U4306 ; P3_U6345
g4525 nand P3_ADD_344_U75 P3_U2362 ; P3_U6346
g4526 nand P3_ADD_371_1212_U17 P3_U2360 ; P3_U6347
g4527 nand P3_U3921 P3_U6330 P3_U3922 P3_U3924 P3_U3929 ; P3_U6348
g4528 nand P3_U2402 P3_REIP_REG_29__SCAN_IN ; P3_U6349
g4529 nand P3_U4318 P3_U6348 ; P3_U6350
g4530 nand P3_U5631 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_U6351
g4531 nand P3_ADD_360_1242_U77 P3_U2395 ; P3_U6352
g4532 nand P3_SUB_357_1258_U77 P3_U2393 ; P3_U6353
g4533 nand P3_ADD_558_U73 P3_U3220 ; P3_U6354
g4534 nand P3_ADD_553_U73 P3_U4298 ; P3_U6355
g4535 nand P3_ADD_547_U73 P3_U4299 ; P3_U6356
g4536 nand P3_ADD_541_U70 P3_U4300 ; P3_U6357
g4537 nand P3_ADD_536_U70 P3_U4301 ; P3_U6358
g4538 nand P3_ADD_531_U73 P3_U2354 ; P3_U6359
g4539 nand P3_ADD_526_U59 P3_U2355 ; P3_U6360
g4540 nand P3_ADD_515_U70 P3_U4302 ; P3_U6361
g4541 nand P3_ADD_494_U70 P3_U2356 ; P3_U6362
g4542 nand P3_ADD_476_U70 P3_U4303 ; P3_U6363
g4543 nand P3_ADD_441_U70 P3_U4304 ; P3_U6364
g4544 nand P3_ADD_405_U70 P3_U4305 ; P3_U6365
g4545 nand P3_ADD_394_U70 P3_U2357 ; P3_U6366
g4546 nand P3_ADD_385_U73 P3_U2358 ; P3_U6367
g4547 nand P3_ADD_380_U73 P3_U2359 ; P3_U6368
g4548 nand P3_ADD_349_U73 P3_U4306 ; P3_U6369
g4549 nand P3_ADD_344_U73 P3_U2362 ; P3_U6370
g4550 nand P3_ADD_371_1212_U79 P3_U2360 ; P3_U6371
g4551 nand P3_U3930 P3_U6354 P3_U3931 P3_U3933 P3_U3938 ; P3_U6372
g4552 nand P3_U2402 P3_REIP_REG_30__SCAN_IN ; P3_U6373
g4553 nand P3_U4318 P3_U6372 ; P3_U6374
g4554 nand P3_U5631 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_U6375
g4555 nand P3_ADD_360_1242_U90 P3_U2395 ; P3_U6376
g4556 nand P3_SUB_357_1258_U20 P3_U2393 ; P3_U6377
g4557 nand P3_ADD_558_U72 P3_U3220 ; P3_U6378
g4558 nand P3_ADD_553_U72 P3_U4298 ; P3_U6379
g4559 nand P3_ADD_547_U72 P3_U4299 ; P3_U6380
g4560 nand P3_ADD_541_U69 P3_U4300 ; P3_U6381
g4561 nand P3_ADD_536_U69 P3_U4301 ; P3_U6382
g4562 nand P3_ADD_531_U72 P3_U2354 ; P3_U6383
g4563 nand P3_ADD_526_U58 P3_U2355 ; P3_U6384
g4564 nand P3_ADD_515_U69 P3_U4302 ; P3_U6385
g4565 nand P3_ADD_494_U69 P3_U2356 ; P3_U6386
g4566 nand P3_ADD_476_U69 P3_U4303 ; P3_U6387
g4567 nand P3_ADD_441_U69 P3_U4304 ; P3_U6388
g4568 nand P3_ADD_405_U69 P3_U4305 ; P3_U6389
g4569 nand P3_ADD_394_U69 P3_U2357 ; P3_U6390
g4570 nand P3_ADD_385_U72 P3_U2358 ; P3_U6391
g4571 nand P3_ADD_380_U72 P3_U2359 ; P3_U6392
g4572 nand P3_ADD_349_U72 P3_U4306 ; P3_U6393
g4573 nand P3_ADD_344_U72 P3_U2362 ; P3_U6394
g4574 nand P3_ADD_371_1212_U92 P3_U2360 ; P3_U6395
g4575 nand P3_U3950 P3_U3945 ; P3_U6396
g4576 nand P3_U2402 P3_REIP_REG_31__SCAN_IN ; P3_U6397
g4577 nand P3_U5631 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_U6398
g4578 nand P3_GTE_355_U6 P3_U2361 ; P3_U6399
g4579 nand P3_GTE_370_U6 P3_U2360 ; P3_U6400
g4580 nand P3_U6400 P3_U6399 ; P3_U6401
g4581 nand P3_U2390 P3_U6401 ; P3_U6402
g4582 nand P3_U3234 P3_U3121 ; P3_U6403
g4583 not P3_U3249 ; P3_U6404
g4584 nand P3_U2398 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U6405
g4585 nand P3_U2397 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U6406
g4586 nand P3_U2396 P3_ADD_360_1242_U85 ; P3_U6407
g4587 nand P3_U2394 P3_SUB_357_1258_U69 ; P3_U6408
g4588 nand P3_U2389 P3_REIP_REG_0__SCAN_IN ; P3_U6409
g4589 nand P3_U2388 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U6410
g4590 nand P3_U2387 P3_ADD_371_1212_U87 ; P3_U6411
g4591 nand P3_U6404 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U6412
g4592 nand P3_ADD_318_U4 P3_U2398 ; P3_U6413
g4593 nand P3_U2397 P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_U6414
g4594 nand P3_U2396 P3_ADD_360_1242_U19 ; P3_U6415
g4595 nand P3_U2394 P3_SUB_357_1258_U21 ; P3_U6416
g4596 nand P3_U2389 P3_REIP_REG_1__SCAN_IN ; P3_U6417
g4597 nand P3_ADD_339_U4 P3_U2388 ; P3_U6418
g4598 nand P3_U2387 P3_ADD_371_1212_U20 ; P3_U6419
g4599 nand P3_U6404 P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_U6420
g4600 nand P3_ADD_318_U71 P3_U2398 ; P3_U6421
g4601 nand P3_ADD_315_U4 P3_U2397 ; P3_U6422
g4602 nand P3_U2396 P3_ADD_360_1242_U91 ; P3_U6423
g4603 nand P3_U2394 P3_SUB_357_1258_U78 ; P3_U6424
g4604 nand P3_U2389 P3_REIP_REG_2__SCAN_IN ; P3_U6425
g4605 nand P3_ADD_339_U71 P3_U2388 ; P3_U6426
g4606 nand P3_U2387 P3_ADD_371_1212_U93 ; P3_U6427
g4607 nand P3_U6404 P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_U6428
g4608 nand P3_ADD_318_U68 P3_U2398 ; P3_U6429
g4609 nand P3_ADD_315_U66 P3_U2397 ; P3_U6430
g4610 nand P3_U2396 P3_ADD_360_1242_U17 ; P3_U6431
g4611 nand P3_U2394 P3_SUB_357_1258_U76 ; P3_U6432
g4612 nand P3_U2389 P3_REIP_REG_3__SCAN_IN ; P3_U6433
g4613 nand P3_ADD_339_U68 P3_U2388 ; P3_U6434
g4614 nand P3_U2387 P3_ADD_371_1212_U18 ; P3_U6435
g4615 nand P3_U6404 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_U6436
g4616 nand P3_ADD_318_U67 P3_U2398 ; P3_U6437
g4617 nand P3_ADD_315_U65 P3_U2397 ; P3_U6438
g4618 nand P3_U2396 P3_ADD_360_1242_U18 ; P3_U6439
g4619 nand P3_U2394 P3_SUB_357_1258_U75 ; P3_U6440
g4620 nand P3_U2389 P3_REIP_REG_4__SCAN_IN ; P3_U6441
g4621 nand P3_ADD_339_U67 P3_U2388 ; P3_U6442
g4622 nand P3_U2387 P3_ADD_371_1212_U91 ; P3_U6443
g4623 nand P3_U6404 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_U6444
g4624 nand P3_ADD_318_U66 P3_U2398 ; P3_U6445
g4625 nand P3_ADD_315_U64 P3_U2397 ; P3_U6446
g4626 nand P3_U2396 P3_ADD_360_1242_U89 ; P3_U6447
g4627 nand P3_U2394 P3_SUB_357_1258_U74 ; P3_U6448
g4628 nand P3_U2389 P3_REIP_REG_5__SCAN_IN ; P3_U6449
g4629 nand P3_ADD_339_U66 P3_U2388 ; P3_U6450
g4630 nand P3_U2387 P3_ADD_371_1212_U19 ; P3_U6451
g4631 nand P3_U6404 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_U6452
g4632 nand P3_ADD_318_U65 P3_U2398 ; P3_U6453
g4633 nand P3_ADD_315_U63 P3_U2397 ; P3_U6454
g4634 nand P3_U2396 P3_ADD_360_1242_U88 ; P3_U6455
g4635 nand P3_U2394 P3_SUB_357_1258_U73 ; P3_U6456
g4636 nand P3_U2389 P3_REIP_REG_6__SCAN_IN ; P3_U6457
g4637 nand P3_ADD_339_U65 P3_U2388 ; P3_U6458
g4638 nand P3_U2387 P3_ADD_371_1212_U90 ; P3_U6459
g4639 nand P3_U6404 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_U6460
g4640 nand P3_ADD_318_U64 P3_U2398 ; P3_U6461
g4641 nand P3_ADD_315_U62 P3_U2397 ; P3_U6462
g4642 nand P3_U2396 P3_ADD_360_1242_U87 ; P3_U6463
g4643 nand P3_U2394 P3_SUB_357_1258_U72 ; P3_U6464
g4644 nand P3_U2389 P3_REIP_REG_7__SCAN_IN ; P3_U6465
g4645 nand P3_ADD_339_U64 P3_U2388 ; P3_U6466
g4646 nand P3_U2387 P3_ADD_371_1212_U89 ; P3_U6467
g4647 nand P3_U6404 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_U6468
g4648 nand P3_ADD_318_U63 P3_U2398 ; P3_U6469
g4649 nand P3_ADD_315_U61 P3_U2397 ; P3_U6470
g4650 nand P3_U2396 P3_ADD_360_1242_U86 ; P3_U6471
g4651 nand P3_U2394 P3_SUB_357_1258_U71 ; P3_U6472
g4652 nand P3_U2389 P3_REIP_REG_8__SCAN_IN ; P3_U6473
g4653 nand P3_ADD_339_U63 P3_U2388 ; P3_U6474
g4654 nand P3_U2387 P3_ADD_371_1212_U88 ; P3_U6475
g4655 nand P3_U6404 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_U6476
g4656 nand P3_ADD_318_U62 P3_U2398 ; P3_U6477
g4657 nand P3_ADD_315_U60 P3_U2397 ; P3_U6478
g4658 nand P3_U2396 P3_ADD_360_1242_U106 ; P3_U6479
g4659 nand P3_U2394 P3_SUB_357_1258_U70 ; P3_U6480
g4660 nand P3_U2389 P3_REIP_REG_9__SCAN_IN ; P3_U6481
g4661 nand P3_ADD_339_U62 P3_U2388 ; P3_U6482
g4662 nand P3_U2387 P3_ADD_371_1212_U109 ; P3_U6483
g4663 nand P3_U6404 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_U6484
g4664 nand P3_ADD_318_U91 P3_U2398 ; P3_U6485
g4665 nand P3_ADD_315_U88 P3_U2397 ; P3_U6486
g4666 nand P3_U2396 P3_ADD_360_1242_U4 ; P3_U6487
g4667 nand P3_U2394 P3_SUB_357_1258_U93 ; P3_U6488
g4668 nand P3_U2389 P3_REIP_REG_10__SCAN_IN ; P3_U6489
g4669 nand P3_ADD_339_U91 P3_U2388 ; P3_U6490
g4670 nand P3_U2387 P3_ADD_371_1212_U5 ; P3_U6491
g4671 nand P3_U6404 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_U6492
g4672 nand P3_ADD_318_U90 P3_U2398 ; P3_U6493
g4673 nand P3_ADD_315_U87 P3_U2397 ; P3_U6494
g4674 nand P3_U2396 P3_ADD_360_1242_U84 ; P3_U6495
g4675 nand P3_U2394 P3_SUB_357_1258_U92 ; P3_U6496
g4676 nand P3_U2389 P3_REIP_REG_11__SCAN_IN ; P3_U6497
g4677 nand P3_ADD_339_U90 P3_U2388 ; P3_U6498
g4678 nand P3_U2387 P3_ADD_371_1212_U86 ; P3_U6499
g4679 nand P3_U6404 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_U6500
g4680 nand P3_ADD_318_U89 P3_U2398 ; P3_U6501
g4681 nand P3_ADD_315_U86 P3_U2397 ; P3_U6502
g4682 nand P3_U2396 P3_ADD_360_1242_U5 ; P3_U6503
g4683 nand P3_U2394 P3_SUB_357_1258_U91 ; P3_U6504
g4684 nand P3_U2389 P3_REIP_REG_12__SCAN_IN ; P3_U6505
g4685 nand P3_ADD_339_U89 P3_U2388 ; P3_U6506
g4686 nand P3_U2387 P3_ADD_371_1212_U6 ; P3_U6507
g4687 nand P3_U6404 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_U6508
g4688 nand P3_ADD_318_U88 P3_U2398 ; P3_U6509
g4689 nand P3_ADD_315_U85 P3_U2397 ; P3_U6510
g4690 nand P3_U2396 P3_ADD_360_1242_U6 ; P3_U6511
g4691 nand P3_U2394 P3_SUB_357_1258_U15 ; P3_U6512
g4692 nand P3_U2389 P3_REIP_REG_13__SCAN_IN ; P3_U6513
g4693 nand P3_ADD_339_U88 P3_U2388 ; P3_U6514
g4694 nand P3_U2387 P3_ADD_371_1212_U7 ; P3_U6515
g4695 nand P3_U6404 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_U6516
g4696 nand P3_ADD_318_U87 P3_U2398 ; P3_U6517
g4697 nand P3_ADD_315_U84 P3_U2397 ; P3_U6518
g4698 nand P3_U2396 P3_ADD_360_1242_U83 ; P3_U6519
g4699 nand P3_U2394 P3_SUB_357_1258_U90 ; P3_U6520
g4700 nand P3_U2389 P3_REIP_REG_14__SCAN_IN ; P3_U6521
g4701 nand P3_ADD_339_U87 P3_U2388 ; P3_U6522
g4702 nand P3_U2387 P3_ADD_371_1212_U85 ; P3_U6523
g4703 nand P3_U6404 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_U6524
g4704 nand P3_ADD_318_U86 P3_U2398 ; P3_U6525
g4705 nand P3_ADD_315_U83 P3_U2397 ; P3_U6526
g4706 nand P3_U2396 P3_ADD_360_1242_U7 ; P3_U6527
g4707 nand P3_U2394 P3_SUB_357_1258_U89 ; P3_U6528
g4708 nand P3_U2389 P3_REIP_REG_15__SCAN_IN ; P3_U6529
g4709 nand P3_ADD_339_U86 P3_U2388 ; P3_U6530
g4710 nand P3_U2387 P3_ADD_371_1212_U8 ; P3_U6531
g4711 nand P3_U6404 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_U6532
g4712 nand P3_ADD_318_U85 P3_U2398 ; P3_U6533
g4713 nand P3_ADD_315_U82 P3_U2397 ; P3_U6534
g4714 nand P3_U2396 P3_ADD_360_1242_U82 ; P3_U6535
g4715 nand P3_U2394 P3_SUB_357_1258_U88 ; P3_U6536
g4716 nand P3_U2389 P3_REIP_REG_16__SCAN_IN ; P3_U6537
g4717 nand P3_ADD_339_U85 P3_U2388 ; P3_U6538
g4718 nand P3_U2387 P3_ADD_371_1212_U84 ; P3_U6539
g4719 nand P3_U6404 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_U6540
g4720 nand P3_ADD_318_U84 P3_U2398 ; P3_U6541
g4721 nand P3_ADD_315_U81 P3_U2397 ; P3_U6542
g4722 nand P3_U2396 P3_ADD_360_1242_U8 ; P3_U6543
g4723 nand P3_U2394 P3_SUB_357_1258_U16 ; P3_U6544
g4724 nand P3_U2389 P3_REIP_REG_17__SCAN_IN ; P3_U6545
g4725 nand P3_ADD_339_U84 P3_U2388 ; P3_U6546
g4726 nand P3_U2387 P3_ADD_371_1212_U9 ; P3_U6547
g4727 nand P3_U6404 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_U6548
g4728 nand P3_ADD_318_U83 P3_U2398 ; P3_U6549
g4729 nand P3_ADD_315_U80 P3_U2397 ; P3_U6550
g4730 nand P3_U2396 P3_ADD_360_1242_U81 ; P3_U6551
g4731 nand P3_U2394 P3_SUB_357_1258_U87 ; P3_U6552
g4732 nand P3_U2389 P3_REIP_REG_18__SCAN_IN ; P3_U6553
g4733 nand P3_ADD_339_U83 P3_U2388 ; P3_U6554
g4734 nand P3_U2387 P3_ADD_371_1212_U83 ; P3_U6555
g4735 nand P3_U6404 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_U6556
g4736 nand P3_ADD_318_U82 P3_U2398 ; P3_U6557
g4737 nand P3_ADD_315_U79 P3_U2397 ; P3_U6558
g4738 nand P3_U2396 P3_ADD_360_1242_U9 ; P3_U6559
g4739 nand P3_U2394 P3_SUB_357_1258_U86 ; P3_U6560
g4740 nand P3_U2389 P3_REIP_REG_19__SCAN_IN ; P3_U6561
g4741 nand P3_ADD_339_U82 P3_U2388 ; P3_U6562
g4742 nand P3_U2387 P3_ADD_371_1212_U10 ; P3_U6563
g4743 nand P3_U6404 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_U6564
g4744 nand P3_ADD_318_U81 P3_U2398 ; P3_U6565
g4745 nand P3_ADD_315_U78 P3_U2397 ; P3_U6566
g4746 nand P3_U2396 P3_ADD_360_1242_U10 ; P3_U6567
g4747 nand P3_U2394 P3_SUB_357_1258_U17 ; P3_U6568
g4748 nand P3_U2389 P3_REIP_REG_20__SCAN_IN ; P3_U6569
g4749 nand P3_ADD_339_U81 P3_U2388 ; P3_U6570
g4750 nand P3_U2387 P3_ADD_371_1212_U11 ; P3_U6571
g4751 nand P3_U6404 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_U6572
g4752 nand P3_ADD_318_U80 P3_U2398 ; P3_U6573
g4753 nand P3_ADD_315_U77 P3_U2397 ; P3_U6574
g4754 nand P3_U2396 P3_ADD_360_1242_U11 ; P3_U6575
g4755 nand P3_U2394 P3_SUB_357_1258_U85 ; P3_U6576
g4756 nand P3_U2389 P3_REIP_REG_21__SCAN_IN ; P3_U6577
g4757 nand P3_ADD_339_U80 P3_U2388 ; P3_U6578
g4758 nand P3_U2387 P3_ADD_371_1212_U12 ; P3_U6579
g4759 nand P3_U6404 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_U6580
g4760 nand P3_ADD_318_U79 P3_U2398 ; P3_U6581
g4761 nand P3_ADD_315_U76 P3_U2397 ; P3_U6582
g4762 nand P3_U2396 P3_ADD_360_1242_U80 ; P3_U6583
g4763 nand P3_U2394 P3_SUB_357_1258_U84 ; P3_U6584
g4764 nand P3_U2389 P3_REIP_REG_22__SCAN_IN ; P3_U6585
g4765 nand P3_ADD_339_U79 P3_U2388 ; P3_U6586
g4766 nand P3_U2387 P3_ADD_371_1212_U82 ; P3_U6587
g4767 nand P3_U6404 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_U6588
g4768 nand P3_ADD_318_U78 P3_U2398 ; P3_U6589
g4769 nand P3_ADD_315_U75 P3_U2397 ; P3_U6590
g4770 nand P3_U2396 P3_ADD_360_1242_U12 ; P3_U6591
g4771 nand P3_U2394 P3_SUB_357_1258_U83 ; P3_U6592
g4772 nand P3_U2389 P3_REIP_REG_23__SCAN_IN ; P3_U6593
g4773 nand P3_ADD_339_U78 P3_U2388 ; P3_U6594
g4774 nand P3_U2387 P3_ADD_371_1212_U13 ; P3_U6595
g4775 nand P3_U6404 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_U6596
g4776 nand P3_ADD_318_U77 P3_U2398 ; P3_U6597
g4777 nand P3_ADD_315_U74 P3_U2397 ; P3_U6598
g4778 nand P3_U2396 P3_ADD_360_1242_U79 ; P3_U6599
g4779 nand P3_U2394 P3_SUB_357_1258_U82 ; P3_U6600
g4780 nand P3_U2389 P3_REIP_REG_24__SCAN_IN ; P3_U6601
g4781 nand P3_ADD_339_U77 P3_U2388 ; P3_U6602
g4782 nand P3_U2387 P3_ADD_371_1212_U81 ; P3_U6603
g4783 nand P3_U6404 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_U6604
g4784 nand P3_ADD_318_U76 P3_U2398 ; P3_U6605
g4785 nand P3_ADD_315_U73 P3_U2397 ; P3_U6606
g4786 nand P3_U2396 P3_ADD_360_1242_U13 ; P3_U6607
g4787 nand P3_U2394 P3_SUB_357_1258_U81 ; P3_U6608
g4788 nand P3_U2389 P3_REIP_REG_25__SCAN_IN ; P3_U6609
g4789 nand P3_ADD_339_U76 P3_U2388 ; P3_U6610
g4790 nand P3_U2387 P3_ADD_371_1212_U14 ; P3_U6611
g4791 nand P3_U6404 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_U6612
g4792 nand P3_ADD_318_U75 P3_U2398 ; P3_U6613
g4793 nand P3_ADD_315_U72 P3_U2397 ; P3_U6614
g4794 nand P3_U2396 P3_ADD_360_1242_U14 ; P3_U6615
g4795 nand P3_U2394 P3_SUB_357_1258_U18 ; P3_U6616
g4796 nand P3_U2389 P3_REIP_REG_26__SCAN_IN ; P3_U6617
g4797 nand P3_ADD_339_U75 P3_U2388 ; P3_U6618
g4798 nand P3_U2387 P3_ADD_371_1212_U15 ; P3_U6619
g4799 nand P3_U6404 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_U6620
g4800 nand P3_ADD_318_U74 P3_U2398 ; P3_U6621
g4801 nand P3_ADD_315_U71 P3_U2397 ; P3_U6622
g4802 nand P3_U2396 P3_ADD_360_1242_U78 ; P3_U6623
g4803 nand P3_U2394 P3_SUB_357_1258_U80 ; P3_U6624
g4804 nand P3_U2389 P3_REIP_REG_27__SCAN_IN ; P3_U6625
g4805 nand P3_ADD_339_U74 P3_U2388 ; P3_U6626
g4806 nand P3_U2387 P3_ADD_371_1212_U80 ; P3_U6627
g4807 nand P3_U6404 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_U6628
g4808 nand P3_ADD_318_U73 P3_U2398 ; P3_U6629
g4809 nand P3_ADD_315_U70 P3_U2397 ; P3_U6630
g4810 nand P3_U2396 P3_ADD_360_1242_U15 ; P3_U6631
g4811 nand P3_U2394 P3_SUB_357_1258_U19 ; P3_U6632
g4812 nand P3_U2389 P3_REIP_REG_28__SCAN_IN ; P3_U6633
g4813 nand P3_ADD_339_U73 P3_U2388 ; P3_U6634
g4814 nand P3_U2387 P3_ADD_371_1212_U16 ; P3_U6635
g4815 nand P3_U6404 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_U6636
g4816 nand P3_ADD_318_U72 P3_U2398 ; P3_U6637
g4817 nand P3_ADD_315_U69 P3_U2397 ; P3_U6638
g4818 nand P3_U2396 P3_ADD_360_1242_U16 ; P3_U6639
g4819 nand P3_U2394 P3_SUB_357_1258_U79 ; P3_U6640
g4820 nand P3_U2389 P3_REIP_REG_29__SCAN_IN ; P3_U6641
g4821 nand P3_ADD_339_U72 P3_U2388 ; P3_U6642
g4822 nand P3_U2387 P3_ADD_371_1212_U17 ; P3_U6643
g4823 nand P3_U6404 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_U6644
g4824 nand P3_ADD_318_U70 P3_U2398 ; P3_U6645
g4825 nand P3_ADD_315_U68 P3_U2397 ; P3_U6646
g4826 nand P3_U2396 P3_ADD_360_1242_U77 ; P3_U6647
g4827 nand P3_U2394 P3_SUB_357_1258_U77 ; P3_U6648
g4828 nand P3_U2389 P3_REIP_REG_30__SCAN_IN ; P3_U6649
g4829 nand P3_ADD_339_U70 P3_U2388 ; P3_U6650
g4830 nand P3_U2387 P3_ADD_371_1212_U79 ; P3_U6651
g4831 nand P3_U6404 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_U6652
g4832 nand P3_ADD_318_U69 P3_U2398 ; P3_U6653
g4833 nand P3_ADD_315_U67 P3_U2397 ; P3_U6654
g4834 nand P3_U2396 P3_ADD_360_1242_U90 ; P3_U6655
g4835 nand P3_U2394 P3_SUB_357_1258_U20 ; P3_U6656
g4836 nand P3_U2389 P3_REIP_REG_31__SCAN_IN ; P3_U6657
g4837 nand P3_ADD_339_U69 P3_U2388 ; P3_U6658
g4838 nand P3_U2387 P3_ADD_371_1212_U92 ; P3_U6659
g4839 nand P3_U6404 P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_U6660
g4840 nand P3_U4304 P3_U2630 P3_GTE_412_U6 ; P3_U6661
g4841 nand P3_GTE_450_U6 P3_U4303 ; P3_U6662
g4842 nand P3_U6662 P3_U6661 ; P3_U6663
g4843 nand P3_U2407 P3_EAX_REG_15__SCAN_IN ; P3_U6664
g4844 nand P3_U2406 BUF2_REG_15__SCAN_IN ; P3_U6665
g4845 nand P3_U3250 P3_LWORD_REG_15__SCAN_IN ; P3_U6666
g4846 nand P3_U2407 P3_EAX_REG_14__SCAN_IN ; P3_U6667
g4847 nand P3_U2406 BUF2_REG_14__SCAN_IN ; P3_U6668
g4848 nand P3_U3250 P3_LWORD_REG_14__SCAN_IN ; P3_U6669
g4849 nand P3_U2407 P3_EAX_REG_13__SCAN_IN ; P3_U6670
g4850 nand P3_U2406 BUF2_REG_13__SCAN_IN ; P3_U6671
g4851 nand P3_U3250 P3_LWORD_REG_13__SCAN_IN ; P3_U6672
g4852 nand P3_U2407 P3_EAX_REG_12__SCAN_IN ; P3_U6673
g4853 nand P3_U2406 BUF2_REG_12__SCAN_IN ; P3_U6674
g4854 nand P3_U3250 P3_LWORD_REG_12__SCAN_IN ; P3_U6675
g4855 nand P3_U2407 P3_EAX_REG_11__SCAN_IN ; P3_U6676
g4856 nand P3_U2406 BUF2_REG_11__SCAN_IN ; P3_U6677
g4857 nand P3_U3250 P3_LWORD_REG_11__SCAN_IN ; P3_U6678
g4858 nand P3_U2407 P3_EAX_REG_10__SCAN_IN ; P3_U6679
g4859 nand P3_U2406 BUF2_REG_10__SCAN_IN ; P3_U6680
g4860 nand P3_U3250 P3_LWORD_REG_10__SCAN_IN ; P3_U6681
g4861 nand P3_U2407 P3_EAX_REG_9__SCAN_IN ; P3_U6682
g4862 nand P3_U2406 BUF2_REG_9__SCAN_IN ; P3_U6683
g4863 nand P3_U3250 P3_LWORD_REG_9__SCAN_IN ; P3_U6684
g4864 nand P3_U2407 P3_EAX_REG_8__SCAN_IN ; P3_U6685
g4865 nand P3_U2406 BUF2_REG_8__SCAN_IN ; P3_U6686
g4866 nand P3_U3250 P3_LWORD_REG_8__SCAN_IN ; P3_U6687
g4867 nand P3_U2407 P3_EAX_REG_7__SCAN_IN ; P3_U6688
g4868 nand P3_U2406 BUF2_REG_7__SCAN_IN ; P3_U6689
g4869 nand P3_U3250 P3_LWORD_REG_7__SCAN_IN ; P3_U6690
g4870 nand P3_U2407 P3_EAX_REG_6__SCAN_IN ; P3_U6691
g4871 nand P3_U2406 BUF2_REG_6__SCAN_IN ; P3_U6692
g4872 nand P3_U3250 P3_LWORD_REG_6__SCAN_IN ; P3_U6693
g4873 nand P3_U2407 P3_EAX_REG_5__SCAN_IN ; P3_U6694
g4874 nand P3_U2406 BUF2_REG_5__SCAN_IN ; P3_U6695
g4875 nand P3_U3250 P3_LWORD_REG_5__SCAN_IN ; P3_U6696
g4876 nand P3_U2407 P3_EAX_REG_4__SCAN_IN ; P3_U6697
g4877 nand P3_U2406 BUF2_REG_4__SCAN_IN ; P3_U6698
g4878 nand P3_U3250 P3_LWORD_REG_4__SCAN_IN ; P3_U6699
g4879 nand P3_U2407 P3_EAX_REG_3__SCAN_IN ; P3_U6700
g4880 nand P3_U2406 BUF2_REG_3__SCAN_IN ; P3_U6701
g4881 nand P3_U3250 P3_LWORD_REG_3__SCAN_IN ; P3_U6702
g4882 nand P3_U2407 P3_EAX_REG_2__SCAN_IN ; P3_U6703
g4883 nand P3_U2406 BUF2_REG_2__SCAN_IN ; P3_U6704
g4884 nand P3_U3250 P3_LWORD_REG_2__SCAN_IN ; P3_U6705
g4885 nand P3_U2407 P3_EAX_REG_1__SCAN_IN ; P3_U6706
g4886 nand P3_U2406 BUF2_REG_1__SCAN_IN ; P3_U6707
g4887 nand P3_U3250 P3_LWORD_REG_1__SCAN_IN ; P3_U6708
g4888 nand P3_U2407 P3_EAX_REG_0__SCAN_IN ; P3_U6709
g4889 nand P3_U2406 BUF2_REG_0__SCAN_IN ; P3_U6710
g4890 nand P3_U3250 P3_LWORD_REG_0__SCAN_IN ; P3_U6711
g4891 nand P3_U2407 P3_EAX_REG_30__SCAN_IN ; P3_U6712
g4892 nand P3_U2406 BUF2_REG_14__SCAN_IN ; P3_U6713
g4893 nand P3_U3250 P3_UWORD_REG_14__SCAN_IN ; P3_U6714
g4894 nand P3_U2407 P3_EAX_REG_29__SCAN_IN ; P3_U6715
g4895 nand P3_U2406 BUF2_REG_13__SCAN_IN ; P3_U6716
g4896 nand P3_U3250 P3_UWORD_REG_13__SCAN_IN ; P3_U6717
g4897 nand P3_U2407 P3_EAX_REG_28__SCAN_IN ; P3_U6718
g4898 nand P3_U2406 BUF2_REG_12__SCAN_IN ; P3_U6719
g4899 nand P3_U3250 P3_UWORD_REG_12__SCAN_IN ; P3_U6720
g4900 nand P3_U2407 P3_EAX_REG_27__SCAN_IN ; P3_U6721
g4901 nand P3_U2406 BUF2_REG_11__SCAN_IN ; P3_U6722
g4902 nand P3_U3250 P3_UWORD_REG_11__SCAN_IN ; P3_U6723
g4903 nand P3_U2407 P3_EAX_REG_26__SCAN_IN ; P3_U6724
g4904 nand P3_U2406 BUF2_REG_10__SCAN_IN ; P3_U6725
g4905 nand P3_U3250 P3_UWORD_REG_10__SCAN_IN ; P3_U6726
g4906 nand P3_U2407 P3_EAX_REG_25__SCAN_IN ; P3_U6727
g4907 nand P3_U2406 BUF2_REG_9__SCAN_IN ; P3_U6728
g4908 nand P3_U3250 P3_UWORD_REG_9__SCAN_IN ; P3_U6729
g4909 nand P3_U2407 P3_EAX_REG_24__SCAN_IN ; P3_U6730
g4910 nand P3_U2406 BUF2_REG_8__SCAN_IN ; P3_U6731
g4911 nand P3_U3250 P3_UWORD_REG_8__SCAN_IN ; P3_U6732
g4912 nand P3_U2407 P3_EAX_REG_23__SCAN_IN ; P3_U6733
g4913 nand P3_U2406 BUF2_REG_7__SCAN_IN ; P3_U6734
g4914 nand P3_U3250 P3_UWORD_REG_7__SCAN_IN ; P3_U6735
g4915 nand P3_U2407 P3_EAX_REG_22__SCAN_IN ; P3_U6736
g4916 nand P3_U2406 BUF2_REG_6__SCAN_IN ; P3_U6737
g4917 nand P3_U3250 P3_UWORD_REG_6__SCAN_IN ; P3_U6738
g4918 nand P3_U2407 P3_EAX_REG_21__SCAN_IN ; P3_U6739
g4919 nand P3_U2406 BUF2_REG_5__SCAN_IN ; P3_U6740
g4920 nand P3_U3250 P3_UWORD_REG_5__SCAN_IN ; P3_U6741
g4921 nand P3_U2407 P3_EAX_REG_20__SCAN_IN ; P3_U6742
g4922 nand P3_U2406 BUF2_REG_4__SCAN_IN ; P3_U6743
g4923 nand P3_U3250 P3_UWORD_REG_4__SCAN_IN ; P3_U6744
g4924 nand P3_U2407 P3_EAX_REG_19__SCAN_IN ; P3_U6745
g4925 nand P3_U2406 BUF2_REG_3__SCAN_IN ; P3_U6746
g4926 nand P3_U3250 P3_UWORD_REG_3__SCAN_IN ; P3_U6747
g4927 nand P3_U2407 P3_EAX_REG_18__SCAN_IN ; P3_U6748
g4928 nand P3_U2406 BUF2_REG_2__SCAN_IN ; P3_U6749
g4929 nand P3_U3250 P3_UWORD_REG_2__SCAN_IN ; P3_U6750
g4930 nand P3_U2407 P3_EAX_REG_17__SCAN_IN ; P3_U6751
g4931 nand P3_U2406 BUF2_REG_1__SCAN_IN ; P3_U6752
g4932 nand P3_U3250 P3_UWORD_REG_1__SCAN_IN ; P3_U6753
g4933 nand P3_U2407 P3_EAX_REG_16__SCAN_IN ; P3_U6754
g4934 nand P3_U2406 BUF2_REG_0__SCAN_IN ; P3_U6755
g4935 nand P3_U3250 P3_UWORD_REG_0__SCAN_IN ; P3_U6756
g4936 nand P3_U3986 P3_U3255 ; P3_U6757
g4937 nand P3_U2453 P3_U3121 ; P3_U6758
g4938 not P3_U3251 ; P3_U6759
g4939 nand P3_U2410 P3_LWORD_REG_0__SCAN_IN ; P3_U6760
g4940 nand P3_U2409 P3_EAX_REG_0__SCAN_IN ; P3_U6761
g4941 nand P3_U6759 P3_DATAO_REG_0__SCAN_IN ; P3_U6762
g4942 nand P3_U2410 P3_LWORD_REG_1__SCAN_IN ; P3_U6763
g4943 nand P3_U2409 P3_EAX_REG_1__SCAN_IN ; P3_U6764
g4944 nand P3_U6759 P3_DATAO_REG_1__SCAN_IN ; P3_U6765
g4945 nand P3_U2410 P3_LWORD_REG_2__SCAN_IN ; P3_U6766
g4946 nand P3_U2409 P3_EAX_REG_2__SCAN_IN ; P3_U6767
g4947 nand P3_U6759 P3_DATAO_REG_2__SCAN_IN ; P3_U6768
g4948 nand P3_U2410 P3_LWORD_REG_3__SCAN_IN ; P3_U6769
g4949 nand P3_U2409 P3_EAX_REG_3__SCAN_IN ; P3_U6770
g4950 nand P3_U6759 P3_DATAO_REG_3__SCAN_IN ; P3_U6771
g4951 nand P3_U2410 P3_LWORD_REG_4__SCAN_IN ; P3_U6772
g4952 nand P3_U2409 P3_EAX_REG_4__SCAN_IN ; P3_U6773
g4953 nand P3_U6759 P3_DATAO_REG_4__SCAN_IN ; P3_U6774
g4954 nand P3_U2410 P3_LWORD_REG_5__SCAN_IN ; P3_U6775
g4955 nand P3_U2409 P3_EAX_REG_5__SCAN_IN ; P3_U6776
g4956 nand P3_U6759 P3_DATAO_REG_5__SCAN_IN ; P3_U6777
g4957 nand P3_U2410 P3_LWORD_REG_6__SCAN_IN ; P3_U6778
g4958 nand P3_U2409 P3_EAX_REG_6__SCAN_IN ; P3_U6779
g4959 nand P3_U6759 P3_DATAO_REG_6__SCAN_IN ; P3_U6780
g4960 nand P3_U2410 P3_LWORD_REG_7__SCAN_IN ; P3_U6781
g4961 nand P3_U2409 P3_EAX_REG_7__SCAN_IN ; P3_U6782
g4962 nand P3_U6759 P3_DATAO_REG_7__SCAN_IN ; P3_U6783
g4963 nand P3_U2410 P3_LWORD_REG_8__SCAN_IN ; P3_U6784
g4964 nand P3_U2409 P3_EAX_REG_8__SCAN_IN ; P3_U6785
g4965 nand P3_U6759 P3_DATAO_REG_8__SCAN_IN ; P3_U6786
g4966 nand P3_U2410 P3_LWORD_REG_9__SCAN_IN ; P3_U6787
g4967 nand P3_U2409 P3_EAX_REG_9__SCAN_IN ; P3_U6788
g4968 nand P3_U6759 P3_DATAO_REG_9__SCAN_IN ; P3_U6789
g4969 nand P3_U2410 P3_LWORD_REG_10__SCAN_IN ; P3_U6790
g4970 nand P3_U2409 P3_EAX_REG_10__SCAN_IN ; P3_U6791
g4971 nand P3_U6759 P3_DATAO_REG_10__SCAN_IN ; P3_U6792
g4972 nand P3_U2410 P3_LWORD_REG_11__SCAN_IN ; P3_U6793
g4973 nand P3_U2409 P3_EAX_REG_11__SCAN_IN ; P3_U6794
g4974 nand P3_U6759 P3_DATAO_REG_11__SCAN_IN ; P3_U6795
g4975 nand P3_U2410 P3_LWORD_REG_12__SCAN_IN ; P3_U6796
g4976 nand P3_U2409 P3_EAX_REG_12__SCAN_IN ; P3_U6797
g4977 nand P3_U6759 P3_DATAO_REG_12__SCAN_IN ; P3_U6798
g4978 nand P3_U2410 P3_LWORD_REG_13__SCAN_IN ; P3_U6799
g4979 nand P3_U2409 P3_EAX_REG_13__SCAN_IN ; P3_U6800
g4980 nand P3_U6759 P3_DATAO_REG_13__SCAN_IN ; P3_U6801
g4981 nand P3_U2410 P3_LWORD_REG_14__SCAN_IN ; P3_U6802
g4982 nand P3_U2409 P3_EAX_REG_14__SCAN_IN ; P3_U6803
g4983 nand P3_U6759 P3_DATAO_REG_14__SCAN_IN ; P3_U6804
g4984 nand P3_U2410 P3_LWORD_REG_15__SCAN_IN ; P3_U6805
g4985 nand P3_U2409 P3_EAX_REG_15__SCAN_IN ; P3_U6806
g4986 nand P3_U6759 P3_DATAO_REG_15__SCAN_IN ; P3_U6807
g4987 nand P3_U2447 P3_EAX_REG_16__SCAN_IN ; P3_U6808
g4988 nand P3_U2410 P3_UWORD_REG_0__SCAN_IN ; P3_U6809
g4989 nand P3_U6759 P3_DATAO_REG_16__SCAN_IN ; P3_U6810
g4990 nand P3_U2447 P3_EAX_REG_17__SCAN_IN ; P3_U6811
g4991 nand P3_U2410 P3_UWORD_REG_1__SCAN_IN ; P3_U6812
g4992 nand P3_U6759 P3_DATAO_REG_17__SCAN_IN ; P3_U6813
g4993 nand P3_U2447 P3_EAX_REG_18__SCAN_IN ; P3_U6814
g4994 nand P3_U2410 P3_UWORD_REG_2__SCAN_IN ; P3_U6815
g4995 nand P3_U6759 P3_DATAO_REG_18__SCAN_IN ; P3_U6816
g4996 nand P3_U2447 P3_EAX_REG_19__SCAN_IN ; P3_U6817
g4997 nand P3_U2410 P3_UWORD_REG_3__SCAN_IN ; P3_U6818
g4998 nand P3_U6759 P3_DATAO_REG_19__SCAN_IN ; P3_U6819
g4999 nand P3_U2447 P3_EAX_REG_20__SCAN_IN ; P3_U6820
g5000 nand P3_U2410 P3_UWORD_REG_4__SCAN_IN ; P3_U6821
g5001 nand P3_U6759 P3_DATAO_REG_20__SCAN_IN ; P3_U6822
g5002 nand P3_U2447 P3_EAX_REG_21__SCAN_IN ; P3_U6823
g5003 nand P3_U2410 P3_UWORD_REG_5__SCAN_IN ; P3_U6824
g5004 nand P3_U6759 P3_DATAO_REG_21__SCAN_IN ; P3_U6825
g5005 nand P3_U2447 P3_EAX_REG_22__SCAN_IN ; P3_U6826
g5006 nand P3_U2410 P3_UWORD_REG_6__SCAN_IN ; P3_U6827
g5007 nand P3_U6759 P3_DATAO_REG_22__SCAN_IN ; P3_U6828
g5008 nand P3_U2447 P3_EAX_REG_23__SCAN_IN ; P3_U6829
g5009 nand P3_U2410 P3_UWORD_REG_7__SCAN_IN ; P3_U6830
g5010 nand P3_U6759 P3_DATAO_REG_23__SCAN_IN ; P3_U6831
g5011 nand P3_U2447 P3_EAX_REG_24__SCAN_IN ; P3_U6832
g5012 nand P3_U2410 P3_UWORD_REG_8__SCAN_IN ; P3_U6833
g5013 nand P3_U6759 P3_DATAO_REG_24__SCAN_IN ; P3_U6834
g5014 nand P3_U2447 P3_EAX_REG_25__SCAN_IN ; P3_U6835
g5015 nand P3_U2410 P3_UWORD_REG_9__SCAN_IN ; P3_U6836
g5016 nand P3_U6759 P3_DATAO_REG_25__SCAN_IN ; P3_U6837
g5017 nand P3_U2447 P3_EAX_REG_26__SCAN_IN ; P3_U6838
g5018 nand P3_U2410 P3_UWORD_REG_10__SCAN_IN ; P3_U6839
g5019 nand P3_U6759 P3_DATAO_REG_26__SCAN_IN ; P3_U6840
g5020 nand P3_U2447 P3_EAX_REG_27__SCAN_IN ; P3_U6841
g5021 nand P3_U2410 P3_UWORD_REG_11__SCAN_IN ; P3_U6842
g5022 nand P3_U6759 P3_DATAO_REG_27__SCAN_IN ; P3_U6843
g5023 nand P3_U2447 P3_EAX_REG_28__SCAN_IN ; P3_U6844
g5024 nand P3_U2410 P3_UWORD_REG_12__SCAN_IN ; P3_U6845
g5025 nand P3_U6759 P3_DATAO_REG_28__SCAN_IN ; P3_U6846
g5026 nand P3_U2447 P3_EAX_REG_29__SCAN_IN ; P3_U6847
g5027 nand P3_U2410 P3_UWORD_REG_13__SCAN_IN ; P3_U6848
g5028 nand P3_U6759 P3_DATAO_REG_29__SCAN_IN ; P3_U6849
g5029 nand P3_U2447 P3_EAX_REG_30__SCAN_IN ; P3_U6850
g5030 nand P3_U2410 P3_UWORD_REG_14__SCAN_IN ; P3_U6851
g5031 nand P3_U6759 P3_DATAO_REG_30__SCAN_IN ; P3_U6852
g5032 nand P3_U2516 P3_U3243 ; P3_U6853
g5033 nand P3_U2446 BUF2_REG_0__SCAN_IN ; P3_U6854
g5034 nand P3_U2621 P3_U2411 ; P3_U6855
g5035 nand P3_ADD_546_U5 P3_U2400 ; P3_U6856
g5036 nand P3_U3252 P3_EAX_REG_0__SCAN_IN ; P3_U6857
g5037 nand P3_U2446 BUF2_REG_1__SCAN_IN ; P3_U6858
g5038 nand P3_U2622 P3_U2411 ; P3_U6859
g5039 nand P3_ADD_546_U71 P3_U2400 ; P3_U6860
g5040 nand P3_U3252 P3_EAX_REG_1__SCAN_IN ; P3_U6861
g5041 nand P3_U2446 BUF2_REG_2__SCAN_IN ; P3_U6862
g5042 nand P3_U2623 P3_U2411 ; P3_U6863
g5043 nand P3_ADD_546_U60 P3_U2400 ; P3_U6864
g5044 nand P3_U3252 P3_EAX_REG_2__SCAN_IN ; P3_U6865
g5045 nand P3_U2446 BUF2_REG_3__SCAN_IN ; P3_U6866
g5046 nand P3_U2624 P3_U2411 ; P3_U6867
g5047 nand P3_ADD_546_U57 P3_U2400 ; P3_U6868
g5048 nand P3_U3252 P3_EAX_REG_3__SCAN_IN ; P3_U6869
g5049 nand P3_U2446 BUF2_REG_4__SCAN_IN ; P3_U6870
g5050 nand P3_U2625 P3_U2411 ; P3_U6871
g5051 nand P3_ADD_546_U56 P3_U2400 ; P3_U6872
g5052 nand P3_U3252 P3_EAX_REG_4__SCAN_IN ; P3_U6873
g5053 nand P3_U2446 BUF2_REG_5__SCAN_IN ; P3_U6874
g5054 nand P3_U2626 P3_U2411 ; P3_U6875
g5055 nand P3_ADD_546_U55 P3_U2400 ; P3_U6876
g5056 nand P3_U3252 P3_EAX_REG_5__SCAN_IN ; P3_U6877
g5057 nand P3_U2446 BUF2_REG_6__SCAN_IN ; P3_U6878
g5058 nand P3_U2627 P3_U2411 ; P3_U6879
g5059 nand P3_ADD_546_U54 P3_U2400 ; P3_U6880
g5060 nand P3_U3252 P3_EAX_REG_6__SCAN_IN ; P3_U6881
g5061 nand P3_U2446 BUF2_REG_7__SCAN_IN ; P3_U6882
g5062 nand P3_U2628 P3_U2411 ; P3_U6883
g5063 nand P3_ADD_546_U53 P3_U2400 ; P3_U6884
g5064 nand P3_U3252 P3_EAX_REG_7__SCAN_IN ; P3_U6885
g5065 nand P3_U2446 BUF2_REG_8__SCAN_IN ; P3_U6886
g5066 nand P3_U2605 P3_U2411 ; P3_U6887
g5067 nand P3_ADD_546_U52 P3_U2400 ; P3_U6888
g5068 nand P3_U3252 P3_EAX_REG_8__SCAN_IN ; P3_U6889
g5069 nand P3_U2446 BUF2_REG_9__SCAN_IN ; P3_U6890
g5070 nand P3_U2606 P3_U2411 ; P3_U6891
g5071 nand P3_ADD_546_U51 P3_U2400 ; P3_U6892
g5072 nand P3_U3252 P3_EAX_REG_9__SCAN_IN ; P3_U6893
g5073 nand P3_U2446 BUF2_REG_10__SCAN_IN ; P3_U6894
g5074 nand P3_U2607 P3_U2411 ; P3_U6895
g5075 nand P3_ADD_546_U81 P3_U2400 ; P3_U6896
g5076 nand P3_U3252 P3_EAX_REG_10__SCAN_IN ; P3_U6897
g5077 nand P3_U2446 BUF2_REG_11__SCAN_IN ; P3_U6898
g5078 nand P3_U2608 P3_U2411 ; P3_U6899
g5079 nand P3_ADD_546_U80 P3_U2400 ; P3_U6900
g5080 nand P3_U3252 P3_EAX_REG_11__SCAN_IN ; P3_U6901
g5081 nand P3_U2446 BUF2_REG_12__SCAN_IN ; P3_U6902
g5082 nand P3_U2609 P3_U2411 ; P3_U6903
g5083 nand P3_ADD_546_U79 P3_U2400 ; P3_U6904
g5084 nand P3_U3252 P3_EAX_REG_12__SCAN_IN ; P3_U6905
g5085 nand P3_U2446 BUF2_REG_13__SCAN_IN ; P3_U6906
g5086 nand P3_U2610 P3_U2411 ; P3_U6907
g5087 nand P3_ADD_546_U78 P3_U2400 ; P3_U6908
g5088 nand P3_U3252 P3_EAX_REG_13__SCAN_IN ; P3_U6909
g5089 nand P3_U2446 BUF2_REG_14__SCAN_IN ; P3_U6910
g5090 nand P3_U2611 P3_U2411 ; P3_U6911
g5091 nand P3_ADD_546_U77 P3_U2400 ; P3_U6912
g5092 nand P3_U3252 P3_EAX_REG_14__SCAN_IN ; P3_U6913
g5093 nand P3_U2446 BUF2_REG_15__SCAN_IN ; P3_U6914
g5094 nand P3_U2612 P3_U2411 ; P3_U6915
g5095 nand P3_ADD_546_U76 P3_U2400 ; P3_U6916
g5096 nand P3_U3252 P3_EAX_REG_15__SCAN_IN ; P3_U6917
g5097 nand P3_U2448 BUF2_REG_0__SCAN_IN ; P3_U6918
g5098 nand P3_U2444 BUF2_REG_16__SCAN_IN ; P3_U6919
g5099 nand P3_U3062 P3_U2411 ; P3_U6920
g5100 nand P3_ADD_546_U75 P3_U2400 ; P3_U6921
g5101 nand P3_U3252 P3_EAX_REG_16__SCAN_IN ; P3_U6922
g5102 nand P3_U2448 BUF2_REG_1__SCAN_IN ; P3_U6923
g5103 nand P3_U2444 BUF2_REG_17__SCAN_IN ; P3_U6924
g5104 nand P3_U3063 P3_U2411 ; P3_U6925
g5105 nand P3_ADD_546_U74 P3_U2400 ; P3_U6926
g5106 nand P3_U3252 P3_EAX_REG_17__SCAN_IN ; P3_U6927
g5107 nand P3_U2448 BUF2_REG_2__SCAN_IN ; P3_U6928
g5108 nand P3_U2444 BUF2_REG_18__SCAN_IN ; P3_U6929
g5109 nand P3_U3064 P3_U2411 ; P3_U6930
g5110 nand P3_ADD_546_U73 P3_U2400 ; P3_U6931
g5111 nand P3_U3252 P3_EAX_REG_18__SCAN_IN ; P3_U6932
g5112 nand P3_U2448 BUF2_REG_3__SCAN_IN ; P3_U6933
g5113 nand P3_U2444 BUF2_REG_19__SCAN_IN ; P3_U6934
g5114 nand P3_U3065 P3_U2411 ; P3_U6935
g5115 nand P3_ADD_546_U72 P3_U2400 ; P3_U6936
g5116 nand P3_U3252 P3_EAX_REG_19__SCAN_IN ; P3_U6937
g5117 nand P3_U2448 BUF2_REG_4__SCAN_IN ; P3_U6938
g5118 nand P3_U2444 BUF2_REG_20__SCAN_IN ; P3_U6939
g5119 nand P3_U3066 P3_U2411 ; P3_U6940
g5120 nand P3_ADD_546_U70 P3_U2400 ; P3_U6941
g5121 nand P3_U3252 P3_EAX_REG_20__SCAN_IN ; P3_U6942
g5122 nand P3_U2448 BUF2_REG_5__SCAN_IN ; P3_U6943
g5123 nand P3_U2444 BUF2_REG_21__SCAN_IN ; P3_U6944
g5124 nand P3_U3067 P3_U2411 ; P3_U6945
g5125 nand P3_ADD_546_U69 P3_U2400 ; P3_U6946
g5126 nand P3_U3252 P3_EAX_REG_21__SCAN_IN ; P3_U6947
g5127 nand P3_U2448 BUF2_REG_6__SCAN_IN ; P3_U6948
g5128 nand P3_U2444 BUF2_REG_22__SCAN_IN ; P3_U6949
g5129 nand P3_U3068 P3_U2411 ; P3_U6950
g5130 nand P3_ADD_546_U68 P3_U2400 ; P3_U6951
g5131 nand P3_U3252 P3_EAX_REG_22__SCAN_IN ; P3_U6952
g5132 nand P3_U2448 BUF2_REG_7__SCAN_IN ; P3_U6953
g5133 nand P3_U2444 BUF2_REG_23__SCAN_IN ; P3_U6954
g5134 nand P3_ADD_391_1180_U25 P3_U2411 ; P3_U6955
g5135 nand P3_ADD_546_U67 P3_U2400 ; P3_U6956
g5136 nand P3_U3252 P3_EAX_REG_23__SCAN_IN ; P3_U6957
g5137 nand P3_U2448 BUF2_REG_8__SCAN_IN ; P3_U6958
g5138 nand P3_U2444 BUF2_REG_24__SCAN_IN ; P3_U6959
g5139 nand P3_ADD_391_1180_U24 P3_U2411 ; P3_U6960
g5140 nand P3_ADD_546_U66 P3_U2400 ; P3_U6961
g5141 nand P3_U3252 P3_EAX_REG_24__SCAN_IN ; P3_U6962
g5142 nand P3_U2448 BUF2_REG_9__SCAN_IN ; P3_U6963
g5143 nand P3_U2444 BUF2_REG_25__SCAN_IN ; P3_U6964
g5144 nand P3_ADD_391_1180_U23 P3_U2411 ; P3_U6965
g5145 nand P3_ADD_546_U65 P3_U2400 ; P3_U6966
g5146 nand P3_U3252 P3_EAX_REG_25__SCAN_IN ; P3_U6967
g5147 nand P3_U2448 BUF2_REG_10__SCAN_IN ; P3_U6968
g5148 nand P3_U2444 BUF2_REG_26__SCAN_IN ; P3_U6969
g5149 nand P3_ADD_391_1180_U22 P3_U2411 ; P3_U6970
g5150 nand P3_ADD_546_U64 P3_U2400 ; P3_U6971
g5151 nand P3_U3252 P3_EAX_REG_26__SCAN_IN ; P3_U6972
g5152 nand P3_U2448 BUF2_REG_11__SCAN_IN ; P3_U6973
g5153 nand P3_U2444 BUF2_REG_27__SCAN_IN ; P3_U6974
g5154 nand P3_ADD_391_1180_U21 P3_U2411 ; P3_U6975
g5155 nand P3_ADD_546_U63 P3_U2400 ; P3_U6976
g5156 nand P3_U3252 P3_EAX_REG_27__SCAN_IN ; P3_U6977
g5157 nand P3_U2448 BUF2_REG_12__SCAN_IN ; P3_U6978
g5158 nand P3_U2444 BUF2_REG_28__SCAN_IN ; P3_U6979
g5159 nand P3_ADD_391_1180_U20 P3_U2411 ; P3_U6980
g5160 nand P3_ADD_546_U62 P3_U2400 ; P3_U6981
g5161 nand P3_U3252 P3_EAX_REG_28__SCAN_IN ; P3_U6982
g5162 nand P3_U2448 BUF2_REG_13__SCAN_IN ; P3_U6983
g5163 nand P3_U2444 BUF2_REG_29__SCAN_IN ; P3_U6984
g5164 nand P3_ADD_391_1180_U19 P3_U2411 ; P3_U6985
g5165 nand P3_ADD_546_U61 P3_U2400 ; P3_U6986
g5166 nand P3_U3252 P3_EAX_REG_29__SCAN_IN ; P3_U6987
g5167 nand P3_U2448 BUF2_REG_14__SCAN_IN ; P3_U6988
g5168 nand P3_U2444 BUF2_REG_30__SCAN_IN ; P3_U6989
g5169 nand P3_ADD_391_1180_U18 P3_U2411 ; P3_U6990
g5170 nand P3_ADD_546_U59 P3_U2400 ; P3_U6991
g5171 nand P3_U3252 P3_EAX_REG_30__SCAN_IN ; P3_U6992
g5172 nand P3_U2444 BUF2_REG_31__SCAN_IN ; P3_U6993
g5173 nand P3_ADD_546_U58 P3_U2400 ; P3_U6994
g5174 nand P3_U3252 P3_EAX_REG_31__SCAN_IN ; P3_U6995
g5175 nand P3_GTE_401_U6 P3_U4305 ; P3_U6996
g5176 nand P3_U3242 P3_U6996 ; P3_U6997
g5177 nand P3_U2408 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U6998
g5178 nand P3_ADD_552_U5 P3_U2399 ; P3_U6999
g5179 nand P3_U3253 P3_EBX_REG_0__SCAN_IN ; P3_U7000
g5180 nand P3_U2408 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U7001
g5181 nand P3_ADD_552_U71 P3_U2399 ; P3_U7002
g5182 nand P3_U3253 P3_EBX_REG_1__SCAN_IN ; P3_U7003
g5183 nand P3_U2408 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U7004
g5184 nand P3_ADD_552_U60 P3_U2399 ; P3_U7005
g5185 nand P3_U3253 P3_EBX_REG_2__SCAN_IN ; P3_U7006
g5186 nand P3_U2408 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U7007
g5187 nand P3_ADD_552_U57 P3_U2399 ; P3_U7008
g5188 nand P3_U3253 P3_EBX_REG_3__SCAN_IN ; P3_U7009
g5189 nand P3_U2408 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U7010
g5190 nand P3_ADD_552_U56 P3_U2399 ; P3_U7011
g5191 nand P3_U3253 P3_EBX_REG_4__SCAN_IN ; P3_U7012
g5192 nand P3_U2408 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U7013
g5193 nand P3_ADD_552_U55 P3_U2399 ; P3_U7014
g5194 nand P3_U3253 P3_EBX_REG_5__SCAN_IN ; P3_U7015
g5195 nand P3_U2408 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U7016
g5196 nand P3_ADD_552_U54 P3_U2399 ; P3_U7017
g5197 nand P3_U3253 P3_EBX_REG_6__SCAN_IN ; P3_U7018
g5198 nand P3_U2408 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U7019
g5199 nand P3_ADD_552_U53 P3_U2399 ; P3_U7020
g5200 nand P3_U3253 P3_EBX_REG_7__SCAN_IN ; P3_U7021
g5201 nand P3_U2605 P3_U2408 ; P3_U7022
g5202 nand P3_ADD_552_U52 P3_U2399 ; P3_U7023
g5203 nand P3_U3253 P3_EBX_REG_8__SCAN_IN ; P3_U7024
g5204 nand P3_U2606 P3_U2408 ; P3_U7025
g5205 nand P3_ADD_552_U51 P3_U2399 ; P3_U7026
g5206 nand P3_U3253 P3_EBX_REG_9__SCAN_IN ; P3_U7027
g5207 nand P3_U2607 P3_U2408 ; P3_U7028
g5208 nand P3_ADD_552_U81 P3_U2399 ; P3_U7029
g5209 nand P3_U3253 P3_EBX_REG_10__SCAN_IN ; P3_U7030
g5210 nand P3_U2608 P3_U2408 ; P3_U7031
g5211 nand P3_ADD_552_U80 P3_U2399 ; P3_U7032
g5212 nand P3_U3253 P3_EBX_REG_11__SCAN_IN ; P3_U7033
g5213 nand P3_U2609 P3_U2408 ; P3_U7034
g5214 nand P3_ADD_552_U79 P3_U2399 ; P3_U7035
g5215 nand P3_U3253 P3_EBX_REG_12__SCAN_IN ; P3_U7036
g5216 nand P3_U2610 P3_U2408 ; P3_U7037
g5217 nand P3_ADD_552_U78 P3_U2399 ; P3_U7038
g5218 nand P3_U3253 P3_EBX_REG_13__SCAN_IN ; P3_U7039
g5219 nand P3_U2611 P3_U2408 ; P3_U7040
g5220 nand P3_ADD_552_U77 P3_U2399 ; P3_U7041
g5221 nand P3_U3253 P3_EBX_REG_14__SCAN_IN ; P3_U7042
g5222 nand P3_U2612 P3_U2408 ; P3_U7043
g5223 nand P3_ADD_552_U76 P3_U2399 ; P3_U7044
g5224 nand P3_U3253 P3_EBX_REG_15__SCAN_IN ; P3_U7045
g5225 nand P3_U3062 P3_U2408 ; P3_U7046
g5226 nand P3_ADD_552_U75 P3_U2399 ; P3_U7047
g5227 nand P3_U3253 P3_EBX_REG_16__SCAN_IN ; P3_U7048
g5228 nand P3_U3063 P3_U2408 ; P3_U7049
g5229 nand P3_ADD_552_U74 P3_U2399 ; P3_U7050
g5230 nand P3_U3253 P3_EBX_REG_17__SCAN_IN ; P3_U7051
g5231 nand P3_U3064 P3_U2408 ; P3_U7052
g5232 nand P3_ADD_552_U73 P3_U2399 ; P3_U7053
g5233 nand P3_U3253 P3_EBX_REG_18__SCAN_IN ; P3_U7054
g5234 nand P3_U3065 P3_U2408 ; P3_U7055
g5235 nand P3_ADD_552_U72 P3_U2399 ; P3_U7056
g5236 nand P3_U3253 P3_EBX_REG_19__SCAN_IN ; P3_U7057
g5237 nand P3_U3066 P3_U2408 ; P3_U7058
g5238 nand P3_ADD_552_U70 P3_U2399 ; P3_U7059
g5239 nand P3_U3253 P3_EBX_REG_20__SCAN_IN ; P3_U7060
g5240 nand P3_U3067 P3_U2408 ; P3_U7061
g5241 nand P3_ADD_552_U69 P3_U2399 ; P3_U7062
g5242 nand P3_U3253 P3_EBX_REG_21__SCAN_IN ; P3_U7063
g5243 nand P3_U3068 P3_U2408 ; P3_U7064
g5244 nand P3_ADD_552_U68 P3_U2399 ; P3_U7065
g5245 nand P3_U3253 P3_EBX_REG_22__SCAN_IN ; P3_U7066
g5246 nand P3_ADD_402_1132_U25 P3_U2408 ; P3_U7067
g5247 nand P3_ADD_552_U67 P3_U2399 ; P3_U7068
g5248 nand P3_U3253 P3_EBX_REG_23__SCAN_IN ; P3_U7069
g5249 nand P3_ADD_402_1132_U24 P3_U2408 ; P3_U7070
g5250 nand P3_ADD_552_U66 P3_U2399 ; P3_U7071
g5251 nand P3_U3253 P3_EBX_REG_24__SCAN_IN ; P3_U7072
g5252 nand P3_ADD_402_1132_U23 P3_U2408 ; P3_U7073
g5253 nand P3_ADD_552_U65 P3_U2399 ; P3_U7074
g5254 nand P3_U3253 P3_EBX_REG_25__SCAN_IN ; P3_U7075
g5255 nand P3_ADD_402_1132_U22 P3_U2408 ; P3_U7076
g5256 nand P3_ADD_552_U64 P3_U2399 ; P3_U7077
g5257 nand P3_U3253 P3_EBX_REG_26__SCAN_IN ; P3_U7078
g5258 nand P3_ADD_402_1132_U21 P3_U2408 ; P3_U7079
g5259 nand P3_ADD_552_U63 P3_U2399 ; P3_U7080
g5260 nand P3_U3253 P3_EBX_REG_27__SCAN_IN ; P3_U7081
g5261 nand P3_ADD_402_1132_U20 P3_U2408 ; P3_U7082
g5262 nand P3_ADD_552_U62 P3_U2399 ; P3_U7083
g5263 nand P3_U3253 P3_EBX_REG_28__SCAN_IN ; P3_U7084
g5264 nand P3_ADD_402_1132_U19 P3_U2408 ; P3_U7085
g5265 nand P3_ADD_552_U61 P3_U2399 ; P3_U7086
g5266 nand P3_U3253 P3_EBX_REG_29__SCAN_IN ; P3_U7087
g5267 nand P3_ADD_402_1132_U18 P3_U2408 ; P3_U7088
g5268 nand P3_ADD_552_U59 P3_U2399 ; P3_U7089
g5269 nand P3_U3253 P3_EBX_REG_30__SCAN_IN ; P3_U7090
g5270 nand P3_ADD_552_U58 P3_U2399 ; P3_U7091
g5271 nand P3_U3253 P3_EBX_REG_31__SCAN_IN ; P3_U7092
g5272 nand P3_U5488 P3_U5491 ; P3_U7093
g5273 not P3_U3260 ; P3_U7094
g5274 not P3_U3257 ; P3_U7095
g5275 or U209 P3_STATEBS16_REG_SCAN_IN ; P3_U7096
g5276 nand P3_U2602 P3_EBX_REG_0__SCAN_IN ; P3_U7097
g5277 nand P3_U2601 P3_REIP_REG_0__SCAN_IN ; P3_U7098
g5278 nand P3_U7910 P3_EBX_REG_0__SCAN_IN ; P3_U7099
g5279 nand P3_ADD_505_U5 P3_U2455 ; P3_U7100
g5280 nand P3_ADD_486_U5 P3_U2454 ; P3_U7101
g5281 nand P3_U2405 P3_REIP_REG_0__SCAN_IN ; P3_U7102
g5282 nand P3_U2403 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U7103
g5283 nand P3_U4319 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U7104
g5284 nand P3_U2401 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_U7105
g5285 nand P3_U7094 P3_REIP_REG_0__SCAN_IN ; P3_U7106
g5286 nand P3_SUB_414_U50 P3_U2602 ; P3_U7107
g5287 nand P3_ADD_467_U4 P3_U2601 ; P3_U7108
g5288 nand P3_U7910 P3_EBX_REG_1__SCAN_IN ; P3_U7109
g5289 nand P3_ADD_505_U17 P3_U2455 ; P3_U7110
g5290 nand P3_ADD_486_U17 P3_U2454 ; P3_U7111
g5291 nand P3_ADD_430_U4 P3_U2405 ; P3_U7112
g5292 nand P3_U2403 P3_ADD_318_U4 ; P3_U7113
g5293 nand P3_SUB_320_U50 P3_U4319 ; P3_U7114
g5294 nand P3_U2401 P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_U7115
g5295 nand P3_U7094 P3_REIP_REG_1__SCAN_IN ; P3_U7116
g5296 nand P3_SUB_414_U17 P3_U2602 ; P3_U7117
g5297 nand P3_ADD_467_U71 P3_U2601 ; P3_U7118
g5298 nand P3_U7910 P3_EBX_REG_2__SCAN_IN ; P3_U7119
g5299 nand P3_ADD_505_U16 P3_U2455 ; P3_U7120
g5300 nand P3_ADD_486_U16 P3_U2454 ; P3_U7121
g5301 nand P3_ADD_430_U71 P3_U2405 ; P3_U7122
g5302 nand P3_U2403 P3_ADD_318_U71 ; P3_U7123
g5303 nand P3_SUB_320_U17 P3_U4319 ; P3_U7124
g5304 nand P3_U2401 P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_U7125
g5305 nand P3_U7094 P3_REIP_REG_2__SCAN_IN ; P3_U7126
g5306 nand P3_SUB_414_U59 P3_U2602 ; P3_U7127
g5307 nand P3_ADD_467_U68 P3_U2601 ; P3_U7128
g5308 nand P3_U7910 P3_EBX_REG_3__SCAN_IN ; P3_U7129
g5309 nand P3_ADD_505_U15 P3_U2455 ; P3_U7130
g5310 nand P3_ADD_486_U15 P3_U2454 ; P3_U7131
g5311 nand P3_ADD_430_U68 P3_U2405 ; P3_U7132
g5312 nand P3_U2403 P3_ADD_318_U68 ; P3_U7133
g5313 nand P3_SUB_320_U59 P3_U4319 ; P3_U7134
g5314 nand P3_U2401 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_U7135
g5315 nand P3_U7094 P3_REIP_REG_3__SCAN_IN ; P3_U7136
g5316 nand P3_SUB_414_U18 P3_U2602 ; P3_U7137
g5317 nand P3_ADD_467_U67 P3_U2601 ; P3_U7138
g5318 nand P3_U7910 P3_EBX_REG_4__SCAN_IN ; P3_U7139
g5319 nand P3_ADD_505_U14 P3_U2455 ; P3_U7140
g5320 nand P3_ADD_486_U14 P3_U2454 ; P3_U7141
g5321 nand P3_ADD_430_U67 P3_U2405 ; P3_U7142
g5322 nand P3_U2403 P3_ADD_318_U67 ; P3_U7143
g5323 nand P3_SUB_320_U18 P3_U4319 ; P3_U7144
g5324 nand P3_U2401 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_U7145
g5325 nand P3_U7094 P3_REIP_REG_4__SCAN_IN ; P3_U7146
g5326 nand P3_SUB_414_U57 P3_U2602 ; P3_U7147
g5327 nand P3_ADD_467_U66 P3_U2601 ; P3_U7148
g5328 nand P3_U7910 P3_EBX_REG_5__SCAN_IN ; P3_U7149
g5329 nand P3_ADD_505_U6 P3_U2455 ; P3_U7150
g5330 nand P3_ADD_486_U6 P3_U2454 ; P3_U7151
g5331 nand P3_ADD_430_U66 P3_U2405 ; P3_U7152
g5332 nand P3_U2403 P3_ADD_318_U66 ; P3_U7153
g5333 nand P3_SUB_320_U57 P3_U4319 ; P3_U7154
g5334 nand P3_U2401 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_U7155
g5335 nand P3_U7094 P3_REIP_REG_5__SCAN_IN ; P3_U7156
g5336 nand P3_SUB_414_U19 P3_U2602 ; P3_U7157
g5337 nand P3_ADD_467_U65 P3_U2601 ; P3_U7158
g5338 nand P3_U7910 P3_EBX_REG_6__SCAN_IN ; P3_U7159
g5339 nand P3_ADD_430_U65 P3_U2405 ; P3_U7160
g5340 nand P3_U2403 P3_ADD_318_U65 ; P3_U7161
g5341 nand P3_SUB_320_U19 P3_U4319 ; P3_U7162
g5342 nand P3_U2401 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_U7163
g5343 nand P3_U7094 P3_REIP_REG_6__SCAN_IN ; P3_U7164
g5344 nand P3_SUB_414_U55 P3_U2602 ; P3_U7165
g5345 nand P3_ADD_467_U64 P3_U2601 ; P3_U7166
g5346 nand P3_U7910 P3_EBX_REG_7__SCAN_IN ; P3_U7167
g5347 nand P3_ADD_430_U64 P3_U2405 ; P3_U7168
g5348 nand P3_U2403 P3_ADD_318_U64 ; P3_U7169
g5349 nand P3_SUB_320_U55 P3_U4319 ; P3_U7170
g5350 nand P3_U2401 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_U7171
g5351 nand P3_U7094 P3_REIP_REG_7__SCAN_IN ; P3_U7172
g5352 nand P3_SUB_414_U20 P3_U2602 ; P3_U7173
g5353 nand P3_ADD_467_U63 P3_U2601 ; P3_U7174
g5354 nand P3_U7910 P3_EBX_REG_8__SCAN_IN ; P3_U7175
g5355 nand P3_ADD_430_U63 P3_U2405 ; P3_U7176
g5356 nand P3_U2403 P3_ADD_318_U63 ; P3_U7177
g5357 nand P3_SUB_320_U20 P3_U4319 ; P3_U7178
g5358 nand P3_U2401 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_U7179
g5359 nand P3_U7094 P3_REIP_REG_8__SCAN_IN ; P3_U7180
g5360 nand P3_SUB_414_U53 P3_U2602 ; P3_U7181
g5361 nand P3_ADD_467_U62 P3_U2601 ; P3_U7182
g5362 nand P3_U7910 P3_EBX_REG_9__SCAN_IN ; P3_U7183
g5363 nand P3_ADD_430_U62 P3_U2405 ; P3_U7184
g5364 nand P3_U2403 P3_ADD_318_U62 ; P3_U7185
g5365 nand P3_SUB_320_U53 P3_U4319 ; P3_U7186
g5366 nand P3_U2401 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_U7187
g5367 nand P3_U7094 P3_REIP_REG_9__SCAN_IN ; P3_U7188
g5368 nand P3_SUB_414_U6 P3_U2602 ; P3_U7189
g5369 nand P3_ADD_467_U91 P3_U2601 ; P3_U7190
g5370 nand P3_U7910 P3_EBX_REG_10__SCAN_IN ; P3_U7191
g5371 nand P3_ADD_430_U91 P3_U2405 ; P3_U7192
g5372 nand P3_U2403 P3_ADD_318_U91 ; P3_U7193
g5373 nand P3_SUB_320_U6 P3_U4319 ; P3_U7194
g5374 nand P3_U2401 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_U7195
g5375 nand P3_U7094 P3_REIP_REG_10__SCAN_IN ; P3_U7196
g5376 nand P3_SUB_414_U82 P3_U2602 ; P3_U7197
g5377 nand P3_ADD_467_U90 P3_U2601 ; P3_U7198
g5378 nand P3_U7910 P3_EBX_REG_11__SCAN_IN ; P3_U7199
g5379 nand P3_ADD_430_U90 P3_U2405 ; P3_U7200
g5380 nand P3_U2403 P3_ADD_318_U90 ; P3_U7201
g5381 nand P3_SUB_320_U82 P3_U4319 ; P3_U7202
g5382 nand P3_U2401 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_U7203
g5383 nand P3_U7094 P3_REIP_REG_11__SCAN_IN ; P3_U7204
g5384 nand P3_SUB_414_U7 P3_U2602 ; P3_U7205
g5385 nand P3_ADD_467_U89 P3_U2601 ; P3_U7206
g5386 nand P3_U7910 P3_EBX_REG_12__SCAN_IN ; P3_U7207
g5387 nand P3_ADD_430_U89 P3_U2405 ; P3_U7208
g5388 nand P3_U2403 P3_ADD_318_U89 ; P3_U7209
g5389 nand P3_SUB_320_U7 P3_U4319 ; P3_U7210
g5390 nand P3_U2401 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_U7211
g5391 nand P3_U7094 P3_REIP_REG_12__SCAN_IN ; P3_U7212
g5392 nand P3_SUB_414_U80 P3_U2602 ; P3_U7213
g5393 nand P3_ADD_467_U88 P3_U2601 ; P3_U7214
g5394 nand P3_U7910 P3_EBX_REG_13__SCAN_IN ; P3_U7215
g5395 nand P3_ADD_430_U88 P3_U2405 ; P3_U7216
g5396 nand P3_U2403 P3_ADD_318_U88 ; P3_U7217
g5397 nand P3_SUB_320_U80 P3_U4319 ; P3_U7218
g5398 nand P3_U2401 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_U7219
g5399 nand P3_U7094 P3_REIP_REG_13__SCAN_IN ; P3_U7220
g5400 nand P3_SUB_414_U8 P3_U2602 ; P3_U7221
g5401 nand P3_ADD_467_U87 P3_U2601 ; P3_U7222
g5402 nand P3_U7910 P3_EBX_REG_14__SCAN_IN ; P3_U7223
g5403 nand P3_ADD_430_U87 P3_U2405 ; P3_U7224
g5404 nand P3_U2403 P3_ADD_318_U87 ; P3_U7225
g5405 nand P3_SUB_320_U8 P3_U4319 ; P3_U7226
g5406 nand P3_U2401 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_U7227
g5407 nand P3_U7094 P3_REIP_REG_14__SCAN_IN ; P3_U7228
g5408 nand P3_SUB_414_U78 P3_U2602 ; P3_U7229
g5409 nand P3_ADD_467_U86 P3_U2601 ; P3_U7230
g5410 nand P3_U7910 P3_EBX_REG_15__SCAN_IN ; P3_U7231
g5411 nand P3_ADD_430_U86 P3_U2405 ; P3_U7232
g5412 nand P3_U2403 P3_ADD_318_U86 ; P3_U7233
g5413 nand P3_SUB_320_U78 P3_U4319 ; P3_U7234
g5414 nand P3_U2401 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_U7235
g5415 nand P3_U7094 P3_REIP_REG_15__SCAN_IN ; P3_U7236
g5416 nand P3_SUB_414_U9 P3_U2602 ; P3_U7237
g5417 nand P3_ADD_467_U85 P3_U2601 ; P3_U7238
g5418 nand P3_U7910 P3_EBX_REG_16__SCAN_IN ; P3_U7239
g5419 nand P3_ADD_430_U85 P3_U2405 ; P3_U7240
g5420 nand P3_U2403 P3_ADD_318_U85 ; P3_U7241
g5421 nand P3_SUB_320_U9 P3_U4319 ; P3_U7242
g5422 nand P3_U2401 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_U7243
g5423 nand P3_U7094 P3_REIP_REG_16__SCAN_IN ; P3_U7244
g5424 nand P3_SUB_414_U76 P3_U2602 ; P3_U7245
g5425 nand P3_ADD_467_U84 P3_U2601 ; P3_U7246
g5426 nand P3_U7910 P3_EBX_REG_17__SCAN_IN ; P3_U7247
g5427 nand P3_ADD_430_U84 P3_U2405 ; P3_U7248
g5428 nand P3_U2403 P3_ADD_318_U84 ; P3_U7249
g5429 nand P3_SUB_320_U76 P3_U4319 ; P3_U7250
g5430 nand P3_U2401 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_U7251
g5431 nand P3_U7094 P3_REIP_REG_17__SCAN_IN ; P3_U7252
g5432 nand P3_SUB_414_U10 P3_U2602 ; P3_U7253
g5433 nand P3_ADD_467_U83 P3_U2601 ; P3_U7254
g5434 nand P3_U7910 P3_EBX_REG_18__SCAN_IN ; P3_U7255
g5435 nand P3_ADD_430_U83 P3_U2405 ; P3_U7256
g5436 nand P3_U2403 P3_ADD_318_U83 ; P3_U7257
g5437 nand P3_SUB_320_U10 P3_U4319 ; P3_U7258
g5438 nand P3_U2401 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_U7259
g5439 nand P3_U7094 P3_REIP_REG_18__SCAN_IN ; P3_U7260
g5440 nand P3_SUB_414_U74 P3_U2602 ; P3_U7261
g5441 nand P3_ADD_467_U82 P3_U2601 ; P3_U7262
g5442 nand P3_U7910 P3_EBX_REG_19__SCAN_IN ; P3_U7263
g5443 nand P3_ADD_430_U82 P3_U2405 ; P3_U7264
g5444 nand P3_U2403 P3_ADD_318_U82 ; P3_U7265
g5445 nand P3_SUB_320_U74 P3_U4319 ; P3_U7266
g5446 nand P3_U2401 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_U7267
g5447 nand P3_U7094 P3_REIP_REG_19__SCAN_IN ; P3_U7268
g5448 nand P3_SUB_414_U11 P3_U2602 ; P3_U7269
g5449 nand P3_ADD_467_U81 P3_U2601 ; P3_U7270
g5450 nand P3_U7910 P3_EBX_REG_20__SCAN_IN ; P3_U7271
g5451 nand P3_ADD_430_U81 P3_U2405 ; P3_U7272
g5452 nand P3_U2403 P3_ADD_318_U81 ; P3_U7273
g5453 nand P3_SUB_320_U11 P3_U4319 ; P3_U7274
g5454 nand P3_U2401 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_U7275
g5455 nand P3_U7094 P3_REIP_REG_20__SCAN_IN ; P3_U7276
g5456 nand P3_SUB_414_U70 P3_U2602 ; P3_U7277
g5457 nand P3_ADD_467_U80 P3_U2601 ; P3_U7278
g5458 nand P3_U7910 P3_EBX_REG_21__SCAN_IN ; P3_U7279
g5459 nand P3_ADD_430_U80 P3_U2405 ; P3_U7280
g5460 nand P3_U2403 P3_ADD_318_U80 ; P3_U7281
g5461 nand P3_SUB_320_U70 P3_U4319 ; P3_U7282
g5462 nand P3_U2401 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_U7283
g5463 nand P3_U7094 P3_REIP_REG_21__SCAN_IN ; P3_U7284
g5464 nand P3_SUB_414_U12 P3_U2602 ; P3_U7285
g5465 nand P3_ADD_467_U79 P3_U2601 ; P3_U7286
g5466 nand P3_U7910 P3_EBX_REG_22__SCAN_IN ; P3_U7287
g5467 nand P3_ADD_430_U79 P3_U2405 ; P3_U7288
g5468 nand P3_U2403 P3_ADD_318_U79 ; P3_U7289
g5469 nand P3_SUB_320_U12 P3_U4319 ; P3_U7290
g5470 nand P3_U2401 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_U7291
g5471 nand P3_U7094 P3_REIP_REG_22__SCAN_IN ; P3_U7292
g5472 nand P3_SUB_414_U68 P3_U2602 ; P3_U7293
g5473 nand P3_ADD_467_U78 P3_U2601 ; P3_U7294
g5474 nand P3_U7910 P3_EBX_REG_23__SCAN_IN ; P3_U7295
g5475 nand P3_ADD_430_U78 P3_U2405 ; P3_U7296
g5476 nand P3_U2403 P3_ADD_318_U78 ; P3_U7297
g5477 nand P3_SUB_320_U68 P3_U4319 ; P3_U7298
g5478 nand P3_U2401 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_U7299
g5479 nand P3_U7094 P3_REIP_REG_23__SCAN_IN ; P3_U7300
g5480 nand P3_SUB_414_U13 P3_U2602 ; P3_U7301
g5481 nand P3_ADD_467_U77 P3_U2601 ; P3_U7302
g5482 nand P3_U7910 P3_EBX_REG_24__SCAN_IN ; P3_U7303
g5483 nand P3_ADD_430_U77 P3_U2405 ; P3_U7304
g5484 nand P3_U2403 P3_ADD_318_U77 ; P3_U7305
g5485 nand P3_SUB_320_U13 P3_U4319 ; P3_U7306
g5486 nand P3_U2401 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_U7307
g5487 nand P3_U7094 P3_REIP_REG_24__SCAN_IN ; P3_U7308
g5488 nand P3_SUB_414_U66 P3_U2602 ; P3_U7309
g5489 nand P3_ADD_467_U76 P3_U2601 ; P3_U7310
g5490 nand P3_U7910 P3_EBX_REG_25__SCAN_IN ; P3_U7311
g5491 nand P3_ADD_430_U76 P3_U2405 ; P3_U7312
g5492 nand P3_U2403 P3_ADD_318_U76 ; P3_U7313
g5493 nand P3_SUB_320_U66 P3_U4319 ; P3_U7314
g5494 nand P3_U2401 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_U7315
g5495 nand P3_U7094 P3_REIP_REG_25__SCAN_IN ; P3_U7316
g5496 nand P3_SUB_414_U14 P3_U2602 ; P3_U7317
g5497 nand P3_ADD_467_U75 P3_U2601 ; P3_U7318
g5498 nand P3_U7910 P3_EBX_REG_26__SCAN_IN ; P3_U7319
g5499 nand P3_ADD_430_U75 P3_U2405 ; P3_U7320
g5500 nand P3_U2403 P3_ADD_318_U75 ; P3_U7321
g5501 nand P3_SUB_320_U14 P3_U4319 ; P3_U7322
g5502 nand P3_U2401 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_U7323
g5503 nand P3_U7094 P3_REIP_REG_26__SCAN_IN ; P3_U7324
g5504 nand P3_SUB_414_U64 P3_U2602 ; P3_U7325
g5505 nand P3_ADD_467_U74 P3_U2601 ; P3_U7326
g5506 nand P3_U7910 P3_EBX_REG_27__SCAN_IN ; P3_U7327
g5507 nand P3_ADD_430_U74 P3_U2405 ; P3_U7328
g5508 nand P3_U2403 P3_ADD_318_U74 ; P3_U7329
g5509 nand P3_SUB_320_U64 P3_U4319 ; P3_U7330
g5510 nand P3_U2401 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_U7331
g5511 nand P3_U7094 P3_REIP_REG_27__SCAN_IN ; P3_U7332
g5512 nand P3_SUB_414_U15 P3_U2602 ; P3_U7333
g5513 nand P3_ADD_467_U73 P3_U2601 ; P3_U7334
g5514 nand P3_U7910 P3_EBX_REG_28__SCAN_IN ; P3_U7335
g5515 nand P3_ADD_430_U73 P3_U2405 ; P3_U7336
g5516 nand P3_U2403 P3_ADD_318_U73 ; P3_U7337
g5517 nand P3_SUB_320_U15 P3_U4319 ; P3_U7338
g5518 nand P3_U2401 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_U7339
g5519 nand P3_U7094 P3_REIP_REG_28__SCAN_IN ; P3_U7340
g5520 nand P3_SUB_414_U16 P3_U2602 ; P3_U7341
g5521 nand P3_ADD_467_U72 P3_U2601 ; P3_U7342
g5522 nand P3_U7910 P3_EBX_REG_29__SCAN_IN ; P3_U7343
g5523 nand P3_ADD_430_U72 P3_U2405 ; P3_U7344
g5524 nand P3_U2403 P3_ADD_318_U72 ; P3_U7345
g5525 nand P3_SUB_320_U16 P3_U4319 ; P3_U7346
g5526 nand P3_U2401 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_U7347
g5527 nand P3_U7094 P3_REIP_REG_29__SCAN_IN ; P3_U7348
g5528 nand P3_SUB_414_U62 P3_U2602 ; P3_U7349
g5529 nand P3_ADD_467_U70 P3_U2601 ; P3_U7350
g5530 nand P3_U7910 P3_EBX_REG_30__SCAN_IN ; P3_U7351
g5531 nand P3_ADD_430_U70 P3_U2405 ; P3_U7352
g5532 nand P3_U2403 P3_ADD_318_U70 ; P3_U7353
g5533 nand P3_SUB_320_U62 P3_U4319 ; P3_U7354
g5534 nand P3_U2401 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_U7355
g5535 nand P3_U7094 P3_REIP_REG_30__SCAN_IN ; P3_U7356
g5536 nand P3_U4135 P3_U2603 ; P3_U7357
g5537 nand P3_SUB_414_U51 P3_U2602 ; P3_U7358
g5538 nand P3_ADD_467_U69 P3_U2601 ; P3_U7359
g5539 nand P3_U7910 P3_EBX_REG_31__SCAN_IN ; P3_U7360
g5540 nand P3_ADD_430_U69 P3_U2405 ; P3_U7361
g5541 nand P3_U2403 P3_ADD_318_U69 ; P3_U7362
g5542 not P3_U7362 ; P3_U7363
g5543 nand P3_U2401 P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_U7364
g5544 nand P3_U7094 P3_REIP_REG_31__SCAN_IN ; P3_U7365
g5545 nand P3_DATAWIDTH_REG_0__SCAN_IN P3_DATAWIDTH_REG_1__SCAN_IN ; P3_U7366
g5546 or P3_REIP_REG_0__SCAN_IN P3_REIP_REG_1__SCAN_IN ; P3_U7367
g5547 not P3_U4285 ; P3_U7368
g5548 nand P3_U4285 P3_FLUSH_REG_SCAN_IN ; P3_U7369
g5549 nand P3_U4623 P3_U2390 ; P3_U7370
g5550 nand P3_U2453 P3_U2630 ; P3_U7371
g5551 nand P3_U3123 P3_U7371 ; P3_U7372
g5552 nand P3_U7372 P3_U3121 ; P3_U7373
g5553 not P3_U4287 ; P3_U7374
g5554 nand P3_U4296 P3_U2631 ; P3_U7375
g5555 nand P3_U3112 P3_U3118 ; P3_U7376
g5556 nand P3_U7919 P3_U4150 P3_STATE2_REG_2__SCAN_IN ; P3_U7377
g5557 nand P3_U7377 P3_STATE2_REG_0__SCAN_IN ; P3_U7378
g5558 nand P3_U3125 P3_U7378 ; P3_U7379
g5559 nand P3_U2390 P3_U2604 ; P3_U7380
g5560 nand P3_U7380 P3_CODEFETCH_REG_SCAN_IN ; P3_U7381
g5561 nand P3_U4347 P3_STATE2_REG_0__SCAN_IN ; P3_U7382
g5562 nand P3_STATE_REG_0__SCAN_IN P3_ADS_N_REG_SCAN_IN ; P3_U7383
g5563 not P3_U4288 ; P3_U7384
g5564 nand P3_U3111 P3_U3114 P3_STATE2_REG_2__SCAN_IN ; P3_U7385
g5565 nand P3_U4488 P3_STATE2_REG_2__SCAN_IN ; P3_U7386
g5566 nand P3_U2542 P3_INSTQUEUE_REG_15__7__SCAN_IN ; P3_U7387
g5567 nand P3_U2541 P3_INSTQUEUE_REG_14__7__SCAN_IN ; P3_U7388
g5568 nand P3_U2540 P3_INSTQUEUE_REG_13__7__SCAN_IN ; P3_U7389
g5569 nand P3_U2539 P3_INSTQUEUE_REG_12__7__SCAN_IN ; P3_U7390
g5570 nand P3_U2537 P3_INSTQUEUE_REG_11__7__SCAN_IN ; P3_U7391
g5571 nand P3_U2536 P3_INSTQUEUE_REG_10__7__SCAN_IN ; P3_U7392
g5572 nand P3_U2535 P3_INSTQUEUE_REG_9__7__SCAN_IN ; P3_U7393
g5573 nand P3_U2534 P3_INSTQUEUE_REG_8__7__SCAN_IN ; P3_U7394
g5574 nand P3_U2532 P3_INSTQUEUE_REG_7__7__SCAN_IN ; P3_U7395
g5575 nand P3_U2531 P3_INSTQUEUE_REG_6__7__SCAN_IN ; P3_U7396
g5576 nand P3_U2530 P3_INSTQUEUE_REG_5__7__SCAN_IN ; P3_U7397
g5577 nand P3_U2529 P3_INSTQUEUE_REG_4__7__SCAN_IN ; P3_U7398
g5578 nand P3_U2527 P3_INSTQUEUE_REG_3__7__SCAN_IN ; P3_U7399
g5579 nand P3_U2525 P3_INSTQUEUE_REG_2__7__SCAN_IN ; P3_U7400
g5580 nand P3_U2523 P3_INSTQUEUE_REG_1__7__SCAN_IN ; P3_U7401
g5581 nand P3_U2521 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U7402
g5582 nand P3_U2542 P3_INSTQUEUE_REG_15__6__SCAN_IN ; P3_U7403
g5583 nand P3_U2541 P3_INSTQUEUE_REG_14__6__SCAN_IN ; P3_U7404
g5584 nand P3_U2540 P3_INSTQUEUE_REG_13__6__SCAN_IN ; P3_U7405
g5585 nand P3_U2539 P3_INSTQUEUE_REG_12__6__SCAN_IN ; P3_U7406
g5586 nand P3_U2537 P3_INSTQUEUE_REG_11__6__SCAN_IN ; P3_U7407
g5587 nand P3_U2536 P3_INSTQUEUE_REG_10__6__SCAN_IN ; P3_U7408
g5588 nand P3_U2535 P3_INSTQUEUE_REG_9__6__SCAN_IN ; P3_U7409
g5589 nand P3_U2534 P3_INSTQUEUE_REG_8__6__SCAN_IN ; P3_U7410
g5590 nand P3_U2532 P3_INSTQUEUE_REG_7__6__SCAN_IN ; P3_U7411
g5591 nand P3_U2531 P3_INSTQUEUE_REG_6__6__SCAN_IN ; P3_U7412
g5592 nand P3_U2530 P3_INSTQUEUE_REG_5__6__SCAN_IN ; P3_U7413
g5593 nand P3_U2529 P3_INSTQUEUE_REG_4__6__SCAN_IN ; P3_U7414
g5594 nand P3_U2527 P3_INSTQUEUE_REG_3__6__SCAN_IN ; P3_U7415
g5595 nand P3_U2525 P3_INSTQUEUE_REG_2__6__SCAN_IN ; P3_U7416
g5596 nand P3_U2523 P3_INSTQUEUE_REG_1__6__SCAN_IN ; P3_U7417
g5597 nand P3_U2521 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U7418
g5598 nand P3_U2542 P3_INSTQUEUE_REG_15__5__SCAN_IN ; P3_U7419
g5599 nand P3_U2541 P3_INSTQUEUE_REG_14__5__SCAN_IN ; P3_U7420
g5600 nand P3_U2540 P3_INSTQUEUE_REG_13__5__SCAN_IN ; P3_U7421
g5601 nand P3_U2539 P3_INSTQUEUE_REG_12__5__SCAN_IN ; P3_U7422
g5602 nand P3_U2537 P3_INSTQUEUE_REG_11__5__SCAN_IN ; P3_U7423
g5603 nand P3_U2536 P3_INSTQUEUE_REG_10__5__SCAN_IN ; P3_U7424
g5604 nand P3_U2535 P3_INSTQUEUE_REG_9__5__SCAN_IN ; P3_U7425
g5605 nand P3_U2534 P3_INSTQUEUE_REG_8__5__SCAN_IN ; P3_U7426
g5606 nand P3_U2532 P3_INSTQUEUE_REG_7__5__SCAN_IN ; P3_U7427
g5607 nand P3_U2531 P3_INSTQUEUE_REG_6__5__SCAN_IN ; P3_U7428
g5608 nand P3_U2530 P3_INSTQUEUE_REG_5__5__SCAN_IN ; P3_U7429
g5609 nand P3_U2529 P3_INSTQUEUE_REG_4__5__SCAN_IN ; P3_U7430
g5610 nand P3_U2527 P3_INSTQUEUE_REG_3__5__SCAN_IN ; P3_U7431
g5611 nand P3_U2525 P3_INSTQUEUE_REG_2__5__SCAN_IN ; P3_U7432
g5612 nand P3_U2523 P3_INSTQUEUE_REG_1__5__SCAN_IN ; P3_U7433
g5613 nand P3_U2521 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U7434
g5614 nand P3_U2542 P3_INSTQUEUE_REG_15__4__SCAN_IN ; P3_U7435
g5615 nand P3_U2541 P3_INSTQUEUE_REG_14__4__SCAN_IN ; P3_U7436
g5616 nand P3_U2540 P3_INSTQUEUE_REG_13__4__SCAN_IN ; P3_U7437
g5617 nand P3_U2539 P3_INSTQUEUE_REG_12__4__SCAN_IN ; P3_U7438
g5618 nand P3_U2537 P3_INSTQUEUE_REG_11__4__SCAN_IN ; P3_U7439
g5619 nand P3_U2536 P3_INSTQUEUE_REG_10__4__SCAN_IN ; P3_U7440
g5620 nand P3_U2535 P3_INSTQUEUE_REG_9__4__SCAN_IN ; P3_U7441
g5621 nand P3_U2534 P3_INSTQUEUE_REG_8__4__SCAN_IN ; P3_U7442
g5622 nand P3_U2532 P3_INSTQUEUE_REG_7__4__SCAN_IN ; P3_U7443
g5623 nand P3_U2531 P3_INSTQUEUE_REG_6__4__SCAN_IN ; P3_U7444
g5624 nand P3_U2530 P3_INSTQUEUE_REG_5__4__SCAN_IN ; P3_U7445
g5625 nand P3_U2529 P3_INSTQUEUE_REG_4__4__SCAN_IN ; P3_U7446
g5626 nand P3_U2527 P3_INSTQUEUE_REG_3__4__SCAN_IN ; P3_U7447
g5627 nand P3_U2525 P3_INSTQUEUE_REG_2__4__SCAN_IN ; P3_U7448
g5628 nand P3_U2523 P3_INSTQUEUE_REG_1__4__SCAN_IN ; P3_U7449
g5629 nand P3_U2521 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U7450
g5630 nand P3_U2542 P3_INSTQUEUE_REG_15__3__SCAN_IN ; P3_U7451
g5631 nand P3_U2541 P3_INSTQUEUE_REG_14__3__SCAN_IN ; P3_U7452
g5632 nand P3_U2540 P3_INSTQUEUE_REG_13__3__SCAN_IN ; P3_U7453
g5633 nand P3_U2539 P3_INSTQUEUE_REG_12__3__SCAN_IN ; P3_U7454
g5634 nand P3_U2537 P3_INSTQUEUE_REG_11__3__SCAN_IN ; P3_U7455
g5635 nand P3_U2536 P3_INSTQUEUE_REG_10__3__SCAN_IN ; P3_U7456
g5636 nand P3_U2535 P3_INSTQUEUE_REG_9__3__SCAN_IN ; P3_U7457
g5637 nand P3_U2534 P3_INSTQUEUE_REG_8__3__SCAN_IN ; P3_U7458
g5638 nand P3_U2532 P3_INSTQUEUE_REG_7__3__SCAN_IN ; P3_U7459
g5639 nand P3_U2531 P3_INSTQUEUE_REG_6__3__SCAN_IN ; P3_U7460
g5640 nand P3_U2530 P3_INSTQUEUE_REG_5__3__SCAN_IN ; P3_U7461
g5641 nand P3_U2529 P3_INSTQUEUE_REG_4__3__SCAN_IN ; P3_U7462
g5642 nand P3_U2527 P3_INSTQUEUE_REG_3__3__SCAN_IN ; P3_U7463
g5643 nand P3_U2525 P3_INSTQUEUE_REG_2__3__SCAN_IN ; P3_U7464
g5644 nand P3_U2523 P3_INSTQUEUE_REG_1__3__SCAN_IN ; P3_U7465
g5645 nand P3_U2521 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U7466
g5646 nand P3_U2542 P3_INSTQUEUE_REG_15__2__SCAN_IN ; P3_U7467
g5647 nand P3_U2541 P3_INSTQUEUE_REG_14__2__SCAN_IN ; P3_U7468
g5648 nand P3_U2540 P3_INSTQUEUE_REG_13__2__SCAN_IN ; P3_U7469
g5649 nand P3_U2539 P3_INSTQUEUE_REG_12__2__SCAN_IN ; P3_U7470
g5650 nand P3_U2537 P3_INSTQUEUE_REG_11__2__SCAN_IN ; P3_U7471
g5651 nand P3_U2536 P3_INSTQUEUE_REG_10__2__SCAN_IN ; P3_U7472
g5652 nand P3_U2535 P3_INSTQUEUE_REG_9__2__SCAN_IN ; P3_U7473
g5653 nand P3_U2534 P3_INSTQUEUE_REG_8__2__SCAN_IN ; P3_U7474
g5654 nand P3_U2532 P3_INSTQUEUE_REG_7__2__SCAN_IN ; P3_U7475
g5655 nand P3_U2531 P3_INSTQUEUE_REG_6__2__SCAN_IN ; P3_U7476
g5656 nand P3_U2530 P3_INSTQUEUE_REG_5__2__SCAN_IN ; P3_U7477
g5657 nand P3_U2529 P3_INSTQUEUE_REG_4__2__SCAN_IN ; P3_U7478
g5658 nand P3_U2527 P3_INSTQUEUE_REG_3__2__SCAN_IN ; P3_U7479
g5659 nand P3_U2525 P3_INSTQUEUE_REG_2__2__SCAN_IN ; P3_U7480
g5660 nand P3_U2523 P3_INSTQUEUE_REG_1__2__SCAN_IN ; P3_U7481
g5661 nand P3_U2521 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U7482
g5662 nand P3_U2542 P3_INSTQUEUE_REG_15__1__SCAN_IN ; P3_U7483
g5663 nand P3_U2541 P3_INSTQUEUE_REG_14__1__SCAN_IN ; P3_U7484
g5664 nand P3_U2540 P3_INSTQUEUE_REG_13__1__SCAN_IN ; P3_U7485
g5665 nand P3_U2539 P3_INSTQUEUE_REG_12__1__SCAN_IN ; P3_U7486
g5666 nand P3_U2537 P3_INSTQUEUE_REG_11__1__SCAN_IN ; P3_U7487
g5667 nand P3_U2536 P3_INSTQUEUE_REG_10__1__SCAN_IN ; P3_U7488
g5668 nand P3_U2535 P3_INSTQUEUE_REG_9__1__SCAN_IN ; P3_U7489
g5669 nand P3_U2534 P3_INSTQUEUE_REG_8__1__SCAN_IN ; P3_U7490
g5670 nand P3_U2532 P3_INSTQUEUE_REG_7__1__SCAN_IN ; P3_U7491
g5671 nand P3_U2531 P3_INSTQUEUE_REG_6__1__SCAN_IN ; P3_U7492
g5672 nand P3_U2530 P3_INSTQUEUE_REG_5__1__SCAN_IN ; P3_U7493
g5673 nand P3_U2529 P3_INSTQUEUE_REG_4__1__SCAN_IN ; P3_U7494
g5674 nand P3_U2527 P3_INSTQUEUE_REG_3__1__SCAN_IN ; P3_U7495
g5675 nand P3_U2525 P3_INSTQUEUE_REG_2__1__SCAN_IN ; P3_U7496
g5676 nand P3_U2523 P3_INSTQUEUE_REG_1__1__SCAN_IN ; P3_U7497
g5677 nand P3_U2521 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U7498
g5678 nand P3_U2542 P3_INSTQUEUE_REG_15__0__SCAN_IN ; P3_U7499
g5679 nand P3_U2541 P3_INSTQUEUE_REG_14__0__SCAN_IN ; P3_U7500
g5680 nand P3_U2540 P3_INSTQUEUE_REG_13__0__SCAN_IN ; P3_U7501
g5681 nand P3_U2539 P3_INSTQUEUE_REG_12__0__SCAN_IN ; P3_U7502
g5682 nand P3_U2537 P3_INSTQUEUE_REG_11__0__SCAN_IN ; P3_U7503
g5683 nand P3_U2536 P3_INSTQUEUE_REG_10__0__SCAN_IN ; P3_U7504
g5684 nand P3_U2535 P3_INSTQUEUE_REG_9__0__SCAN_IN ; P3_U7505
g5685 nand P3_U2534 P3_INSTQUEUE_REG_8__0__SCAN_IN ; P3_U7506
g5686 nand P3_U2532 P3_INSTQUEUE_REG_7__0__SCAN_IN ; P3_U7507
g5687 nand P3_U2531 P3_INSTQUEUE_REG_6__0__SCAN_IN ; P3_U7508
g5688 nand P3_U2530 P3_INSTQUEUE_REG_5__0__SCAN_IN ; P3_U7509
g5689 nand P3_U2529 P3_INSTQUEUE_REG_4__0__SCAN_IN ; P3_U7510
g5690 nand P3_U2527 P3_INSTQUEUE_REG_3__0__SCAN_IN ; P3_U7511
g5691 nand P3_U2525 P3_INSTQUEUE_REG_2__0__SCAN_IN ; P3_U7512
g5692 nand P3_U2523 P3_INSTQUEUE_REG_1__0__SCAN_IN ; P3_U7513
g5693 nand P3_U2521 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U7514
g5694 nand P3_U4470 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U7515
g5695 not P3_U3266 ; P3_U7516
g5696 nand P3_U2562 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U7517
g5697 nand P3_U2561 P3_INSTQUEUE_REG_1__7__SCAN_IN ; P3_U7518
g5698 nand P3_U2560 P3_INSTQUEUE_REG_2__7__SCAN_IN ; P3_U7519
g5699 nand P3_U2559 P3_INSTQUEUE_REG_3__7__SCAN_IN ; P3_U7520
g5700 nand P3_U2557 P3_INSTQUEUE_REG_4__7__SCAN_IN ; P3_U7521
g5701 nand P3_U2556 P3_INSTQUEUE_REG_5__7__SCAN_IN ; P3_U7522
g5702 nand P3_U2555 P3_INSTQUEUE_REG_6__7__SCAN_IN ; P3_U7523
g5703 nand P3_U2554 P3_INSTQUEUE_REG_7__7__SCAN_IN ; P3_U7524
g5704 nand P3_U2552 P3_INSTQUEUE_REG_8__7__SCAN_IN ; P3_U7525
g5705 nand P3_U2551 P3_INSTQUEUE_REG_9__7__SCAN_IN ; P3_U7526
g5706 nand P3_U2550 P3_INSTQUEUE_REG_10__7__SCAN_IN ; P3_U7527
g5707 nand P3_U2549 P3_INSTQUEUE_REG_11__7__SCAN_IN ; P3_U7528
g5708 nand P3_U2547 P3_INSTQUEUE_REG_12__7__SCAN_IN ; P3_U7529
g5709 nand P3_U2546 P3_INSTQUEUE_REG_13__7__SCAN_IN ; P3_U7530
g5710 nand P3_U2545 P3_INSTQUEUE_REG_14__7__SCAN_IN ; P3_U7531
g5711 nand P3_U2544 P3_INSTQUEUE_REG_15__7__SCAN_IN ; P3_U7532
g5712 nand P3_U2562 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U7533
g5713 nand P3_U2561 P3_INSTQUEUE_REG_1__6__SCAN_IN ; P3_U7534
g5714 nand P3_U2560 P3_INSTQUEUE_REG_2__6__SCAN_IN ; P3_U7535
g5715 nand P3_U2559 P3_INSTQUEUE_REG_3__6__SCAN_IN ; P3_U7536
g5716 nand P3_U2557 P3_INSTQUEUE_REG_4__6__SCAN_IN ; P3_U7537
g5717 nand P3_U2556 P3_INSTQUEUE_REG_5__6__SCAN_IN ; P3_U7538
g5718 nand P3_U2555 P3_INSTQUEUE_REG_6__6__SCAN_IN ; P3_U7539
g5719 nand P3_U2554 P3_INSTQUEUE_REG_7__6__SCAN_IN ; P3_U7540
g5720 nand P3_U2552 P3_INSTQUEUE_REG_8__6__SCAN_IN ; P3_U7541
g5721 nand P3_U2551 P3_INSTQUEUE_REG_9__6__SCAN_IN ; P3_U7542
g5722 nand P3_U2550 P3_INSTQUEUE_REG_10__6__SCAN_IN ; P3_U7543
g5723 nand P3_U2549 P3_INSTQUEUE_REG_11__6__SCAN_IN ; P3_U7544
g5724 nand P3_U2547 P3_INSTQUEUE_REG_12__6__SCAN_IN ; P3_U7545
g5725 nand P3_U2546 P3_INSTQUEUE_REG_13__6__SCAN_IN ; P3_U7546
g5726 nand P3_U2545 P3_INSTQUEUE_REG_14__6__SCAN_IN ; P3_U7547
g5727 nand P3_U2544 P3_INSTQUEUE_REG_15__6__SCAN_IN ; P3_U7548
g5728 nand P3_U2562 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U7549
g5729 nand P3_U2561 P3_INSTQUEUE_REG_1__5__SCAN_IN ; P3_U7550
g5730 nand P3_U2560 P3_INSTQUEUE_REG_2__5__SCAN_IN ; P3_U7551
g5731 nand P3_U2559 P3_INSTQUEUE_REG_3__5__SCAN_IN ; P3_U7552
g5732 nand P3_U2557 P3_INSTQUEUE_REG_4__5__SCAN_IN ; P3_U7553
g5733 nand P3_U2556 P3_INSTQUEUE_REG_5__5__SCAN_IN ; P3_U7554
g5734 nand P3_U2555 P3_INSTQUEUE_REG_6__5__SCAN_IN ; P3_U7555
g5735 nand P3_U2554 P3_INSTQUEUE_REG_7__5__SCAN_IN ; P3_U7556
g5736 nand P3_U2552 P3_INSTQUEUE_REG_8__5__SCAN_IN ; P3_U7557
g5737 nand P3_U2551 P3_INSTQUEUE_REG_9__5__SCAN_IN ; P3_U7558
g5738 nand P3_U2550 P3_INSTQUEUE_REG_10__5__SCAN_IN ; P3_U7559
g5739 nand P3_U2549 P3_INSTQUEUE_REG_11__5__SCAN_IN ; P3_U7560
g5740 nand P3_U2547 P3_INSTQUEUE_REG_12__5__SCAN_IN ; P3_U7561
g5741 nand P3_U2546 P3_INSTQUEUE_REG_13__5__SCAN_IN ; P3_U7562
g5742 nand P3_U2545 P3_INSTQUEUE_REG_14__5__SCAN_IN ; P3_U7563
g5743 nand P3_U2544 P3_INSTQUEUE_REG_15__5__SCAN_IN ; P3_U7564
g5744 nand P3_U2562 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U7565
g5745 nand P3_U2561 P3_INSTQUEUE_REG_1__4__SCAN_IN ; P3_U7566
g5746 nand P3_U2560 P3_INSTQUEUE_REG_2__4__SCAN_IN ; P3_U7567
g5747 nand P3_U2559 P3_INSTQUEUE_REG_3__4__SCAN_IN ; P3_U7568
g5748 nand P3_U2557 P3_INSTQUEUE_REG_4__4__SCAN_IN ; P3_U7569
g5749 nand P3_U2556 P3_INSTQUEUE_REG_5__4__SCAN_IN ; P3_U7570
g5750 nand P3_U2555 P3_INSTQUEUE_REG_6__4__SCAN_IN ; P3_U7571
g5751 nand P3_U2554 P3_INSTQUEUE_REG_7__4__SCAN_IN ; P3_U7572
g5752 nand P3_U2552 P3_INSTQUEUE_REG_8__4__SCAN_IN ; P3_U7573
g5753 nand P3_U2551 P3_INSTQUEUE_REG_9__4__SCAN_IN ; P3_U7574
g5754 nand P3_U2550 P3_INSTQUEUE_REG_10__4__SCAN_IN ; P3_U7575
g5755 nand P3_U2549 P3_INSTQUEUE_REG_11__4__SCAN_IN ; P3_U7576
g5756 nand P3_U2547 P3_INSTQUEUE_REG_12__4__SCAN_IN ; P3_U7577
g5757 nand P3_U2546 P3_INSTQUEUE_REG_13__4__SCAN_IN ; P3_U7578
g5758 nand P3_U2545 P3_INSTQUEUE_REG_14__4__SCAN_IN ; P3_U7579
g5759 nand P3_U2544 P3_INSTQUEUE_REG_15__4__SCAN_IN ; P3_U7580
g5760 nand P3_U2562 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U7581
g5761 nand P3_U2561 P3_INSTQUEUE_REG_1__3__SCAN_IN ; P3_U7582
g5762 nand P3_U2560 P3_INSTQUEUE_REG_2__3__SCAN_IN ; P3_U7583
g5763 nand P3_U2559 P3_INSTQUEUE_REG_3__3__SCAN_IN ; P3_U7584
g5764 nand P3_U2557 P3_INSTQUEUE_REG_4__3__SCAN_IN ; P3_U7585
g5765 nand P3_U2556 P3_INSTQUEUE_REG_5__3__SCAN_IN ; P3_U7586
g5766 nand P3_U2555 P3_INSTQUEUE_REG_6__3__SCAN_IN ; P3_U7587
g5767 nand P3_U2554 P3_INSTQUEUE_REG_7__3__SCAN_IN ; P3_U7588
g5768 nand P3_U2552 P3_INSTQUEUE_REG_8__3__SCAN_IN ; P3_U7589
g5769 nand P3_U2551 P3_INSTQUEUE_REG_9__3__SCAN_IN ; P3_U7590
g5770 nand P3_U2550 P3_INSTQUEUE_REG_10__3__SCAN_IN ; P3_U7591
g5771 nand P3_U2549 P3_INSTQUEUE_REG_11__3__SCAN_IN ; P3_U7592
g5772 nand P3_U2547 P3_INSTQUEUE_REG_12__3__SCAN_IN ; P3_U7593
g5773 nand P3_U2546 P3_INSTQUEUE_REG_13__3__SCAN_IN ; P3_U7594
g5774 nand P3_U2545 P3_INSTQUEUE_REG_14__3__SCAN_IN ; P3_U7595
g5775 nand P3_U2544 P3_INSTQUEUE_REG_15__3__SCAN_IN ; P3_U7596
g5776 nand P3_U2562 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U7597
g5777 nand P3_U2561 P3_INSTQUEUE_REG_1__2__SCAN_IN ; P3_U7598
g5778 nand P3_U2560 P3_INSTQUEUE_REG_2__2__SCAN_IN ; P3_U7599
g5779 nand P3_U2559 P3_INSTQUEUE_REG_3__2__SCAN_IN ; P3_U7600
g5780 nand P3_U2557 P3_INSTQUEUE_REG_4__2__SCAN_IN ; P3_U7601
g5781 nand P3_U2556 P3_INSTQUEUE_REG_5__2__SCAN_IN ; P3_U7602
g5782 nand P3_U2555 P3_INSTQUEUE_REG_6__2__SCAN_IN ; P3_U7603
g5783 nand P3_U2554 P3_INSTQUEUE_REG_7__2__SCAN_IN ; P3_U7604
g5784 nand P3_U2552 P3_INSTQUEUE_REG_8__2__SCAN_IN ; P3_U7605
g5785 nand P3_U2551 P3_INSTQUEUE_REG_9__2__SCAN_IN ; P3_U7606
g5786 nand P3_U2550 P3_INSTQUEUE_REG_10__2__SCAN_IN ; P3_U7607
g5787 nand P3_U2549 P3_INSTQUEUE_REG_11__2__SCAN_IN ; P3_U7608
g5788 nand P3_U2547 P3_INSTQUEUE_REG_12__2__SCAN_IN ; P3_U7609
g5789 nand P3_U2546 P3_INSTQUEUE_REG_13__2__SCAN_IN ; P3_U7610
g5790 nand P3_U2545 P3_INSTQUEUE_REG_14__2__SCAN_IN ; P3_U7611
g5791 nand P3_U2544 P3_INSTQUEUE_REG_15__2__SCAN_IN ; P3_U7612
g5792 nand P3_U2562 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U7613
g5793 nand P3_U2561 P3_INSTQUEUE_REG_1__1__SCAN_IN ; P3_U7614
g5794 nand P3_U2560 P3_INSTQUEUE_REG_2__1__SCAN_IN ; P3_U7615
g5795 nand P3_U2559 P3_INSTQUEUE_REG_3__1__SCAN_IN ; P3_U7616
g5796 nand P3_U2557 P3_INSTQUEUE_REG_4__1__SCAN_IN ; P3_U7617
g5797 nand P3_U2556 P3_INSTQUEUE_REG_5__1__SCAN_IN ; P3_U7618
g5798 nand P3_U2555 P3_INSTQUEUE_REG_6__1__SCAN_IN ; P3_U7619
g5799 nand P3_U2554 P3_INSTQUEUE_REG_7__1__SCAN_IN ; P3_U7620
g5800 nand P3_U2552 P3_INSTQUEUE_REG_8__1__SCAN_IN ; P3_U7621
g5801 nand P3_U2551 P3_INSTQUEUE_REG_9__1__SCAN_IN ; P3_U7622
g5802 nand P3_U2550 P3_INSTQUEUE_REG_10__1__SCAN_IN ; P3_U7623
g5803 nand P3_U2549 P3_INSTQUEUE_REG_11__1__SCAN_IN ; P3_U7624
g5804 nand P3_U2547 P3_INSTQUEUE_REG_12__1__SCAN_IN ; P3_U7625
g5805 nand P3_U2546 P3_INSTQUEUE_REG_13__1__SCAN_IN ; P3_U7626
g5806 nand P3_U2545 P3_INSTQUEUE_REG_14__1__SCAN_IN ; P3_U7627
g5807 nand P3_U2544 P3_INSTQUEUE_REG_15__1__SCAN_IN ; P3_U7628
g5808 nand P3_U2562 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U7629
g5809 nand P3_U2561 P3_INSTQUEUE_REG_1__0__SCAN_IN ; P3_U7630
g5810 nand P3_U2560 P3_INSTQUEUE_REG_2__0__SCAN_IN ; P3_U7631
g5811 nand P3_U2559 P3_INSTQUEUE_REG_3__0__SCAN_IN ; P3_U7632
g5812 nand P3_U2557 P3_INSTQUEUE_REG_4__0__SCAN_IN ; P3_U7633
g5813 nand P3_U2556 P3_INSTQUEUE_REG_5__0__SCAN_IN ; P3_U7634
g5814 nand P3_U2555 P3_INSTQUEUE_REG_6__0__SCAN_IN ; P3_U7635
g5815 nand P3_U2554 P3_INSTQUEUE_REG_7__0__SCAN_IN ; P3_U7636
g5816 nand P3_U2552 P3_INSTQUEUE_REG_8__0__SCAN_IN ; P3_U7637
g5817 nand P3_U2551 P3_INSTQUEUE_REG_9__0__SCAN_IN ; P3_U7638
g5818 nand P3_U2550 P3_INSTQUEUE_REG_10__0__SCAN_IN ; P3_U7639
g5819 nand P3_U2549 P3_INSTQUEUE_REG_11__0__SCAN_IN ; P3_U7640
g5820 nand P3_U2547 P3_INSTQUEUE_REG_12__0__SCAN_IN ; P3_U7641
g5821 nand P3_U2546 P3_INSTQUEUE_REG_13__0__SCAN_IN ; P3_U7642
g5822 nand P3_U2545 P3_INSTQUEUE_REG_14__0__SCAN_IN ; P3_U7643
g5823 nand P3_U2544 P3_INSTQUEUE_REG_15__0__SCAN_IN ; P3_U7644
g5824 not P3_U4289 ; P3_U7645
g5825 nand P3_U2582 P3_INSTQUEUE_REG_8__7__SCAN_IN ; P3_U7646
g5826 nand P3_U2581 P3_INSTQUEUE_REG_9__7__SCAN_IN ; P3_U7647
g5827 nand P3_U2580 P3_INSTQUEUE_REG_10__7__SCAN_IN ; P3_U7648
g5828 nand P3_U2579 P3_INSTQUEUE_REG_11__7__SCAN_IN ; P3_U7649
g5829 nand P3_U2577 P3_INSTQUEUE_REG_12__7__SCAN_IN ; P3_U7650
g5830 nand P3_U2576 P3_INSTQUEUE_REG_13__7__SCAN_IN ; P3_U7651
g5831 nand P3_U2575 P3_INSTQUEUE_REG_14__7__SCAN_IN ; P3_U7652
g5832 nand P3_U2574 P3_INSTQUEUE_REG_15__7__SCAN_IN ; P3_U7653
g5833 nand P3_U2572 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U7654
g5834 nand P3_U2571 P3_INSTQUEUE_REG_1__7__SCAN_IN ; P3_U7655
g5835 nand P3_U2570 P3_INSTQUEUE_REG_2__7__SCAN_IN ; P3_U7656
g5836 nand P3_U2569 P3_INSTQUEUE_REG_3__7__SCAN_IN ; P3_U7657
g5837 nand P3_U2567 P3_INSTQUEUE_REG_4__7__SCAN_IN ; P3_U7658
g5838 nand P3_U2566 P3_INSTQUEUE_REG_5__7__SCAN_IN ; P3_U7659
g5839 nand P3_U2565 P3_INSTQUEUE_REG_6__7__SCAN_IN ; P3_U7660
g5840 nand P3_U2564 P3_INSTQUEUE_REG_7__7__SCAN_IN ; P3_U7661
g5841 nand P3_U2582 P3_INSTQUEUE_REG_8__6__SCAN_IN ; P3_U7662
g5842 nand P3_U2581 P3_INSTQUEUE_REG_9__6__SCAN_IN ; P3_U7663
g5843 nand P3_U2580 P3_INSTQUEUE_REG_10__6__SCAN_IN ; P3_U7664
g5844 nand P3_U2579 P3_INSTQUEUE_REG_11__6__SCAN_IN ; P3_U7665
g5845 nand P3_U2577 P3_INSTQUEUE_REG_12__6__SCAN_IN ; P3_U7666
g5846 nand P3_U2576 P3_INSTQUEUE_REG_13__6__SCAN_IN ; P3_U7667
g5847 nand P3_U2575 P3_INSTQUEUE_REG_14__6__SCAN_IN ; P3_U7668
g5848 nand P3_U2574 P3_INSTQUEUE_REG_15__6__SCAN_IN ; P3_U7669
g5849 nand P3_U2572 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U7670
g5850 nand P3_U2571 P3_INSTQUEUE_REG_1__6__SCAN_IN ; P3_U7671
g5851 nand P3_U2570 P3_INSTQUEUE_REG_2__6__SCAN_IN ; P3_U7672
g5852 nand P3_U2569 P3_INSTQUEUE_REG_3__6__SCAN_IN ; P3_U7673
g5853 nand P3_U2567 P3_INSTQUEUE_REG_4__6__SCAN_IN ; P3_U7674
g5854 nand P3_U2566 P3_INSTQUEUE_REG_5__6__SCAN_IN ; P3_U7675
g5855 nand P3_U2565 P3_INSTQUEUE_REG_6__6__SCAN_IN ; P3_U7676
g5856 nand P3_U2564 P3_INSTQUEUE_REG_7__6__SCAN_IN ; P3_U7677
g5857 nand P3_U2582 P3_INSTQUEUE_REG_8__5__SCAN_IN ; P3_U7678
g5858 nand P3_U2581 P3_INSTQUEUE_REG_9__5__SCAN_IN ; P3_U7679
g5859 nand P3_U2580 P3_INSTQUEUE_REG_10__5__SCAN_IN ; P3_U7680
g5860 nand P3_U2579 P3_INSTQUEUE_REG_11__5__SCAN_IN ; P3_U7681
g5861 nand P3_U2577 P3_INSTQUEUE_REG_12__5__SCAN_IN ; P3_U7682
g5862 nand P3_U2576 P3_INSTQUEUE_REG_13__5__SCAN_IN ; P3_U7683
g5863 nand P3_U2575 P3_INSTQUEUE_REG_14__5__SCAN_IN ; P3_U7684
g5864 nand P3_U2574 P3_INSTQUEUE_REG_15__5__SCAN_IN ; P3_U7685
g5865 nand P3_U2572 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U7686
g5866 nand P3_U2571 P3_INSTQUEUE_REG_1__5__SCAN_IN ; P3_U7687
g5867 nand P3_U2570 P3_INSTQUEUE_REG_2__5__SCAN_IN ; P3_U7688
g5868 nand P3_U2569 P3_INSTQUEUE_REG_3__5__SCAN_IN ; P3_U7689
g5869 nand P3_U2567 P3_INSTQUEUE_REG_4__5__SCAN_IN ; P3_U7690
g5870 nand P3_U2566 P3_INSTQUEUE_REG_5__5__SCAN_IN ; P3_U7691
g5871 nand P3_U2565 P3_INSTQUEUE_REG_6__5__SCAN_IN ; P3_U7692
g5872 nand P3_U2564 P3_INSTQUEUE_REG_7__5__SCAN_IN ; P3_U7693
g5873 nand P3_U2582 P3_INSTQUEUE_REG_8__4__SCAN_IN ; P3_U7694
g5874 nand P3_U2581 P3_INSTQUEUE_REG_9__4__SCAN_IN ; P3_U7695
g5875 nand P3_U2580 P3_INSTQUEUE_REG_10__4__SCAN_IN ; P3_U7696
g5876 nand P3_U2579 P3_INSTQUEUE_REG_11__4__SCAN_IN ; P3_U7697
g5877 nand P3_U2577 P3_INSTQUEUE_REG_12__4__SCAN_IN ; P3_U7698
g5878 nand P3_U2576 P3_INSTQUEUE_REG_13__4__SCAN_IN ; P3_U7699
g5879 nand P3_U2575 P3_INSTQUEUE_REG_14__4__SCAN_IN ; P3_U7700
g5880 nand P3_U2574 P3_INSTQUEUE_REG_15__4__SCAN_IN ; P3_U7701
g5881 nand P3_U2572 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U7702
g5882 nand P3_U2571 P3_INSTQUEUE_REG_1__4__SCAN_IN ; P3_U7703
g5883 nand P3_U2570 P3_INSTQUEUE_REG_2__4__SCAN_IN ; P3_U7704
g5884 nand P3_U2569 P3_INSTQUEUE_REG_3__4__SCAN_IN ; P3_U7705
g5885 nand P3_U2567 P3_INSTQUEUE_REG_4__4__SCAN_IN ; P3_U7706
g5886 nand P3_U2566 P3_INSTQUEUE_REG_5__4__SCAN_IN ; P3_U7707
g5887 nand P3_U2565 P3_INSTQUEUE_REG_6__4__SCAN_IN ; P3_U7708
g5888 nand P3_U2564 P3_INSTQUEUE_REG_7__4__SCAN_IN ; P3_U7709
g5889 nand P3_U2582 P3_INSTQUEUE_REG_8__3__SCAN_IN ; P3_U7710
g5890 nand P3_U2581 P3_INSTQUEUE_REG_9__3__SCAN_IN ; P3_U7711
g5891 nand P3_U2580 P3_INSTQUEUE_REG_10__3__SCAN_IN ; P3_U7712
g5892 nand P3_U2579 P3_INSTQUEUE_REG_11__3__SCAN_IN ; P3_U7713
g5893 nand P3_U2577 P3_INSTQUEUE_REG_12__3__SCAN_IN ; P3_U7714
g5894 nand P3_U2576 P3_INSTQUEUE_REG_13__3__SCAN_IN ; P3_U7715
g5895 nand P3_U2575 P3_INSTQUEUE_REG_14__3__SCAN_IN ; P3_U7716
g5896 nand P3_U2574 P3_INSTQUEUE_REG_15__3__SCAN_IN ; P3_U7717
g5897 nand P3_U2572 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U7718
g5898 nand P3_U2571 P3_INSTQUEUE_REG_1__3__SCAN_IN ; P3_U7719
g5899 nand P3_U2570 P3_INSTQUEUE_REG_2__3__SCAN_IN ; P3_U7720
g5900 nand P3_U2569 P3_INSTQUEUE_REG_3__3__SCAN_IN ; P3_U7721
g5901 nand P3_U2567 P3_INSTQUEUE_REG_4__3__SCAN_IN ; P3_U7722
g5902 nand P3_U2566 P3_INSTQUEUE_REG_5__3__SCAN_IN ; P3_U7723
g5903 nand P3_U2565 P3_INSTQUEUE_REG_6__3__SCAN_IN ; P3_U7724
g5904 nand P3_U2564 P3_INSTQUEUE_REG_7__3__SCAN_IN ; P3_U7725
g5905 nand P3_U2582 P3_INSTQUEUE_REG_8__2__SCAN_IN ; P3_U7726
g5906 nand P3_U2581 P3_INSTQUEUE_REG_9__2__SCAN_IN ; P3_U7727
g5907 nand P3_U2580 P3_INSTQUEUE_REG_10__2__SCAN_IN ; P3_U7728
g5908 nand P3_U2579 P3_INSTQUEUE_REG_11__2__SCAN_IN ; P3_U7729
g5909 nand P3_U2577 P3_INSTQUEUE_REG_12__2__SCAN_IN ; P3_U7730
g5910 nand P3_U2576 P3_INSTQUEUE_REG_13__2__SCAN_IN ; P3_U7731
g5911 nand P3_U2575 P3_INSTQUEUE_REG_14__2__SCAN_IN ; P3_U7732
g5912 nand P3_U2574 P3_INSTQUEUE_REG_15__2__SCAN_IN ; P3_U7733
g5913 nand P3_U2572 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U7734
g5914 nand P3_U2571 P3_INSTQUEUE_REG_1__2__SCAN_IN ; P3_U7735
g5915 nand P3_U2570 P3_INSTQUEUE_REG_2__2__SCAN_IN ; P3_U7736
g5916 nand P3_U2569 P3_INSTQUEUE_REG_3__2__SCAN_IN ; P3_U7737
g5917 nand P3_U2567 P3_INSTQUEUE_REG_4__2__SCAN_IN ; P3_U7738
g5918 nand P3_U2566 P3_INSTQUEUE_REG_5__2__SCAN_IN ; P3_U7739
g5919 nand P3_U2565 P3_INSTQUEUE_REG_6__2__SCAN_IN ; P3_U7740
g5920 nand P3_U2564 P3_INSTQUEUE_REG_7__2__SCAN_IN ; P3_U7741
g5921 nand P3_U2582 P3_INSTQUEUE_REG_8__1__SCAN_IN ; P3_U7742
g5922 nand P3_U2581 P3_INSTQUEUE_REG_9__1__SCAN_IN ; P3_U7743
g5923 nand P3_U2580 P3_INSTQUEUE_REG_10__1__SCAN_IN ; P3_U7744
g5924 nand P3_U2579 P3_INSTQUEUE_REG_11__1__SCAN_IN ; P3_U7745
g5925 nand P3_U2577 P3_INSTQUEUE_REG_12__1__SCAN_IN ; P3_U7746
g5926 nand P3_U2576 P3_INSTQUEUE_REG_13__1__SCAN_IN ; P3_U7747
g5927 nand P3_U2575 P3_INSTQUEUE_REG_14__1__SCAN_IN ; P3_U7748
g5928 nand P3_U2574 P3_INSTQUEUE_REG_15__1__SCAN_IN ; P3_U7749
g5929 nand P3_U2572 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U7750
g5930 nand P3_U2571 P3_INSTQUEUE_REG_1__1__SCAN_IN ; P3_U7751
g5931 nand P3_U2570 P3_INSTQUEUE_REG_2__1__SCAN_IN ; P3_U7752
g5932 nand P3_U2569 P3_INSTQUEUE_REG_3__1__SCAN_IN ; P3_U7753
g5933 nand P3_U2567 P3_INSTQUEUE_REG_4__1__SCAN_IN ; P3_U7754
g5934 nand P3_U2566 P3_INSTQUEUE_REG_5__1__SCAN_IN ; P3_U7755
g5935 nand P3_U2565 P3_INSTQUEUE_REG_6__1__SCAN_IN ; P3_U7756
g5936 nand P3_U2564 P3_INSTQUEUE_REG_7__1__SCAN_IN ; P3_U7757
g5937 nand P3_U2582 P3_INSTQUEUE_REG_8__0__SCAN_IN ; P3_U7758
g5938 nand P3_U2581 P3_INSTQUEUE_REG_9__0__SCAN_IN ; P3_U7759
g5939 nand P3_U2580 P3_INSTQUEUE_REG_10__0__SCAN_IN ; P3_U7760
g5940 nand P3_U2579 P3_INSTQUEUE_REG_11__0__SCAN_IN ; P3_U7761
g5941 nand P3_U2577 P3_INSTQUEUE_REG_12__0__SCAN_IN ; P3_U7762
g5942 nand P3_U2576 P3_INSTQUEUE_REG_13__0__SCAN_IN ; P3_U7763
g5943 nand P3_U2575 P3_INSTQUEUE_REG_14__0__SCAN_IN ; P3_U7764
g5944 nand P3_U2574 P3_INSTQUEUE_REG_15__0__SCAN_IN ; P3_U7765
g5945 nand P3_U2572 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U7766
g5946 nand P3_U2571 P3_INSTQUEUE_REG_1__0__SCAN_IN ; P3_U7767
g5947 nand P3_U2570 P3_INSTQUEUE_REG_2__0__SCAN_IN ; P3_U7768
g5948 nand P3_U2569 P3_INSTQUEUE_REG_3__0__SCAN_IN ; P3_U7769
g5949 nand P3_U2567 P3_INSTQUEUE_REG_4__0__SCAN_IN ; P3_U7770
g5950 nand P3_U2566 P3_INSTQUEUE_REG_5__0__SCAN_IN ; P3_U7771
g5951 nand P3_U2565 P3_INSTQUEUE_REG_6__0__SCAN_IN ; P3_U7772
g5952 nand P3_U2564 P3_INSTQUEUE_REG_7__0__SCAN_IN ; P3_U7773
g5953 nand P3_U3097 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U7774
g5954 not P3_U3268 ; P3_U7775
g5955 nand P3_U2600 P3_INSTQUEUE_REG_8__7__SCAN_IN ; P3_U7776
g5956 nand P3_U2599 P3_INSTQUEUE_REG_9__7__SCAN_IN ; P3_U7777
g5957 nand P3_U2598 P3_INSTQUEUE_REG_10__7__SCAN_IN ; P3_U7778
g5958 nand P3_U2597 P3_INSTQUEUE_REG_11__7__SCAN_IN ; P3_U7779
g5959 nand P3_U2595 P3_INSTQUEUE_REG_12__7__SCAN_IN ; P3_U7780
g5960 nand P3_U2594 P3_INSTQUEUE_REG_13__7__SCAN_IN ; P3_U7781
g5961 nand P3_U2593 P3_INSTQUEUE_REG_14__7__SCAN_IN ; P3_U7782
g5962 nand P3_U2592 P3_INSTQUEUE_REG_15__7__SCAN_IN ; P3_U7783
g5963 nand P3_U2591 P3_INSTQUEUE_REG_0__7__SCAN_IN ; P3_U7784
g5964 nand P3_U2590 P3_INSTQUEUE_REG_1__7__SCAN_IN ; P3_U7785
g5965 nand P3_U2589 P3_INSTQUEUE_REG_2__7__SCAN_IN ; P3_U7786
g5966 nand P3_U2588 P3_INSTQUEUE_REG_3__7__SCAN_IN ; P3_U7787
g5967 nand P3_U2586 P3_INSTQUEUE_REG_4__7__SCAN_IN ; P3_U7788
g5968 nand P3_U2585 P3_INSTQUEUE_REG_5__7__SCAN_IN ; P3_U7789
g5969 nand P3_U2584 P3_INSTQUEUE_REG_6__7__SCAN_IN ; P3_U7790
g5970 nand P3_U2583 P3_INSTQUEUE_REG_7__7__SCAN_IN ; P3_U7791
g5971 nand P3_U2600 P3_INSTQUEUE_REG_8__6__SCAN_IN ; P3_U7792
g5972 nand P3_U2599 P3_INSTQUEUE_REG_9__6__SCAN_IN ; P3_U7793
g5973 nand P3_U2598 P3_INSTQUEUE_REG_10__6__SCAN_IN ; P3_U7794
g5974 nand P3_U2597 P3_INSTQUEUE_REG_11__6__SCAN_IN ; P3_U7795
g5975 nand P3_U2595 P3_INSTQUEUE_REG_12__6__SCAN_IN ; P3_U7796
g5976 nand P3_U2594 P3_INSTQUEUE_REG_13__6__SCAN_IN ; P3_U7797
g5977 nand P3_U2593 P3_INSTQUEUE_REG_14__6__SCAN_IN ; P3_U7798
g5978 nand P3_U2592 P3_INSTQUEUE_REG_15__6__SCAN_IN ; P3_U7799
g5979 nand P3_U2591 P3_INSTQUEUE_REG_0__6__SCAN_IN ; P3_U7800
g5980 nand P3_U2590 P3_INSTQUEUE_REG_1__6__SCAN_IN ; P3_U7801
g5981 nand P3_U2589 P3_INSTQUEUE_REG_2__6__SCAN_IN ; P3_U7802
g5982 nand P3_U2588 P3_INSTQUEUE_REG_3__6__SCAN_IN ; P3_U7803
g5983 nand P3_U2586 P3_INSTQUEUE_REG_4__6__SCAN_IN ; P3_U7804
g5984 nand P3_U2585 P3_INSTQUEUE_REG_5__6__SCAN_IN ; P3_U7805
g5985 nand P3_U2584 P3_INSTQUEUE_REG_6__6__SCAN_IN ; P3_U7806
g5986 nand P3_U2583 P3_INSTQUEUE_REG_7__6__SCAN_IN ; P3_U7807
g5987 nand P3_U2600 P3_INSTQUEUE_REG_8__5__SCAN_IN ; P3_U7808
g5988 nand P3_U2599 P3_INSTQUEUE_REG_9__5__SCAN_IN ; P3_U7809
g5989 nand P3_U2598 P3_INSTQUEUE_REG_10__5__SCAN_IN ; P3_U7810
g5990 nand P3_U2597 P3_INSTQUEUE_REG_11__5__SCAN_IN ; P3_U7811
g5991 nand P3_U2595 P3_INSTQUEUE_REG_12__5__SCAN_IN ; P3_U7812
g5992 nand P3_U2594 P3_INSTQUEUE_REG_13__5__SCAN_IN ; P3_U7813
g5993 nand P3_U2593 P3_INSTQUEUE_REG_14__5__SCAN_IN ; P3_U7814
g5994 nand P3_U2592 P3_INSTQUEUE_REG_15__5__SCAN_IN ; P3_U7815
g5995 nand P3_U2591 P3_INSTQUEUE_REG_0__5__SCAN_IN ; P3_U7816
g5996 nand P3_U2590 P3_INSTQUEUE_REG_1__5__SCAN_IN ; P3_U7817
g5997 nand P3_U2589 P3_INSTQUEUE_REG_2__5__SCAN_IN ; P3_U7818
g5998 nand P3_U2588 P3_INSTQUEUE_REG_3__5__SCAN_IN ; P3_U7819
g5999 nand P3_U2586 P3_INSTQUEUE_REG_4__5__SCAN_IN ; P3_U7820
g6000 nand P3_U2585 P3_INSTQUEUE_REG_5__5__SCAN_IN ; P3_U7821
g6001 nand P3_U2584 P3_INSTQUEUE_REG_6__5__SCAN_IN ; P3_U7822
g6002 nand P3_U2583 P3_INSTQUEUE_REG_7__5__SCAN_IN ; P3_U7823
g6003 nand P3_U2600 P3_INSTQUEUE_REG_8__4__SCAN_IN ; P3_U7824
g6004 nand P3_U2599 P3_INSTQUEUE_REG_9__4__SCAN_IN ; P3_U7825
g6005 nand P3_U2598 P3_INSTQUEUE_REG_10__4__SCAN_IN ; P3_U7826
g6006 nand P3_U2597 P3_INSTQUEUE_REG_11__4__SCAN_IN ; P3_U7827
g6007 nand P3_U2595 P3_INSTQUEUE_REG_12__4__SCAN_IN ; P3_U7828
g6008 nand P3_U2594 P3_INSTQUEUE_REG_13__4__SCAN_IN ; P3_U7829
g6009 nand P3_U2593 P3_INSTQUEUE_REG_14__4__SCAN_IN ; P3_U7830
g6010 nand P3_U2592 P3_INSTQUEUE_REG_15__4__SCAN_IN ; P3_U7831
g6011 nand P3_U2591 P3_INSTQUEUE_REG_0__4__SCAN_IN ; P3_U7832
g6012 nand P3_U2590 P3_INSTQUEUE_REG_1__4__SCAN_IN ; P3_U7833
g6013 nand P3_U2589 P3_INSTQUEUE_REG_2__4__SCAN_IN ; P3_U7834
g6014 nand P3_U2588 P3_INSTQUEUE_REG_3__4__SCAN_IN ; P3_U7835
g6015 nand P3_U2586 P3_INSTQUEUE_REG_4__4__SCAN_IN ; P3_U7836
g6016 nand P3_U2585 P3_INSTQUEUE_REG_5__4__SCAN_IN ; P3_U7837
g6017 nand P3_U2584 P3_INSTQUEUE_REG_6__4__SCAN_IN ; P3_U7838
g6018 nand P3_U2583 P3_INSTQUEUE_REG_7__4__SCAN_IN ; P3_U7839
g6019 nand P3_U2600 P3_INSTQUEUE_REG_8__3__SCAN_IN ; P3_U7840
g6020 nand P3_U2599 P3_INSTQUEUE_REG_9__3__SCAN_IN ; P3_U7841
g6021 nand P3_U2598 P3_INSTQUEUE_REG_10__3__SCAN_IN ; P3_U7842
g6022 nand P3_U2597 P3_INSTQUEUE_REG_11__3__SCAN_IN ; P3_U7843
g6023 nand P3_U2595 P3_INSTQUEUE_REG_12__3__SCAN_IN ; P3_U7844
g6024 nand P3_U2594 P3_INSTQUEUE_REG_13__3__SCAN_IN ; P3_U7845
g6025 nand P3_U2593 P3_INSTQUEUE_REG_14__3__SCAN_IN ; P3_U7846
g6026 nand P3_U2592 P3_INSTQUEUE_REG_15__3__SCAN_IN ; P3_U7847
g6027 nand P3_U2591 P3_INSTQUEUE_REG_0__3__SCAN_IN ; P3_U7848
g6028 nand P3_U2590 P3_INSTQUEUE_REG_1__3__SCAN_IN ; P3_U7849
g6029 nand P3_U2589 P3_INSTQUEUE_REG_2__3__SCAN_IN ; P3_U7850
g6030 nand P3_U2588 P3_INSTQUEUE_REG_3__3__SCAN_IN ; P3_U7851
g6031 nand P3_U2586 P3_INSTQUEUE_REG_4__3__SCAN_IN ; P3_U7852
g6032 nand P3_U2585 P3_INSTQUEUE_REG_5__3__SCAN_IN ; P3_U7853
g6033 nand P3_U2584 P3_INSTQUEUE_REG_6__3__SCAN_IN ; P3_U7854
g6034 nand P3_U2583 P3_INSTQUEUE_REG_7__3__SCAN_IN ; P3_U7855
g6035 nand P3_U2600 P3_INSTQUEUE_REG_8__2__SCAN_IN ; P3_U7856
g6036 nand P3_U2599 P3_INSTQUEUE_REG_9__2__SCAN_IN ; P3_U7857
g6037 nand P3_U2598 P3_INSTQUEUE_REG_10__2__SCAN_IN ; P3_U7858
g6038 nand P3_U2597 P3_INSTQUEUE_REG_11__2__SCAN_IN ; P3_U7859
g6039 nand P3_U2595 P3_INSTQUEUE_REG_12__2__SCAN_IN ; P3_U7860
g6040 nand P3_U2594 P3_INSTQUEUE_REG_13__2__SCAN_IN ; P3_U7861
g6041 nand P3_U2593 P3_INSTQUEUE_REG_14__2__SCAN_IN ; P3_U7862
g6042 nand P3_U2592 P3_INSTQUEUE_REG_15__2__SCAN_IN ; P3_U7863
g6043 nand P3_U2591 P3_INSTQUEUE_REG_0__2__SCAN_IN ; P3_U7864
g6044 nand P3_U2590 P3_INSTQUEUE_REG_1__2__SCAN_IN ; P3_U7865
g6045 nand P3_U2589 P3_INSTQUEUE_REG_2__2__SCAN_IN ; P3_U7866
g6046 nand P3_U2588 P3_INSTQUEUE_REG_3__2__SCAN_IN ; P3_U7867
g6047 nand P3_U2586 P3_INSTQUEUE_REG_4__2__SCAN_IN ; P3_U7868
g6048 nand P3_U2585 P3_INSTQUEUE_REG_5__2__SCAN_IN ; P3_U7869
g6049 nand P3_U2584 P3_INSTQUEUE_REG_6__2__SCAN_IN ; P3_U7870
g6050 nand P3_U2583 P3_INSTQUEUE_REG_7__2__SCAN_IN ; P3_U7871
g6051 nand P3_U2600 P3_INSTQUEUE_REG_8__1__SCAN_IN ; P3_U7872
g6052 nand P3_U2599 P3_INSTQUEUE_REG_9__1__SCAN_IN ; P3_U7873
g6053 nand P3_U2598 P3_INSTQUEUE_REG_10__1__SCAN_IN ; P3_U7874
g6054 nand P3_U2597 P3_INSTQUEUE_REG_11__1__SCAN_IN ; P3_U7875
g6055 nand P3_U2595 P3_INSTQUEUE_REG_12__1__SCAN_IN ; P3_U7876
g6056 nand P3_U2594 P3_INSTQUEUE_REG_13__1__SCAN_IN ; P3_U7877
g6057 nand P3_U2593 P3_INSTQUEUE_REG_14__1__SCAN_IN ; P3_U7878
g6058 nand P3_U2592 P3_INSTQUEUE_REG_15__1__SCAN_IN ; P3_U7879
g6059 nand P3_U2591 P3_INSTQUEUE_REG_0__1__SCAN_IN ; P3_U7880
g6060 nand P3_U2590 P3_INSTQUEUE_REG_1__1__SCAN_IN ; P3_U7881
g6061 nand P3_U2589 P3_INSTQUEUE_REG_2__1__SCAN_IN ; P3_U7882
g6062 nand P3_U2588 P3_INSTQUEUE_REG_3__1__SCAN_IN ; P3_U7883
g6063 nand P3_U2586 P3_INSTQUEUE_REG_4__1__SCAN_IN ; P3_U7884
g6064 nand P3_U2585 P3_INSTQUEUE_REG_5__1__SCAN_IN ; P3_U7885
g6065 nand P3_U2584 P3_INSTQUEUE_REG_6__1__SCAN_IN ; P3_U7886
g6066 nand P3_U2583 P3_INSTQUEUE_REG_7__1__SCAN_IN ; P3_U7887
g6067 nand P3_U2600 P3_INSTQUEUE_REG_8__0__SCAN_IN ; P3_U7888
g6068 nand P3_U2599 P3_INSTQUEUE_REG_9__0__SCAN_IN ; P3_U7889
g6069 nand P3_U2598 P3_INSTQUEUE_REG_10__0__SCAN_IN ; P3_U7890
g6070 nand P3_U2597 P3_INSTQUEUE_REG_11__0__SCAN_IN ; P3_U7891
g6071 nand P3_U2595 P3_INSTQUEUE_REG_12__0__SCAN_IN ; P3_U7892
g6072 nand P3_U2594 P3_INSTQUEUE_REG_13__0__SCAN_IN ; P3_U7893
g6073 nand P3_U2593 P3_INSTQUEUE_REG_14__0__SCAN_IN ; P3_U7894
g6074 nand P3_U2592 P3_INSTQUEUE_REG_15__0__SCAN_IN ; P3_U7895
g6075 nand P3_U2591 P3_INSTQUEUE_REG_0__0__SCAN_IN ; P3_U7896
g6076 nand P3_U2590 P3_INSTQUEUE_REG_1__0__SCAN_IN ; P3_U7897
g6077 nand P3_U2589 P3_INSTQUEUE_REG_2__0__SCAN_IN ; P3_U7898
g6078 nand P3_U2588 P3_INSTQUEUE_REG_3__0__SCAN_IN ; P3_U7899
g6079 nand P3_U2586 P3_INSTQUEUE_REG_4__0__SCAN_IN ; P3_U7900
g6080 nand P3_U2585 P3_INSTQUEUE_REG_5__0__SCAN_IN ; P3_U7901
g6081 nand P3_U2584 P3_INSTQUEUE_REG_6__0__SCAN_IN ; P3_U7902
g6082 nand P3_U2583 P3_INSTQUEUE_REG_7__0__SCAN_IN ; P3_U7903
g6083 nand P3_U4292 P3_STATE_REG_0__SCAN_IN ; P3_U7904
g6084 or U209 P3_STATE2_REG_2__SCAN_IN ; P3_U7905
g6085 nand P3_U3939 P3_U6397 ; P3_U7906
g6086 nand P3_U4134 P3_U2603 ; P3_U7907
g6087 nand P3_U2404 P3_U3256 ; P3_U7908
g6088 nand P3_U2392 P3_U7096 ; P3_U7909
g6089 nand P3_U7908 P3_U4317 P3_U7909 ; P3_U7910
g6090 not P3_U3086 ; P3_U7911
g6091 nand P3_U7911 P3_U3088 ; P3_U7912
g6092 nand P3_U4449 P3_U4446 P3_STATE_REG_1__SCAN_IN ; P3_U7913
g6093 nand P3_U7904 P3_STATE_REG_2__SCAN_IN ; P3_U7914
g6094 nand P3_U4446 P3_STATE_REG_1__SCAN_IN ; P3_U7915
g6095 nand P3_U4505 P3_U3106 ; P3_U7916
g6096 nand P3_U4488 P3_U4522 ; P3_U7917
g6097 nand P3_U3208 P3_U3219 ; P3_U7918
g6098 nand P3_U7376 P3_U3105 ; P3_U7919
g6099 nand P3_U3077 P3_BE_N_REG_3__SCAN_IN ; P3_U7920
g6100 nand P3_U4308 P3_BYTEENABLE_REG_3__SCAN_IN ; P3_U7921
g6101 nand P3_U3077 P3_BE_N_REG_2__SCAN_IN ; P3_U7922
g6102 nand P3_U4308 P3_BYTEENABLE_REG_2__SCAN_IN ; P3_U7923
g6103 nand P3_U3077 P3_BE_N_REG_1__SCAN_IN ; P3_U7924
g6104 nand P3_U4308 P3_BYTEENABLE_REG_1__SCAN_IN ; P3_U7925
g6105 nand P3_U3077 P3_BE_N_REG_0__SCAN_IN ; P3_U7926
g6106 nand P3_U4308 P3_BYTEENABLE_REG_0__SCAN_IN ; P3_U7927
g6107 nand P3_U3079 P3_STATE_REG_0__SCAN_IN P3_REQUESTPENDING_REG_SCAN_IN ; P3_U7928
g6108 nand P3_U3086 P3_STATE_REG_2__SCAN_IN ; P3_U7929
g6109 nand P3_U7929 P3_U7928 ; P3_U7930
g6110 nand P3_U7914 P3_U4449 P3_STATE_REG_1__SCAN_IN ; P3_U7931
g6111 nand P3_U7930 P3_U3076 ; P3_U7932
g6112 nand P3_U3087 P3_STATE_REG_2__SCAN_IN P3_STATE_REG_0__SCAN_IN ; P3_U7933
g6113 nand P3_U4459 P3_U3079 ; P3_U7934
g6114 or P3_STATE_REG_1__SCAN_IN P3_STATE_REG_0__SCAN_IN ; P3_U7935
g6115 nand P3_U4346 P3_STATE_REG_0__SCAN_IN ; P3_U7936
g6116 not P3_U3278 ; P3_U7937
g6117 nand P3_U7937 P3_DATAWIDTH_REG_0__SCAN_IN ; P3_U7938
g6118 nand P3_U3279 P3_U3278 ; P3_U7939
g6119 nand P3_U3278 P3_U4464 ; P3_U7940
g6120 nand P3_U7937 P3_DATAWIDTH_REG_1__SCAN_IN ; P3_U7941
g6121 nand P3_U4505 P3_U3211 ; P3_U7942
g6122 nand P3_U3104 P3_U3214 ; P3_U7943
g6123 nand P3_U4505 P3_U3213 ; P3_U7944
g6124 nand P3_U3104 P3_U3210 ; P3_U7945
g6125 nand P3_U4539 P3_U4618 ; P3_U7946
g6126 nand P3_U4620 P3_U3101 ; P3_U7947
g6127 nand P3_U4281 P3_U4617 ; P3_U7948
g6128 nand P3_U4622 P3_U4624 ; P3_U7949
g6129 nand P3_U4505 P3_U3237 ; P3_U7950
g6130 nand P3_U3104 P3_U3238 ; P3_U7951
g6131 nand P3_U4627 P3_STATE2_REG_0__SCAN_IN ; P3_U7952
g6132 nand P3_U4628 P3_U3121 ; P3_U7953
g6133 nand P3_U3122 P3_STATE2_REG_3__SCAN_IN ; P3_U7954
g6134 nand P3_U2453 P3_U4630 ; P3_U7955
g6135 or P3_STATE2_REG_0__SCAN_IN P3_STATEBS16_REG_SCAN_IN ; P3_U7956
g6136 nand P3_U7905 P3_STATE2_REG_0__SCAN_IN ; P3_U7957
g6137 nand P3_U4638 P3_STATE2_REG_0__SCAN_IN ; P3_U7958
g6138 nand P3_U4637 P3_U4629 P3_U3121 ; P3_U7959
g6139 nand P3_U3130 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_U7960
g6140 nand P3_U4648 P3_U3131 ; P3_U7961
g6141 not P3_U3269 ; P3_U7962
g6142 nand P3_U7962 P3_U4653 ; P3_U7963
g6143 nand P3_U3269 P3_U3138 ; P3_U7964
g6144 not P3_U3270 ; P3_U7965
g6145 nand P3_U7965 P3_U4657 ; P3_U7966
g6146 nand P3_U3270 P3_U3140 ; P3_U7967
g6147 not P3_U3271 ; P3_U7968
g6148 nand P3_U3109 P3_U3101 ; P3_U7969
g6149 nand P3_U4539 P3_U5483 ; P3_U7970
g6150 nand P3_U3283 P3_U4283 ; P3_U7971
g6151 nand P3_U5499 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_U7972
g6152 nand P3_U3218 P3_U3107 ; P3_U7973
g6153 nand P3_U4573 P3_U4590 ; P3_U7974
g6154 nand P3_U4539 P3_U5512 ; P3_U7975
g6155 nand P3_U5515 P3_U3101 ; P3_U7976
g6156 nand P3_U4556 P3_U5517 P3_U3110 ; P3_U7977
g6157 nand P3_U5513 P3_U3107 P3_U4590 ; P3_U7978
g6158 nand P3_U5499 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U7979
g6159 nand P3_U5546 P3_U4283 ; P3_U7980
g6160 nand P3_U3221 P3_U3094 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U7981
g6161 nand P3_U5531 P3_U3097 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U7982
g6162 nand P3_U4284 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_U7983
g6163 nand P3_SUB_580_U6 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_U7984
g6164 not P3_U3287 ; P3_U7985
g6165 nand P3_U4284 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_U7986
g6166 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_U7987
g6167 not P3_U3286 ; P3_U7988
g6168 nand P3_U5499 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U7989
g6169 nand P3_U5557 P3_U4283 ; P3_U7990
g6170 nand P3_U5499 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U7991
g6171 nand P3_U5570 P3_U4283 ; P3_U7992
g6172 nand P3_U3221 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U7993
g6173 nand P3_U5571 P3_U3093 ; P3_U7994
g6174 nand P3_U5499 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U7995
g6175 nand P3_U5577 P3_U4283 ; P3_U7996
g6176 nand P3_U7968 P3_U4647 ; P3_U7997
g6177 nand P3_U3271 P3_U3143 ; P3_U7998
g6178 nand P3_U7998 P3_U7997 ; P3_U7999
g6179 nand P3_U5622 P3_U3104 ; P3_U8000
g6180 nand P3_U4505 P3_U5619 ; P3_U8001
g6181 nand P3_U3261 P3_BYTEENABLE_REG_3__SCAN_IN ; P3_U8002
g6182 nand P3_U3291 P3_U4307 ; P3_U8003
g6183 or P3_DATAWIDTH_REG_0__SCAN_IN P3_DATAWIDTH_REG_1__SCAN_IN ; P3_U8004
g6184 nand P3_U3240 P3_DATAWIDTH_REG_0__SCAN_IN ; P3_U8005
g6185 nand P3_U8005 P3_U8004 ; P3_U8006
g6186 nand P3_U8006 P3_U3081 ; P3_U8007
g6187 nand P3_REIP_REG_0__SCAN_IN P3_REIP_REG_1__SCAN_IN ; P3_U8008
g6188 nand P3_U8008 P3_U8007 ; P3_U8009
g6189 nand P3_U3261 P3_BYTEENABLE_REG_2__SCAN_IN ; P3_U8010
g6190 nand P3_U8009 P3_U4307 ; P3_U8011
g6191 nand P3_U3261 P3_BYTEENABLE_REG_1__SCAN_IN ; P3_U8012
g6192 nand P3_U4307 P3_REIP_REG_1__SCAN_IN ; P3_U8013
g6193 nand P3_U3261 P3_BYTEENABLE_REG_0__SCAN_IN ; P3_U8014
g6194 nand P3_U4307 P3_U7367 ; P3_U8015
g6195 nand P3_U4308 P3_U3264 ; P3_U8016
g6196 nand P3_U3077 P3_W_R_N_REG_SCAN_IN ; P3_U8017
g6197 nand P3_U7368 P3_U4617 ; P3_U8018
g6198 nand P3_U4285 P3_MORE_REG_SCAN_IN ; P3_U8019
g6199 nand P3_U7937 P3_STATEBS16_REG_SCAN_IN ; P3_U8020
g6200 nand BS16 P3_U3278 ; P3_U8021
g6201 nand P3_U7374 P3_REQUESTPENDING_REG_SCAN_IN ; P3_U8022
g6202 nand P3_U7379 P3_U4287 ; P3_U8023
g6203 nand P3_U4308 P3_U3263 ; P3_U8024
g6204 nand P3_U3077 P3_D_C_N_REG_SCAN_IN ; P3_U8025
g6205 nand P3_U3077 P3_M_IO_N_REG_SCAN_IN ; P3_U8026
g6206 nand P3_U4308 P3_MEMORYFETCH_REG_SCAN_IN ; P3_U8027
g6207 nand P3_U7384 P3_READREQUEST_REG_SCAN_IN ; P3_U8028
g6208 nand P3_U7385 P3_U4288 ; P3_U8029
g6209 nand P3_U7384 P3_MEMORYFETCH_REG_SCAN_IN ; P3_U8030
g6210 nand P3_U7386 P3_U4288 ; P3_U8031
g6211 nand P3_U3097 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U8032
g6212 nand P3_U3094 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U8033
g6213 not P3_U3272 ; P3_U8034
g6214 nand P3_U4289 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U8035
g6215 nand P3_U7645 P3_U3100 ; P3_U8036
g6216 not P3_U3273 ; P3_U8037
g6217 nand P3_U3207 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U8038
g6218 nand P3_U3287 P3_U3286 P3_FLUSH_REG_SCAN_IN ; P3_U8039
g6219 nand P3_U3207 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U8040
g6220 nand P3_U3286 P3_U7985 P3_FLUSH_REG_SCAN_IN ; P3_U8041
g6221 nand P3_U3207 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U8042
g6222 nand P3_U7988 P3_FLUSH_REG_SCAN_IN ; P3_U8043
g6223 nand P3_U3303 P3_U4290 ; P3_U8044
g6224 nand P3_U5496 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_U8045
g6225 nand P3_U5496 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_U8046
g6226 nand P3_U5542 P3_U4290 ; P3_U8047
g6227 nand P3_U5496 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_U8048
g6228 nand P3_U5553 P3_U4290 ; P3_U8049
g6229 nand P3_U5496 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_U8050
g6230 nand P3_U5566 P3_U4290 ; P3_U8051
g6231 nand P3_U5496 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_U8052
g6232 nand P3_U5573 P3_U4290 ; P3_U8053
g6233 and P2_U2617 P2_U3300 P2_U7873 ; P2_U2352
g6234 and P2_U4343 P2_U2439 ; P2_U2353
g6235 and P2_U7861 P2_U7873 P2_STATE2_REG_0__SCAN_IN ; P2_U2354
g6236 and P2_U2447 P2_U7861 ; P2_U2355
g6237 and P2_U3253 P2_STATE2_REG_0__SCAN_IN ; P2_U2356
g6238 and P2_U3712 P2_U2458 ; P2_U2357
g6239 and P2_U4431 P2_STATE2_REG_0__SCAN_IN ; P2_U2358
g6240 and P2_U4411 P2_U3265 ; P2_U2359
g6241 nor U211 P2_STATEBS16_REG_SCAN_IN ; P2_U2360
g6242 and P2_R2238_U6 P2_U2356 ; P2_U2361
g6243 and P2_U2398 P2_U4443 ; P2_U2362
g6244 and P2_U3535 P2_STATE2_REG_2__SCAN_IN ; P2_U2363
g6245 and P2_U3546 P2_STATE2_REG_2__SCAN_IN ; P2_U2364
g6246 and P2_U4443 P2_STATE2_REG_3__SCAN_IN ; P2_U2365
g6247 and P2_U3546 P2_STATE2_REG_1__SCAN_IN ; P2_U2366
g6248 and P2_U2364 P2_U4417 ; P2_U2367
g6249 and P2_U2363 P2_U4420 ; P2_U2368
g6250 and P2_U2364 P2_U4428 ; P2_U2369
g6251 and P2_U2447 P2_U3537 ; P2_U2370
g6252 and P2_U3990 P2_U3537 ; P2_U2371
g6253 and P2_U3989 P2_U3537 ; P2_U2372
g6254 and P2_U4419 P2_U3537 ; P2_U2373
g6255 and P2_U4468 P2_STATE2_REG_0__SCAN_IN ; P2_U2374
g6256 and P2_U4441 P2_U3521 ; P2_U2375
g6257 and P2_U3873 P2_U2436 ; P2_U2376
g6258 and P2_U2367 P2_U4411 ; P2_U2377
g6259 and P2_U3546 P2_STATE2_REG_3__SCAN_IN ; P2_U2378
g6260 and P2_U4440 P2_U7865 ; P2_U2379
g6261 and P2_U4441 P2_U7865 ; P2_U2380
g6262 and P2_U3535 P2_U3270 ; P2_U2381
g6263 and P2_U2366 P2_U3647 ; P2_U2382
g6264 and P2_U2366 P2_U3528 ; P2_U2383
g6265 and P2_U2368 P2_U4417 ; P2_U2384
g6266 and P2_U2368 P2_U4428 ; P2_U2385
g6267 and P2_U2363 P2_U4436 ; P2_U2386
g6268 and P2_U5940 P2_U3537 ; P2_U2387
g6269 and P2_U2363 P2_U5675 ; P2_U2388
g6270 and P2_U2363 P2_U5677 ; P2_U2389
g6271 and P2_U2363 P2_U5679 ; P2_U2390
g6272 and P2_U2369 P2_U3545 ; P2_U2391
g6273 and P2_U6571 P2_U2369 ; P2_U2392
g6274 and P2_U4440 P2_U3521 ; P2_U2393
g6275 and P2_U4442 P2_U2616 ; P2_U2394
g6276 and P2_U4442 P2_U7873 ; P2_U2395
g6277 and P2_U3541 P2_U3284 ; P2_U2396
g6278 and P2_U4441 P2_U4601 ; P2_U2397
g6279 and P2_U4430 P2_STATEBS16_REG_SCAN_IN ; P2_U2398
g6280 and U314 P2_U4443 ; P2_U2399
g6281 and U303 P2_U4443 ; P2_U2400
g6282 and U292 P2_U4443 ; P2_U2401
g6283 and U289 P2_U4443 ; P2_U2402
g6284 and U288 P2_U4443 ; P2_U2403
g6285 and U287 P2_U4443 ; P2_U2404
g6286 and U286 P2_U4443 ; P2_U2405
g6287 and U285 P2_U4443 ; P2_U2406
g6288 and U298 P2_U2362 ; P2_U2407
g6289 and U307 P2_U2362 ; P2_U2408
g6290 and U297 P2_U2362 ; P2_U2409
g6291 and U306 P2_U2362 ; P2_U2410
g6292 and U296 P2_U2362 ; P2_U2411
g6293 and U305 P2_U2362 ; P2_U2412
g6294 and U295 P2_U2362 ; P2_U2413
g6295 and U304 P2_U2362 ; P2_U2414
g6296 and U294 P2_U2362 ; P2_U2415
g6297 and U302 P2_U2362 ; P2_U2416
g6298 and U293 P2_U2362 ; P2_U2417
g6299 and U301 P2_U2362 ; P2_U2418
g6300 and U291 P2_U2362 ; P2_U2419
g6301 and U300 P2_U2362 ; P2_U2420
g6302 and U290 P2_U2362 ; P2_U2421
g6303 and U299 P2_U2362 ; P2_U2422
g6304 and P2_U2365 P2_U3255 ; P2_U2423
g6305 and P2_U2365 P2_U3278 ; P2_U2424
g6306 and P2_U2365 P2_U3521 ; P2_U2425
g6307 and P2_U2365 P2_U3279 ; P2_U2426
g6308 and P2_U2375 P2_U3279 ; P2_U2427
g6309 and P2_U2365 P2_U2616 ; P2_U2428
g6310 and P2_U2365 P2_U2617 ; P2_U2429
g6311 and P2_U3541 P2_STATE2_REG_0__SCAN_IN ; P2_U2430
g6312 and P2_U2365 P2_U3253 ; P2_U2431
g6313 and P2_U2365 P2_U3280 ; P2_U2432
g6314 and P2_U2375 P2_U3295 ; P2_U2433
g6315 and P2_U2375 P2_U7869 ; P2_U2434
g6316 and P2_U2356 P2_U3541 ; P2_U2435
g6317 and P2_U7859 P2_U7867 ; P2_U2436
g6318 and P2_U2364 P2_U7871 ; P2_U2437
g6319 and P2_U7859 P2_U3278 ; P2_U2438
g6320 and P2_U4339 P2_U3521 ; P2_U2439
g6321 and P2_U3580 P2_U3428 ; P2_U2440
g6322 and P2_U4647 P2_U3580 ; P2_U2441
g6323 and P2_U8067 P2_U3428 ; P2_U2442
g6324 and P2_U4647 P2_U8067 ; P2_U2443
g6325 and P2_U3243 P2_U3307 ; P2_U2444
g6326 and P2_U4650 P2_U3307 ; P2_U2445
g6327 and P2_R2088_U6 P2_U4424 ; P2_U2446
g6328 and P2_U2616 P2_STATE2_REG_0__SCAN_IN ; P2_U2447
g6329 and P2_STATE2_REG_2__SCAN_IN P2_STATE2_REG_1__SCAN_IN ; P2_U2448
g6330 and P2_U3278 P2_U3521 ; P2_U2449
g6331 and P2_U2354 P2_U7871 ; P2_U2450
g6332 and P2_U4601 P2_U2457 P2_U2438 ; P2_U2451
g6333 and P2_U3272 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U2452
g6334 and P2_U3271 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2453
g6335 and P2_U3271 P2_U3272 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U2454
g6336 and P2_U3276 P2_U3272 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U2455
g6337 and P2_U3276 P2_U3271 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2456
g6338 and P2_U3521 P2_U3255 ; P2_U2457
g6339 and P2_U2617 P2_U3279 P2_U7863 ; P2_U2458
g6340 and P2_U8053 P2_U8052 P2_U4393 ; P2_U2459
g6341 and P2_R2182_U40 P2_U3317 ; P2_U2460
g6342 and P2_U3579 P2_U3426 ; P2_U2461
g6343 and P2_R2182_U76 P2_R2182_U40 ; P2_U2462
g6344 and P2_U4637 P2_U2462 ; P2_U2463
g6345 and P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U2464
g6346 and P2_U3309 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U2465
g6347 and P2_R2099_U96 P2_R2099_U95 ; P2_U2466
g6348 and P2_R2099_U5 P2_R2099_U94 ; P2_U2467
g6349 and P2_U3320 P2_U4657 ; P2_U2468
g6350 and P2_U4633 P2_U2462 ; P2_U2469
g6351 and P2_R2099_U5 P2_U3323 ; P2_U2470
g6352 and P2_U3339 P2_U4715 ; P2_U2471
g6353 and P2_U4634 P2_U2462 ; P2_U2472
g6354 and P2_R2099_U94 P2_U3324 ; P2_U2473
g6355 and P2_U3354 P2_U4774 ; P2_U2474
g6356 and P2_U4635 P2_R2182_U69 ; P2_U2475
g6357 nor P2_R2182_U69 P2_R2182_U68 ; P2_U2476
g6358 and P2_U2476 P2_U2462 ; P2_U2477
g6359 nor P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U2478
g6360 nor P2_R2099_U94 P2_R2099_U5 ; P2_U2479
g6361 and P2_U3366 P2_U4831 ; P2_U2480
g6362 and P2_U8064 P2_U3426 ; P2_U2481
g6363 and P2_U4638 P2_U4637 ; P2_U2482
g6364 and P2_R2099_U95 P2_U3322 ; P2_U2483
g6365 and P2_U3379 P2_U4889 ; P2_U2484
g6366 and P2_U4638 P2_U4633 ; P2_U2485
g6367 and P2_U3391 P2_U4946 ; P2_U2486
g6368 and P2_U4638 P2_U4634 ; P2_U2487
g6369 and P2_U3402 P2_U5004 ; P2_U2488
g6370 and P2_U4638 P2_U2476 ; P2_U2489
g6371 and P2_U3414 P2_U5061 ; P2_U2490
g6372 and P2_U4640 P2_U3579 ; P2_U2491
g6373 and P2_R2099_U96 P2_U3321 ; P2_U2492
g6374 and P2_U3427 P2_U3425 ; P2_U2493
g6375 and P2_U4633 P2_U2460 ; P2_U2494
g6376 and P2_U3440 P2_U5174 ; P2_U2495
g6377 and P2_U4634 P2_U2460 ; P2_U2496
g6378 and P2_U3451 P2_U5232 ; P2_U2497
g6379 and P2_U2476 P2_U2460 ; P2_U2498
g6380 and P2_U3463 P2_U5289 ; P2_U2499
g6381 and P2_U4640 P2_U8064 ; P2_U2500
g6382 nor P2_R2182_U40 P2_R2182_U76 ; P2_U2501
g6383 and P2_U2501 P2_U4637 ; P2_U2502
g6384 nor P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U2503
g6385 nor P2_R2099_U95 P2_R2099_U96 ; P2_U2504
g6386 and P2_U3474 P2_U5347 ; P2_U2505
g6387 and P2_U2501 P2_U4633 ; P2_U2506
g6388 and P2_U3486 P2_U5404 ; P2_U2507
g6389 and P2_U2501 P2_U4634 ; P2_U2508
g6390 and P2_U3497 P2_U5462 ; P2_U2509
g6391 and P2_U2501 P2_U2476 ; P2_U2510
g6392 and P2_U3509 P2_U5519 ; P2_U2511
g6393 and P2_U8069 P2_U8068 P2_U3869 ; P2_U2512
g6394 and P2_U5580 P2_U5579 ; P2_U2513
g6395 and P2_U3881 P2_U7896 P2_U3882 ; P2_U2514
g6396 and P2_U8082 P2_U8100 ; P2_U2515
g6397 and P2_U5616 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2516
g6398 and P2_U2515 P2_U2516 ; P2_U2517
g6399 and P2_U5616 P2_U3272 ; P2_U2518
g6400 and P2_U2515 P2_U2518 ; P2_U2519
g6401 and P2_U8082 P2_U3582 ; P2_U2520
g6402 and P2_U2520 P2_U2516 ; P2_U2521
g6403 and P2_U2520 P2_U2518 ; P2_U2522
g6404 and P2_U3530 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2523
g6405 and P2_U2515 P2_U2523 ; P2_U2524
g6406 and P2_U3272 P2_U3530 ; P2_U2525
g6407 and P2_U2515 P2_U2525 ; P2_U2526
g6408 and P2_U2520 P2_U2523 ; P2_U2527
g6409 and P2_U2520 P2_U2525 ; P2_U2528
g6410 and P2_U3582 P2_U3581 ; P2_U2529
g6411 and P2_U2525 P2_U2529 ; P2_U2530
g6412 and P2_U2523 P2_U2529 ; P2_U2531
g6413 and P2_U8100 P2_U3581 ; P2_U2532
g6414 and P2_U2525 P2_U2532 ; P2_U2533
g6415 and P2_U2523 P2_U2532 ; P2_U2534
g6416 and P2_U2529 P2_U2518 ; P2_U2535
g6417 and P2_U2529 P2_U2516 ; P2_U2536
g6418 and P2_U2518 P2_U2532 ; P2_U2537
g6419 and P2_U2516 P2_U2532 ; P2_U2538
g6420 nor P2_R2147_U8 P2_R2147_U4 ; P2_U2539
g6421 nor P2_R2147_U9 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2540
g6422 and P2_U2539 P2_U2540 ; P2_U2541
g6423 and P2_U3529 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2542
g6424 and P2_U2539 P2_U2542 ; P2_U2543
g6425 and P2_R2147_U4 P2_U3526 ; P2_U2544
g6426 and P2_U2544 P2_U2540 ; P2_U2545
g6427 and P2_U2544 P2_U2542 ; P2_U2546
g6428 and P2_R2147_U9 P2_U3532 ; P2_U2547
g6429 and P2_U2539 P2_U2547 ; P2_U2548
g6430 and P2_R2147_U9 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2549
g6431 and P2_U2539 P2_U2549 ; P2_U2550
g6432 and P2_U2544 P2_U2547 ; P2_U2551
g6433 and P2_U2544 P2_U2549 ; P2_U2552
g6434 and P2_R2147_U8 P2_U3531 ; P2_U2553
g6435 and P2_U2540 P2_U2553 ; P2_U2554
g6436 and P2_U2542 P2_U2553 ; P2_U2555
g6437 and P2_R2147_U4 P2_R2147_U8 ; P2_U2556
g6438 and P2_U2540 P2_U2556 ; P2_U2557
g6439 and P2_U2542 P2_U2556 ; P2_U2558
g6440 and P2_U2553 P2_U2547 ; P2_U2559
g6441 and P2_U2553 P2_U2549 ; P2_U2560
g6442 and P2_U2547 P2_U2556 ; P2_U2561
g6443 and P2_U2549 P2_U2556 ; P2_U2562
g6444 and P2_U8100 P2_U3272 ; P2_U2563
g6445 and P2_U4409 P2_U3583 ; P2_U2564
g6446 and P2_U2564 P2_U2563 ; P2_U2565
g6447 and P2_U8100 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2566
g6448 and P2_U2564 P2_U2566 ; P2_U2567
g6449 and P2_U3582 P2_U3272 ; P2_U2568
g6450 and P2_U2564 P2_U2568 ; P2_U2569
g6451 and P2_U3582 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U2570
g6452 and P2_U2564 P2_U2570 ; P2_U2571
g6453 and P2_U3583 P2_U3553 ; P2_U2572
g6454 and P2_U2572 P2_U2563 ; P2_U2573
g6455 and P2_U2572 P2_U2566 ; P2_U2574
g6456 and P2_U2572 P2_U2568 ; P2_U2575
g6457 and P2_U2572 P2_U2570 ; P2_U2576
g6458 and P2_U4409 P2_U8149 ; P2_U2577
g6459 and P2_U2577 P2_U2563 ; P2_U2578
g6460 and P2_U2577 P2_U2566 ; P2_U2579
g6461 and P2_U2577 P2_U2568 ; P2_U2580
g6462 and P2_U2577 P2_U2570 ; P2_U2581
g6463 and P2_U8149 P2_U3553 ; P2_U2582
g6464 and P2_U2563 P2_U2582 ; P2_U2583
g6465 and P2_U2566 P2_U2582 ; P2_U2584
g6466 and P2_U2568 P2_U2582 ; P2_U2585
g6467 and P2_U2570 P2_U2582 ; P2_U2586
g6468 and P2_U2391 P2_EBX_REG_31__SCAN_IN ; P2_U2587
g6469 and P2_U2377 P2_U2360 ; P2_U2588
g6470 and P2_U7581 P2_U3550 P2_U4457 P2_U3549 ; P2_U2589
g6471 and P2_U5590 P2_U2436 ; P2_U2590
g6472 nand P2_U4274 P2_U4273 ; P2_U2591
g6473 nand P2_U4272 P2_U4271 ; P2_U2592
g6474 nand P2_U4270 P2_U4269 ; P2_U2593
g6475 nand P2_U4268 P2_U4267 ; P2_U2594
g6476 nand P2_U4266 P2_U4265 ; P2_U2595
g6477 nand P2_U4264 P2_U4263 ; P2_U2596
g6478 nand P2_U4262 P2_U4261 ; P2_U2597
g6479 nand P2_U4260 P2_U4259 ; P2_U2598
g6480 nand P2_U4258 P2_U4257 P2_U4256 P2_U4255 ; P2_U2599
g6481 nand P2_U4254 P2_U4253 P2_U4252 P2_U4251 ; P2_U2600
g6482 nand P2_U4250 P2_U4249 P2_U4248 P2_U4247 ; P2_U2601
g6483 nand P2_U4246 P2_U4245 P2_U4244 P2_U4243 ; P2_U2602
g6484 nand P2_U4242 P2_U4241 P2_U4240 P2_U4239 ; P2_U2603
g6485 nand P2_U4238 P2_U4237 P2_U4236 P2_U4235 ; P2_U2604
g6486 nand P2_U4234 P2_U4233 P2_U4232 P2_U4231 ; P2_U2605
g6487 nand P2_U4230 P2_U4229 P2_U4228 P2_U4227 ; P2_U2606
g6488 nand P2_U4226 P2_U4225 P2_U4224 P2_U4223 ; P2_U2607
g6489 nand P2_U4222 P2_U4221 P2_U4220 P2_U4219 ; P2_U2608
g6490 nand P2_U4218 P2_U4217 P2_U4216 P2_U4215 ; P2_U2609
g6491 nand P2_U4214 P2_U4213 P2_U4212 P2_U4211 ; P2_U2610
g6492 nand P2_U4210 P2_U4209 P2_U4208 P2_U4207 ; P2_U2611
g6493 nand P2_U4206 P2_U4205 P2_U4204 P2_U4203 ; P2_U2612
g6494 nand P2_U4202 P2_U4201 P2_U4200 P2_U4199 ; P2_U2613
g6495 nand P2_U4198 P2_U4197 P2_U4196 P2_U4195 ; P2_U2614
g6496 and P2_U3519 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U2615
g6497 nand P2_U3706 P2_U3705 ; P2_U2616
g6498 nand P2_U3694 P2_U3693 ; P2_U2617
g6499 nand P2_U4350 P2_U7453 ; P2_U2618
g6500 nand P2_U4351 P2_U7456 ; P2_U2619
g6501 nand P2_U4353 P2_U7462 ; P2_U2620
g6502 nand P2_U4354 P2_U7465 ; P2_U2621
g6503 nand P2_U4355 P2_U7468 ; P2_U2622
g6504 nand P2_U4356 P2_U7471 ; P2_U2623
g6505 nand P2_U4357 P2_U7474 ; P2_U2624
g6506 nand P2_U4358 P2_U7477 ; P2_U2625
g6507 nand P2_U4359 P2_U7480 ; P2_U2626
g6508 nand P2_U4360 P2_U7483 ; P2_U2627
g6509 nand P2_U4361 P2_U7486 ; P2_U2628
g6510 nand P2_U4362 P2_U7489 ; P2_U2629
g6511 nand P2_U4364 P2_U7495 ; P2_U2630
g6512 nand P2_U4365 P2_U7498 ; P2_U2631
g6513 nand P2_U4366 P2_U7501 ; P2_U2632
g6514 nand P2_U4367 P2_U7504 ; P2_U2633
g6515 nand P2_U7508 P2_U7507 P2_U4368 ; P2_U2634
g6516 nand P2_U7512 P2_U7511 P2_U4369 ; P2_U2635
g6517 nand P2_U7516 P2_U7515 P2_U4370 ; P2_U2636
g6518 nand P2_U7520 P2_U7519 P2_U4371 ; P2_U2637
g6519 nand P2_U7524 P2_U7523 P2_U4372 ; P2_U2638
g6520 nand P2_U7528 P2_U7527 P2_U4373 ; P2_U2639
g6521 nand P2_U7434 P2_U7433 P2_U4344 ; P2_U2640
g6522 nand P2_U7438 P2_U7437 P2_U4345 ; P2_U2641
g6523 nand P2_U4346 P2_U7441 ; P2_U2642
g6524 nand P2_U4347 P2_U7444 ; P2_U2643
g6525 nand P2_U4348 P2_U7447 ; P2_U2644
g6526 nand P2_U4349 P2_U7450 ; P2_U2645
g6527 nand P2_U4352 P2_U7459 ; P2_U2646
g6528 nand P2_U4363 P2_U7492 ; P2_U2647
g6529 nand P2_U4374 P2_U7531 ; P2_U2648
g6530 nand P2_U7534 P2_U3300 P2_U4375 ; P2_U2649
g6531 and P2_U2352 P2_U3242 ; P2_U2650
g6532 and P2_U2352 P2_U7217 ; P2_U2651
g6533 and P2_U2352 P2_U7251 ; P2_U2652
g6534 and P2_U2352 P2_U7285 ; P2_U2653
g6535 nand P2_U7423 P2_U7422 ; P2_U2654
g6536 nand P2_U4338 P2_U7424 ; P2_U2655
g6537 nand P2_U4340 P2_U7427 ; P2_U2656
g6538 nand P2_U4342 P2_U7429 ; P2_U2657
g6539 and P2_U2354 P2_U2598 ; P2_U2658
g6540 and P2_U2354 P2_U2597 ; P2_U2659
g6541 and P2_U2354 P2_U2596 ; P2_U2660
g6542 and P2_U2354 P2_U2595 ; P2_U2661
g6543 and P2_U2354 P2_U2594 ; P2_U2662
g6544 and P2_U2354 P2_U2593 ; P2_U2663
g6545 and P2_U2354 P2_U2592 ; P2_U2664
g6546 and P2_U2354 P2_U2591 ; P2_U2665
g6547 and P2_U2614 P2_U2355 ; P2_U2666
g6548 and P2_U2613 P2_U2355 ; P2_U2667
g6549 and P2_U2612 P2_U2355 ; P2_U2668
g6550 and P2_U2611 P2_U2355 ; P2_U2669
g6551 and P2_U2610 P2_U2355 ; P2_U2670
g6552 and P2_U2609 P2_U2355 ; P2_U2671
g6553 and P2_U2608 P2_U2355 ; P2_U2672
g6554 and P2_U2607 P2_U2355 ; P2_U2673
g6555 and P2_U2355 P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U2674
g6556 and P2_U2355 P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U2675
g6557 and P2_U2355 P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U2676
g6558 and P2_U2355 P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U2677
g6559 and P2_U2355 P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U2678
g6560 and P2_U2355 P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U2679
g6561 and P2_U2355 P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U2680
g6562 nand P2_U7166 P2_U4275 ; P2_U2681
g6563 and P2_U2355 P2_ADD_402_1132_U18 ; P2_U2682
g6564 and P2_ADD_402_1132_U19 P2_U2355 ; P2_U2683
g6565 and P2_ADD_402_1132_U24 P2_U2355 ; P2_U2684
g6566 and P2_ADD_402_1132_U22 P2_U2355 ; P2_U2685
g6567 and P2_ADD_402_1132_U21 P2_U2355 ; P2_U2686
g6568 and P2_ADD_402_1132_U25 P2_U2355 ; P2_U2687
g6569 and P2_ADD_402_1132_U20 P2_U2355 ; P2_U2688
g6570 nand P2_U7142 P2_U7141 ; P2_U2689
g6571 nand P2_U7144 P2_U7143 ; P2_U2690
g6572 nand P2_U7146 P2_U7145 ; P2_U2691
g6573 nand P2_U7148 P2_U7147 ; P2_U2692
g6574 nand P2_U7153 P2_U7152 ; P2_U2693
g6575 nand P2_U7155 P2_U7154 ; P2_U2694
g6576 nand P2_U7157 P2_U7156 ; P2_U2695
g6577 nand P2_U7159 P2_U7158 ; P2_U2696
g6578 and P2_U3554 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U2698
g6579 nand P2_U7139 P2_U7140 P2_U7138 ; P2_U2699
g6580 nand P2_U7150 P2_U7151 P2_U7149 ; P2_U2700
g6581 nand P2_U7161 P2_U7162 P2_U7160 ; P2_U2701
g6582 nand P2_U7164 P2_U7165 P2_U7163 ; P2_U2702
g6583 nand P2_U7727 P2_U7726 ; P2_U2703
g6584 nand P2_U7729 P2_U7728 ; P2_U2704
g6585 nand P2_U4390 P2_U7730 ; P2_U2705
g6586 nand P2_U7732 P2_U7733 P2_U3550 ; P2_U2706
g6587 nand P2_U4391 P2_U7734 ; P2_U2707
g6588 and P2_R2219_U25 P2_U7723 ; P2_U2708
g6589 and P2_R2219_U26 P2_U7723 ; P2_U2709
g6590 and P2_R2219_U27 P2_U7723 ; P2_U2710
g6591 nand P2_U7724 P2_STATE2_REG_0__SCAN_IN ; P2_U2711
g6592 nand P2_U7871 P2_U4407 P2_STATE2_REG_0__SCAN_IN ; P2_U2712
g6593 nand P2_U7725 P2_STATE2_REG_0__SCAN_IN ; P2_U2713
g6594 nand P2_U7871 P2_U4408 P2_STATE2_REG_0__SCAN_IN ; P2_U2714
g6595 nand P2_U2356 P2_U2616 ; P2_U2715
g6596 nand P2_U7620 P2_U7619 P2_U7618 P2_U7617 ; P2_U2716
g6597 nand P2_U7624 P2_U7623 P2_U7622 P2_U7621 ; P2_U2717
g6598 nand P2_U7632 P2_U7631 P2_U7630 P2_U7629 ; P2_U2718
g6599 nand P2_U7636 P2_U7635 P2_U7634 P2_U7633 ; P2_U2719
g6600 nand P2_U7640 P2_U7639 P2_U7638 P2_U7637 ; P2_U2720
g6601 nand P2_U7644 P2_U7643 P2_U7642 P2_U7641 ; P2_U2721
g6602 nand P2_U7648 P2_U7647 P2_U7646 P2_U7645 ; P2_U2722
g6603 nand P2_U7652 P2_U7651 P2_U7650 P2_U7649 ; P2_U2723
g6604 nand P2_U7656 P2_U7655 P2_U7654 P2_U7653 ; P2_U2724
g6605 nand P2_U7660 P2_U7659 P2_U7658 P2_U7657 ; P2_U2725
g6606 nand P2_U7664 P2_U7663 P2_U7662 P2_U7661 ; P2_U2726
g6607 nand P2_U7668 P2_U7667 P2_U7666 P2_U7665 ; P2_U2727
g6608 nand P2_U7676 P2_U7675 P2_U7674 P2_U7673 ; P2_U2728
g6609 nand P2_U7680 P2_U7679 P2_U7678 P2_U7677 ; P2_U2729
g6610 nand P2_U7684 P2_U7683 P2_U7682 P2_U7681 ; P2_U2730
g6611 nand P2_U7688 P2_U7687 P2_U7686 P2_U7685 ; P2_U2731
g6612 nand P2_U7692 P2_U7691 P2_U7690 P2_U7689 ; P2_U2732
g6613 nand P2_U7696 P2_U7695 P2_U7694 P2_U7693 ; P2_U2733
g6614 nand P2_U7700 P2_U7699 P2_U7698 P2_U7697 ; P2_U2734
g6615 nand P2_U7704 P2_U7703 P2_U7702 P2_U7701 ; P2_U2735
g6616 nand P2_U7708 P2_U7707 P2_U7706 P2_U7705 ; P2_U2736
g6617 nand P2_U7712 P2_U7711 P2_U7710 P2_U7709 ; P2_U2737
g6618 nand P2_U7596 P2_U7595 P2_U7594 P2_U7593 ; P2_U2738
g6619 nand P2_U7600 P2_U7599 P2_U7598 P2_U7597 ; P2_U2739
g6620 nand P2_U7604 P2_U7603 P2_U7602 P2_U7601 ; P2_U2740
g6621 nand P2_U7608 P2_U7607 P2_U7606 P2_U7605 ; P2_U2741
g6622 nand P2_U7612 P2_U7611 P2_U7610 P2_U7609 ; P2_U2742
g6623 nand P2_U7616 P2_U7615 P2_U7614 P2_U7613 ; P2_U2743
g6624 nand P2_U7628 P2_U7627 P2_U7626 P2_U7625 ; P2_U2744
g6625 nand P2_U7672 P2_U7671 P2_U7670 P2_U7669 ; P2_U2745
g6626 nand P2_U7716 P2_U7715 P2_U7714 P2_U7713 ; P2_U2746
g6627 nand P2_U7886 P2_U7721 P2_U4389 P2_U4388 P2_U7717 ; P2_U2747
g6628 nand P2_U7583 P2_U7582 ; P2_U2748
g6629 nand P2_U4380 P2_U7584 ; P2_U2749
g6630 nand P2_U4382 P2_U7588 ; P2_U2750
g6631 and P2_U7888 P2_U7737 ; P2_U2751
g6632 and P2_U3280 P2_U7873 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U2752
g6633 nand P2_U3286 P2_U7572 ; P2_U2753
g6634 nand P2_U3286 P2_U7573 ; P2_U2754
g6635 nand P2_U3286 P2_U7574 ; P2_U2755
g6636 nand P2_U3286 P2_U7575 ; P2_U2756
g6637 nand P2_U3286 P2_U7576 ; P2_U2757
g6638 and P2_U4428 P2_U3242 ; P2_U2758
g6639 and P2_U4428 P2_U7217 ; P2_U2759
g6640 and P2_U4428 P2_U7251 ; P2_U2760
g6641 nand P2_U7563 P2_U7562 ; P2_U2761
g6642 nand P2_U7565 P2_U7564 ; P2_U2762
g6643 nand P2_U7567 P2_U7566 ; P2_U2763
g6644 nand P2_U7569 P2_U7568 ; P2_U2764
g6645 nand P2_U7571 P2_U7570 ; P2_U2765
g6646 nand P2_U4447 P2_U7539 ; P2_U2766
g6647 nand P2_U4447 P2_U7540 ; P2_U2767
g6648 nand P2_U4447 P2_U7541 ; P2_U2768
g6649 nand P2_U4447 P2_U7542 ; P2_U2769
g6650 nand P2_U4447 P2_U7543 ; P2_U2770
g6651 nand P2_U4447 P2_U7544 ; P2_U2771
g6652 nand P2_U4447 P2_U7545 ; P2_U2772
g6653 nand P2_U4447 P2_U7546 ; P2_U2773
g6654 nand P2_U4447 P2_U7547 ; P2_U2774
g6655 nand P2_U4447 P2_U7548 ; P2_U2775
g6656 nand P2_U4447 P2_U7549 ; P2_U2776
g6657 nand P2_U4447 P2_U7550 ; P2_U2777
g6658 nand P2_U4447 P2_U7551 ; P2_U2778
g6659 nand P2_U4447 P2_U7552 ; P2_U2779
g6660 nand P2_U4447 P2_U7553 ; P2_U2780
g6661 nand P2_U4447 P2_U7554 ; P2_U2781
g6662 nand P2_U4447 P2_U7555 ; P2_U2782
g6663 nand P2_U4447 P2_U7556 ; P2_U2783
g6664 nand P2_U4447 P2_U7557 ; P2_U2784
g6665 nand P2_U4447 P2_U7558 ; P2_U2785
g6666 nand P2_U4447 P2_U7559 ; P2_U2786
g6667 nand P2_U4447 P2_U7560 ; P2_U2787
g6668 nand P2_U4447 P2_U7537 ; P2_U2788
g6669 nand P2_U4447 P2_U7538 ; P2_U2789
g6670 and P2_U3242 P2_R2267_U63 ; P2_U2790
g6671 and P2_U3242 P2_R2267_U16 ; P2_U2791
g6672 and P2_U3242 P2_R2267_U15 ; P2_U2792
g6673 and P2_U3242 P2_R2267_U67 ; P2_U2793
g6674 and P2_U3242 P2_R2267_U14 ; P2_U2794
g6675 and P2_U3242 P2_R2267_U69 ; P2_U2795
g6676 and P2_U3242 P2_R2267_U13 ; P2_U2796
g6677 and P2_U3242 P2_R2267_U71 ; P2_U2797
g6678 and P2_U3242 P2_R2267_U12 ; P2_U2798
g6679 and P2_U3242 P2_R2267_U73 ; P2_U2799
g6680 and P2_U3242 P2_R2267_U11 ; P2_U2800
g6681 and P2_U3242 P2_R2267_U75 ; P2_U2801
g6682 and P2_U3242 P2_R2267_U10 ; P2_U2802
g6683 and P2_U3242 P2_R2267_U79 ; P2_U2803
g6684 and P2_U3242 P2_R2267_U9 ; P2_U2804
g6685 and P2_U3242 P2_R2267_U81 ; P2_U2805
g6686 and P2_U3242 P2_R2267_U8 ; P2_U2806
g6687 and P2_U3242 P2_R2267_U83 ; P2_U2807
g6688 and P2_U3242 P2_R2267_U7 ; P2_U2808
g6689 and P2_U3242 P2_R2267_U85 ; P2_U2809
g6690 and P2_U3242 P2_R2267_U6 ; P2_U2810
g6691 and P2_U3242 P2_R2267_U87 ; P2_U2811
g6692 and P2_U3242 P2_R2267_U20 ; P2_U2812
g6693 and P2_U3519 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U2813
g6694 nand P2_U4190 P2_U6861 ; P2_U2814
g6695 nand P2_U7917 P2_U6856 ; P2_U2815
g6696 nand P2_U6855 P2_U6854 ; P2_U2816
g6697 nand P2_U8140 P2_U8139 P2_U4463 ; P2_U2817
g6698 nand P2_U8136 P2_U8135 P2_U4463 ; P2_U2818
g6699 nand P2_U6840 P2_U6839 ; P2_U2819
g6700 nand P2_U8128 P2_U8127 P2_U3548 ; P2_U2820
g6701 nand P2_U3548 P2_U4452 P2_U6837 ; P2_U2821
g6702 nand P2_U4398 P2_U6836 ; P2_U2822
g6703 nand P2_U8124 P2_U8123 P2_U4452 ; P2_U2823
g6704 nand P2_U6827 P2_U6829 P2_U4168 P2_U6830 P2_U6828 ; P2_U2824
g6705 nand P2_U6819 P2_U6821 P2_U4166 P2_U6822 P2_U6820 ; P2_U2825
g6706 nand P2_U6811 P2_U6813 P2_U4164 P2_U6814 P2_U6812 ; P2_U2826
g6707 nand P2_U6803 P2_U6805 P2_U4162 P2_U6806 P2_U6804 ; P2_U2827
g6708 nand P2_U6795 P2_U6797 P2_U4160 P2_U6798 P2_U6796 ; P2_U2828
g6709 nand P2_U6787 P2_U6789 P2_U4158 P2_U6790 P2_U6788 ; P2_U2829
g6710 nand P2_U6779 P2_U6781 P2_U6782 P2_U4156 P2_U6780 ; P2_U2830
g6711 nand P2_U6772 P2_U4152 ; P2_U2831
g6712 nand P2_U6764 P2_U4149 ; P2_U2832
g6713 nand P2_U6755 P2_U6757 P2_U6758 P2_U6756 P2_U4148 ; P2_U2833
g6714 nand P2_U4146 P2_U4144 ; P2_U2834
g6715 nand P2_U4143 P2_U4141 ; P2_U2835
g6716 nand P2_U4140 P2_U4138 ; P2_U2836
g6717 nand P2_U4136 P2_U4134 ; P2_U2837
g6718 nand P2_U4132 P2_U4130 ; P2_U2838
g6719 nand P2_U4128 P2_U4126 ; P2_U2839
g6720 nand P2_U4124 P2_U4122 ; P2_U2840
g6721 nand P2_U6693 P2_U4118 P2_U6692 P2_U6696 P2_U4119 ; P2_U2841
g6722 nand P2_U6685 P2_U4115 P2_U6684 P2_U6688 P2_U4116 ; P2_U2842
g6723 nand P2_U6677 P2_U4112 P2_U6676 P2_U6680 P2_U4113 ; P2_U2843
g6724 nand P2_U6670 P2_U6669 P2_U4109 P2_U6672 P2_U4110 ; P2_U2844
g6725 nand P2_U6662 P2_U6661 P2_U4106 P2_U6664 P2_U4107 ; P2_U2845
g6726 nand P2_U6654 P2_U6653 P2_U4103 P2_U6656 P2_U4104 ; P2_U2846
g6727 nand P2_U6646 P2_U6645 P2_U4100 P2_U6648 P2_U4101 ; P2_U2847
g6728 nand P2_U6638 P2_U6637 P2_U4097 P2_U6640 P2_U4098 ; P2_U2848
g6729 nand P2_U6630 P2_U6629 P2_U4094 P2_U6632 P2_U4095 ; P2_U2849
g6730 nand P2_U4093 P2_U4091 ; P2_U2850
g6731 nand P2_U4089 P2_U4087 ; P2_U2851
g6732 nand P2_U6602 P2_U4082 P2_U6606 P2_U4084 ; P2_U2852
g6733 nand P2_U6593 P2_U4078 P2_U6597 P2_U4080 ; P2_U2853
g6734 nand P2_U6584 P2_U4074 P2_U6588 P2_U4076 ; P2_U2854
g6735 nand P2_U6575 P2_U4070 P2_U6579 P2_U4072 ; P2_U2855
g6736 nand P2_U6565 P2_U6564 ; P2_U2856
g6737 nand P2_U6562 P2_U6563 P2_U6561 ; P2_U2857
g6738 nand P2_U6559 P2_U6560 P2_U6558 ; P2_U2858
g6739 nand P2_U6556 P2_U6557 P2_U6555 ; P2_U2859
g6740 nand P2_U6553 P2_U6554 P2_U6552 ; P2_U2860
g6741 nand P2_U6550 P2_U6551 P2_U6549 ; P2_U2861
g6742 nand P2_U6547 P2_U6548 P2_U6546 ; P2_U2862
g6743 nand P2_U6544 P2_U6545 P2_U6543 ; P2_U2863
g6744 nand P2_U6541 P2_U6542 P2_U6540 ; P2_U2864
g6745 nand P2_U6538 P2_U6539 P2_U6537 ; P2_U2865
g6746 nand P2_U6535 P2_U6536 P2_U6534 ; P2_U2866
g6747 nand P2_U6532 P2_U6533 P2_U6531 ; P2_U2867
g6748 nand P2_U6529 P2_U6530 P2_U6528 ; P2_U2868
g6749 nand P2_U6526 P2_U6527 P2_U6525 ; P2_U2869
g6750 nand P2_U6523 P2_U6524 P2_U6522 ; P2_U2870
g6751 nand P2_U6520 P2_U6521 P2_U6519 ; P2_U2871
g6752 nand P2_U6517 P2_U6518 P2_U6516 ; P2_U2872
g6753 nand P2_U6514 P2_U6515 P2_U6513 ; P2_U2873
g6754 nand P2_U6511 P2_U6512 P2_U6510 ; P2_U2874
g6755 nand P2_U6508 P2_U6509 P2_U6507 ; P2_U2875
g6756 nand P2_U6505 P2_U6506 P2_U6504 ; P2_U2876
g6757 nand P2_U6502 P2_U6503 P2_U6501 ; P2_U2877
g6758 nand P2_U6499 P2_U6500 P2_U6498 ; P2_U2878
g6759 nand P2_U6496 P2_U6497 P2_U6495 ; P2_U2879
g6760 nand P2_U6493 P2_U6492 P2_U6494 ; P2_U2880
g6761 nand P2_U6490 P2_U6489 P2_U6491 ; P2_U2881
g6762 nand P2_U6487 P2_U6486 P2_U6488 ; P2_U2882
g6763 nand P2_U6484 P2_U6483 P2_U6485 ; P2_U2883
g6764 nand P2_U6481 P2_U6480 P2_U6482 ; P2_U2884
g6765 nand P2_U6478 P2_U6477 P2_U6479 ; P2_U2885
g6766 nand P2_U6475 P2_U6474 P2_U6476 ; P2_U2886
g6767 nand P2_U6472 P2_U6471 P2_U6473 ; P2_U2887
g6768 nand P2_U6468 P2_U6466 P2_U6467 ; P2_U2888
g6769 nand P2_U6462 P2_U6461 P2_U6465 P2_U6464 P2_U6463 ; P2_U2889
g6770 nand P2_U6457 P2_U6456 P2_U6460 P2_U6459 P2_U6458 ; P2_U2890
g6771 nand P2_U6452 P2_U6451 P2_U6455 P2_U6454 P2_U6453 ; P2_U2891
g6772 nand P2_U6447 P2_U6446 P2_U6450 P2_U6449 P2_U6448 ; P2_U2892
g6773 nand P2_U6442 P2_U6441 P2_U6445 P2_U6444 P2_U6443 ; P2_U2893
g6774 nand P2_U6437 P2_U6436 P2_U6440 P2_U6439 P2_U6438 ; P2_U2894
g6775 nand P2_U6432 P2_U6431 P2_U6435 P2_U6434 P2_U6433 ; P2_U2895
g6776 nand P2_U6427 P2_U6426 P2_U6430 P2_U6429 P2_U6428 ; P2_U2896
g6777 nand P2_U6422 P2_U6421 P2_U6425 P2_U6424 P2_U6423 ; P2_U2897
g6778 nand P2_U6417 P2_U6416 P2_U6420 P2_U6419 P2_U6418 ; P2_U2898
g6779 nand P2_U6412 P2_U6411 P2_U6415 P2_U6414 P2_U6413 ; P2_U2899
g6780 nand P2_U6407 P2_U6406 P2_U6410 P2_U6409 P2_U6408 ; P2_U2900
g6781 nand P2_U6402 P2_U6401 P2_U6405 P2_U6404 P2_U6403 ; P2_U2901
g6782 nand P2_U6397 P2_U6396 P2_U6400 P2_U6399 P2_U6398 ; P2_U2902
g6783 nand P2_U6392 P2_U6391 P2_U6395 P2_U6394 P2_U6393 ; P2_U2903
g6784 nand P2_U6390 P2_U6387 P2_U6389 P2_U6388 ; P2_U2904
g6785 nand P2_U6386 P2_U6383 P2_U6385 P2_U6384 ; P2_U2905
g6786 nand P2_U6382 P2_U6379 P2_U6381 P2_U6380 ; P2_U2906
g6787 nand P2_U6378 P2_U6375 P2_U6377 P2_U6376 ; P2_U2907
g6788 nand P2_U6374 P2_U6371 P2_U6373 P2_U6372 ; P2_U2908
g6789 nand P2_U6370 P2_U6367 P2_U6369 P2_U6368 ; P2_U2909
g6790 nand P2_U4068 P2_U6363 P2_U6364 ; P2_U2910
g6791 nand P2_U4067 P2_U6359 P2_U6360 ; P2_U2911
g6792 nand P2_U4066 P2_U6355 P2_U6356 ; P2_U2912
g6793 nand P2_U6352 P2_U6351 P2_U4065 ; P2_U2913
g6794 nand P2_U6348 P2_U6347 P2_U4064 ; P2_U2914
g6795 nand P2_U6344 P2_U6343 P2_U4063 ; P2_U2915
g6796 nand P2_U6340 P2_U6339 P2_U4062 ; P2_U2916
g6797 nand P2_U6336 P2_U6335 P2_U4061 ; P2_U2917
g6798 nand P2_U6332 P2_U6331 P2_U4060 ; P2_U2918
g6799 nand P2_U6328 P2_U6327 P2_U4059 ; P2_U2919
g6800 and P2_U6232 P2_DATAO_REG_31__SCAN_IN ; P2_U2920
g6801 nand P2_U6324 P2_U6323 P2_U6325 ; P2_U2921
g6802 nand P2_U6321 P2_U6320 P2_U6322 ; P2_U2922
g6803 nand P2_U6318 P2_U6317 P2_U6319 ; P2_U2923
g6804 nand P2_U6315 P2_U6314 P2_U6316 ; P2_U2924
g6805 nand P2_U6312 P2_U6311 P2_U6313 ; P2_U2925
g6806 nand P2_U6309 P2_U6308 P2_U6310 ; P2_U2926
g6807 nand P2_U6306 P2_U6305 P2_U6307 ; P2_U2927
g6808 nand P2_U6303 P2_U6302 P2_U6304 ; P2_U2928
g6809 nand P2_U6300 P2_U6299 P2_U6301 ; P2_U2929
g6810 nand P2_U6297 P2_U6296 P2_U6298 ; P2_U2930
g6811 nand P2_U6294 P2_U6293 P2_U6295 ; P2_U2931
g6812 nand P2_U6291 P2_U6290 P2_U6292 ; P2_U2932
g6813 nand P2_U6288 P2_U6287 P2_U6289 ; P2_U2933
g6814 nand P2_U6285 P2_U6284 P2_U6286 ; P2_U2934
g6815 nand P2_U6282 P2_U6281 P2_U6283 ; P2_U2935
g6816 nand P2_U6279 P2_U6278 P2_U6280 ; P2_U2936
g6817 nand P2_U6276 P2_U6275 P2_U6277 ; P2_U2937
g6818 nand P2_U6273 P2_U6272 P2_U6274 ; P2_U2938
g6819 nand P2_U6270 P2_U6269 P2_U6271 ; P2_U2939
g6820 nand P2_U6267 P2_U6266 P2_U6268 ; P2_U2940
g6821 nand P2_U6264 P2_U6263 P2_U6265 ; P2_U2941
g6822 nand P2_U6261 P2_U6260 P2_U6262 ; P2_U2942
g6823 nand P2_U6258 P2_U6257 P2_U6259 ; P2_U2943
g6824 nand P2_U6255 P2_U6254 P2_U6256 ; P2_U2944
g6825 nand P2_U6252 P2_U6251 P2_U6253 ; P2_U2945
g6826 nand P2_U6249 P2_U6248 P2_U6250 ; P2_U2946
g6827 nand P2_U6246 P2_U6245 P2_U6247 ; P2_U2947
g6828 nand P2_U6243 P2_U6242 P2_U6244 ; P2_U2948
g6829 nand P2_U6240 P2_U6239 P2_U6241 ; P2_U2949
g6830 nand P2_U6237 P2_U6236 P2_U6238 ; P2_U2950
g6831 nand P2_U6234 P2_U6233 P2_U6235 ; P2_U2951
g6832 nand P2_U6225 P2_U6224 P2_U6226 ; P2_U2952
g6833 nand P2_U6222 P2_U6221 P2_U6223 ; P2_U2953
g6834 nand P2_U6219 P2_U6218 P2_U6220 ; P2_U2954
g6835 nand P2_U6216 P2_U6215 P2_U6217 ; P2_U2955
g6836 nand P2_U6213 P2_U6212 P2_U6214 ; P2_U2956
g6837 nand P2_U6210 P2_U6209 P2_U6211 ; P2_U2957
g6838 nand P2_U6207 P2_U6206 P2_U6208 ; P2_U2958
g6839 nand P2_U6204 P2_U6203 P2_U6205 ; P2_U2959
g6840 nand P2_U6201 P2_U6200 P2_U6202 ; P2_U2960
g6841 nand P2_U6198 P2_U6197 P2_U6199 ; P2_U2961
g6842 nand P2_U6195 P2_U6194 P2_U6196 ; P2_U2962
g6843 nand P2_U6192 P2_U6191 P2_U6193 ; P2_U2963
g6844 nand P2_U6189 P2_U6188 P2_U6190 ; P2_U2964
g6845 nand P2_U6186 P2_U6185 P2_U6187 ; P2_U2965
g6846 nand P2_U6183 P2_U6182 P2_U6184 ; P2_U2966
g6847 nand P2_U6180 P2_U6179 P2_U6181 ; P2_U2967
g6848 nand P2_U6177 P2_U6176 P2_U6178 ; P2_U2968
g6849 nand P2_U6174 P2_U6173 P2_U6175 ; P2_U2969
g6850 nand P2_U6171 P2_U6170 P2_U6172 ; P2_U2970
g6851 nand P2_U6168 P2_U6167 P2_U6169 ; P2_U2971
g6852 nand P2_U6165 P2_U6164 P2_U6166 ; P2_U2972
g6853 nand P2_U6162 P2_U6161 P2_U6163 ; P2_U2973
g6854 nand P2_U6159 P2_U6158 P2_U6160 ; P2_U2974
g6855 nand P2_U6156 P2_U6155 P2_U6157 ; P2_U2975
g6856 nand P2_U6153 P2_U6152 P2_U6154 ; P2_U2976
g6857 nand P2_U6150 P2_U6149 P2_U6151 ; P2_U2977
g6858 nand P2_U6147 P2_U6146 P2_U6148 ; P2_U2978
g6859 nand P2_U6144 P2_U6143 P2_U6145 ; P2_U2979
g6860 nand P2_U6141 P2_U6140 P2_U6142 ; P2_U2980
g6861 nand P2_U6138 P2_U6137 P2_U6139 ; P2_U2981
g6862 nand P2_U6135 P2_U6134 P2_U6136 ; P2_U2982
g6863 nand P2_U4054 P2_U4053 ; P2_U2983
g6864 nand P2_U4052 P2_U4051 ; P2_U2984
g6865 nand P2_U4050 P2_U4049 ; P2_U2985
g6866 nand P2_U4048 P2_U4047 ; P2_U2986
g6867 nand P2_U4046 P2_U4045 ; P2_U2987
g6868 nand P2_U4044 P2_U4043 ; P2_U2988
g6869 nand P2_U4042 P2_U4041 ; P2_U2989
g6870 nand P2_U4040 P2_U4039 ; P2_U2990
g6871 nand P2_U4038 P2_U4037 ; P2_U2991
g6872 nand P2_U4036 P2_U4035 ; P2_U2992
g6873 nand P2_U4034 P2_U4033 ; P2_U2993
g6874 nand P2_U4032 P2_U4031 ; P2_U2994
g6875 nand P2_U4030 P2_U4029 ; P2_U2995
g6876 nand P2_U4028 P2_U4027 ; P2_U2996
g6877 nand P2_U4026 P2_U4025 ; P2_U2997
g6878 nand P2_U4024 P2_U4023 ; P2_U2998
g6879 nand P2_U4022 P2_U4021 ; P2_U2999
g6880 nand P2_U4020 P2_U4019 ; P2_U3000
g6881 nand P2_U4018 P2_U4017 ; P2_U3001
g6882 nand P2_U4016 P2_U4015 ; P2_U3002
g6883 nand P2_U4014 P2_U4013 ; P2_U3003
g6884 nand P2_U4012 P2_U4011 ; P2_U3004
g6885 nand P2_U4010 P2_U4009 ; P2_U3005
g6886 nand P2_U4008 P2_U4007 ; P2_U3006
g6887 nand P2_U4006 P2_U4005 ; P2_U3007
g6888 nand P2_U4004 P2_U4003 ; P2_U3008
g6889 nand P2_U4002 P2_U4001 ; P2_U3009
g6890 nand P2_U4000 P2_U3999 ; P2_U3010
g6891 nand P2_U3998 P2_U3997 ; P2_U3011
g6892 nand P2_U3996 P2_U3995 ; P2_U3012
g6893 nand P2_U3994 P2_U3993 ; P2_U3013
g6894 nand P2_U3992 P2_U3991 ; P2_U3014
g6895 nand P2_U5933 P2_U5932 P2_U3988 P2_U3987 P2_U5928 ; P2_U3015
g6896 nand P2_U5925 P2_U5924 P2_U3986 P2_U3985 P2_U5920 ; P2_U3016
g6897 nand P2_U5917 P2_U5916 P2_U3984 P2_U3983 ; P2_U3017
g6898 nand P2_U5909 P2_U5908 P2_U3982 P2_U3981 P2_U3980 ; P2_U3018
g6899 nand P2_U5901 P2_U5900 P2_U3979 P2_U3978 P2_U3977 ; P2_U3019
g6900 nand P2_U5893 P2_U5892 P2_U3976 P2_U3975 P2_U3974 ; P2_U3020
g6901 nand P2_U5885 P2_U5884 P2_U3973 P2_U3972 P2_U3971 ; P2_U3021
g6902 nand P2_U5877 P2_U5876 P2_U3970 P2_U3969 P2_U3968 ; P2_U3022
g6903 nand P2_U5869 P2_U5868 P2_U3967 P2_U3966 P2_U3965 ; P2_U3023
g6904 nand P2_U5861 P2_U5860 P2_U3964 P2_U3963 P2_U3962 ; P2_U3024
g6905 nand P2_U5853 P2_U5852 P2_U3961 P2_U3960 P2_U3959 ; P2_U3025
g6906 nand P2_U5845 P2_U5844 P2_U3958 P2_U3957 P2_U3956 ; P2_U3026
g6907 nand P2_U5837 P2_U5836 P2_U3955 P2_U3954 P2_U3953 ; P2_U3027
g6908 nand P2_U5829 P2_U5828 P2_U3952 P2_U3951 P2_U3950 ; P2_U3028
g6909 nand P2_U5821 P2_U5820 P2_U3949 P2_U3948 P2_U3947 ; P2_U3029
g6910 nand P2_U5813 P2_U5812 P2_U3946 P2_U3945 P2_U3944 ; P2_U3030
g6911 nand P2_U5805 P2_U5804 P2_U3943 P2_U3942 P2_U3941 ; P2_U3031
g6912 nand P2_U5797 P2_U5796 P2_U3940 P2_U3939 P2_U3938 ; P2_U3032
g6913 nand P2_U5789 P2_U5788 P2_U3937 P2_U3936 P2_U3935 ; P2_U3033
g6914 nand P2_U5781 P2_U5780 P2_U3934 P2_U3933 P2_U3932 ; P2_U3034
g6915 nand P2_U5773 P2_U5772 P2_U3931 P2_U3930 P2_U3929 ; P2_U3035
g6916 nand P2_U5765 P2_U5764 P2_U3928 P2_U3927 P2_U3926 ; P2_U3036
g6917 nand P2_U5757 P2_U5756 P2_U3925 P2_U3924 P2_U3923 ; P2_U3037
g6918 nand P2_U5749 P2_U5748 P2_U3922 P2_U3921 P2_U3920 ; P2_U3038
g6919 nand P2_U5741 P2_U5740 P2_U3919 P2_U3918 P2_U3917 ; P2_U3039
g6920 nand P2_U5733 P2_U5732 P2_U3916 P2_U3915 P2_U3914 ; P2_U3040
g6921 nand P2_U5725 P2_U5724 P2_U3913 P2_U3912 P2_U3911 ; P2_U3041
g6922 nand P2_U5717 P2_U5716 P2_U3910 P2_U3909 P2_U3908 ; P2_U3042
g6923 nand P2_U5709 P2_U5708 P2_U3907 P2_U3906 P2_U3905 ; P2_U3043
g6924 nand P2_U5701 P2_U5700 P2_U3904 P2_U3903 P2_U3902 ; P2_U3044
g6925 nand P2_U5693 P2_U5692 P2_U3901 P2_U3900 P2_U3899 ; P2_U3045
g6926 nand P2_U5685 P2_U5684 P2_U3898 P2_U3897 P2_U3896 ; P2_U3046
g6927 and P2_U5643 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_U3047
g6928 nand P2_U5570 P2_U5569 P2_U3865 ; P2_U3048
g6929 nand P2_U5565 P2_U5564 P2_U3864 ; P2_U3049
g6930 nand P2_U5560 P2_U5559 P2_U3863 ; P2_U3050
g6931 nand P2_U5555 P2_U5554 P2_U3862 ; P2_U3051
g6932 nand P2_U5550 P2_U5549 P2_U3861 ; P2_U3052
g6933 nand P2_U5545 P2_U5544 P2_U3860 ; P2_U3053
g6934 nand P2_U5540 P2_U5539 P2_U3859 ; P2_U3054
g6935 nand P2_U5535 P2_U5534 P2_U3858 ; P2_U3055
g6936 nand P2_U5513 P2_U5512 P2_U3856 ; P2_U3056
g6937 nand P2_U5508 P2_U5507 P2_U3855 ; P2_U3057
g6938 nand P2_U5503 P2_U5502 P2_U3854 ; P2_U3058
g6939 nand P2_U5498 P2_U5497 P2_U3853 ; P2_U3059
g6940 nand P2_U5493 P2_U5492 P2_U3852 ; P2_U3060
g6941 nand P2_U5488 P2_U5487 P2_U3851 ; P2_U3061
g6942 nand P2_U5483 P2_U5482 P2_U3850 ; P2_U3062
g6943 nand P2_U5478 P2_U5477 P2_U3849 ; P2_U3063
g6944 nand P2_U5455 P2_U5454 P2_U3847 ; P2_U3064
g6945 nand P2_U5450 P2_U5449 P2_U3846 ; P2_U3065
g6946 nand P2_U5445 P2_U5444 P2_U3845 ; P2_U3066
g6947 nand P2_U5440 P2_U5439 P2_U3844 ; P2_U3067
g6948 nand P2_U5435 P2_U5434 P2_U3843 ; P2_U3068
g6949 nand P2_U5430 P2_U5429 P2_U3842 ; P2_U3069
g6950 nand P2_U5425 P2_U5424 P2_U3841 ; P2_U3070
g6951 nand P2_U5420 P2_U5419 P2_U3840 ; P2_U3071
g6952 nand P2_U5398 P2_U5397 P2_U3838 ; P2_U3072
g6953 nand P2_U5393 P2_U5392 P2_U3837 ; P2_U3073
g6954 nand P2_U5388 P2_U5387 P2_U3836 ; P2_U3074
g6955 nand P2_U5383 P2_U5382 P2_U3835 ; P2_U3075
g6956 nand P2_U5378 P2_U5377 P2_U3834 ; P2_U3076
g6957 nand P2_U5373 P2_U5372 P2_U3833 ; P2_U3077
g6958 nand P2_U5368 P2_U5367 P2_U3832 ; P2_U3078
g6959 nand P2_U5363 P2_U5362 P2_U3831 ; P2_U3079
g6960 nand P2_U5340 P2_U5339 P2_U3829 ; P2_U3080
g6961 nand P2_U5335 P2_U5334 P2_U3828 ; P2_U3081
g6962 nand P2_U5330 P2_U5329 P2_U3827 ; P2_U3082
g6963 nand P2_U5325 P2_U5324 P2_U3826 ; P2_U3083
g6964 nand P2_U5320 P2_U5319 P2_U3825 ; P2_U3084
g6965 nand P2_U5315 P2_U5314 P2_U3824 ; P2_U3085
g6966 nand P2_U5310 P2_U5309 P2_U3823 ; P2_U3086
g6967 nand P2_U5305 P2_U5304 P2_U3822 ; P2_U3087
g6968 nand P2_U5283 P2_U5282 P2_U3820 ; P2_U3088
g6969 nand P2_U5278 P2_U5277 P2_U3819 ; P2_U3089
g6970 nand P2_U5273 P2_U5272 P2_U3818 ; P2_U3090
g6971 nand P2_U5268 P2_U5267 P2_U3817 ; P2_U3091
g6972 nand P2_U5263 P2_U5262 P2_U3816 ; P2_U3092
g6973 nand P2_U5258 P2_U5257 P2_U3815 ; P2_U3093
g6974 nand P2_U5253 P2_U5252 P2_U3814 ; P2_U3094
g6975 nand P2_U5248 P2_U5247 P2_U3813 ; P2_U3095
g6976 nand P2_U5225 P2_U5224 P2_U3811 ; P2_U3096
g6977 nand P2_U5220 P2_U5219 P2_U3810 ; P2_U3097
g6978 nand P2_U5215 P2_U5214 P2_U3809 ; P2_U3098
g6979 nand P2_U5210 P2_U5209 P2_U3808 ; P2_U3099
g6980 nand P2_U5205 P2_U5204 P2_U3807 ; P2_U3100
g6981 nand P2_U5200 P2_U5199 P2_U3806 ; P2_U3101
g6982 nand P2_U5195 P2_U5194 P2_U3805 ; P2_U3102
g6983 nand P2_U5190 P2_U5189 P2_U3804 ; P2_U3103
g6984 nand P2_U5168 P2_U5167 P2_U3802 ; P2_U3104
g6985 nand P2_U5163 P2_U5162 P2_U3801 ; P2_U3105
g6986 nand P2_U5158 P2_U5157 P2_U3800 ; P2_U3106
g6987 nand P2_U5153 P2_U5152 P2_U3799 ; P2_U3107
g6988 nand P2_U5148 P2_U5147 P2_U3798 ; P2_U3108
g6989 nand P2_U5143 P2_U5142 P2_U3797 ; P2_U3109
g6990 nand P2_U5138 P2_U5137 P2_U3796 ; P2_U3110
g6991 nand P2_U5133 P2_U5132 P2_U3795 ; P2_U3111
g6992 nand P2_U5112 P2_U5111 P2_U3793 ; P2_U3112
g6993 nand P2_U5107 P2_U5106 P2_U3792 ; P2_U3113
g6994 nand P2_U5102 P2_U5101 P2_U3791 ; P2_U3114
g6995 nand P2_U5097 P2_U5096 P2_U3790 ; P2_U3115
g6996 nand P2_U5092 P2_U5091 P2_U3789 ; P2_U3116
g6997 nand P2_U5087 P2_U5086 P2_U3788 ; P2_U3117
g6998 nand P2_U5082 P2_U5081 P2_U3787 ; P2_U3118
g6999 nand P2_U5077 P2_U5076 P2_U3786 ; P2_U3119
g7000 nand P2_U5055 P2_U5054 P2_U3784 ; P2_U3120
g7001 nand P2_U5050 P2_U5049 P2_U3783 ; P2_U3121
g7002 nand P2_U5045 P2_U5044 P2_U3782 ; P2_U3122
g7003 nand P2_U5040 P2_U5039 P2_U3781 ; P2_U3123
g7004 nand P2_U5035 P2_U5034 P2_U3780 ; P2_U3124
g7005 nand P2_U5030 P2_U5029 P2_U3779 ; P2_U3125
g7006 nand P2_U5025 P2_U5024 P2_U3778 ; P2_U3126
g7007 nand P2_U5020 P2_U5019 P2_U3777 ; P2_U3127
g7008 nand P2_U4997 P2_U4996 P2_U3775 ; P2_U3128
g7009 nand P2_U4992 P2_U4991 P2_U3774 ; P2_U3129
g7010 nand P2_U4987 P2_U4986 P2_U3773 ; P2_U3130
g7011 nand P2_U4982 P2_U4981 P2_U3772 ; P2_U3131
g7012 nand P2_U4977 P2_U4976 P2_U3771 ; P2_U3132
g7013 nand P2_U4972 P2_U4971 P2_U3770 ; P2_U3133
g7014 nand P2_U4967 P2_U4966 P2_U3769 ; P2_U3134
g7015 nand P2_U4962 P2_U4961 P2_U3768 ; P2_U3135
g7016 nand P2_U4940 P2_U4939 P2_U3766 ; P2_U3136
g7017 nand P2_U4935 P2_U4934 P2_U3765 ; P2_U3137
g7018 nand P2_U4930 P2_U4929 P2_U3764 ; P2_U3138
g7019 nand P2_U4925 P2_U4924 P2_U3763 ; P2_U3139
g7020 nand P2_U4920 P2_U4919 P2_U3762 ; P2_U3140
g7021 nand P2_U4915 P2_U4914 P2_U3761 ; P2_U3141
g7022 nand P2_U4910 P2_U4909 P2_U3760 ; P2_U3142
g7023 nand P2_U4905 P2_U4904 P2_U3759 ; P2_U3143
g7024 nand P2_U4882 P2_U4881 P2_U3757 ; P2_U3144
g7025 nand P2_U4877 P2_U4876 P2_U3756 ; P2_U3145
g7026 nand P2_U4872 P2_U4871 P2_U3755 ; P2_U3146
g7027 nand P2_U4867 P2_U4866 P2_U3754 ; P2_U3147
g7028 nand P2_U4862 P2_U4861 P2_U3753 ; P2_U3148
g7029 nand P2_U4857 P2_U4856 P2_U3752 ; P2_U3149
g7030 nand P2_U4852 P2_U4851 P2_U3751 ; P2_U3150
g7031 nand P2_U4847 P2_U4846 P2_U3750 ; P2_U3151
g7032 nand P2_U4825 P2_U4824 P2_U3748 ; P2_U3152
g7033 nand P2_U4820 P2_U4819 P2_U3747 ; P2_U3153
g7034 nand P2_U4815 P2_U4814 P2_U3746 ; P2_U3154
g7035 nand P2_U4810 P2_U4809 P2_U3745 ; P2_U3155
g7036 nand P2_U4805 P2_U4804 P2_U3744 ; P2_U3156
g7037 nand P2_U4800 P2_U4799 P2_U3743 ; P2_U3157
g7038 nand P2_U4795 P2_U4794 P2_U3742 ; P2_U3158
g7039 nand P2_U4790 P2_U4789 P2_U3741 ; P2_U3159
g7040 nand P2_U4766 P2_U4765 P2_U3739 ; P2_U3160
g7041 nand P2_U4761 P2_U4760 P2_U3738 ; P2_U3161
g7042 nand P2_U4756 P2_U4755 P2_U3737 ; P2_U3162
g7043 nand P2_U4751 P2_U4750 P2_U3736 ; P2_U3163
g7044 nand P2_U4746 P2_U4745 P2_U3735 ; P2_U3164
g7045 nand P2_U4741 P2_U4740 P2_U3734 ; P2_U3165
g7046 nand P2_U4736 P2_U4735 P2_U3733 ; P2_U3166
g7047 nand P2_U4731 P2_U4730 P2_U3732 ; P2_U3167
g7048 nand P2_U4708 P2_U4707 P2_U3730 ; P2_U3168
g7049 nand P2_U4703 P2_U4702 P2_U3729 ; P2_U3169
g7050 nand P2_U4698 P2_U4697 P2_U3728 ; P2_U3170
g7051 nand P2_U4693 P2_U4692 P2_U3727 ; P2_U3171
g7052 nand P2_U4688 P2_U4687 P2_U3726 ; P2_U3172
g7053 nand P2_U4683 P2_U4682 P2_U3725 ; P2_U3173
g7054 nand P2_U4678 P2_U4677 P2_U3724 ; P2_U3174
g7055 nand P2_U4673 P2_U4672 P2_U3723 ; P2_U3175
g7056 nand P2_U8061 P2_U8060 P2_U3721 ; P2_U3176
g7057 nand P2_U4629 P2_U4628 P2_U4627 P2_U4454 ; P2_U3177
g7058 nand P2_U3716 P2_U4625 ; P2_U3178
g7059 and P2_U7917 P2_DATAWIDTH_REG_31__SCAN_IN ; P2_U3179
g7060 and P2_U7917 P2_DATAWIDTH_REG_30__SCAN_IN ; P2_U3180
g7061 and P2_U7917 P2_DATAWIDTH_REG_29__SCAN_IN ; P2_U3181
g7062 and P2_U7917 P2_DATAWIDTH_REG_28__SCAN_IN ; P2_U3182
g7063 and P2_U7917 P2_DATAWIDTH_REG_27__SCAN_IN ; P2_U3183
g7064 and P2_U7917 P2_DATAWIDTH_REG_26__SCAN_IN ; P2_U3184
g7065 and P2_U7917 P2_DATAWIDTH_REG_25__SCAN_IN ; P2_U3185
g7066 and P2_U7917 P2_DATAWIDTH_REG_24__SCAN_IN ; P2_U3186
g7067 and P2_U7917 P2_DATAWIDTH_REG_23__SCAN_IN ; P2_U3187
g7068 and P2_U7917 P2_DATAWIDTH_REG_22__SCAN_IN ; P2_U3188
g7069 and P2_U7917 P2_DATAWIDTH_REG_21__SCAN_IN ; P2_U3189
g7070 and P2_U7917 P2_DATAWIDTH_REG_20__SCAN_IN ; P2_U3190
g7071 and P2_U7917 P2_DATAWIDTH_REG_19__SCAN_IN ; P2_U3191
g7072 and P2_U7917 P2_DATAWIDTH_REG_18__SCAN_IN ; P2_U3192
g7073 and P2_U7917 P2_DATAWIDTH_REG_17__SCAN_IN ; P2_U3193
g7074 and P2_U7917 P2_DATAWIDTH_REG_16__SCAN_IN ; P2_U3194
g7075 and P2_U7917 P2_DATAWIDTH_REG_15__SCAN_IN ; P2_U3195
g7076 and P2_U7917 P2_DATAWIDTH_REG_14__SCAN_IN ; P2_U3196
g7077 and P2_U7917 P2_DATAWIDTH_REG_13__SCAN_IN ; P2_U3197
g7078 and P2_U7917 P2_DATAWIDTH_REG_12__SCAN_IN ; P2_U3198
g7079 and P2_U7917 P2_DATAWIDTH_REG_11__SCAN_IN ; P2_U3199
g7080 and P2_U7917 P2_DATAWIDTH_REG_10__SCAN_IN ; P2_U3200
g7081 and P2_U7917 P2_DATAWIDTH_REG_9__SCAN_IN ; P2_U3201
g7082 and P2_U7917 P2_DATAWIDTH_REG_8__SCAN_IN ; P2_U3202
g7083 and P2_U7917 P2_DATAWIDTH_REG_7__SCAN_IN ; P2_U3203
g7084 and P2_U7917 P2_DATAWIDTH_REG_6__SCAN_IN ; P2_U3204
g7085 and P2_U7917 P2_DATAWIDTH_REG_5__SCAN_IN ; P2_U3205
g7086 and P2_U7917 P2_DATAWIDTH_REG_4__SCAN_IN ; P2_U3206
g7087 and P2_U7917 P2_DATAWIDTH_REG_3__SCAN_IN ; P2_U3207
g7088 and P2_U7917 P2_DATAWIDTH_REG_2__SCAN_IN ; P2_U3208
g7089 nand P2_U7914 P2_U7913 P2_U4588 ; P2_U3209
g7090 nand P2_U7912 P2_U7911 P2_U3691 ; P2_U3210
g7091 nand P2_U3690 P2_U4579 ; P2_U3211
g7092 nand P2_U4566 P2_U4565 P2_U4567 ; P2_U3212
g7093 nand P2_U4563 P2_U4562 P2_U4564 ; P2_U3213
g7094 nand P2_U4560 P2_U4559 P2_U4561 ; P2_U3214
g7095 nand P2_U4557 P2_U4556 P2_U4558 ; P2_U3215
g7096 nand P2_U4554 P2_U4553 P2_U4555 ; P2_U3216
g7097 nand P2_U4551 P2_U4550 P2_U4552 ; P2_U3217
g7098 nand P2_U4548 P2_U4547 P2_U4549 ; P2_U3218
g7099 nand P2_U4545 P2_U4544 P2_U4546 ; P2_U3219
g7100 nand P2_U4542 P2_U4541 P2_U4543 ; P2_U3220
g7101 nand P2_U4539 P2_U4538 P2_U4540 ; P2_U3221
g7102 nand P2_U4536 P2_U4535 P2_U4537 ; P2_U3222
g7103 nand P2_U4533 P2_U4532 P2_U4534 ; P2_U3223
g7104 nand P2_U4530 P2_U4529 P2_U4531 ; P2_U3224
g7105 nand P2_U4527 P2_U4526 P2_U4528 ; P2_U3225
g7106 nand P2_U4524 P2_U4523 P2_U4525 ; P2_U3226
g7107 nand P2_U4521 P2_U4520 P2_U4522 ; P2_U3227
g7108 nand P2_U4518 P2_U4517 P2_U4519 ; P2_U3228
g7109 nand P2_U4515 P2_U4514 P2_U4516 ; P2_U3229
g7110 nand P2_U4512 P2_U4511 P2_U4513 ; P2_U3230
g7111 nand P2_U4509 P2_U4508 P2_U4510 ; P2_U3231
g7112 nand P2_U4506 P2_U4505 P2_U4507 ; P2_U3232
g7113 nand P2_U4503 P2_U4502 P2_U4504 ; P2_U3233
g7114 nand P2_U4500 P2_U4499 P2_U4501 ; P2_U3234
g7115 nand P2_U4497 P2_U4496 P2_U4498 ; P2_U3235
g7116 nand P2_U4494 P2_U4493 P2_U4495 ; P2_U3236
g7117 nand P2_U4491 P2_U4490 P2_U4492 ; P2_U3237
g7118 nand P2_U4488 P2_U4487 P2_U4489 ; P2_U3238
g7119 nand P2_U4485 P2_U4484 P2_U4486 ; P2_U3239
g7120 nand P2_U4482 P2_U4481 P2_U4483 ; P2_U3240
g7121 nand P2_U4479 P2_U4478 P2_U4480 ; P2_U3241
g7122 nand P2_U4194 P2_U4193 P2_U4192 P2_U4191 ; P2_U3242
g7123 nand P2_U3349 P2_U3335 ; P2_U3243
g7124 not P2_STATE_REG_2__SCAN_IN ; P2_U3244
g7125 nand P2_U2440 P2_U3243 ; P2_U3245
g7126 nand P2_U2440 P2_U4650 ; P2_U3246
g7127 nand P2_U2442 P2_U3243 ; P2_U3247
g7128 nand P2_U2442 P2_U4650 ; P2_U3248
g7129 nand P2_U2441 P2_U3243 ; P2_U3249
g7130 nand P2_U2441 P2_U4650 ; P2_U3250
g7131 nand P2_U2443 P2_U3243 ; P2_U3251
g7132 nand P2_U2443 P2_U4650 ; P2_U3252
g7133 nand P2_U3708 P2_U3707 ; P2_U3253
g7134 nand P2_U2590 P2_U4429 ; P2_U3254
g7135 nand P2_U3696 P2_U3695 ; P2_U3255
g7136 not P2_REQUESTPENDING_REG_SCAN_IN ; P2_U3256
g7137 nand P2_U8051 P2_U8050 P2_U4609 P2_U4608 ; P2_U3257
g7138 not P2_STATE_REG_1__SCAN_IN ; P2_U3258
g7139 nand P2_U3266 P2_STATE_REG_1__SCAN_IN ; P2_U3259
g7140 nand P2_U4439 P2_U3244 ; P2_U3260
g7141 nand P2_U4439 P2_STATE_REG_2__SCAN_IN ; P2_U3261
g7142 nand P2_U3244 P2_STATE_REG_1__SCAN_IN ; P2_U3262
g7143 or P2_STATE_REG_2__SCAN_IN P2_STATE_REG_1__SCAN_IN ; P2_U3263
g7144 not HOLD ; P2_U3264
g7145 not U211 ; P2_U3265
g7146 not P2_STATE_REG_0__SCAN_IN ; P2_U3266
g7147 nand P2_U3264 P2_REQUESTPENDING_REG_SCAN_IN ; P2_U3267
g7148 or HOLD P2_REQUESTPENDING_REG_SCAN_IN ; P2_U3268
g7149 not P2_STATE2_REG_1__SCAN_IN ; P2_U3269
g7150 not P2_STATE2_REG_2__SCAN_IN ; P2_U3270
g7151 not P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U3271
g7152 not P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U3272
g7153 not P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U3273
g7154 nand P2_U3276 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U3274
g7155 or P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U3275
g7156 not P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U3276
g7157 nand P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U3277
g7158 nand P2_U3700 P2_U3699 ; P2_U3278
g7159 nand P2_U3702 P2_U3701 ; P2_U3279
g7160 nand P2_U3704 P2_U3703 ; P2_U3280
g7161 nand P2_U7861 P2_U7863 P2_U7859 ; P2_U3281
g7162 nand P2_U2457 P2_U7869 P2_U4476 ; P2_U3282
g7163 nand P2_U3253 P2_U7873 ; P2_U3283
g7164 not P2_STATE2_REG_0__SCAN_IN ; P2_U3284
g7165 nand P2_U4424 P2_U3709 ; P2_U3285
g7166 nand P2_U3253 P2_U2616 ; P2_U3286
g7167 not P2_GTE_370_U6 ; P2_U3287
g7168 nand P2_U2457 P2_U7859 P2_U2458 ; P2_U3288
g7169 nand P2_U2616 P2_U7871 ; P2_U3289
g7170 nand P2_U4595 P2_U3266 ; P2_U3290
g7171 nand P2_U3713 P2_U2459 ; P2_U3291
g7172 not P2_R2243_U8 ; P2_U3292
g7173 nand P2_U2357 P2_U3280 ; P2_U3293
g7174 nand P2_U7871 P2_U7873 ; P2_U3294
g7175 nand P2_U7861 P2_U2617 ; P2_U3295
g7176 nand P2_U2451 P2_U4428 ; P2_U3296
g7177 not P2_R2167_U6 ; P2_U3297
g7178 nand P2_U7894 P2_U4444 P2_LT_563_U6 P2_U4614 P2_U4610 ; P2_U3298
g7179 nand P2_U4619 P2_STATE2_REG_0__SCAN_IN ; P2_U3299
g7180 not P2_STATE2_REG_3__SCAN_IN ; P2_U3300
g7181 nand P2_U3270 P2_STATE2_REG_0__SCAN_IN ; P2_U3301
g7182 not P2_STATEBS16_REG_SCAN_IN ; P2_U3302
g7183 or P2_STATE2_REG_3__SCAN_IN P2_STATE2_REG_1__SCAN_IN ; P2_U3303
g7184 nand P2_U3269 P2_STATE2_REG_2__SCAN_IN ; P2_U3304
g7185 nand P2_R2167_U6 P2_STATE2_REG_3__SCAN_IN ; P2_U3305
g7186 nand P2_U4656 P2_U3284 ; P2_U3306
g7187 not P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U3307
g7188 not P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_U3308
g7189 not P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U3309
g7190 not P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U3310
g7191 nand P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U3311
g7192 nand P2_U4642 P2_U2464 ; P2_U3312
g7193 or P2_STATE2_REG_3__SCAN_IN P2_STATE2_REG_2__SCAN_IN ; P2_U3313
g7194 not P2_R2182_U69 ; P2_U3314
g7195 not P2_R2182_U68 ; P2_U3315
g7196 not P2_R2182_U40 ; P2_U3316
g7197 not P2_R2182_U76 ; P2_U3317
g7198 nand P2_R2182_U68 P2_R2182_U69 ; P2_U3318
g7199 nand P2_U3352 P2_U3314 ; P2_U3319
g7200 nand P2_U4636 P2_U2461 ; P2_U3320
g7201 not P2_R2099_U95 ; P2_U3321
g7202 not P2_R2099_U96 ; P2_U3322
g7203 not P2_R2099_U94 ; P2_U3323
g7204 not P2_R2099_U5 ; P2_U3324
g7205 nand P2_U3312 P2_U4651 ; P2_U3325
g7206 nand P2_U3570 P2_U3312 ; P2_U3326
g7207 not P2_INSTQUEUE_REG_15__7__SCAN_IN ; P2_U3327
g7208 not P2_INSTQUEUE_REG_15__6__SCAN_IN ; P2_U3328
g7209 not P2_INSTQUEUE_REG_15__5__SCAN_IN ; P2_U3329
g7210 not P2_INSTQUEUE_REG_15__4__SCAN_IN ; P2_U3330
g7211 not P2_INSTQUEUE_REG_15__3__SCAN_IN ; P2_U3331
g7212 not P2_INSTQUEUE_REG_15__2__SCAN_IN ; P2_U3332
g7213 not P2_INSTQUEUE_REG_15__1__SCAN_IN ; P2_U3333
g7214 not P2_INSTQUEUE_REG_15__0__SCAN_IN ; P2_U3334
g7215 nand P2_U3307 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_U3335
g7216 nand P2_U4649 P2_U2464 ; P2_U3336
g7217 nand P2_R2182_U68 P2_U3314 ; P2_U3337
g7218 nand P2_R2182_U69 P2_U3352 ; P2_U3338
g7219 nand P2_U4709 P2_U2461 ; P2_U3339
g7220 nand P2_U3569 P2_U3336 ; P2_U3340
g7221 not P2_INSTQUEUE_REG_14__7__SCAN_IN ; P2_U3341
g7222 not P2_INSTQUEUE_REG_14__6__SCAN_IN ; P2_U3342
g7223 not P2_INSTQUEUE_REG_14__5__SCAN_IN ; P2_U3343
g7224 not P2_INSTQUEUE_REG_14__4__SCAN_IN ; P2_U3344
g7225 not P2_INSTQUEUE_REG_14__3__SCAN_IN ; P2_U3345
g7226 not P2_INSTQUEUE_REG_14__2__SCAN_IN ; P2_U3346
g7227 not P2_INSTQUEUE_REG_14__1__SCAN_IN ; P2_U3347
g7228 not P2_INSTQUEUE_REG_14__0__SCAN_IN ; P2_U3348
g7229 nand P2_U3308 P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U3349
g7230 nand P2_U4648 P2_U2464 ; P2_U3350
g7231 nand P2_R2182_U69 P2_U3315 ; P2_U3351
g7232 nand P2_U3337 P2_U3351 ; P2_U3352
g7233 nand P2_U4635 P2_U3314 ; P2_U3353
g7234 nand P2_U4767 P2_U2461 ; P2_U3354
g7235 nand P2_U3350 P2_U4770 ; P2_U3355
g7236 nand P2_U3568 P2_U3350 ; P2_U3356
g7237 not P2_INSTQUEUE_REG_13__7__SCAN_IN ; P2_U3357
g7238 not P2_INSTQUEUE_REG_13__6__SCAN_IN ; P2_U3358
g7239 not P2_INSTQUEUE_REG_13__5__SCAN_IN ; P2_U3359
g7240 not P2_INSTQUEUE_REG_13__4__SCAN_IN ; P2_U3360
g7241 not P2_INSTQUEUE_REG_13__3__SCAN_IN ; P2_U3361
g7242 not P2_INSTQUEUE_REG_13__2__SCAN_IN ; P2_U3362
g7243 not P2_INSTQUEUE_REG_13__1__SCAN_IN ; P2_U3363
g7244 not P2_INSTQUEUE_REG_13__0__SCAN_IN ; P2_U3364
g7245 nand P2_U2478 P2_U2464 ; P2_U3365
g7246 nand P2_U2475 P2_U2461 ; P2_U3366
g7247 nand P2_U3567 P2_U3365 ; P2_U3367
g7248 not P2_INSTQUEUE_REG_12__7__SCAN_IN ; P2_U3368
g7249 not P2_INSTQUEUE_REG_12__6__SCAN_IN ; P2_U3369
g7250 not P2_INSTQUEUE_REG_12__5__SCAN_IN ; P2_U3370
g7251 not P2_INSTQUEUE_REG_12__4__SCAN_IN ; P2_U3371
g7252 not P2_INSTQUEUE_REG_12__3__SCAN_IN ; P2_U3372
g7253 not P2_INSTQUEUE_REG_12__2__SCAN_IN ; P2_U3373
g7254 not P2_INSTQUEUE_REG_12__1__SCAN_IN ; P2_U3374
g7255 not P2_INSTQUEUE_REG_12__0__SCAN_IN ; P2_U3375
g7256 nand P2_U3310 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U3376
g7257 nand P2_U4645 P2_U4642 ; P2_U3377
g7258 nand P2_R2182_U76 P2_U3316 ; P2_U3378
g7259 nand P2_U2481 P2_U4636 ; P2_U3379
g7260 nand P2_U3377 P2_U4885 ; P2_U3380
g7261 nand P2_U3566 P2_U3377 ; P2_U3381
g7262 not P2_INSTQUEUE_REG_11__7__SCAN_IN ; P2_U3382
g7263 not P2_INSTQUEUE_REG_11__6__SCAN_IN ; P2_U3383
g7264 not P2_INSTQUEUE_REG_11__5__SCAN_IN ; P2_U3384
g7265 not P2_INSTQUEUE_REG_11__4__SCAN_IN ; P2_U3385
g7266 not P2_INSTQUEUE_REG_11__3__SCAN_IN ; P2_U3386
g7267 not P2_INSTQUEUE_REG_11__2__SCAN_IN ; P2_U3387
g7268 not P2_INSTQUEUE_REG_11__1__SCAN_IN ; P2_U3388
g7269 not P2_INSTQUEUE_REG_11__0__SCAN_IN ; P2_U3389
g7270 nand P2_U4645 P2_U4649 ; P2_U3390
g7271 nand P2_U2481 P2_U4709 ; P2_U3391
g7272 nand P2_U3565 P2_U3390 ; P2_U3392
g7273 not P2_INSTQUEUE_REG_10__7__SCAN_IN ; P2_U3393
g7274 not P2_INSTQUEUE_REG_10__6__SCAN_IN ; P2_U3394
g7275 not P2_INSTQUEUE_REG_10__5__SCAN_IN ; P2_U3395
g7276 not P2_INSTQUEUE_REG_10__4__SCAN_IN ; P2_U3396
g7277 not P2_INSTQUEUE_REG_10__3__SCAN_IN ; P2_U3397
g7278 not P2_INSTQUEUE_REG_10__2__SCAN_IN ; P2_U3398
g7279 not P2_INSTQUEUE_REG_10__1__SCAN_IN ; P2_U3399
g7280 not P2_INSTQUEUE_REG_10__0__SCAN_IN ; P2_U3400
g7281 nand P2_U4645 P2_U4648 ; P2_U3401
g7282 nand P2_U2481 P2_U4767 ; P2_U3402
g7283 nand P2_U3401 P2_U5000 ; P2_U3403
g7284 nand P2_U3564 P2_U3401 ; P2_U3404
g7285 not P2_INSTQUEUE_REG_9__7__SCAN_IN ; P2_U3405
g7286 not P2_INSTQUEUE_REG_9__6__SCAN_IN ; P2_U3406
g7287 not P2_INSTQUEUE_REG_9__5__SCAN_IN ; P2_U3407
g7288 not P2_INSTQUEUE_REG_9__4__SCAN_IN ; P2_U3408
g7289 not P2_INSTQUEUE_REG_9__3__SCAN_IN ; P2_U3409
g7290 not P2_INSTQUEUE_REG_9__2__SCAN_IN ; P2_U3410
g7291 not P2_INSTQUEUE_REG_9__1__SCAN_IN ; P2_U3411
g7292 not P2_INSTQUEUE_REG_9__0__SCAN_IN ; P2_U3412
g7293 nand P2_U4645 P2_U2478 ; P2_U3413
g7294 nand P2_U2481 P2_U2475 ; P2_U3414
g7295 nand P2_U3563 P2_U3413 ; P2_U3415
g7296 not P2_INSTQUEUE_REG_8__7__SCAN_IN ; P2_U3416
g7297 not P2_INSTQUEUE_REG_8__6__SCAN_IN ; P2_U3417
g7298 not P2_INSTQUEUE_REG_8__5__SCAN_IN ; P2_U3418
g7299 not P2_INSTQUEUE_REG_8__4__SCAN_IN ; P2_U3419
g7300 not P2_INSTQUEUE_REG_8__3__SCAN_IN ; P2_U3420
g7301 not P2_INSTQUEUE_REG_8__2__SCAN_IN ; P2_U3421
g7302 not P2_INSTQUEUE_REG_8__1__SCAN_IN ; P2_U3422
g7303 not P2_INSTQUEUE_REG_8__0__SCAN_IN ; P2_U3423
g7304 nand P2_U2465 P2_U4642 ; P2_U3424
g7305 nand P2_U2460 P2_U4637 ; P2_U3425
g7306 nand P2_U3378 P2_U4639 P2_U3425 ; P2_U3426
g7307 nand P2_U2491 P2_U4636 ; P2_U3427
g7308 nand P2_U3376 P2_U4646 P2_U3424 ; P2_U3428
g7309 nand P2_U3424 P2_U5114 ; P2_U3429
g7310 nand P2_U3562 P2_U3424 ; P2_U3430
g7311 not P2_INSTQUEUE_REG_7__7__SCAN_IN ; P2_U3431
g7312 not P2_INSTQUEUE_REG_7__6__SCAN_IN ; P2_U3432
g7313 not P2_INSTQUEUE_REG_7__5__SCAN_IN ; P2_U3433
g7314 not P2_INSTQUEUE_REG_7__4__SCAN_IN ; P2_U3434
g7315 not P2_INSTQUEUE_REG_7__3__SCAN_IN ; P2_U3435
g7316 not P2_INSTQUEUE_REG_7__2__SCAN_IN ; P2_U3436
g7317 not P2_INSTQUEUE_REG_7__1__SCAN_IN ; P2_U3437
g7318 not P2_INSTQUEUE_REG_7__0__SCAN_IN ; P2_U3438
g7319 nand P2_U4649 P2_U2465 ; P2_U3439
g7320 nand P2_U2491 P2_U4709 ; P2_U3440
g7321 nand P2_U3561 P2_U3439 ; P2_U3441
g7322 not P2_INSTQUEUE_REG_6__7__SCAN_IN ; P2_U3442
g7323 not P2_INSTQUEUE_REG_6__6__SCAN_IN ; P2_U3443
g7324 not P2_INSTQUEUE_REG_6__5__SCAN_IN ; P2_U3444
g7325 not P2_INSTQUEUE_REG_6__4__SCAN_IN ; P2_U3445
g7326 not P2_INSTQUEUE_REG_6__3__SCAN_IN ; P2_U3446
g7327 not P2_INSTQUEUE_REG_6__2__SCAN_IN ; P2_U3447
g7328 not P2_INSTQUEUE_REG_6__1__SCAN_IN ; P2_U3448
g7329 not P2_INSTQUEUE_REG_6__0__SCAN_IN ; P2_U3449
g7330 nand P2_U4648 P2_U2465 ; P2_U3450
g7331 nand P2_U2491 P2_U4767 ; P2_U3451
g7332 nand P2_U3450 P2_U5228 ; P2_U3452
g7333 nand P2_U3560 P2_U3450 ; P2_U3453
g7334 not P2_INSTQUEUE_REG_5__7__SCAN_IN ; P2_U3454
g7335 not P2_INSTQUEUE_REG_5__6__SCAN_IN ; P2_U3455
g7336 not P2_INSTQUEUE_REG_5__5__SCAN_IN ; P2_U3456
g7337 not P2_INSTQUEUE_REG_5__4__SCAN_IN ; P2_U3457
g7338 not P2_INSTQUEUE_REG_5__3__SCAN_IN ; P2_U3458
g7339 not P2_INSTQUEUE_REG_5__2__SCAN_IN ; P2_U3459
g7340 not P2_INSTQUEUE_REG_5__1__SCAN_IN ; P2_U3460
g7341 not P2_INSTQUEUE_REG_5__0__SCAN_IN ; P2_U3461
g7342 nand P2_U2478 P2_U2465 ; P2_U3462
g7343 nand P2_U2491 P2_U2475 ; P2_U3463
g7344 nand P2_U3559 P2_U3462 ; P2_U3464
g7345 not P2_INSTQUEUE_REG_4__7__SCAN_IN ; P2_U3465
g7346 not P2_INSTQUEUE_REG_4__6__SCAN_IN ; P2_U3466
g7347 not P2_INSTQUEUE_REG_4__5__SCAN_IN ; P2_U3467
g7348 not P2_INSTQUEUE_REG_4__4__SCAN_IN ; P2_U3468
g7349 not P2_INSTQUEUE_REG_4__3__SCAN_IN ; P2_U3469
g7350 not P2_INSTQUEUE_REG_4__2__SCAN_IN ; P2_U3470
g7351 not P2_INSTQUEUE_REG_4__1__SCAN_IN ; P2_U3471
g7352 not P2_INSTQUEUE_REG_4__0__SCAN_IN ; P2_U3472
g7353 nand P2_U2503 P2_U4642 ; P2_U3473
g7354 nand P2_U2500 P2_U4636 ; P2_U3474
g7355 nand P2_U3473 P2_U5343 ; P2_U3475
g7356 nand P2_U3558 P2_U3473 ; P2_U3476
g7357 not P2_INSTQUEUE_REG_3__7__SCAN_IN ; P2_U3477
g7358 not P2_INSTQUEUE_REG_3__6__SCAN_IN ; P2_U3478
g7359 not P2_INSTQUEUE_REG_3__5__SCAN_IN ; P2_U3479
g7360 not P2_INSTQUEUE_REG_3__4__SCAN_IN ; P2_U3480
g7361 not P2_INSTQUEUE_REG_3__3__SCAN_IN ; P2_U3481
g7362 not P2_INSTQUEUE_REG_3__2__SCAN_IN ; P2_U3482
g7363 not P2_INSTQUEUE_REG_3__1__SCAN_IN ; P2_U3483
g7364 not P2_INSTQUEUE_REG_3__0__SCAN_IN ; P2_U3484
g7365 nand P2_U2503 P2_U4649 ; P2_U3485
g7366 nand P2_U2500 P2_U4709 ; P2_U3486
g7367 nand P2_U3557 P2_U3485 ; P2_U3487
g7368 not P2_INSTQUEUE_REG_2__7__SCAN_IN ; P2_U3488
g7369 not P2_INSTQUEUE_REG_2__6__SCAN_IN ; P2_U3489
g7370 not P2_INSTQUEUE_REG_2__5__SCAN_IN ; P2_U3490
g7371 not P2_INSTQUEUE_REG_2__4__SCAN_IN ; P2_U3491
g7372 not P2_INSTQUEUE_REG_2__3__SCAN_IN ; P2_U3492
g7373 not P2_INSTQUEUE_REG_2__2__SCAN_IN ; P2_U3493
g7374 not P2_INSTQUEUE_REG_2__1__SCAN_IN ; P2_U3494
g7375 not P2_INSTQUEUE_REG_2__0__SCAN_IN ; P2_U3495
g7376 nand P2_U2503 P2_U4648 ; P2_U3496
g7377 nand P2_U2500 P2_U4767 ; P2_U3497
g7378 nand P2_U3496 P2_U5458 ; P2_U3498
g7379 nand P2_U3556 P2_U3496 ; P2_U3499
g7380 not P2_INSTQUEUE_REG_1__7__SCAN_IN ; P2_U3500
g7381 not P2_INSTQUEUE_REG_1__6__SCAN_IN ; P2_U3501
g7382 not P2_INSTQUEUE_REG_1__5__SCAN_IN ; P2_U3502
g7383 not P2_INSTQUEUE_REG_1__4__SCAN_IN ; P2_U3503
g7384 not P2_INSTQUEUE_REG_1__3__SCAN_IN ; P2_U3504
g7385 not P2_INSTQUEUE_REG_1__2__SCAN_IN ; P2_U3505
g7386 not P2_INSTQUEUE_REG_1__1__SCAN_IN ; P2_U3506
g7387 not P2_INSTQUEUE_REG_1__0__SCAN_IN ; P2_U3507
g7388 nand P2_U2503 P2_U2478 ; P2_U3508
g7389 nand P2_U2500 P2_U2475 ; P2_U3509
g7390 nand P2_U3555 P2_U3508 ; P2_U3510
g7391 not P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U3511
g7392 not P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U3512
g7393 not P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U3513
g7394 not P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U3514
g7395 not P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U3515
g7396 not P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U3516
g7397 not P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U3517
g7398 not P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U3518
g7399 not P2_FLUSH_REG_SCAN_IN ; P2_U3519
g7400 not P2_R2088_U6 ; P2_U3520
g7401 nand P2_U3698 P2_U3697 ; P2_U3521
g7402 nand P2_U2451 P2_U4429 ; P2_U3522
g7403 nand P2_U4475 P2_U4427 ; P2_U3523
g7404 nand P2_U4429 P2_U4475 ; P2_U3524
g7405 nand P2_U7865 P2_U7863 P2_U3279 P2_U7869 ; P2_U3525
g7406 not P2_R2147_U8 ; P2_U3526
g7407 nand P2_U3283 P2_U3289 ; P2_U3527
g7408 not P2_U3647 ; P2_U3528
g7409 not P2_R2147_U9 ; P2_U3529
g7410 nand P2_U3274 P2_U5615 ; P2_U3530
g7411 not P2_R2147_U4 ; P2_U3531
g7412 not P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U3532
g7413 nand P2_U4455 P2_U3306 P2_U5642 ; P2_U3533
g7414 nand P2_U4430 P2_U3269 ; P2_U3534
g7415 nand P2_U5672 P2_U5671 ; P2_U3535
g7416 nand P2_U7873 P2_STATE2_REG_0__SCAN_IN ; P2_U3536
g7417 nand P2_U5937 P2_U5936 ; P2_U3537
g7418 nand P2_U4055 P2_U2446 ; P2_U3538
g7419 nand P2_U4056 P2_U2357 ; P2_U3539
g7420 nand P2_U3284 P2_STATE2_REG_2__SCAN_IN ; P2_U3540
g7421 nand P2_U6231 P2_U6230 ; P2_U3541
g7422 nand P2_U2374 P2_U6326 ; P2_U3542
g7423 nand P2_U2374 P2_U6470 ; P2_U3543
g7424 not P2_EBX_REG_31__SCAN_IN ; P2_U3544
g7425 or U211 P2_STATEBS16_REG_SCAN_IN ; P2_U3545
g7426 nand P2_U4069 P2_U4462 ; P2_U3546
g7427 nand P2_U4181 P2_U4177 P2_U4174 P2_U4171 ; P2_U3547
g7428 nand P2_U4438 P2_REIP_REG_1__SCAN_IN ; P2_U3548
g7429 nand P2_U2356 P2_U4420 ; P2_U3549
g7430 nand P2_U4427 P2_STATE2_REG_0__SCAN_IN ; P2_U3550
g7431 not P2_CODEFETCH_REG_SCAN_IN ; P2_U3551
g7432 not P2_READREQUEST_REG_SCAN_IN ; P2_U3552
g7433 nand P2_U4405 P2_U3275 ; P2_U3553
g7434 nand P2_U4415 P2_U3576 ; P2_U3554
g7435 nand P2_U2504 P2_U2479 ; P2_U3555
g7436 nand P2_U2504 P2_U2473 ; P2_U3556
g7437 nand P2_U2504 P2_U2470 ; P2_U3557
g7438 nand P2_U2504 P2_U2467 ; P2_U3558
g7439 nand P2_U2492 P2_U2479 ; P2_U3559
g7440 nand P2_U2492 P2_U2473 ; P2_U3560
g7441 nand P2_U2492 P2_U2470 ; P2_U3561
g7442 nand P2_U2492 P2_U2467 ; P2_U3562
g7443 nand P2_U2483 P2_U2479 ; P2_U3563
g7444 nand P2_U2483 P2_U2473 ; P2_U3564
g7445 nand P2_U2483 P2_U2470 ; P2_U3565
g7446 nand P2_U2483 P2_U2467 ; P2_U3566
g7447 nand P2_U2479 P2_U2466 ; P2_U3567
g7448 nand P2_U2473 P2_U2466 ; P2_U3568
g7449 nand P2_U2470 P2_U2466 ; P2_U3569
g7450 nand P2_U2466 P2_U2467 ; P2_U3570
g7451 nand P2_U7865 P2_U3300 ; P2_U3571
g7452 not P2_U3242 ; P2_U3572
g7453 or P2_STATE2_REG_1__SCAN_IN P2_STATE2_REG_0__SCAN_IN ; P2_U3573
g7454 nand P2_U5571 P2_U3295 P2_U3521 ; P2_U3574
g7455 nand P2_U4419 P2_U7871 ; P2_U3575
g7456 nand P2_U4419 P2_U3279 ; P2_U3576
g7457 nand P2_U4424 P2_U6845 ; P2_U3577
g7458 nand P2_U2590 P2_U4428 ; P2_U3578
g7459 nand P2_U8063 P2_U8062 ; P2_U3579
g7460 nand P2_U8066 P2_U8065 ; P2_U3580
g7461 nand P2_U8081 P2_U8080 ; P2_U3581
g7462 nand P2_U8099 P2_U8098 ; P2_U3582
g7463 nand P2_U8148 P2_U8147 ; P2_U3583
g7464 nand P2_U8151 P2_U8150 ; P2_U3584
g7465 nand P2_U7900 P2_U7899 ; P2_U3585
g7466 nand P2_U7902 P2_U7901 ; P2_U3586
g7467 nand P2_U7904 P2_U7903 ; P2_U3587
g7468 nand P2_U7906 P2_U7905 ; P2_U3588
g7469 nand P2_U7916 P2_U7915 ; P2_U3589
g7470 and P2_U3263 P2_U4401 ; P2_U3590
g7471 nand P2_U7919 P2_U7918 ; P2_U3591
g7472 nand P2_U7921 P2_U7920 ; P2_U3592
g7473 nand P2_U8059 P2_U8058 ; P2_U3593
g7474 and P2_U3866 P2_U4434 ; P2_U3594
g7475 nand P2_U8073 P2_U8072 ; P2_U3595
g7476 nand P2_U8084 P2_U8083 ; P2_U3596
g7477 nand P2_U8086 P2_U8085 ; P2_U3597
g7478 nand P2_U8089 P2_U8088 ; P2_U3598
g7479 nand P2_U8094 P2_U8093 ; P2_U3599
g7480 nand P2_U8102 P2_U8101 ; P2_U3600
g7481 nand P2_U8104 P2_U8103 ; P2_U3601
g7482 nand P2_U8106 P2_U8105 ; P2_U3602
g7483 nand P2_U8111 P2_U8110 ; P2_U3603
g7484 nand P2_U8113 P2_U8112 ; P2_U3604
g7485 nand P2_U8115 P2_U8114 ; P2_U3605
g7486 nor P2_DATAWIDTH_REG_1__SCAN_IN P2_REIP_REG_1__SCAN_IN ; P2_U3606
g7487 and P2_U4183 P2_U7898 ; P2_U3607
g7488 nand P2_U8130 P2_U8129 ; P2_U3608
g7489 nand P2_U8134 P2_U8133 ; P2_U3609
g7490 nand P2_U8138 P2_U8137 ; P2_U3610
g7491 nand P2_U8142 P2_U8141 ; P2_U3611
g7492 nand P2_U8144 P2_U8143 ; P2_U3612
g7493 nand P2_U8282 P2_U8281 ; P2_U3613
g7494 nand P2_U8284 P2_U8283 ; P2_U3614
g7495 nand P2_U8286 P2_U8285 ; P2_U3615
g7496 and P2_U4434 P2_R2147_U7 ; P2_U3616
g7497 nand P2_U8288 P2_U8287 ; P2_U3617
g7498 nand P2_U8290 P2_U8289 ; P2_U3618
g7499 nand P2_U8292 P2_U8291 ; P2_U3619
g7500 nand P2_U8294 P2_U8293 ; P2_U3620
g7501 nand P2_U8296 P2_U8295 ; P2_U3621
g7502 nand P2_U8298 P2_U8297 ; P2_U3622
g7503 nand P2_U8300 P2_U8299 ; P2_U3623
g7504 nand P2_U8302 P2_U8301 ; P2_U3624
g7505 nand P2_U8304 P2_U8303 ; P2_U3625
g7506 nand P2_U8306 P2_U8305 ; P2_U3626
g7507 nand P2_U8308 P2_U8307 ; P2_U3627
g7508 nand P2_U8310 P2_U8309 ; P2_U3628
g7509 nand P2_U8312 P2_U8311 ; P2_U3629
g7510 nand P2_U8314 P2_U8313 ; P2_U3630
g7511 nand P2_U8316 P2_U8315 ; P2_U3631
g7512 nand P2_U8318 P2_U8317 ; P2_U3632
g7513 nand P2_U8320 P2_U8319 ; P2_U3633
g7514 nand P2_U8322 P2_U8321 ; P2_U3634
g7515 nand P2_U8324 P2_U8323 ; P2_U3635
g7516 nand P2_U8326 P2_U8325 ; P2_U3636
g7517 nand P2_U8328 P2_U8327 ; P2_U3637
g7518 nand P2_U8330 P2_U8329 ; P2_U3638
g7519 nand P2_U8332 P2_U8331 ; P2_U3639
g7520 nand P2_U8334 P2_U8333 ; P2_U3640
g7521 nand P2_U8336 P2_U8335 ; P2_U3641
g7522 nand P2_U8338 P2_U8337 ; P2_U3642
g7523 nand P2_U8340 P2_U8339 ; P2_U3643
g7524 nand P2_U8342 P2_U8341 ; P2_U3644
g7525 nand P2_U8344 P2_U8343 ; P2_U3645
g7526 nand P2_U8346 P2_U8345 ; P2_U3646
g7527 nand P2_U8350 P2_U8349 ; P2_U3647
g7528 nand P2_U8352 P2_U8351 ; P2_U3648
g7529 nand P2_U8354 P2_U8353 ; P2_U3649
g7530 nand P2_U8356 P2_U8355 ; P2_U3650
g7531 nand P2_U8358 P2_U8357 ; P2_U3651
g7532 nand P2_U8360 P2_U8359 ; P2_U3652
g7533 nand P2_U8362 P2_U8361 ; P2_U3653
g7534 nand P2_U8364 P2_U8363 ; P2_U3654
g7535 nand P2_U8366 P2_U8365 ; P2_U3655
g7536 nand P2_U8368 P2_U8367 ; P2_U3656
g7537 nand P2_U8370 P2_U8369 ; P2_U3657
g7538 nand P2_U8372 P2_U8371 ; P2_U3658
g7539 nand P2_U8374 P2_U8373 ; P2_U3659
g7540 nand P2_U8376 P2_U8375 ; P2_U3660
g7541 nand P2_U8378 P2_U8377 ; P2_U3661
g7542 nand P2_U8380 P2_U8379 ; P2_U3662
g7543 nand P2_U8382 P2_U8381 ; P2_U3663
g7544 nand P2_U8384 P2_U8383 ; P2_U3664
g7545 nand P2_U8386 P2_U8385 ; P2_U3665
g7546 nand P2_U8388 P2_U8387 ; P2_U3666
g7547 nand P2_U8390 P2_U8389 ; P2_U3667
g7548 nand P2_U8392 P2_U8391 ; P2_U3668
g7549 nand P2_U8394 P2_U8393 ; P2_U3669
g7550 nand P2_U8396 P2_U8395 ; P2_U3670
g7551 nand P2_U8398 P2_U8397 ; P2_U3671
g7552 nand P2_U8400 P2_U8399 ; P2_U3672
g7553 nand P2_U8402 P2_U8401 ; P2_U3673
g7554 nand P2_U8404 P2_U8403 ; P2_U3674
g7555 nand P2_U8406 P2_U8405 ; P2_U3675
g7556 nand P2_U8408 P2_U8407 ; P2_U3676
g7557 nand P2_U8410 P2_U8409 ; P2_U3677
g7558 nand P2_U8412 P2_U8411 ; P2_U3678
g7559 nand P2_U8414 P2_U8413 ; P2_U3679
g7560 nand P2_U8416 P2_U8415 ; P2_U3680
g7561 nand P2_U8418 P2_U8417 ; P2_U3681
g7562 nand P2_U8420 P2_U8419 ; P2_U3682
g7563 nand P2_U8422 P2_U8421 ; P2_U3683
g7564 nand P2_U8424 P2_U8423 ; P2_U3684
g7565 nand P2_U8426 P2_U8425 ; P2_U3685
g7566 nand P2_U8428 P2_U8427 ; P2_U3686
g7567 nand P2_U8430 P2_U8429 ; P2_U3687
g7568 nand P2_U8432 P2_U8431 ; P2_U3688
g7569 nand P2_U8434 P2_U8433 ; P2_U3689
g7570 and P2_U4578 P2_U3261 ; P2_U3690
g7571 and P2_U4583 P2_U3260 ; P2_U3691
g7572 and P2_STATE_REG_0__SCAN_IN P2_REQUESTPENDING_REG_SCAN_IN ; P2_U3692
g7573 and P2_U7799 P2_U7783 P2_U7767 P2_U7751 ; P2_U3693
g7574 and P2_U7868 P2_U7847 P2_U7831 P2_U7815 ; P2_U3694
g7575 and P2_U7798 P2_U7782 P2_U7766 P2_U7750 ; P2_U3695
g7576 and P2_U7866 P2_U7846 P2_U7830 P2_U7814 ; P2_U3696
g7577 and P2_U7797 P2_U7781 P2_U7765 P2_U7749 ; P2_U3697
g7578 and P2_U7864 P2_U7845 P2_U7829 P2_U7813 ; P2_U3698
g7579 and P2_U7796 P2_U7780 P2_U7764 P2_U7748 ; P2_U3699
g7580 and P2_U7862 P2_U7844 P2_U7828 P2_U7812 ; P2_U3700
g7581 and P2_U7795 P2_U7779 P2_U7763 P2_U7747 ; P2_U3701
g7582 and P2_U7860 P2_U7843 P2_U7827 P2_U7811 ; P2_U3702
g7583 and P2_U7794 P2_U7778 P2_U7762 P2_U7746 ; P2_U3703
g7584 and P2_U7858 P2_U7842 P2_U7826 P2_U7810 ; P2_U3704
g7585 and P2_U7801 P2_U7785 P2_U7769 P2_U7753 ; P2_U3705
g7586 and P2_U7872 P2_U7849 P2_U7833 P2_U7817 ; P2_U3706
g7587 and P2_U7800 P2_U7784 P2_U7768 P2_U7752 ; P2_U3707
g7588 and P2_U7870 P2_U7848 P2_U7832 P2_U7816 ; P2_U3708
g7589 and P2_U3710 P2_U4417 ; P2_U3709
g7590 and P2_U4595 P2_STATE2_REG_0__SCAN_IN ; P2_U3710
g7591 and P2_U2360 P2_U3266 ; P2_U3711
g7592 and P2_U3521 P2_U7867 ; P2_U3712
g7593 and P2_U4599 P2_U4598 ; P2_U3713
g7594 and P2_U3573 P2_STATE2_REG_2__SCAN_IN ; P2_U3714
g7595 and P2_U3714 P2_U4618 ; P2_U3715
g7596 and P2_U4624 P2_U3304 ; P2_U3716
g7597 and P2_U4466 P2_U3265 ; P2_U3717
g7598 and P2_U3269 P2_STATE2_REG_3__SCAN_IN ; P2_U3718
g7599 nor P2_STATE2_REG_2__SCAN_IN P2_STATE2_REG_1__SCAN_IN ; P2_U3719
g7600 and P2_U4465 P2_U4453 ; P2_U3720
g7601 and P2_U3720 P2_U4632 ; P2_U3721
g7602 and P2_U4661 P2_U4662 P2_U4443 ; P2_U3722
g7603 and P2_U4670 P2_U4669 P2_U4671 ; P2_U3723
g7604 and P2_U4675 P2_U4674 P2_U4676 ; P2_U3724
g7605 and P2_U4680 P2_U4679 P2_U4681 ; P2_U3725
g7606 and P2_U4685 P2_U4684 P2_U4686 ; P2_U3726
g7607 and P2_U4690 P2_U4689 P2_U4691 ; P2_U3727
g7608 and P2_U4695 P2_U4694 P2_U4696 ; P2_U3728
g7609 and P2_U4700 P2_U4699 P2_U4701 ; P2_U3729
g7610 and P2_U4705 P2_U4704 P2_U4706 ; P2_U3730
g7611 and P2_U4719 P2_U4720 P2_U4443 ; P2_U3731
g7612 and P2_U4728 P2_U4727 P2_U4729 ; P2_U3732
g7613 and P2_U4733 P2_U4732 P2_U4734 ; P2_U3733
g7614 and P2_U4738 P2_U4737 P2_U4739 ; P2_U3734
g7615 and P2_U4743 P2_U4742 P2_U4744 ; P2_U3735
g7616 and P2_U4748 P2_U4747 P2_U4749 ; P2_U3736
g7617 and P2_U4753 P2_U4752 P2_U4754 ; P2_U3737
g7618 and P2_U4758 P2_U4757 P2_U4759 ; P2_U3738
g7619 and P2_U4763 P2_U4762 P2_U4764 ; P2_U3739
g7620 and P2_U4778 P2_U4779 P2_U4443 ; P2_U3740
g7621 and P2_U4787 P2_U4786 P2_U4788 ; P2_U3741
g7622 and P2_U4792 P2_U4791 P2_U4793 ; P2_U3742
g7623 and P2_U4797 P2_U4796 P2_U4798 ; P2_U3743
g7624 and P2_U4802 P2_U4801 P2_U4803 ; P2_U3744
g7625 and P2_U4807 P2_U4806 P2_U4808 ; P2_U3745
g7626 and P2_U4812 P2_U4811 P2_U4813 ; P2_U3746
g7627 and P2_U4817 P2_U4816 P2_U4818 ; P2_U3747
g7628 and P2_U4822 P2_U4821 P2_U4823 ; P2_U3748
g7629 and P2_U4835 P2_U4836 P2_U4443 ; P2_U3749
g7630 and P2_U4844 P2_U4843 P2_U4845 ; P2_U3750
g7631 and P2_U4849 P2_U4848 P2_U4850 ; P2_U3751
g7632 and P2_U4854 P2_U4853 P2_U4855 ; P2_U3752
g7633 and P2_U4859 P2_U4858 P2_U4860 ; P2_U3753
g7634 and P2_U4864 P2_U4863 P2_U4865 ; P2_U3754
g7635 and P2_U4869 P2_U4868 P2_U4870 ; P2_U3755
g7636 and P2_U4874 P2_U4873 P2_U4875 ; P2_U3756
g7637 and P2_U4879 P2_U4878 P2_U4880 ; P2_U3757
g7638 and P2_U4893 P2_U4894 P2_U4443 ; P2_U3758
g7639 and P2_U4902 P2_U4901 P2_U4903 ; P2_U3759
g7640 and P2_U4907 P2_U4906 P2_U4908 ; P2_U3760
g7641 and P2_U4912 P2_U4911 P2_U4913 ; P2_U3761
g7642 and P2_U4917 P2_U4916 P2_U4918 ; P2_U3762
g7643 and P2_U4922 P2_U4921 P2_U4923 ; P2_U3763
g7644 and P2_U4927 P2_U4926 P2_U4928 ; P2_U3764
g7645 and P2_U4932 P2_U4931 P2_U4933 ; P2_U3765
g7646 and P2_U4937 P2_U4936 P2_U4938 ; P2_U3766
g7647 and P2_U4950 P2_U4951 P2_U4443 ; P2_U3767
g7648 and P2_U4959 P2_U4958 P2_U4960 ; P2_U3768
g7649 and P2_U4964 P2_U4963 P2_U4965 ; P2_U3769
g7650 and P2_U4969 P2_U4968 P2_U4970 ; P2_U3770
g7651 and P2_U4974 P2_U4973 P2_U4975 ; P2_U3771
g7652 and P2_U4979 P2_U4978 P2_U4980 ; P2_U3772
g7653 and P2_U4984 P2_U4983 P2_U4985 ; P2_U3773
g7654 and P2_U4989 P2_U4988 P2_U4990 ; P2_U3774
g7655 and P2_U4994 P2_U4993 P2_U4995 ; P2_U3775
g7656 and P2_U5008 P2_U5009 P2_U4443 ; P2_U3776
g7657 and P2_U5017 P2_U5016 P2_U5018 ; P2_U3777
g7658 and P2_U5022 P2_U5021 P2_U5023 ; P2_U3778
g7659 and P2_U5027 P2_U5026 P2_U5028 ; P2_U3779
g7660 and P2_U5032 P2_U5031 P2_U5033 ; P2_U3780
g7661 and P2_U5037 P2_U5036 P2_U5038 ; P2_U3781
g7662 and P2_U5042 P2_U5041 P2_U5043 ; P2_U3782
g7663 and P2_U5047 P2_U5046 P2_U5048 ; P2_U3783
g7664 and P2_U5052 P2_U5051 P2_U5053 ; P2_U3784
g7665 and P2_U5065 P2_U5066 P2_U4443 ; P2_U3785
g7666 and P2_U5074 P2_U5073 P2_U5075 ; P2_U3786
g7667 and P2_U5079 P2_U5078 P2_U5080 ; P2_U3787
g7668 and P2_U5084 P2_U5083 P2_U5085 ; P2_U3788
g7669 and P2_U5089 P2_U5088 P2_U5090 ; P2_U3789
g7670 and P2_U5094 P2_U5093 P2_U5095 ; P2_U3790
g7671 and P2_U5099 P2_U5098 P2_U5100 ; P2_U3791
g7672 and P2_U5104 P2_U5103 P2_U5105 ; P2_U3792
g7673 and P2_U5109 P2_U5108 P2_U5110 ; P2_U3793
g7674 and P2_U5121 P2_U5122 P2_U4443 ; P2_U3794
g7675 and P2_U5130 P2_U5129 P2_U5131 ; P2_U3795
g7676 and P2_U5135 P2_U5134 P2_U5136 ; P2_U3796
g7677 and P2_U5140 P2_U5139 P2_U5141 ; P2_U3797
g7678 and P2_U5145 P2_U5144 P2_U5146 ; P2_U3798
g7679 and P2_U5150 P2_U5149 P2_U5151 ; P2_U3799
g7680 and P2_U5155 P2_U5154 P2_U5156 ; P2_U3800
g7681 and P2_U5160 P2_U5159 P2_U5161 ; P2_U3801
g7682 and P2_U5165 P2_U5164 P2_U5166 ; P2_U3802
g7683 and P2_U5178 P2_U5179 P2_U4443 ; P2_U3803
g7684 and P2_U5187 P2_U5186 P2_U5188 ; P2_U3804
g7685 and P2_U5192 P2_U5191 P2_U5193 ; P2_U3805
g7686 and P2_U5197 P2_U5196 P2_U5198 ; P2_U3806
g7687 and P2_U5202 P2_U5201 P2_U5203 ; P2_U3807
g7688 and P2_U5207 P2_U5206 P2_U5208 ; P2_U3808
g7689 and P2_U5212 P2_U5211 P2_U5213 ; P2_U3809
g7690 and P2_U5217 P2_U5216 P2_U5218 ; P2_U3810
g7691 and P2_U5222 P2_U5221 P2_U5223 ; P2_U3811
g7692 and P2_U5236 P2_U5237 P2_U4443 ; P2_U3812
g7693 and P2_U5245 P2_U5244 P2_U5246 ; P2_U3813
g7694 and P2_U5250 P2_U5249 P2_U5251 ; P2_U3814
g7695 and P2_U5255 P2_U5254 P2_U5256 ; P2_U3815
g7696 and P2_U5260 P2_U5259 P2_U5261 ; P2_U3816
g7697 and P2_U5265 P2_U5264 P2_U5266 ; P2_U3817
g7698 and P2_U5270 P2_U5269 P2_U5271 ; P2_U3818
g7699 and P2_U5275 P2_U5274 P2_U5276 ; P2_U3819
g7700 and P2_U5280 P2_U5279 P2_U5281 ; P2_U3820
g7701 and P2_U5293 P2_U5294 P2_U4443 ; P2_U3821
g7702 and P2_U5302 P2_U5301 P2_U5303 ; P2_U3822
g7703 and P2_U5307 P2_U5306 P2_U5308 ; P2_U3823
g7704 and P2_U5312 P2_U5311 P2_U5313 ; P2_U3824
g7705 and P2_U5317 P2_U5316 P2_U5318 ; P2_U3825
g7706 and P2_U5322 P2_U5321 P2_U5323 ; P2_U3826
g7707 and P2_U5327 P2_U5326 P2_U5328 ; P2_U3827
g7708 and P2_U5332 P2_U5331 P2_U5333 ; P2_U3828
g7709 and P2_U5337 P2_U5336 P2_U5338 ; P2_U3829
g7710 and P2_U5351 P2_U5352 P2_U4443 ; P2_U3830
g7711 and P2_U5360 P2_U5359 P2_U5361 ; P2_U3831
g7712 and P2_U5365 P2_U5364 P2_U5366 ; P2_U3832
g7713 and P2_U5370 P2_U5369 P2_U5371 ; P2_U3833
g7714 and P2_U5375 P2_U5374 P2_U5376 ; P2_U3834
g7715 and P2_U5380 P2_U5379 P2_U5381 ; P2_U3835
g7716 and P2_U5385 P2_U5384 P2_U5386 ; P2_U3836
g7717 and P2_U5390 P2_U5389 P2_U5391 ; P2_U3837
g7718 and P2_U5395 P2_U5394 P2_U5396 ; P2_U3838
g7719 and P2_U5408 P2_U5409 P2_U4443 ; P2_U3839
g7720 and P2_U5417 P2_U5416 P2_U5418 ; P2_U3840
g7721 and P2_U5422 P2_U5421 P2_U5423 ; P2_U3841
g7722 and P2_U5427 P2_U5426 P2_U5428 ; P2_U3842
g7723 and P2_U5432 P2_U5431 P2_U5433 ; P2_U3843
g7724 and P2_U5437 P2_U5436 P2_U5438 ; P2_U3844
g7725 and P2_U5442 P2_U5441 P2_U5443 ; P2_U3845
g7726 and P2_U5447 P2_U5446 P2_U5448 ; P2_U3846
g7727 and P2_U5452 P2_U5451 P2_U5453 ; P2_U3847
g7728 and P2_U5466 P2_U5467 P2_U4443 ; P2_U3848
g7729 and P2_U5475 P2_U5474 P2_U5476 ; P2_U3849
g7730 and P2_U5480 P2_U5479 P2_U5481 ; P2_U3850
g7731 and P2_U5485 P2_U5484 P2_U5486 ; P2_U3851
g7732 and P2_U5490 P2_U5489 P2_U5491 ; P2_U3852
g7733 and P2_U5495 P2_U5494 P2_U5496 ; P2_U3853
g7734 and P2_U5500 P2_U5499 P2_U5501 ; P2_U3854
g7735 and P2_U5505 P2_U5504 P2_U5506 ; P2_U3855
g7736 and P2_U5510 P2_U5509 P2_U5511 ; P2_U3856
g7737 and P2_U5523 P2_U5524 P2_U4443 ; P2_U3857
g7738 and P2_U5532 P2_U5531 P2_U5533 ; P2_U3858
g7739 and P2_U5537 P2_U5536 P2_U5538 ; P2_U3859
g7740 and P2_U5542 P2_U5541 P2_U5543 ; P2_U3860
g7741 and P2_U5547 P2_U5546 P2_U5548 ; P2_U3861
g7742 and P2_U5552 P2_U5551 P2_U5553 ; P2_U3862
g7743 and P2_U5557 P2_U5556 P2_U5558 ; P2_U3863
g7744 and P2_U5562 P2_U5561 P2_U5563 ; P2_U3864
g7745 and P2_U5567 P2_U5566 P2_U5568 ; P2_U3865
g7746 and P2_R2147_U7 P2_U4466 ; P2_U3866
g7747 and P2_STATE2_REG_0__SCAN_IN P2_FLUSH_REG_SCAN_IN ; P2_U3867
g7748 and P2_U5573 P2_U5571 ; P2_U3868
g7749 and P2_U3868 P2_U5576 ; P2_U3869
g7750 and P2_U4460 P2_U4456 ; P2_U3870
g7751 and P2_U8071 P2_U8070 P2_U3870 P2_U2512 ; P2_U3871
g7752 and P2_U5583 P2_U4455 ; P2_U3872
g7753 and P2_U3521 P2_U7869 ; P2_U3873
g7754 and P2_U7861 P2_U3278 ; P2_U3874
g7755 and P2_U3874 P2_U4429 ; P2_U3875
g7756 and P2_U4429 P2_U3279 ; P2_U3876
g7757 and P2_U7859 P2_U5593 ; P2_U3877
g7758 and P2_U7863 P2_U3521 ; P2_U3878
g7759 and P2_U5587 P2_U5588 P2_U3281 ; P2_U3879
g7760 and P2_U5599 P2_U3254 ; P2_U3880
g7761 and P2_U5601 P2_U5600 P2_U3880 ; P2_U3881
g7762 and P2_U7897 P2_U5602 ; P2_U3882
g7763 and P2_U5608 P2_U5607 ; P2_U3883
g7764 and P2_U3883 P2_U5609 ; P2_U3884
g7765 and P2_U4396 P2_U5617 ; P2_U3885
g7766 and P2_U4601 P2_U2449 ; P2_U3886
g7767 and P2_U3582 P2_U7859 ; P2_U3887
g7768 and P2_U5627 P2_U5626 ; P2_U3888
g7769 and P2_U7859 P2_U3272 ; P2_U3889
g7770 and P2_U5635 P2_U5634 ; P2_U3890
g7771 and P2_U5649 P2_U5650 ; P2_U3891
g7772 and P2_U5653 P2_U5654 ; P2_U3892
g7773 and P2_U5658 P2_U5659 ; P2_U3893
g7774 and P2_U4460 P2_U5668 P2_U4456 ; P2_U3894
g7775 and P2_U5674 P2_U3578 ; P2_U3895
g7776 and P2_U5681 P2_U5680 ; P2_U3896
g7777 and P2_U5683 P2_U5682 ; P2_U3897
g7778 and P2_U5687 P2_U5686 ; P2_U3898
g7779 and P2_U5689 P2_U5688 ; P2_U3899
g7780 and P2_U5691 P2_U5690 ; P2_U3900
g7781 and P2_U5695 P2_U5694 ; P2_U3901
g7782 and P2_U5697 P2_U5696 ; P2_U3902
g7783 and P2_U5699 P2_U5698 ; P2_U3903
g7784 and P2_U5703 P2_U5702 ; P2_U3904
g7785 and P2_U5705 P2_U5704 ; P2_U3905
g7786 and P2_U5707 P2_U5706 ; P2_U3906
g7787 and P2_U5711 P2_U5710 ; P2_U3907
g7788 and P2_U5713 P2_U5712 ; P2_U3908
g7789 and P2_U5715 P2_U5714 ; P2_U3909
g7790 and P2_U5719 P2_U5718 ; P2_U3910
g7791 and P2_U5721 P2_U5720 ; P2_U3911
g7792 and P2_U5723 P2_U5722 ; P2_U3912
g7793 and P2_U5727 P2_U5726 ; P2_U3913
g7794 and P2_U5729 P2_U5728 ; P2_U3914
g7795 and P2_U5731 P2_U5730 ; P2_U3915
g7796 and P2_U5735 P2_U5734 ; P2_U3916
g7797 and P2_U5737 P2_U5736 ; P2_U3917
g7798 and P2_U5739 P2_U5738 ; P2_U3918
g7799 and P2_U5743 P2_U5742 ; P2_U3919
g7800 and P2_U5745 P2_U5744 ; P2_U3920
g7801 and P2_U5747 P2_U5746 ; P2_U3921
g7802 and P2_U5751 P2_U5750 ; P2_U3922
g7803 and P2_U5753 P2_U5752 ; P2_U3923
g7804 and P2_U5755 P2_U5754 ; P2_U3924
g7805 and P2_U5759 P2_U5758 ; P2_U3925
g7806 and P2_U5761 P2_U5760 ; P2_U3926
g7807 and P2_U5763 P2_U5762 ; P2_U3927
g7808 and P2_U5767 P2_U5766 ; P2_U3928
g7809 and P2_U5769 P2_U5768 ; P2_U3929
g7810 and P2_U5771 P2_U5770 ; P2_U3930
g7811 and P2_U5775 P2_U5774 ; P2_U3931
g7812 and P2_U5777 P2_U5776 ; P2_U3932
g7813 and P2_U5779 P2_U5778 ; P2_U3933
g7814 and P2_U5783 P2_U5782 ; P2_U3934
g7815 and P2_U5785 P2_U5784 ; P2_U3935
g7816 and P2_U5787 P2_U5786 ; P2_U3936
g7817 and P2_U5791 P2_U5790 ; P2_U3937
g7818 and P2_U5793 P2_U5792 ; P2_U3938
g7819 and P2_U5795 P2_U5794 ; P2_U3939
g7820 and P2_U5799 P2_U5798 ; P2_U3940
g7821 and P2_U5801 P2_U5800 ; P2_U3941
g7822 and P2_U5803 P2_U5802 ; P2_U3942
g7823 and P2_U5807 P2_U5806 ; P2_U3943
g7824 and P2_U5809 P2_U5808 ; P2_U3944
g7825 and P2_U5811 P2_U5810 ; P2_U3945
g7826 and P2_U5815 P2_U5814 ; P2_U3946
g7827 and P2_U5817 P2_U5816 ; P2_U3947
g7828 and P2_U5819 P2_U5818 ; P2_U3948
g7829 and P2_U5823 P2_U5822 ; P2_U3949
g7830 and P2_U5825 P2_U5824 ; P2_U3950
g7831 and P2_U5827 P2_U5826 ; P2_U3951
g7832 and P2_U5831 P2_U5830 ; P2_U3952
g7833 and P2_U5833 P2_U5832 ; P2_U3953
g7834 and P2_U5835 P2_U5834 ; P2_U3954
g7835 and P2_U5839 P2_U5838 ; P2_U3955
g7836 and P2_U5841 P2_U5840 ; P2_U3956
g7837 and P2_U5843 P2_U5842 ; P2_U3957
g7838 and P2_U5847 P2_U5846 ; P2_U3958
g7839 and P2_U5849 P2_U5848 ; P2_U3959
g7840 and P2_U5851 P2_U5850 ; P2_U3960
g7841 and P2_U5855 P2_U5854 ; P2_U3961
g7842 and P2_U5857 P2_U5856 ; P2_U3962
g7843 and P2_U5859 P2_U5858 ; P2_U3963
g7844 and P2_U5863 P2_U5862 ; P2_U3964
g7845 and P2_U5865 P2_U5864 ; P2_U3965
g7846 and P2_U5867 P2_U5866 ; P2_U3966
g7847 and P2_U5871 P2_U5870 ; P2_U3967
g7848 and P2_U5873 P2_U5872 ; P2_U3968
g7849 and P2_U5875 P2_U5874 ; P2_U3969
g7850 and P2_U5879 P2_U5878 ; P2_U3970
g7851 and P2_U5881 P2_U5880 ; P2_U3971
g7852 and P2_U5883 P2_U5882 ; P2_U3972
g7853 and P2_U5887 P2_U5886 ; P2_U3973
g7854 and P2_U5889 P2_U5888 ; P2_U3974
g7855 and P2_U5891 P2_U5890 ; P2_U3975
g7856 and P2_U5895 P2_U5894 ; P2_U3976
g7857 and P2_U5897 P2_U5896 ; P2_U3977
g7858 and P2_U5899 P2_U5898 ; P2_U3978
g7859 and P2_U5903 P2_U5902 ; P2_U3979
g7860 and P2_U5905 P2_U5904 ; P2_U3980
g7861 and P2_U5907 P2_U5906 ; P2_U3981
g7862 and P2_U5911 P2_U5910 ; P2_U3982
g7863 and P2_U5915 P2_U5914 P2_U5913 P2_U5912 ; P2_U3983
g7864 and P2_U5919 P2_U5918 ; P2_U3984
g7865 and P2_U5923 P2_U5922 P2_U5921 ; P2_U3985
g7866 and P2_U5927 P2_U5926 ; P2_U3986
g7867 and P2_U5931 P2_U5930 P2_U5929 ; P2_U3987
g7868 and P2_U5935 P2_U5934 ; P2_U3988
g7869 and P2_STATE2_REG_1__SCAN_IN P2_STATEBS16_REG_SCAN_IN ; P2_U3989
g7870 nor P2_STATE2_REG_2__SCAN_IN P2_STATE2_REG_1__SCAN_IN ; P2_U3990
g7871 and P2_U5942 P2_U5941 P2_U5943 ; P2_U3991
g7872 and P2_U5945 P2_U5944 P2_U5946 ; P2_U3992
g7873 and P2_U5948 P2_U5947 P2_U5949 ; P2_U3993
g7874 and P2_U5951 P2_U5950 P2_U5952 ; P2_U3994
g7875 and P2_U5954 P2_U5953 P2_U5955 ; P2_U3995
g7876 and P2_U5957 P2_U5956 P2_U5958 ; P2_U3996
g7877 and P2_U5960 P2_U5959 P2_U5961 ; P2_U3997
g7878 and P2_U5963 P2_U5962 P2_U5964 ; P2_U3998
g7879 and P2_U5966 P2_U5965 P2_U5967 ; P2_U3999
g7880 and P2_U5969 P2_U5968 P2_U5970 ; P2_U4000
g7881 and P2_U5972 P2_U5971 P2_U5973 ; P2_U4001
g7882 and P2_U5975 P2_U5974 P2_U5976 ; P2_U4002
g7883 and P2_U5978 P2_U5977 P2_U5979 ; P2_U4003
g7884 and P2_U5981 P2_U5980 P2_U5982 ; P2_U4004
g7885 and P2_U5984 P2_U5983 P2_U5985 ; P2_U4005
g7886 and P2_U5987 P2_U5986 P2_U5988 ; P2_U4006
g7887 and P2_U5990 P2_U5989 P2_U5991 ; P2_U4007
g7888 and P2_U5993 P2_U5992 P2_U5994 ; P2_U4008
g7889 and P2_U5996 P2_U5995 P2_U5997 ; P2_U4009
g7890 and P2_U5999 P2_U5998 P2_U6000 ; P2_U4010
g7891 and P2_U6002 P2_U6001 P2_U6003 ; P2_U4011
g7892 and P2_U6005 P2_U6004 P2_U6006 ; P2_U4012
g7893 and P2_U6008 P2_U6007 P2_U6009 ; P2_U4013
g7894 and P2_U6011 P2_U6010 P2_U6012 ; P2_U4014
g7895 and P2_U6014 P2_U6013 P2_U6015 ; P2_U4015
g7896 and P2_U6017 P2_U6016 P2_U6018 ; P2_U4016
g7897 and P2_U6020 P2_U6019 P2_U6021 ; P2_U4017
g7898 and P2_U6023 P2_U6022 P2_U6024 ; P2_U4018
g7899 and P2_U6026 P2_U6025 P2_U6027 ; P2_U4019
g7900 and P2_U6029 P2_U6028 P2_U6030 ; P2_U4020
g7901 and P2_U6032 P2_U6031 P2_U6033 ; P2_U4021
g7902 and P2_U6035 P2_U6034 P2_U6036 ; P2_U4022
g7903 and P2_U6038 P2_U6037 P2_U6039 ; P2_U4023
g7904 and P2_U6041 P2_U6040 P2_U6042 ; P2_U4024
g7905 and P2_U6044 P2_U6043 P2_U6045 ; P2_U4025
g7906 and P2_U6047 P2_U6046 P2_U6048 ; P2_U4026
g7907 and P2_U6050 P2_U6049 P2_U6051 ; P2_U4027
g7908 and P2_U6053 P2_U6052 P2_U6054 ; P2_U4028
g7909 and P2_U6056 P2_U6055 P2_U6057 ; P2_U4029
g7910 and P2_U6059 P2_U6058 P2_U6060 ; P2_U4030
g7911 and P2_U6062 P2_U6061 P2_U6063 ; P2_U4031
g7912 and P2_U6065 P2_U6064 P2_U6066 ; P2_U4032
g7913 and P2_U6068 P2_U6067 P2_U6069 ; P2_U4033
g7914 and P2_U6071 P2_U6070 P2_U6072 ; P2_U4034
g7915 and P2_U6074 P2_U6073 P2_U6075 ; P2_U4035
g7916 and P2_U6077 P2_U6076 P2_U6078 ; P2_U4036
g7917 and P2_U6080 P2_U6079 P2_U6081 ; P2_U4037
g7918 and P2_U6083 P2_U6082 P2_U6084 ; P2_U4038
g7919 and P2_U6086 P2_U6085 P2_U6087 ; P2_U4039
g7920 and P2_U6089 P2_U6088 P2_U6090 ; P2_U4040
g7921 and P2_U6092 P2_U6091 P2_U6093 ; P2_U4041
g7922 and P2_U6095 P2_U6094 P2_U6096 ; P2_U4042
g7923 and P2_U6098 P2_U6097 P2_U6099 ; P2_U4043
g7924 and P2_U6101 P2_U6100 P2_U6102 ; P2_U4044
g7925 and P2_U6104 P2_U6103 P2_U6105 ; P2_U4045
g7926 and P2_U6107 P2_U6106 P2_U6108 ; P2_U4046
g7927 and P2_U6110 P2_U6109 P2_U6111 ; P2_U4047
g7928 and P2_U6113 P2_U6112 P2_U6114 ; P2_U4048
g7929 and P2_U6116 P2_U6115 P2_U6117 ; P2_U4049
g7930 and P2_U6119 P2_U6118 P2_U6120 ; P2_U4050
g7931 and P2_U6122 P2_U6121 P2_U6123 ; P2_U4051
g7932 and P2_U6126 P2_U6124 P2_U6125 ; P2_U4052
g7933 and P2_U6128 P2_U6127 P2_U6129 ; P2_U4053
g7934 and P2_U6131 P2_U6130 P2_U6132 ; P2_U4054
g7935 and P2_U4468 P2_U6133 P2_U2356 ; P2_U4055
g7936 and P2_U3280 P2_U7871 P2_STATE2_REG_0__SCAN_IN ; P2_U4056
g7937 and P2_U2616 P2_U4468 ; P2_U4057
g7938 and P2_U2374 P2_U4417 ; P2_U4058
g7939 and P2_U6330 P2_U6329 ; P2_U4059
g7940 and P2_U6334 P2_U6333 ; P2_U4060
g7941 and P2_U6338 P2_U6337 ; P2_U4061
g7942 and P2_U6342 P2_U6341 ; P2_U4062
g7943 and P2_U6346 P2_U6345 ; P2_U4063
g7944 and P2_U6350 P2_U6349 ; P2_U4064
g7945 and P2_U6354 P2_U6353 ; P2_U4065
g7946 and P2_U6358 P2_U6357 ; P2_U4066
g7947 and P2_U6362 P2_U6361 ; P2_U4067
g7948 and P2_U6366 P2_U6365 ; P2_U4068
g7949 and P2_U4454 P2_U4453 P2_U6569 ; P2_U4069
g7950 and P2_U6574 P2_U6573 P2_U4071 ; P2_U4070
g7951 and P2_U6577 P2_U6576 ; P2_U4071
g7952 and P2_U4073 P2_U6578 ; P2_U4072
g7953 and P2_U6581 P2_U6580 ; P2_U4073
g7954 and P2_U6583 P2_U6582 P2_U4075 ; P2_U4074
g7955 and P2_U6586 P2_U6585 ; P2_U4075
g7956 and P2_U4077 P2_U6587 ; P2_U4076
g7957 and P2_U6590 P2_U6589 ; P2_U4077
g7958 and P2_U6592 P2_U6591 P2_U4079 ; P2_U4078
g7959 and P2_U6595 P2_U6594 ; P2_U4079
g7960 and P2_U4081 P2_U6596 ; P2_U4080
g7961 and P2_U6599 P2_U6598 ; P2_U4081
g7962 and P2_U6601 P2_U6600 P2_U4083 ; P2_U4082
g7963 and P2_U6604 P2_U6603 ; P2_U4083
g7964 and P2_U4085 P2_U6605 ; P2_U4084
g7965 and P2_U6608 P2_U6607 ; P2_U4085
g7966 and P2_U6609 P2_U4446 P2_U6610 ; P2_U4086
g7967 and P2_U4088 P2_U6615 ; P2_U4087
g7968 and P2_U6617 P2_U6616 ; P2_U4088
g7969 and P2_U6612 P2_U6611 P2_U4086 P2_U6613 P2_U6614 ; P2_U4089
g7970 and P2_U6618 P2_U4446 P2_U6619 ; P2_U4090
g7971 and P2_U4092 P2_U6624 ; P2_U4091
g7972 and P2_U6626 P2_U6625 ; P2_U4092
g7973 and P2_U6621 P2_U6620 P2_U4090 P2_U6622 P2_U6623 ; P2_U4093
g7974 and P2_U6627 P2_U4446 P2_U6628 ; P2_U4094
g7975 and P2_U4096 P2_U6631 ; P2_U4095
g7976 and P2_U6634 P2_U6633 ; P2_U4096
g7977 and P2_U6635 P2_U4446 P2_U6636 ; P2_U4097
g7978 and P2_U4099 P2_U6639 ; P2_U4098
g7979 and P2_U6642 P2_U6641 ; P2_U4099
g7980 and P2_U6643 P2_U4446 P2_U6644 ; P2_U4100
g7981 and P2_U4102 P2_U6647 ; P2_U4101
g7982 and P2_U6650 P2_U6649 ; P2_U4102
g7983 and P2_U6651 P2_U4446 P2_U6652 ; P2_U4103
g7984 and P2_U4105 P2_U6655 ; P2_U4104
g7985 and P2_U6658 P2_U6657 ; P2_U4105
g7986 and P2_U6659 P2_U4446 P2_U6660 ; P2_U4106
g7987 and P2_U4108 P2_U6663 ; P2_U4107
g7988 and P2_U6666 P2_U6665 ; P2_U4108
g7989 and P2_U6667 P2_U4446 P2_U6668 ; P2_U4109
g7990 and P2_U4111 P2_U6671 ; P2_U4110
g7991 and P2_U6674 P2_U6673 ; P2_U4111
g7992 and P2_U6675 P2_U4446 P2_U6678 ; P2_U4112
g7993 and P2_U4114 P2_U6679 ; P2_U4113
g7994 and P2_U6682 P2_U6681 ; P2_U4114
g7995 and P2_U6683 P2_U4446 P2_U6686 ; P2_U4115
g7996 and P2_U4117 P2_U6687 ; P2_U4116
g7997 and P2_U6690 P2_U6689 ; P2_U4117
g7998 and P2_U6691 P2_U4446 P2_U6694 ; P2_U4118
g7999 and P2_U4120 P2_U6695 ; P2_U4119
g8000 and P2_U6698 P2_U6697 ; P2_U4120
g8001 and P2_U6699 P2_U4446 ; P2_U4121
g8002 and P2_U4123 P2_U6703 ; P2_U4122
g8003 and P2_U6706 P2_U6705 ; P2_U4123
g8004 and P2_U4121 P2_U6701 P2_U6702 P2_U6700 P2_U6704 ; P2_U4124
g8005 and P2_U6707 P2_U4446 ; P2_U4125
g8006 and P2_U4127 P2_U6711 ; P2_U4126
g8007 and P2_U6714 P2_U6713 ; P2_U4127
g8008 and P2_U4125 P2_U6709 P2_U6710 P2_U6708 P2_U6712 ; P2_U4128
g8009 and P2_U6715 P2_U4446 ; P2_U4129
g8010 and P2_U4131 P2_U6719 ; P2_U4130
g8011 and P2_U6722 P2_U6721 ; P2_U4131
g8012 and P2_U4129 P2_U6717 P2_U6718 P2_U6716 P2_U6720 ; P2_U4132
g8013 and P2_U6723 P2_U4446 ; P2_U4133
g8014 and P2_U4135 P2_U6727 ; P2_U4134
g8015 and P2_U6730 P2_U6729 ; P2_U4135
g8016 and P2_U4133 P2_U6725 P2_U6726 P2_U6724 P2_U6728 ; P2_U4136
g8017 and P2_U6731 P2_U4446 ; P2_U4137
g8018 and P2_U4139 P2_U6735 ; P2_U4138
g8019 and P2_U6738 P2_U6737 ; P2_U4139
g8020 and P2_U4137 P2_U6733 P2_U6734 P2_U6732 P2_U6736 ; P2_U4140
g8021 and P2_U4142 P2_U6743 ; P2_U4141
g8022 and P2_U6746 P2_U6745 ; P2_U4142
g8023 and P2_U6739 P2_U6741 P2_U6742 P2_U6740 P2_U6744 ; P2_U4143
g8024 and P2_U4145 P2_U6751 ; P2_U4144
g8025 and P2_U6754 P2_U6753 ; P2_U4145
g8026 and P2_U6747 P2_U6749 P2_U6750 P2_U6748 P2_U6752 ; P2_U4146
g8027 and P2_U6762 P2_U6761 ; P2_U4147
g8028 and P2_U4147 P2_U6759 P2_U6760 ; P2_U4148
g8029 and P2_U6763 P2_U6765 P2_U6766 P2_U6768 P2_U4150 ; P2_U4149
g8030 and P2_U4151 P2_U6767 ; P2_U4150
g8031 and P2_U6770 P2_U6769 ; P2_U4151
g8032 and P2_U6771 P2_U6773 P2_U6774 P2_U6776 P2_U4153 ; P2_U4152
g8033 and P2_U4154 P2_U6775 ; P2_U4153
g8034 and P2_U6778 P2_U6777 ; P2_U4154
g8035 and P2_U6786 P2_U6785 ; P2_U4155
g8036 and P2_U4155 P2_U6783 P2_U6784 ; P2_U4156
g8037 and P2_U6794 P2_U6793 ; P2_U4157
g8038 and P2_U4157 P2_U6791 P2_U6792 ; P2_U4158
g8039 and P2_U6802 P2_U6801 ; P2_U4159
g8040 and P2_U4159 P2_U6799 P2_U6800 ; P2_U4160
g8041 and P2_U6810 P2_U6809 ; P2_U4161
g8042 and P2_U4161 P2_U6807 P2_U6808 ; P2_U4162
g8043 and P2_U6818 P2_U6817 ; P2_U4163
g8044 and P2_U4163 P2_U6815 P2_U6816 ; P2_U4164
g8045 and P2_U6826 P2_U6825 ; P2_U4165
g8046 and P2_U4165 P2_U6823 P2_U6824 ; P2_U4166
g8047 and P2_U6834 P2_U6833 ; P2_U4167
g8048 and P2_U4167 P2_U6831 P2_U6832 ; P2_U4168
g8049 nor P2_DATAWIDTH_REG_2__SCAN_IN P2_DATAWIDTH_REG_3__SCAN_IN P2_DATAWIDTH_REG_4__SCAN_IN P2_DATAWIDTH_REG_5__SCAN_IN ; P2_U4169
g8050 nor P2_DATAWIDTH_REG_6__SCAN_IN P2_DATAWIDTH_REG_7__SCAN_IN P2_DATAWIDTH_REG_8__SCAN_IN P2_DATAWIDTH_REG_9__SCAN_IN ; P2_U4170
g8051 and P2_U4170 P2_U4169 ; P2_U4171
g8052 nor P2_DATAWIDTH_REG_10__SCAN_IN P2_DATAWIDTH_REG_11__SCAN_IN P2_DATAWIDTH_REG_12__SCAN_IN P2_DATAWIDTH_REG_13__SCAN_IN ; P2_U4172
g8053 nor P2_DATAWIDTH_REG_14__SCAN_IN P2_DATAWIDTH_REG_15__SCAN_IN P2_DATAWIDTH_REG_16__SCAN_IN P2_DATAWIDTH_REG_17__SCAN_IN ; P2_U4173
g8054 and P2_U4173 P2_U4172 ; P2_U4174
g8055 nor P2_DATAWIDTH_REG_18__SCAN_IN P2_DATAWIDTH_REG_19__SCAN_IN P2_DATAWIDTH_REG_20__SCAN_IN P2_DATAWIDTH_REG_21__SCAN_IN ; P2_U4175
g8056 nor P2_DATAWIDTH_REG_22__SCAN_IN P2_DATAWIDTH_REG_23__SCAN_IN P2_DATAWIDTH_REG_24__SCAN_IN P2_DATAWIDTH_REG_25__SCAN_IN ; P2_U4176
g8057 and P2_U4176 P2_U4175 ; P2_U4177
g8058 nor P2_DATAWIDTH_REG_26__SCAN_IN P2_DATAWIDTH_REG_27__SCAN_IN ; P2_U4178
g8059 nor P2_DATAWIDTH_REG_28__SCAN_IN P2_DATAWIDTH_REG_29__SCAN_IN ; P2_U4179
g8060 nor P2_DATAWIDTH_REG_30__SCAN_IN P2_DATAWIDTH_REG_31__SCAN_IN ; P2_U4180
g8061 and P2_U4180 P2_U6835 P2_U4179 P2_U4178 ; P2_U4181
g8062 nor P2_DATAWIDTH_REG_0__SCAN_IN P2_DATAWIDTH_REG_1__SCAN_IN P2_REIP_REG_0__SCAN_IN ; P2_U4182
g8063 nor P2_DATAWIDTH_REG_1__SCAN_IN P2_REIP_REG_1__SCAN_IN ; P2_U4183
g8064 and P2_U6844 P2_U7873 ; P2_U4184
g8065 and P2_U6848 P2_U3301 ; P2_U4185
g8066 and P2_U4185 P2_U6849 ; P2_U4186
g8067 and P2_U3265 P2_STATE2_REG_1__SCAN_IN ; P2_U4187
g8068 and P2_U6842 P2_U3313 P2_U6841 ; P2_U4188
g8069 and P2_U2374 P2_U3253 ; P2_U4189
g8070 and P2_U6860 P2_U3534 ; P2_U4190
g8071 and P2_U6865 P2_U6864 P2_U6863 P2_U6862 ; P2_U4191
g8072 and P2_U6869 P2_U6868 P2_U6867 P2_U6866 ; P2_U4192
g8073 and P2_U6873 P2_U6872 P2_U6871 P2_U6870 ; P2_U4193
g8074 and P2_U6877 P2_U6876 P2_U6875 P2_U6874 ; P2_U4194
g8075 and P2_U6881 P2_U6880 P2_U6879 P2_U6878 ; P2_U4195
g8076 and P2_U6885 P2_U6884 P2_U6883 P2_U6882 ; P2_U4196
g8077 and P2_U6889 P2_U6888 P2_U6887 P2_U6886 ; P2_U4197
g8078 and P2_U6893 P2_U6892 P2_U6891 P2_U6890 ; P2_U4198
g8079 and P2_U6897 P2_U6896 P2_U6895 P2_U6894 ; P2_U4199
g8080 and P2_U6901 P2_U6900 P2_U6899 P2_U6898 ; P2_U4200
g8081 and P2_U6905 P2_U6904 P2_U6903 P2_U6902 ; P2_U4201
g8082 and P2_U6909 P2_U6908 P2_U6907 P2_U6906 ; P2_U4202
g8083 and P2_U6913 P2_U6912 P2_U6911 P2_U6910 ; P2_U4203
g8084 and P2_U6917 P2_U6916 P2_U6915 P2_U6914 ; P2_U4204
g8085 and P2_U6921 P2_U6920 P2_U6919 P2_U6918 ; P2_U4205
g8086 and P2_U6925 P2_U6924 P2_U6923 P2_U6922 ; P2_U4206
g8087 and P2_U6929 P2_U6928 P2_U6927 P2_U6926 ; P2_U4207
g8088 and P2_U6933 P2_U6932 P2_U6931 P2_U6930 ; P2_U4208
g8089 and P2_U6937 P2_U6936 P2_U6935 P2_U6934 ; P2_U4209
g8090 and P2_U6941 P2_U6940 P2_U6939 P2_U6938 ; P2_U4210
g8091 and P2_U6945 P2_U6944 P2_U6943 P2_U6942 ; P2_U4211
g8092 and P2_U6949 P2_U6948 P2_U6947 P2_U6946 ; P2_U4212
g8093 and P2_U6953 P2_U6952 P2_U6951 P2_U6950 ; P2_U4213
g8094 and P2_U6957 P2_U6956 P2_U6955 P2_U6954 ; P2_U4214
g8095 and P2_U6961 P2_U6960 P2_U6959 P2_U6958 ; P2_U4215
g8096 and P2_U6965 P2_U6964 P2_U6963 P2_U6962 ; P2_U4216
g8097 and P2_U6969 P2_U6968 P2_U6967 P2_U6966 ; P2_U4217
g8098 and P2_U6973 P2_U6972 P2_U6971 P2_U6970 ; P2_U4218
g8099 and P2_U6977 P2_U6976 P2_U6975 P2_U6974 ; P2_U4219
g8100 and P2_U6981 P2_U6980 P2_U6979 P2_U6978 ; P2_U4220
g8101 and P2_U6985 P2_U6984 P2_U6983 P2_U6982 ; P2_U4221
g8102 and P2_U6989 P2_U6988 P2_U6987 P2_U6986 ; P2_U4222
g8103 and P2_U6993 P2_U6992 P2_U6991 P2_U6990 ; P2_U4223
g8104 and P2_U6997 P2_U6996 P2_U6995 P2_U6994 ; P2_U4224
g8105 and P2_U7001 P2_U7000 P2_U6999 P2_U6998 ; P2_U4225
g8106 and P2_U7005 P2_U7004 P2_U7003 P2_U7002 ; P2_U4226
g8107 and P2_U7011 P2_U7010 P2_U7009 P2_U7008 ; P2_U4227
g8108 and P2_U7015 P2_U7014 P2_U7013 P2_U7012 ; P2_U4228
g8109 and P2_U7019 P2_U7018 P2_U7017 P2_U7016 ; P2_U4229
g8110 and P2_U7023 P2_U7022 P2_U7021 P2_U7020 ; P2_U4230
g8111 and P2_U7027 P2_U7026 P2_U7025 P2_U7024 ; P2_U4231
g8112 and P2_U7031 P2_U7030 P2_U7029 P2_U7028 ; P2_U4232
g8113 and P2_U7035 P2_U7034 P2_U7033 P2_U7032 ; P2_U4233
g8114 and P2_U7039 P2_U7038 P2_U7037 P2_U7036 ; P2_U4234
g8115 and P2_U7043 P2_U7042 P2_U7041 P2_U7040 ; P2_U4235
g8116 and P2_U7047 P2_U7046 P2_U7045 P2_U7044 ; P2_U4236
g8117 and P2_U7051 P2_U7050 P2_U7049 P2_U7048 ; P2_U4237
g8118 and P2_U7055 P2_U7054 P2_U7053 P2_U7052 ; P2_U4238
g8119 and P2_U7059 P2_U7058 P2_U7057 P2_U7056 ; P2_U4239
g8120 and P2_U7063 P2_U7062 P2_U7061 P2_U7060 ; P2_U4240
g8121 and P2_U7067 P2_U7066 P2_U7065 P2_U7064 ; P2_U4241
g8122 and P2_U7071 P2_U7070 P2_U7069 P2_U7068 ; P2_U4242
g8123 and P2_U7075 P2_U7074 P2_U7073 P2_U7072 ; P2_U4243
g8124 and P2_U7079 P2_U7078 P2_U7077 P2_U7076 ; P2_U4244
g8125 and P2_U7083 P2_U7082 P2_U7081 P2_U7080 ; P2_U4245
g8126 and P2_U7087 P2_U7086 P2_U7085 P2_U7084 ; P2_U4246
g8127 and P2_U7091 P2_U7090 P2_U7089 P2_U7088 ; P2_U4247
g8128 and P2_U7095 P2_U7094 P2_U7093 P2_U7092 ; P2_U4248
g8129 and P2_U7099 P2_U7098 P2_U7097 P2_U7096 ; P2_U4249
g8130 and P2_U7103 P2_U7102 P2_U7101 P2_U7100 ; P2_U4250
g8131 and P2_U7107 P2_U7106 P2_U7105 P2_U7104 ; P2_U4251
g8132 and P2_U7111 P2_U7110 P2_U7109 P2_U7108 ; P2_U4252
g8133 and P2_U7115 P2_U7114 P2_U7113 P2_U7112 ; P2_U4253
g8134 and P2_U7119 P2_U7118 P2_U7117 P2_U7116 ; P2_U4254
g8135 and P2_U7123 P2_U7122 P2_U7121 P2_U7120 ; P2_U4255
g8136 and P2_U7127 P2_U7126 P2_U7125 P2_U7124 ; P2_U4256
g8137 and P2_U7131 P2_U7130 P2_U7129 P2_U7128 ; P2_U4257
g8138 and P2_U7135 P2_U7134 P2_U7133 P2_U7132 ; P2_U4258
g8139 and P2_U7802 P2_U7786 P2_U7770 P2_U7754 ; P2_U4259
g8140 and P2_U7874 P2_U7850 P2_U7834 P2_U7818 ; P2_U4260
g8141 and P2_U7803 P2_U7787 P2_U7771 P2_U7755 ; P2_U4261
g8142 and P2_U7875 P2_U7851 P2_U7835 P2_U7819 ; P2_U4262
g8143 and P2_U7804 P2_U7788 P2_U7772 P2_U7756 ; P2_U4263
g8144 and P2_U7876 P2_U7852 P2_U7836 P2_U7820 ; P2_U4264
g8145 and P2_U7805 P2_U7789 P2_U7773 P2_U7757 ; P2_U4265
g8146 and P2_U7877 P2_U7853 P2_U7837 P2_U7821 ; P2_U4266
g8147 and P2_U7806 P2_U7790 P2_U7774 P2_U7758 ; P2_U4267
g8148 and P2_U7878 P2_U7854 P2_U7838 P2_U7822 ; P2_U4268
g8149 and P2_U7807 P2_U7791 P2_U7775 P2_U7759 ; P2_U4269
g8150 and P2_U7879 P2_U7855 P2_U7839 P2_U7823 ; P2_U4270
g8151 and P2_U7808 P2_U7792 P2_U7776 P2_U7760 ; P2_U4271
g8152 and P2_U7880 P2_U7856 P2_U7840 P2_U7824 ; P2_U4272
g8153 and P2_U7809 P2_U7793 P2_U7777 P2_U7761 ; P2_U4273
g8154 and P2_U7881 P2_U7857 P2_U7841 P2_U7825 ; P2_U4274
g8155 and P2_U7861 P2_U4276 ; P2_U4275
g8156 and P2_U3300 P2_STATE2_REG_2__SCAN_IN P2_STATE2_REG_0__SCAN_IN ; P2_U4276
g8157 and P2_U7170 P2_U7169 P2_U7168 P2_U7167 ; P2_U4277
g8158 and P2_U7174 P2_U7173 P2_U7172 P2_U7171 ; P2_U4278
g8159 and P2_U7178 P2_U7177 P2_U7176 P2_U7175 ; P2_U4279
g8160 and P2_U7182 P2_U7181 P2_U7180 P2_U7179 ; P2_U4280
g8161 and P2_U7187 P2_U7186 P2_U7185 P2_U7184 ; P2_U4281
g8162 and P2_U7191 P2_U7190 P2_U7189 P2_U7188 ; P2_U4282
g8163 and P2_U7195 P2_U7194 P2_U7193 P2_U7192 ; P2_U4283
g8164 and P2_U7199 P2_U7198 P2_U7197 P2_U7196 ; P2_U4284
g8165 and P2_U7204 P2_U7203 P2_U7202 P2_U7201 ; P2_U4285
g8166 and P2_U7208 P2_U7207 P2_U7206 P2_U7205 ; P2_U4286
g8167 and P2_U7212 P2_U7211 P2_U7210 P2_U7209 ; P2_U4287
g8168 and P2_U7216 P2_U7215 P2_U7214 P2_U7213 ; P2_U4288
g8169 and P2_U7221 P2_U7220 P2_U7219 P2_U7218 ; P2_U4289
g8170 and P2_U7225 P2_U7224 P2_U7223 P2_U7222 ; P2_U4290
g8171 and P2_U7229 P2_U7228 P2_U7227 P2_U7226 ; P2_U4291
g8172 and P2_U7233 P2_U7232 P2_U7231 P2_U7230 ; P2_U4292
g8173 and P2_U7238 P2_U7237 P2_U7236 P2_U7235 ; P2_U4293
g8174 and P2_U7242 P2_U7241 P2_U7240 P2_U7239 ; P2_U4294
g8175 and P2_U7246 P2_U7245 P2_U7244 P2_U7243 ; P2_U4295
g8176 and P2_U7250 P2_U7249 P2_U7248 P2_U7247 ; P2_U4296
g8177 and P2_U7255 P2_U7254 P2_U7253 P2_U7252 ; P2_U4297
g8178 and P2_U7259 P2_U7258 P2_U7257 P2_U7256 ; P2_U4298
g8179 and P2_U7263 P2_U7262 P2_U7261 P2_U7260 ; P2_U4299
g8180 and P2_U7267 P2_U7266 P2_U7265 P2_U7264 ; P2_U4300
g8181 and P2_U7272 P2_U7271 P2_U7270 P2_U7269 ; P2_U4301
g8182 and P2_U7276 P2_U7275 P2_U7274 P2_U7273 ; P2_U4302
g8183 and P2_U7280 P2_U7279 P2_U7278 P2_U7277 ; P2_U4303
g8184 and P2_U7284 P2_U7283 P2_U7282 P2_U7281 ; P2_U4304
g8185 and P2_U7289 P2_U7288 P2_U7287 P2_U7286 ; P2_U4305
g8186 and P2_U7293 P2_U7292 P2_U7291 P2_U7290 ; P2_U4306
g8187 and P2_U7297 P2_U7296 P2_U7295 P2_U7294 ; P2_U4307
g8188 and P2_U7301 P2_U7300 P2_U7299 P2_U7298 ; P2_U4308
g8189 and P2_U7306 P2_U7305 P2_U7304 P2_U7303 ; P2_U4309
g8190 and P2_U7310 P2_U7309 P2_U7308 P2_U7307 ; P2_U4310
g8191 and P2_U7314 P2_U7313 P2_U7312 P2_U7311 ; P2_U4311
g8192 and P2_U7318 P2_U7317 P2_U7316 P2_U7315 ; P2_U4312
g8193 and P2_U7323 P2_U7322 P2_U7321 P2_U7320 ; P2_U4313
g8194 and P2_U7327 P2_U7326 P2_U7325 P2_U7324 ; P2_U4314
g8195 and P2_U7331 P2_U7330 P2_U7329 P2_U7328 ; P2_U4315
g8196 and P2_U7335 P2_U7334 P2_U7333 P2_U7332 ; P2_U4316
g8197 and P2_U7340 P2_U7339 P2_U7338 P2_U7337 ; P2_U4317
g8198 and P2_U7344 P2_U7343 P2_U7342 P2_U7341 ; P2_U4318
g8199 and P2_U7348 P2_U7347 P2_U7346 P2_U7345 ; P2_U4319
g8200 and P2_U7352 P2_U7351 P2_U7350 P2_U7349 ; P2_U4320
g8201 and P2_U7357 P2_U7356 P2_U7355 P2_U7354 ; P2_U4321
g8202 and P2_U7361 P2_U7360 P2_U7359 P2_U7358 ; P2_U4322
g8203 and P2_U7365 P2_U7364 P2_U7363 P2_U7362 ; P2_U4323
g8204 and P2_U7369 P2_U7368 P2_U7367 P2_U7366 ; P2_U4324
g8205 and P2_U7374 P2_U7373 P2_U7372 P2_U7371 ; P2_U4325
g8206 and P2_U7378 P2_U7377 P2_U7376 P2_U7375 ; P2_U4326
g8207 and P2_U7382 P2_U7381 P2_U7380 P2_U7379 ; P2_U4327
g8208 and P2_U7386 P2_U7385 P2_U7384 P2_U7383 ; P2_U4328
g8209 and P2_U7391 P2_U7390 P2_U7389 P2_U7388 ; P2_U4329
g8210 and P2_U7395 P2_U7394 P2_U7393 P2_U7392 ; P2_U4330
g8211 and P2_U7399 P2_U7398 P2_U7397 P2_U7396 ; P2_U4331
g8212 and P2_U7403 P2_U7402 P2_U7401 P2_U7400 ; P2_U4332
g8213 and P2_U7408 P2_U7407 P2_U7406 P2_U7405 ; P2_U4333
g8214 and P2_U7412 P2_U7411 P2_U7410 P2_U7409 ; P2_U4334
g8215 and P2_U7416 P2_U7415 P2_U7414 P2_U7413 ; P2_U4335
g8216 and P2_U7420 P2_U7419 P2_U7418 P2_U7417 ; P2_U4336
g8217 and P2_U2616 P2_U3300 ; P2_U4337
g8218 and P2_U7425 P2_U4413 ; P2_U4338
g8219 and P2_U4595 P2_U3300 ; P2_U4339
g8220 and P2_U7426 P2_U4414 P2_U7428 ; P2_U4340
g8221 and P2_U7430 P2_U3571 ; P2_U4341
g8222 and P2_U4413 P2_U4341 ; P2_U4342
g8223 and P2_U7869 P2_U7873 ; P2_U4343
g8224 and P2_U7436 P2_U7435 ; P2_U4344
g8225 and P2_U7440 P2_U7439 ; P2_U4345
g8226 and P2_U7442 P2_U7443 ; P2_U4346
g8227 and P2_U7445 P2_U7446 ; P2_U4347
g8228 and P2_U7448 P2_U7449 ; P2_U4348
g8229 and P2_U7451 P2_U7452 ; P2_U4349
g8230 and P2_U7454 P2_U7455 ; P2_U4350
g8231 and P2_U7457 P2_U7458 ; P2_U4351
g8232 and P2_U7460 P2_U7461 ; P2_U4352
g8233 and P2_U7463 P2_U7464 ; P2_U4353
g8234 and P2_U7466 P2_U7467 ; P2_U4354
g8235 and P2_U7469 P2_U7470 ; P2_U4355
g8236 and P2_U7472 P2_U7473 ; P2_U4356
g8237 and P2_U7475 P2_U7476 ; P2_U4357
g8238 and P2_U7478 P2_U7479 ; P2_U4358
g8239 and P2_U7481 P2_U7482 ; P2_U4359
g8240 and P2_U7484 P2_U7485 ; P2_U4360
g8241 and P2_U7487 P2_U7488 ; P2_U4361
g8242 and P2_U7490 P2_U7491 ; P2_U4362
g8243 and P2_U7493 P2_U7494 ; P2_U4363
g8244 and P2_U7496 P2_U7497 ; P2_U4364
g8245 and P2_U7499 P2_U7500 ; P2_U4365
g8246 and P2_U7502 P2_U7503 ; P2_U4366
g8247 and P2_U7505 P2_U7506 ; P2_U4367
g8248 and P2_U7510 P2_U7509 ; P2_U4368
g8249 and P2_U7514 P2_U7513 ; P2_U4369
g8250 and P2_U7518 P2_U7517 ; P2_U4370
g8251 and P2_U7522 P2_U7521 ; P2_U4371
g8252 and P2_U7526 P2_U7525 ; P2_U4372
g8253 and P2_U7530 P2_U7529 ; P2_U4373
g8254 and P2_U7532 P2_U7533 ; P2_U4374
g8255 and P2_U7536 P2_U7535 ; P2_U4375
g8256 and P2_U3255 P2_U6845 ; P2_U4376
g8257 and P2_U7863 P2_U3255 ; P2_U4377
g8258 and P2_U2356 P2_U7873 ; P2_U4378
g8259 and P2_U7579 P2_U7580 P2_U7578 ; P2_U4379
g8260 and P2_U7585 P2_U3269 ; P2_U4380
g8261 and P2_U2356 P2_U4595 ; P2_U4381
g8262 and P2_U3577 P2_U3539 P2_U4472 P2_U7587 P2_U7586 ; P2_U4382
g8263 and P2_U7579 P2_U4422 ; P2_U4383
g8264 and P2_U4383 P2_U7578 ; P2_U4384
g8265 and P2_U7580 P2_U4458 ; P2_U4385
g8266 and P2_U7590 P2_U7589 ; P2_U4386
g8267 and P2_U7736 P2_STATE2_REG_0__SCAN_IN ; P2_U4387
g8268 and P2_U3573 P2_U4458 P2_U4457 P2_U3549 ; P2_U4388
g8269 and P2_U7719 P2_U7718 ; P2_U4389
g8270 and P2_U7731 P2_U3536 ; P2_U4390
g8271 and P2_U7735 P2_U3536 ; P2_U4391
g8272 and P2_U7908 P2_U7907 ; P2_U4392
g8273 and P2_U8055 P2_U8054 ; P2_U4393
g8274 nand P2_U3872 P2_U5582 ; P2_U4394
g8275 and P2_U8079 P2_U8078 ; P2_U4395
g8276 and P2_U8092 P2_U8091 ; P2_U4396
g8277 and P2_U8120 P2_U8119 ; P2_U4397
g8278 and P2_U8126 P2_U8125 ; P2_U4398
g8279 and P2_U8132 P2_U8131 ; P2_U4399
g8280 nand P2_U2374 P2_U3291 ; P2_U4400
g8281 not BS16 ; P2_U4401
g8282 nand P2_U4462 P2_U4188 ; P2_U4402
g8283 nand P2_U3534 P2_U4462 ; P2_U4403
g8284 and P2_U8146 P2_U8145 ; P2_U4404
g8285 nand P2_U7006 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U4405
g8286 nand P2_U2513 P2_U3871 ; P2_U4406
g8287 not P2_R2219_U29 ; P2_U4407
g8288 not P2_R2219_U8 ; P2_U4408
g8289 not P2_U3553 ; P2_U4409
g8290 nand HOLD P2_U3265 ; P2_U4410
g8291 not P2_U3290 ; P2_U4411
g8292 not P2_U3571 ; P2_U4412
g8293 nand P2_U4337 P2_U4601 ; P2_U4413
g8294 nand P2_U2616 P2_U3300 P2_U7869 ; P2_U4414
g8295 nand P2_U2447 P2_U3279 ; P2_U4415
g8296 not P2_U3576 ; P2_U4416
g8297 not P2_U3283 ; P2_U4417
g8298 not P2_U3550 ; P2_U4418
g8299 not P2_U3536 ; P2_U4419
g8300 not P2_U3288 ; P2_U4420
g8301 not P2_U3539 ; P2_U4421
g8302 nand P2_U2376 P2_U3278 P2_U2450 ; P2_U4422
g8303 not P2_U3577 ; P2_U4423
g8304 not P2_U3282 ; P2_U4424
g8305 not P2_U3285 ; P2_U4425
g8306 not P2_U3549 ; P2_U4426
g8307 not P2_U3289 ; P2_U4427
g8308 not P2_U3286 ; P2_U4428
g8309 not P2_U3294 ; P2_U4429
g8310 not P2_U3313 ; P2_U4430
g8311 not P2_U3578 ; P2_U4431
g8312 not P2_U3254 ; P2_U4432
g8313 not P2_U3523 ; P2_U4433
g8314 not P2_U3524 ; P2_U4434
g8315 not P2_U3296 ; P2_U4435
g8316 not P2_U3522 ; P2_U4436
g8317 nand P2_U3875 P2_U2376 ; P2_U4437
g8318 not P2_U3547 ; P2_U4438
g8319 not P2_U3259 ; P2_U4439
g8320 not P2_U3543 ; P2_U4440
g8321 not P2_U3542 ; P2_U4441
g8322 not P2_U3538 ; P2_U4442
g8323 not P2_U3306 ; P2_U4443
g8324 not P2_LT_563_1260_U6 ; P2_U4444
g8325 nand P2_U4430 P2_U3302 ; P2_U4445
g8326 nand P2_U4461 P2_U3546 ; P2_U4446
g8327 nand P2_R2219_U7 P2_U2617 ; P2_U4447
g8328 nand P2_U2367 P2_U3290 ; P2_U4448
g8329 not P2_U3261 ; P2_U4449
g8330 not P2_U3260 ; P2_U4450
g8331 not P2_U3425 ; P2_U4451
g8332 nand P2_U4182 P2_U4438 ; P2_U4452
g8333 nand P2_U3718 P2_U4474 ; P2_U4453
g8334 nand P2_U3302 P2_U3270 P2_U3284 P2_STATE2_REG_1__SCAN_IN ; P2_U4454
g8335 nand P2_U3867 P2_U2448 ; P2_U4455
g8336 nand P2_U2446 P2_U2359 ; P2_U4456
g8337 nand P2_U2356 P2_U3280 ; P2_U4457
g8338 nand P2_U4378 P2_U7577 ; P2_U4458
g8339 not P2_U3575 ; P2_U4459
g8340 nand P2_U2438 P2_U3295 ; P2_U4460
g8341 not P2_U3534 ; P2_U4461
g8342 nand P2_U2374 P2_U6568 ; P2_U4462
g8343 nand P2_U4574 P2_U3266 ; P2_U4463
g8344 nand P2_U2448 P2_U3292 ; P2_U4464
g8345 nand P2_U4474 U211 ; P2_U4465
g8346 not P2_U3303 ; P2_U4466
g8347 not P2_U3540 ; P2_U4467
g8348 not P2_U3304 ; P2_U4468
g8349 not P2_U3305 ; P2_U4469
g8350 nand P2_U3876 P2_U2376 ; P2_U4470
g8351 not P2_U3573 ; P2_U4471
g8352 nand P2_U2376 P2_U7871 P2_U4416 ; P2_U4472
g8353 not P2_U3262 ; P2_U4473
g8354 not P2_U3301 ; P2_U4474
g8355 not P2_U3293 ; P2_U4475
g8356 not P2_U3281 ; P2_U4476
g8357 not P2_U3548 ; P2_U4477
g8358 nand P2_U4450 P2_REIP_REG_31__SCAN_IN ; P2_U4478
g8359 nand P2_U4449 P2_REIP_REG_30__SCAN_IN ; P2_U4479
g8360 nand P2_U3259 P2_ADDRESS_REG_29__SCAN_IN ; P2_U4480
g8361 nand P2_U4450 P2_REIP_REG_30__SCAN_IN ; P2_U4481
g8362 nand P2_U4449 P2_REIP_REG_29__SCAN_IN ; P2_U4482
g8363 nand P2_U3259 P2_ADDRESS_REG_28__SCAN_IN ; P2_U4483
g8364 nand P2_U4450 P2_REIP_REG_29__SCAN_IN ; P2_U4484
g8365 nand P2_U4449 P2_REIP_REG_28__SCAN_IN ; P2_U4485
g8366 nand P2_U3259 P2_ADDRESS_REG_27__SCAN_IN ; P2_U4486
g8367 nand P2_U4450 P2_REIP_REG_28__SCAN_IN ; P2_U4487
g8368 nand P2_U4449 P2_REIP_REG_27__SCAN_IN ; P2_U4488
g8369 nand P2_U3259 P2_ADDRESS_REG_26__SCAN_IN ; P2_U4489
g8370 nand P2_U4450 P2_REIP_REG_27__SCAN_IN ; P2_U4490
g8371 nand P2_U4449 P2_REIP_REG_26__SCAN_IN ; P2_U4491
g8372 nand P2_U3259 P2_ADDRESS_REG_25__SCAN_IN ; P2_U4492
g8373 nand P2_U4450 P2_REIP_REG_26__SCAN_IN ; P2_U4493
g8374 nand P2_U4449 P2_REIP_REG_25__SCAN_IN ; P2_U4494
g8375 nand P2_U3259 P2_ADDRESS_REG_24__SCAN_IN ; P2_U4495
g8376 nand P2_U4450 P2_REIP_REG_25__SCAN_IN ; P2_U4496
g8377 nand P2_U4449 P2_REIP_REG_24__SCAN_IN ; P2_U4497
g8378 nand P2_U3259 P2_ADDRESS_REG_23__SCAN_IN ; P2_U4498
g8379 nand P2_U4450 P2_REIP_REG_24__SCAN_IN ; P2_U4499
g8380 nand P2_U4449 P2_REIP_REG_23__SCAN_IN ; P2_U4500
g8381 nand P2_U3259 P2_ADDRESS_REG_22__SCAN_IN ; P2_U4501
g8382 nand P2_U4450 P2_REIP_REG_23__SCAN_IN ; P2_U4502
g8383 nand P2_U4449 P2_REIP_REG_22__SCAN_IN ; P2_U4503
g8384 nand P2_U3259 P2_ADDRESS_REG_21__SCAN_IN ; P2_U4504
g8385 nand P2_U4450 P2_REIP_REG_22__SCAN_IN ; P2_U4505
g8386 nand P2_U4449 P2_REIP_REG_21__SCAN_IN ; P2_U4506
g8387 nand P2_U3259 P2_ADDRESS_REG_20__SCAN_IN ; P2_U4507
g8388 nand P2_U4450 P2_REIP_REG_21__SCAN_IN ; P2_U4508
g8389 nand P2_U4449 P2_REIP_REG_20__SCAN_IN ; P2_U4509
g8390 nand P2_U3259 P2_ADDRESS_REG_19__SCAN_IN ; P2_U4510
g8391 nand P2_U4450 P2_REIP_REG_20__SCAN_IN ; P2_U4511
g8392 nand P2_U4449 P2_REIP_REG_19__SCAN_IN ; P2_U4512
g8393 nand P2_U3259 P2_ADDRESS_REG_18__SCAN_IN ; P2_U4513
g8394 nand P2_U4450 P2_REIP_REG_19__SCAN_IN ; P2_U4514
g8395 nand P2_U4449 P2_REIP_REG_18__SCAN_IN ; P2_U4515
g8396 nand P2_U3259 P2_ADDRESS_REG_17__SCAN_IN ; P2_U4516
g8397 nand P2_U4450 P2_REIP_REG_18__SCAN_IN ; P2_U4517
g8398 nand P2_U4449 P2_REIP_REG_17__SCAN_IN ; P2_U4518
g8399 nand P2_U3259 P2_ADDRESS_REG_16__SCAN_IN ; P2_U4519
g8400 nand P2_U4450 P2_REIP_REG_17__SCAN_IN ; P2_U4520
g8401 nand P2_U4449 P2_REIP_REG_16__SCAN_IN ; P2_U4521
g8402 nand P2_U3259 P2_ADDRESS_REG_15__SCAN_IN ; P2_U4522
g8403 nand P2_U4450 P2_REIP_REG_16__SCAN_IN ; P2_U4523
g8404 nand P2_U4449 P2_REIP_REG_15__SCAN_IN ; P2_U4524
g8405 nand P2_U3259 P2_ADDRESS_REG_14__SCAN_IN ; P2_U4525
g8406 nand P2_U4450 P2_REIP_REG_15__SCAN_IN ; P2_U4526
g8407 nand P2_U4449 P2_REIP_REG_14__SCAN_IN ; P2_U4527
g8408 nand P2_U3259 P2_ADDRESS_REG_13__SCAN_IN ; P2_U4528
g8409 nand P2_U4450 P2_REIP_REG_14__SCAN_IN ; P2_U4529
g8410 nand P2_U4449 P2_REIP_REG_13__SCAN_IN ; P2_U4530
g8411 nand P2_U3259 P2_ADDRESS_REG_12__SCAN_IN ; P2_U4531
g8412 nand P2_U4450 P2_REIP_REG_13__SCAN_IN ; P2_U4532
g8413 nand P2_U4449 P2_REIP_REG_12__SCAN_IN ; P2_U4533
g8414 nand P2_U3259 P2_ADDRESS_REG_11__SCAN_IN ; P2_U4534
g8415 nand P2_U4450 P2_REIP_REG_12__SCAN_IN ; P2_U4535
g8416 nand P2_U4449 P2_REIP_REG_11__SCAN_IN ; P2_U4536
g8417 nand P2_U3259 P2_ADDRESS_REG_10__SCAN_IN ; P2_U4537
g8418 nand P2_U4450 P2_REIP_REG_11__SCAN_IN ; P2_U4538
g8419 nand P2_U4449 P2_REIP_REG_10__SCAN_IN ; P2_U4539
g8420 nand P2_U3259 P2_ADDRESS_REG_9__SCAN_IN ; P2_U4540
g8421 nand P2_U4450 P2_REIP_REG_10__SCAN_IN ; P2_U4541
g8422 nand P2_U4449 P2_REIP_REG_9__SCAN_IN ; P2_U4542
g8423 nand P2_U3259 P2_ADDRESS_REG_8__SCAN_IN ; P2_U4543
g8424 nand P2_U4450 P2_REIP_REG_9__SCAN_IN ; P2_U4544
g8425 nand P2_U4449 P2_REIP_REG_8__SCAN_IN ; P2_U4545
g8426 nand P2_U3259 P2_ADDRESS_REG_7__SCAN_IN ; P2_U4546
g8427 nand P2_U4450 P2_REIP_REG_8__SCAN_IN ; P2_U4547
g8428 nand P2_U4449 P2_REIP_REG_7__SCAN_IN ; P2_U4548
g8429 nand P2_U3259 P2_ADDRESS_REG_6__SCAN_IN ; P2_U4549
g8430 nand P2_U4450 P2_REIP_REG_7__SCAN_IN ; P2_U4550
g8431 nand P2_U4449 P2_REIP_REG_6__SCAN_IN ; P2_U4551
g8432 nand P2_U3259 P2_ADDRESS_REG_5__SCAN_IN ; P2_U4552
g8433 nand P2_U4450 P2_REIP_REG_6__SCAN_IN ; P2_U4553
g8434 nand P2_U4449 P2_REIP_REG_5__SCAN_IN ; P2_U4554
g8435 nand P2_U3259 P2_ADDRESS_REG_4__SCAN_IN ; P2_U4555
g8436 nand P2_U4450 P2_REIP_REG_5__SCAN_IN ; P2_U4556
g8437 nand P2_U4449 P2_REIP_REG_4__SCAN_IN ; P2_U4557
g8438 nand P2_U3259 P2_ADDRESS_REG_3__SCAN_IN ; P2_U4558
g8439 nand P2_U4450 P2_REIP_REG_4__SCAN_IN ; P2_U4559
g8440 nand P2_U4449 P2_REIP_REG_3__SCAN_IN ; P2_U4560
g8441 nand P2_U3259 P2_ADDRESS_REG_2__SCAN_IN ; P2_U4561
g8442 nand P2_U4450 P2_REIP_REG_3__SCAN_IN ; P2_U4562
g8443 nand P2_U4449 P2_REIP_REG_2__SCAN_IN ; P2_U4563
g8444 nand P2_U3259 P2_ADDRESS_REG_1__SCAN_IN ; P2_U4564
g8445 nand P2_U4450 P2_REIP_REG_2__SCAN_IN ; P2_U4565
g8446 nand P2_U4449 P2_REIP_REG_1__SCAN_IN ; P2_U4566
g8447 nand P2_U3259 P2_ADDRESS_REG_0__SCAN_IN ; P2_U4567
g8448 not P2_U3267 ; P2_U4568
g8449 nand P2_U4568 P2_U3265 ; P2_U4569
g8450 nand NA P2_U4473 ; P2_U4570
g8451 not P2_U3268 ; P2_U4571
g8452 nand P2_U4571 P2_U3265 ; P2_U4572
g8453 nand P2_U4392 P2_U7891 ; P2_U4573
g8454 not P2_U3263 ; P2_U4574
g8455 nand HOLD P2_U3256 P2_U4574 ; P2_U4575
g8456 nand P2_U3268 U211 P2_STATE_REG_1__SCAN_IN ; P2_U4576
g8457 nand P2_U4576 P2_U4575 ; P2_U4577
g8458 nand P2_U4570 P2_U4577 P2_STATE_REG_0__SCAN_IN ; P2_U4578
g8459 nand P2_U4573 P2_STATE_REG_2__SCAN_IN ; P2_U4579
g8460 nand P2_U4410 P2_STATE_REG_0__SCAN_IN ; P2_U4580
g8461 nand P2_U4580 P2_STATE_REG_2__SCAN_IN ; P2_U4581
g8462 nand P2_U7910 P2_U7909 P2_U7892 ; P2_U4582
g8463 nand U211 P2_U4439 ; P2_U4583
g8464 nand P2_U3692 P2_U7893 ; P2_U4584
g8465 nand P2_U3267 P2_STATE_REG_2__SCAN_IN ; P2_U4585
g8466 nand NA P2_U3266 ; P2_U4586
g8467 nand P2_U4586 P2_U4585 ; P2_U4587
g8468 nand P2_U4587 P2_U3258 ; P2_U4588
g8469 nand P2_U4401 P2_U3263 ; P2_U4589
g8470 not P2_U3277 ; P2_U4590
g8471 nand P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U4591
g8472 not P2_U3274 ; P2_U4592
g8473 not P2_U3275 ; P2_U4593
g8474 nand P2_U3258 P2_STATE_REG_2__SCAN_IN ; P2_U4594
g8475 nand P2_U3262 P2_U4594 ; P2_U4595
g8476 not P2_U3527 ; P2_U4596
g8477 nand P2_U3294 P2_U3286 ; P2_U4597
g8478 nand P2_U4597 P2_U3265 ; P2_U4598
g8479 nand P2_U2359 P2_U3527 ; P2_U4599
g8480 not P2_U3291 ; P2_U4600
g8481 not P2_U3295 ; P2_U4601
g8482 nand P2_U4424 P2_U3253 ; P2_U4602
g8483 nand P2_U3524 P2_U4602 ; P2_U4603
g8484 nand P2_U3523 P2_U3522 ; P2_U4604
g8485 nand P2_R2243_U8 P2_U4428 ; P2_U4605
g8486 nand P2_U4417 P2_U3287 ; P2_U4606
g8487 nand P2_U4606 P2_U4605 ; P2_U4607
g8488 nand P2_U4420 P2_U4607 ; P2_U4608
g8489 nand P2_U4603 P2_U3520 ; P2_U4609
g8490 not P2_U3257 ; P2_U4610
g8491 nand P2_U4428 P2_U3292 ; P2_U4611
g8492 nand P2_GTE_370_U6 P2_U4417 ; P2_U4612
g8493 nand P2_U4612 P2_U4611 ; P2_U4613
g8494 nand P2_U4420 P2_U4613 ; P2_U4614
g8495 or P2_FLUSH_REG_SCAN_IN P2_MORE_REG_SCAN_IN ; P2_U4615
g8496 not P2_U3298 ; P2_U4616
g8497 nand P2_U4616 P2_U3269 ; P2_U4617
g8498 nand P2_U3711 P2_U4425 ; P2_U4618
g8499 nand P2_U8057 P2_U8056 P2_U3715 ; P2_U4619
g8500 not P2_U3299 ; P2_U4620
g8501 nand P2_U4474 P2_U3265 ; P2_U4621
g8502 nand P2_U3284 P2_STATEBS16_REG_SCAN_IN ; P2_U4622
g8503 nand P2_U4622 P2_U4621 ; P2_U4623
g8504 nand P2_U4623 P2_STATE2_REG_1__SCAN_IN ; P2_U4624
g8505 nand P2_U3299 P2_STATE2_REG_2__SCAN_IN ; P2_U4625
g8506 nand P2_U4619 P2_U4465 ; P2_U4626
g8507 nand P2_U3717 P2_U4620 ; P2_U4627
g8508 nand P2_U4626 P2_STATE2_REG_1__SCAN_IN ; P2_U4628
g8509 nand P2_U2374 P2_U4619 ; P2_U4629
g8510 nand P2_U3719 P2_U4469 ; P2_U4630
g8511 nand P2_U4619 P2_U4464 ; P2_U4631
g8512 nand P2_U2374 P2_U3298 ; P2_U4632
g8513 not P2_U3337 ; P2_U4633
g8514 not P2_U3351 ; P2_U4634
g8515 not P2_U3352 ; P2_U4635
g8516 not P2_U3319 ; P2_U4636
g8517 not P2_U3318 ; P2_U4637
g8518 not P2_U3378 ; P2_U4638
g8519 nand P2_R2182_U76 P2_U3318 ; P2_U4639
g8520 not P2_U3426 ; P2_U4640
g8521 not P2_U3320 ; P2_U4641
g8522 not P2_U3311 ; P2_U4642
g8523 not P2_U3312 ; P2_U4643
g8524 not P2_U3424 ; P2_U4644
g8525 not P2_U3376 ; P2_U4645
g8526 nand P2_U3311 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U4646
g8527 not P2_U3428 ; P2_U4647
g8528 not P2_U3349 ; P2_U4648
g8529 not P2_U3335 ; P2_U4649
g8530 not P2_U3243 ; P2_U4650
g8531 nand P2_U2440 P2_U2444 ; P2_U4651
g8532 not P2_U3325 ; P2_U4652
g8533 not P2_U3570 ; P2_U4653
g8534 not P2_U3326 ; P2_U4654
g8535 nand P2_U3270 P2_STATE2_REG_1__SCAN_IN ; P2_U4655
g8536 nand P2_U4655 P2_U3304 P2_U3305 ; P2_U4656
g8537 nand P2_U4637 P2_U2462 ; P2_U4657
g8538 nand P2_U2468 P2_U2362 ; P2_U4658
g8539 nand P2_U4445 P2_U4658 ; P2_U4659
g8540 nand P2_U4652 P2_U4659 ; P2_U4660
g8541 nand P2_U4654 P2_STATE2_REG_2__SCAN_IN ; P2_U4661
g8542 nand P2_U3312 P2_STATE2_REG_3__SCAN_IN ; P2_U4662
g8543 nand P2_U4660 P2_U3722 ; P2_U4663
g8544 nand P2_U2468 P2_U2398 ; P2_U4664
g8545 nand P2_U4445 P2_U4664 ; P2_U4665
g8546 nand P2_U4665 P2_U3325 ; P2_U4666
g8547 nand P2_U3326 P2_STATE2_REG_2__SCAN_IN ; P2_U4667
g8548 nand P2_U4667 P2_U4666 ; P2_U4668
g8549 nand P2_U2425 P2_U4643 ; P2_U4669
g8550 nand P2_U2422 P2_U2463 ; P2_U4670
g8551 nand P2_U2421 P2_U4641 ; P2_U4671
g8552 nand P2_U2406 P2_U4668 ; P2_U4672
g8553 nand P2_U4663 P2_INSTQUEUE_REG_15__7__SCAN_IN ; P2_U4673
g8554 nand P2_U2426 P2_U4643 ; P2_U4674
g8555 nand P2_U2420 P2_U2463 ; P2_U4675
g8556 nand P2_U2419 P2_U4641 ; P2_U4676
g8557 nand P2_U2405 P2_U4668 ; P2_U4677
g8558 nand P2_U4663 P2_INSTQUEUE_REG_15__6__SCAN_IN ; P2_U4678
g8559 nand P2_U2429 P2_U4643 ; P2_U4679
g8560 nand P2_U2418 P2_U2463 ; P2_U4680
g8561 nand P2_U2417 P2_U4641 ; P2_U4681
g8562 nand P2_U2404 P2_U4668 ; P2_U4682
g8563 nand P2_U4663 P2_INSTQUEUE_REG_15__5__SCAN_IN ; P2_U4683
g8564 nand P2_U2424 P2_U4643 ; P2_U4684
g8565 nand P2_U2416 P2_U2463 ; P2_U4685
g8566 nand P2_U2415 P2_U4641 ; P2_U4686
g8567 nand P2_U2403 P2_U4668 ; P2_U4687
g8568 nand P2_U4663 P2_INSTQUEUE_REG_15__4__SCAN_IN ; P2_U4688
g8569 nand P2_U2423 P2_U4643 ; P2_U4689
g8570 nand P2_U2414 P2_U2463 ; P2_U4690
g8571 nand P2_U2413 P2_U4641 ; P2_U4691
g8572 nand P2_U2402 P2_U4668 ; P2_U4692
g8573 nand P2_U4663 P2_INSTQUEUE_REG_15__3__SCAN_IN ; P2_U4693
g8574 nand P2_U2432 P2_U4643 ; P2_U4694
g8575 nand P2_U2412 P2_U2463 ; P2_U4695
g8576 nand P2_U2411 P2_U4641 ; P2_U4696
g8577 nand P2_U2401 P2_U4668 ; P2_U4697
g8578 nand P2_U4663 P2_INSTQUEUE_REG_15__2__SCAN_IN ; P2_U4698
g8579 nand P2_U2428 P2_U4643 ; P2_U4699
g8580 nand P2_U2410 P2_U2463 ; P2_U4700
g8581 nand P2_U2409 P2_U4641 ; P2_U4701
g8582 nand P2_U2400 P2_U4668 ; P2_U4702
g8583 nand P2_U4663 P2_INSTQUEUE_REG_15__1__SCAN_IN ; P2_U4703
g8584 nand P2_U2431 P2_U4643 ; P2_U4704
g8585 nand P2_U2408 P2_U2463 ; P2_U4705
g8586 nand P2_U2407 P2_U4641 ; P2_U4706
g8587 nand P2_U2399 P2_U4668 ; P2_U4707
g8588 nand P2_U4663 P2_INSTQUEUE_REG_15__0__SCAN_IN ; P2_U4708
g8589 not P2_U3338 ; P2_U4709
g8590 not P2_U3339 ; P2_U4710
g8591 not P2_U3336 ; P2_U4711
g8592 not P2_U3245 ; P2_U4712
g8593 not P2_U3569 ; P2_U4713
g8594 not P2_U3340 ; P2_U4714
g8595 nand P2_U4633 P2_U2462 ; P2_U4715
g8596 nand P2_U2471 P2_U2362 ; P2_U4716
g8597 nand P2_U4445 P2_U4716 ; P2_U4717
g8598 nand P2_U4717 P2_U3245 ; P2_U4718
g8599 nand P2_U4714 P2_STATE2_REG_2__SCAN_IN ; P2_U4719
g8600 nand P2_U3336 P2_STATE2_REG_3__SCAN_IN ; P2_U4720
g8601 nand P2_U4718 P2_U3731 ; P2_U4721
g8602 nand P2_U2471 P2_U2398 ; P2_U4722
g8603 nand P2_U4445 P2_U4722 ; P2_U4723
g8604 nand P2_U4723 P2_U4712 ; P2_U4724
g8605 nand P2_U3340 P2_STATE2_REG_2__SCAN_IN ; P2_U4725
g8606 nand P2_U4725 P2_U4724 ; P2_U4726
g8607 nand P2_U4711 P2_U2425 ; P2_U4727
g8608 nand P2_U2469 P2_U2422 ; P2_U4728
g8609 nand P2_U4710 P2_U2421 ; P2_U4729
g8610 nand P2_U2406 P2_U4726 ; P2_U4730
g8611 nand P2_U4721 P2_INSTQUEUE_REG_14__7__SCAN_IN ; P2_U4731
g8612 nand P2_U4711 P2_U2426 ; P2_U4732
g8613 nand P2_U2469 P2_U2420 ; P2_U4733
g8614 nand P2_U4710 P2_U2419 ; P2_U4734
g8615 nand P2_U2405 P2_U4726 ; P2_U4735
g8616 nand P2_U4721 P2_INSTQUEUE_REG_14__6__SCAN_IN ; P2_U4736
g8617 nand P2_U4711 P2_U2429 ; P2_U4737
g8618 nand P2_U2469 P2_U2418 ; P2_U4738
g8619 nand P2_U4710 P2_U2417 ; P2_U4739
g8620 nand P2_U2404 P2_U4726 ; P2_U4740
g8621 nand P2_U4721 P2_INSTQUEUE_REG_14__5__SCAN_IN ; P2_U4741
g8622 nand P2_U4711 P2_U2424 ; P2_U4742
g8623 nand P2_U2469 P2_U2416 ; P2_U4743
g8624 nand P2_U4710 P2_U2415 ; P2_U4744
g8625 nand P2_U2403 P2_U4726 ; P2_U4745
g8626 nand P2_U4721 P2_INSTQUEUE_REG_14__4__SCAN_IN ; P2_U4746
g8627 nand P2_U4711 P2_U2423 ; P2_U4747
g8628 nand P2_U2469 P2_U2414 ; P2_U4748
g8629 nand P2_U4710 P2_U2413 ; P2_U4749
g8630 nand P2_U2402 P2_U4726 ; P2_U4750
g8631 nand P2_U4721 P2_INSTQUEUE_REG_14__3__SCAN_IN ; P2_U4751
g8632 nand P2_U4711 P2_U2432 ; P2_U4752
g8633 nand P2_U2469 P2_U2412 ; P2_U4753
g8634 nand P2_U4710 P2_U2411 ; P2_U4754
g8635 nand P2_U2401 P2_U4726 ; P2_U4755
g8636 nand P2_U4721 P2_INSTQUEUE_REG_14__2__SCAN_IN ; P2_U4756
g8637 nand P2_U4711 P2_U2428 ; P2_U4757
g8638 nand P2_U2469 P2_U2410 ; P2_U4758
g8639 nand P2_U4710 P2_U2409 ; P2_U4759
g8640 nand P2_U2400 P2_U4726 ; P2_U4760
g8641 nand P2_U4721 P2_INSTQUEUE_REG_14__1__SCAN_IN ; P2_U4761
g8642 nand P2_U4711 P2_U2431 ; P2_U4762
g8643 nand P2_U2469 P2_U2408 ; P2_U4763
g8644 nand P2_U4710 P2_U2407 ; P2_U4764
g8645 nand P2_U2399 P2_U4726 ; P2_U4765
g8646 nand P2_U4721 P2_INSTQUEUE_REG_14__0__SCAN_IN ; P2_U4766
g8647 not P2_U3353 ; P2_U4767
g8648 not P2_U3354 ; P2_U4768
g8649 not P2_U3350 ; P2_U4769
g8650 nand P2_U2445 P2_U2440 ; P2_U4770
g8651 not P2_U3355 ; P2_U4771
g8652 not P2_U3568 ; P2_U4772
g8653 not P2_U3356 ; P2_U4773
g8654 nand P2_U4634 P2_U2462 ; P2_U4774
g8655 nand P2_U2474 P2_U2362 ; P2_U4775
g8656 nand P2_U4445 P2_U4775 ; P2_U4776
g8657 nand P2_U4771 P2_U4776 ; P2_U4777
g8658 nand P2_U4773 P2_STATE2_REG_2__SCAN_IN ; P2_U4778
g8659 nand P2_U3350 P2_STATE2_REG_3__SCAN_IN ; P2_U4779
g8660 nand P2_U4777 P2_U3740 ; P2_U4780
g8661 nand P2_U2474 P2_U2398 ; P2_U4781
g8662 nand P2_U4445 P2_U4781 ; P2_U4782
g8663 nand P2_U4782 P2_U3355 ; P2_U4783
g8664 nand P2_U3356 P2_STATE2_REG_2__SCAN_IN ; P2_U4784
g8665 nand P2_U4784 P2_U4783 ; P2_U4785
g8666 nand P2_U4769 P2_U2425 ; P2_U4786
g8667 nand P2_U2472 P2_U2422 ; P2_U4787
g8668 nand P2_U4768 P2_U2421 ; P2_U4788
g8669 nand P2_U2406 P2_U4785 ; P2_U4789
g8670 nand P2_U4780 P2_INSTQUEUE_REG_13__7__SCAN_IN ; P2_U4790
g8671 nand P2_U4769 P2_U2426 ; P2_U4791
g8672 nand P2_U2472 P2_U2420 ; P2_U4792
g8673 nand P2_U4768 P2_U2419 ; P2_U4793
g8674 nand P2_U2405 P2_U4785 ; P2_U4794
g8675 nand P2_U4780 P2_INSTQUEUE_REG_13__6__SCAN_IN ; P2_U4795
g8676 nand P2_U4769 P2_U2429 ; P2_U4796
g8677 nand P2_U2472 P2_U2418 ; P2_U4797
g8678 nand P2_U4768 P2_U2417 ; P2_U4798
g8679 nand P2_U2404 P2_U4785 ; P2_U4799
g8680 nand P2_U4780 P2_INSTQUEUE_REG_13__5__SCAN_IN ; P2_U4800
g8681 nand P2_U4769 P2_U2424 ; P2_U4801
g8682 nand P2_U2472 P2_U2416 ; P2_U4802
g8683 nand P2_U4768 P2_U2415 ; P2_U4803
g8684 nand P2_U2403 P2_U4785 ; P2_U4804
g8685 nand P2_U4780 P2_INSTQUEUE_REG_13__4__SCAN_IN ; P2_U4805
g8686 nand P2_U4769 P2_U2423 ; P2_U4806
g8687 nand P2_U2472 P2_U2414 ; P2_U4807
g8688 nand P2_U4768 P2_U2413 ; P2_U4808
g8689 nand P2_U2402 P2_U4785 ; P2_U4809
g8690 nand P2_U4780 P2_INSTQUEUE_REG_13__3__SCAN_IN ; P2_U4810
g8691 nand P2_U4769 P2_U2432 ; P2_U4811
g8692 nand P2_U2472 P2_U2412 ; P2_U4812
g8693 nand P2_U4768 P2_U2411 ; P2_U4813
g8694 nand P2_U2401 P2_U4785 ; P2_U4814
g8695 nand P2_U4780 P2_INSTQUEUE_REG_13__2__SCAN_IN ; P2_U4815
g8696 nand P2_U4769 P2_U2428 ; P2_U4816
g8697 nand P2_U2472 P2_U2410 ; P2_U4817
g8698 nand P2_U4768 P2_U2409 ; P2_U4818
g8699 nand P2_U2400 P2_U4785 ; P2_U4819
g8700 nand P2_U4780 P2_INSTQUEUE_REG_13__1__SCAN_IN ; P2_U4820
g8701 nand P2_U4769 P2_U2431 ; P2_U4821
g8702 nand P2_U2472 P2_U2408 ; P2_U4822
g8703 nand P2_U4768 P2_U2407 ; P2_U4823
g8704 nand P2_U2399 P2_U4785 ; P2_U4824
g8705 nand P2_U4780 P2_INSTQUEUE_REG_13__0__SCAN_IN ; P2_U4825
g8706 not P2_U3366 ; P2_U4826
g8707 not P2_U3365 ; P2_U4827
g8708 not P2_U3246 ; P2_U4828
g8709 not P2_U3567 ; P2_U4829
g8710 not P2_U3367 ; P2_U4830
g8711 nand P2_U2476 P2_U2462 ; P2_U4831
g8712 nand P2_U2480 P2_U2362 ; P2_U4832
g8713 nand P2_U4445 P2_U4832 ; P2_U4833
g8714 nand P2_U4833 P2_U3246 ; P2_U4834
g8715 nand P2_U4830 P2_STATE2_REG_2__SCAN_IN ; P2_U4835
g8716 nand P2_U3365 P2_STATE2_REG_3__SCAN_IN ; P2_U4836
g8717 nand P2_U4834 P2_U3749 ; P2_U4837
g8718 nand P2_U2480 P2_U2398 ; P2_U4838
g8719 nand P2_U4445 P2_U4838 ; P2_U4839
g8720 nand P2_U4839 P2_U4828 ; P2_U4840
g8721 nand P2_U3367 P2_STATE2_REG_2__SCAN_IN ; P2_U4841
g8722 nand P2_U4841 P2_U4840 ; P2_U4842
g8723 nand P2_U4827 P2_U2425 ; P2_U4843
g8724 nand P2_U2477 P2_U2422 ; P2_U4844
g8725 nand P2_U4826 P2_U2421 ; P2_U4845
g8726 nand P2_U2406 P2_U4842 ; P2_U4846
g8727 nand P2_U4837 P2_INSTQUEUE_REG_12__7__SCAN_IN ; P2_U4847
g8728 nand P2_U4827 P2_U2426 ; P2_U4848
g8729 nand P2_U2477 P2_U2420 ; P2_U4849
g8730 nand P2_U4826 P2_U2419 ; P2_U4850
g8731 nand P2_U2405 P2_U4842 ; P2_U4851
g8732 nand P2_U4837 P2_INSTQUEUE_REG_12__6__SCAN_IN ; P2_U4852
g8733 nand P2_U4827 P2_U2429 ; P2_U4853
g8734 nand P2_U2477 P2_U2418 ; P2_U4854
g8735 nand P2_U4826 P2_U2417 ; P2_U4855
g8736 nand P2_U2404 P2_U4842 ; P2_U4856
g8737 nand P2_U4837 P2_INSTQUEUE_REG_12__5__SCAN_IN ; P2_U4857
g8738 nand P2_U4827 P2_U2424 ; P2_U4858
g8739 nand P2_U2477 P2_U2416 ; P2_U4859
g8740 nand P2_U4826 P2_U2415 ; P2_U4860
g8741 nand P2_U2403 P2_U4842 ; P2_U4861
g8742 nand P2_U4837 P2_INSTQUEUE_REG_12__4__SCAN_IN ; P2_U4862
g8743 nand P2_U4827 P2_U2423 ; P2_U4863
g8744 nand P2_U2477 P2_U2414 ; P2_U4864
g8745 nand P2_U4826 P2_U2413 ; P2_U4865
g8746 nand P2_U2402 P2_U4842 ; P2_U4866
g8747 nand P2_U4837 P2_INSTQUEUE_REG_12__3__SCAN_IN ; P2_U4867
g8748 nand P2_U4827 P2_U2432 ; P2_U4868
g8749 nand P2_U2477 P2_U2412 ; P2_U4869
g8750 nand P2_U4826 P2_U2411 ; P2_U4870
g8751 nand P2_U2401 P2_U4842 ; P2_U4871
g8752 nand P2_U4837 P2_INSTQUEUE_REG_12__2__SCAN_IN ; P2_U4872
g8753 nand P2_U4827 P2_U2428 ; P2_U4873
g8754 nand P2_U2477 P2_U2410 ; P2_U4874
g8755 nand P2_U4826 P2_U2409 ; P2_U4875
g8756 nand P2_U2400 P2_U4842 ; P2_U4876
g8757 nand P2_U4837 P2_INSTQUEUE_REG_12__1__SCAN_IN ; P2_U4877
g8758 nand P2_U4827 P2_U2431 ; P2_U4878
g8759 nand P2_U2477 P2_U2408 ; P2_U4879
g8760 nand P2_U4826 P2_U2407 ; P2_U4880
g8761 nand P2_U2399 P2_U4842 ; P2_U4881
g8762 nand P2_U4837 P2_INSTQUEUE_REG_12__0__SCAN_IN ; P2_U4882
g8763 not P2_U3379 ; P2_U4883
g8764 not P2_U3377 ; P2_U4884
g8765 nand P2_U2442 P2_U2444 ; P2_U4885
g8766 not P2_U3380 ; P2_U4886
g8767 not P2_U3566 ; P2_U4887
g8768 not P2_U3381 ; P2_U4888
g8769 nand P2_U4638 P2_U4637 ; P2_U4889
g8770 nand P2_U2484 P2_U2362 ; P2_U4890
g8771 nand P2_U4445 P2_U4890 ; P2_U4891
g8772 nand P2_U4886 P2_U4891 ; P2_U4892
g8773 nand P2_U4888 P2_STATE2_REG_2__SCAN_IN ; P2_U4893
g8774 nand P2_U3377 P2_STATE2_REG_3__SCAN_IN ; P2_U4894
g8775 nand P2_U4892 P2_U3758 ; P2_U4895
g8776 nand P2_U2484 P2_U2398 ; P2_U4896
g8777 nand P2_U4445 P2_U4896 ; P2_U4897
g8778 nand P2_U4897 P2_U3380 ; P2_U4898
g8779 nand P2_U3381 P2_STATE2_REG_2__SCAN_IN ; P2_U4899
g8780 nand P2_U4899 P2_U4898 ; P2_U4900
g8781 nand P2_U4884 P2_U2425 ; P2_U4901
g8782 nand P2_U2482 P2_U2422 ; P2_U4902
g8783 nand P2_U4883 P2_U2421 ; P2_U4903
g8784 nand P2_U2406 P2_U4900 ; P2_U4904
g8785 nand P2_U4895 P2_INSTQUEUE_REG_11__7__SCAN_IN ; P2_U4905
g8786 nand P2_U4884 P2_U2426 ; P2_U4906
g8787 nand P2_U2482 P2_U2420 ; P2_U4907
g8788 nand P2_U4883 P2_U2419 ; P2_U4908
g8789 nand P2_U2405 P2_U4900 ; P2_U4909
g8790 nand P2_U4895 P2_INSTQUEUE_REG_11__6__SCAN_IN ; P2_U4910
g8791 nand P2_U4884 P2_U2429 ; P2_U4911
g8792 nand P2_U2482 P2_U2418 ; P2_U4912
g8793 nand P2_U4883 P2_U2417 ; P2_U4913
g8794 nand P2_U2404 P2_U4900 ; P2_U4914
g8795 nand P2_U4895 P2_INSTQUEUE_REG_11__5__SCAN_IN ; P2_U4915
g8796 nand P2_U4884 P2_U2424 ; P2_U4916
g8797 nand P2_U2482 P2_U2416 ; P2_U4917
g8798 nand P2_U4883 P2_U2415 ; P2_U4918
g8799 nand P2_U2403 P2_U4900 ; P2_U4919
g8800 nand P2_U4895 P2_INSTQUEUE_REG_11__4__SCAN_IN ; P2_U4920
g8801 nand P2_U4884 P2_U2423 ; P2_U4921
g8802 nand P2_U2482 P2_U2414 ; P2_U4922
g8803 nand P2_U4883 P2_U2413 ; P2_U4923
g8804 nand P2_U2402 P2_U4900 ; P2_U4924
g8805 nand P2_U4895 P2_INSTQUEUE_REG_11__3__SCAN_IN ; P2_U4925
g8806 nand P2_U4884 P2_U2432 ; P2_U4926
g8807 nand P2_U2482 P2_U2412 ; P2_U4927
g8808 nand P2_U4883 P2_U2411 ; P2_U4928
g8809 nand P2_U2401 P2_U4900 ; P2_U4929
g8810 nand P2_U4895 P2_INSTQUEUE_REG_11__2__SCAN_IN ; P2_U4930
g8811 nand P2_U4884 P2_U2428 ; P2_U4931
g8812 nand P2_U2482 P2_U2410 ; P2_U4932
g8813 nand P2_U4883 P2_U2409 ; P2_U4933
g8814 nand P2_U2400 P2_U4900 ; P2_U4934
g8815 nand P2_U4895 P2_INSTQUEUE_REG_11__1__SCAN_IN ; P2_U4935
g8816 nand P2_U4884 P2_U2431 ; P2_U4936
g8817 nand P2_U2482 P2_U2408 ; P2_U4937
g8818 nand P2_U4883 P2_U2407 ; P2_U4938
g8819 nand P2_U2399 P2_U4900 ; P2_U4939
g8820 nand P2_U4895 P2_INSTQUEUE_REG_11__0__SCAN_IN ; P2_U4940
g8821 not P2_U3391 ; P2_U4941
g8822 not P2_U3390 ; P2_U4942
g8823 not P2_U3247 ; P2_U4943
g8824 not P2_U3565 ; P2_U4944
g8825 not P2_U3392 ; P2_U4945
g8826 nand P2_U4638 P2_U4633 ; P2_U4946
g8827 nand P2_U2486 P2_U2362 ; P2_U4947
g8828 nand P2_U4445 P2_U4947 ; P2_U4948
g8829 nand P2_U4948 P2_U3247 ; P2_U4949
g8830 nand P2_U4945 P2_STATE2_REG_2__SCAN_IN ; P2_U4950
g8831 nand P2_U3390 P2_STATE2_REG_3__SCAN_IN ; P2_U4951
g8832 nand P2_U4949 P2_U3767 ; P2_U4952
g8833 nand P2_U2486 P2_U2398 ; P2_U4953
g8834 nand P2_U4445 P2_U4953 ; P2_U4954
g8835 nand P2_U4954 P2_U4943 ; P2_U4955
g8836 nand P2_U3392 P2_STATE2_REG_2__SCAN_IN ; P2_U4956
g8837 nand P2_U4956 P2_U4955 ; P2_U4957
g8838 nand P2_U4942 P2_U2425 ; P2_U4958
g8839 nand P2_U2485 P2_U2422 ; P2_U4959
g8840 nand P2_U4941 P2_U2421 ; P2_U4960
g8841 nand P2_U2406 P2_U4957 ; P2_U4961
g8842 nand P2_U4952 P2_INSTQUEUE_REG_10__7__SCAN_IN ; P2_U4962
g8843 nand P2_U4942 P2_U2426 ; P2_U4963
g8844 nand P2_U2485 P2_U2420 ; P2_U4964
g8845 nand P2_U4941 P2_U2419 ; P2_U4965
g8846 nand P2_U2405 P2_U4957 ; P2_U4966
g8847 nand P2_U4952 P2_INSTQUEUE_REG_10__6__SCAN_IN ; P2_U4967
g8848 nand P2_U4942 P2_U2429 ; P2_U4968
g8849 nand P2_U2485 P2_U2418 ; P2_U4969
g8850 nand P2_U4941 P2_U2417 ; P2_U4970
g8851 nand P2_U2404 P2_U4957 ; P2_U4971
g8852 nand P2_U4952 P2_INSTQUEUE_REG_10__5__SCAN_IN ; P2_U4972
g8853 nand P2_U4942 P2_U2424 ; P2_U4973
g8854 nand P2_U2485 P2_U2416 ; P2_U4974
g8855 nand P2_U4941 P2_U2415 ; P2_U4975
g8856 nand P2_U2403 P2_U4957 ; P2_U4976
g8857 nand P2_U4952 P2_INSTQUEUE_REG_10__4__SCAN_IN ; P2_U4977
g8858 nand P2_U4942 P2_U2423 ; P2_U4978
g8859 nand P2_U2485 P2_U2414 ; P2_U4979
g8860 nand P2_U4941 P2_U2413 ; P2_U4980
g8861 nand P2_U2402 P2_U4957 ; P2_U4981
g8862 nand P2_U4952 P2_INSTQUEUE_REG_10__3__SCAN_IN ; P2_U4982
g8863 nand P2_U4942 P2_U2432 ; P2_U4983
g8864 nand P2_U2485 P2_U2412 ; P2_U4984
g8865 nand P2_U4941 P2_U2411 ; P2_U4985
g8866 nand P2_U2401 P2_U4957 ; P2_U4986
g8867 nand P2_U4952 P2_INSTQUEUE_REG_10__2__SCAN_IN ; P2_U4987
g8868 nand P2_U4942 P2_U2428 ; P2_U4988
g8869 nand P2_U2485 P2_U2410 ; P2_U4989
g8870 nand P2_U4941 P2_U2409 ; P2_U4990
g8871 nand P2_U2400 P2_U4957 ; P2_U4991
g8872 nand P2_U4952 P2_INSTQUEUE_REG_10__1__SCAN_IN ; P2_U4992
g8873 nand P2_U4942 P2_U2431 ; P2_U4993
g8874 nand P2_U2485 P2_U2408 ; P2_U4994
g8875 nand P2_U4941 P2_U2407 ; P2_U4995
g8876 nand P2_U2399 P2_U4957 ; P2_U4996
g8877 nand P2_U4952 P2_INSTQUEUE_REG_10__0__SCAN_IN ; P2_U4997
g8878 not P2_U3402 ; P2_U4998
g8879 not P2_U3401 ; P2_U4999
g8880 nand P2_U2442 P2_U2445 ; P2_U5000
g8881 not P2_U3403 ; P2_U5001
g8882 not P2_U3564 ; P2_U5002
g8883 not P2_U3404 ; P2_U5003
g8884 nand P2_U4638 P2_U4634 ; P2_U5004
g8885 nand P2_U2488 P2_U2362 ; P2_U5005
g8886 nand P2_U4445 P2_U5005 ; P2_U5006
g8887 nand P2_U5001 P2_U5006 ; P2_U5007
g8888 nand P2_U5003 P2_STATE2_REG_2__SCAN_IN ; P2_U5008
g8889 nand P2_U3401 P2_STATE2_REG_3__SCAN_IN ; P2_U5009
g8890 nand P2_U5007 P2_U3776 ; P2_U5010
g8891 nand P2_U2488 P2_U2398 ; P2_U5011
g8892 nand P2_U4445 P2_U5011 ; P2_U5012
g8893 nand P2_U5012 P2_U3403 ; P2_U5013
g8894 nand P2_U3404 P2_STATE2_REG_2__SCAN_IN ; P2_U5014
g8895 nand P2_U5014 P2_U5013 ; P2_U5015
g8896 nand P2_U4999 P2_U2425 ; P2_U5016
g8897 nand P2_U2487 P2_U2422 ; P2_U5017
g8898 nand P2_U4998 P2_U2421 ; P2_U5018
g8899 nand P2_U2406 P2_U5015 ; P2_U5019
g8900 nand P2_U5010 P2_INSTQUEUE_REG_9__7__SCAN_IN ; P2_U5020
g8901 nand P2_U4999 P2_U2426 ; P2_U5021
g8902 nand P2_U2487 P2_U2420 ; P2_U5022
g8903 nand P2_U4998 P2_U2419 ; P2_U5023
g8904 nand P2_U2405 P2_U5015 ; P2_U5024
g8905 nand P2_U5010 P2_INSTQUEUE_REG_9__6__SCAN_IN ; P2_U5025
g8906 nand P2_U4999 P2_U2429 ; P2_U5026
g8907 nand P2_U2487 P2_U2418 ; P2_U5027
g8908 nand P2_U4998 P2_U2417 ; P2_U5028
g8909 nand P2_U2404 P2_U5015 ; P2_U5029
g8910 nand P2_U5010 P2_INSTQUEUE_REG_9__5__SCAN_IN ; P2_U5030
g8911 nand P2_U4999 P2_U2424 ; P2_U5031
g8912 nand P2_U2487 P2_U2416 ; P2_U5032
g8913 nand P2_U4998 P2_U2415 ; P2_U5033
g8914 nand P2_U2403 P2_U5015 ; P2_U5034
g8915 nand P2_U5010 P2_INSTQUEUE_REG_9__4__SCAN_IN ; P2_U5035
g8916 nand P2_U4999 P2_U2423 ; P2_U5036
g8917 nand P2_U2487 P2_U2414 ; P2_U5037
g8918 nand P2_U4998 P2_U2413 ; P2_U5038
g8919 nand P2_U2402 P2_U5015 ; P2_U5039
g8920 nand P2_U5010 P2_INSTQUEUE_REG_9__3__SCAN_IN ; P2_U5040
g8921 nand P2_U4999 P2_U2432 ; P2_U5041
g8922 nand P2_U2487 P2_U2412 ; P2_U5042
g8923 nand P2_U4998 P2_U2411 ; P2_U5043
g8924 nand P2_U2401 P2_U5015 ; P2_U5044
g8925 nand P2_U5010 P2_INSTQUEUE_REG_9__2__SCAN_IN ; P2_U5045
g8926 nand P2_U4999 P2_U2428 ; P2_U5046
g8927 nand P2_U2487 P2_U2410 ; P2_U5047
g8928 nand P2_U4998 P2_U2409 ; P2_U5048
g8929 nand P2_U2400 P2_U5015 ; P2_U5049
g8930 nand P2_U5010 P2_INSTQUEUE_REG_9__1__SCAN_IN ; P2_U5050
g8931 nand P2_U4999 P2_U2431 ; P2_U5051
g8932 nand P2_U2487 P2_U2408 ; P2_U5052
g8933 nand P2_U4998 P2_U2407 ; P2_U5053
g8934 nand P2_U2399 P2_U5015 ; P2_U5054
g8935 nand P2_U5010 P2_INSTQUEUE_REG_9__0__SCAN_IN ; P2_U5055
g8936 not P2_U3414 ; P2_U5056
g8937 not P2_U3413 ; P2_U5057
g8938 not P2_U3248 ; P2_U5058
g8939 not P2_U3563 ; P2_U5059
g8940 not P2_U3415 ; P2_U5060
g8941 nand P2_U4638 P2_U2476 ; P2_U5061
g8942 nand P2_U2490 P2_U2362 ; P2_U5062
g8943 nand P2_U4445 P2_U5062 ; P2_U5063
g8944 nand P2_U5063 P2_U3248 ; P2_U5064
g8945 nand P2_U5060 P2_STATE2_REG_2__SCAN_IN ; P2_U5065
g8946 nand P2_U3413 P2_STATE2_REG_3__SCAN_IN ; P2_U5066
g8947 nand P2_U5064 P2_U3785 ; P2_U5067
g8948 nand P2_U2490 P2_U2398 ; P2_U5068
g8949 nand P2_U4445 P2_U5068 ; P2_U5069
g8950 nand P2_U5069 P2_U5058 ; P2_U5070
g8951 nand P2_U3415 P2_STATE2_REG_2__SCAN_IN ; P2_U5071
g8952 nand P2_U5071 P2_U5070 ; P2_U5072
g8953 nand P2_U5057 P2_U2425 ; P2_U5073
g8954 nand P2_U2489 P2_U2422 ; P2_U5074
g8955 nand P2_U5056 P2_U2421 ; P2_U5075
g8956 nand P2_U2406 P2_U5072 ; P2_U5076
g8957 nand P2_U5067 P2_INSTQUEUE_REG_8__7__SCAN_IN ; P2_U5077
g8958 nand P2_U5057 P2_U2426 ; P2_U5078
g8959 nand P2_U2489 P2_U2420 ; P2_U5079
g8960 nand P2_U5056 P2_U2419 ; P2_U5080
g8961 nand P2_U2405 P2_U5072 ; P2_U5081
g8962 nand P2_U5067 P2_INSTQUEUE_REG_8__6__SCAN_IN ; P2_U5082
g8963 nand P2_U5057 P2_U2429 ; P2_U5083
g8964 nand P2_U2489 P2_U2418 ; P2_U5084
g8965 nand P2_U5056 P2_U2417 ; P2_U5085
g8966 nand P2_U2404 P2_U5072 ; P2_U5086
g8967 nand P2_U5067 P2_INSTQUEUE_REG_8__5__SCAN_IN ; P2_U5087
g8968 nand P2_U5057 P2_U2424 ; P2_U5088
g8969 nand P2_U2489 P2_U2416 ; P2_U5089
g8970 nand P2_U5056 P2_U2415 ; P2_U5090
g8971 nand P2_U2403 P2_U5072 ; P2_U5091
g8972 nand P2_U5067 P2_INSTQUEUE_REG_8__4__SCAN_IN ; P2_U5092
g8973 nand P2_U5057 P2_U2423 ; P2_U5093
g8974 nand P2_U2489 P2_U2414 ; P2_U5094
g8975 nand P2_U5056 P2_U2413 ; P2_U5095
g8976 nand P2_U2402 P2_U5072 ; P2_U5096
g8977 nand P2_U5067 P2_INSTQUEUE_REG_8__3__SCAN_IN ; P2_U5097
g8978 nand P2_U5057 P2_U2432 ; P2_U5098
g8979 nand P2_U2489 P2_U2412 ; P2_U5099
g8980 nand P2_U5056 P2_U2411 ; P2_U5100
g8981 nand P2_U2401 P2_U5072 ; P2_U5101
g8982 nand P2_U5067 P2_INSTQUEUE_REG_8__2__SCAN_IN ; P2_U5102
g8983 nand P2_U5057 P2_U2428 ; P2_U5103
g8984 nand P2_U2489 P2_U2410 ; P2_U5104
g8985 nand P2_U5056 P2_U2409 ; P2_U5105
g8986 nand P2_U2400 P2_U5072 ; P2_U5106
g8987 nand P2_U5067 P2_INSTQUEUE_REG_8__1__SCAN_IN ; P2_U5107
g8988 nand P2_U5057 P2_U2431 ; P2_U5108
g8989 nand P2_U2489 P2_U2408 ; P2_U5109
g8990 nand P2_U5056 P2_U2407 ; P2_U5110
g8991 nand P2_U2399 P2_U5072 ; P2_U5111
g8992 nand P2_U5067 P2_INSTQUEUE_REG_8__0__SCAN_IN ; P2_U5112
g8993 not P2_U3427 ; P2_U5113
g8994 nand P2_U2441 P2_U2444 ; P2_U5114
g8995 not P2_U3429 ; P2_U5115
g8996 not P2_U3562 ; P2_U5116
g8997 not P2_U3430 ; P2_U5117
g8998 nand P2_U2493 P2_U2362 ; P2_U5118
g8999 nand P2_U4445 P2_U5118 ; P2_U5119
g9000 nand P2_U5115 P2_U5119 ; P2_U5120
g9001 nand P2_U5117 P2_STATE2_REG_2__SCAN_IN ; P2_U5121
g9002 nand P2_U3424 P2_STATE2_REG_3__SCAN_IN ; P2_U5122
g9003 nand P2_U5120 P2_U3794 ; P2_U5123
g9004 nand P2_U2493 P2_U2398 ; P2_U5124
g9005 nand P2_U4445 P2_U5124 ; P2_U5125
g9006 nand P2_U5125 P2_U3429 ; P2_U5126
g9007 nand P2_U3430 P2_STATE2_REG_2__SCAN_IN ; P2_U5127
g9008 nand P2_U5127 P2_U5126 ; P2_U5128
g9009 nand P2_U4644 P2_U2425 ; P2_U5129
g9010 nand P2_U4451 P2_U2422 ; P2_U5130
g9011 nand P2_U5113 P2_U2421 ; P2_U5131
g9012 nand P2_U2406 P2_U5128 ; P2_U5132
g9013 nand P2_U5123 P2_INSTQUEUE_REG_7__7__SCAN_IN ; P2_U5133
g9014 nand P2_U4644 P2_U2426 ; P2_U5134
g9015 nand P2_U4451 P2_U2420 ; P2_U5135
g9016 nand P2_U5113 P2_U2419 ; P2_U5136
g9017 nand P2_U2405 P2_U5128 ; P2_U5137
g9018 nand P2_U5123 P2_INSTQUEUE_REG_7__6__SCAN_IN ; P2_U5138
g9019 nand P2_U4644 P2_U2429 ; P2_U5139
g9020 nand P2_U4451 P2_U2418 ; P2_U5140
g9021 nand P2_U5113 P2_U2417 ; P2_U5141
g9022 nand P2_U2404 P2_U5128 ; P2_U5142
g9023 nand P2_U5123 P2_INSTQUEUE_REG_7__5__SCAN_IN ; P2_U5143
g9024 nand P2_U4644 P2_U2424 ; P2_U5144
g9025 nand P2_U4451 P2_U2416 ; P2_U5145
g9026 nand P2_U5113 P2_U2415 ; P2_U5146
g9027 nand P2_U2403 P2_U5128 ; P2_U5147
g9028 nand P2_U5123 P2_INSTQUEUE_REG_7__4__SCAN_IN ; P2_U5148
g9029 nand P2_U4644 P2_U2423 ; P2_U5149
g9030 nand P2_U4451 P2_U2414 ; P2_U5150
g9031 nand P2_U5113 P2_U2413 ; P2_U5151
g9032 nand P2_U2402 P2_U5128 ; P2_U5152
g9033 nand P2_U5123 P2_INSTQUEUE_REG_7__3__SCAN_IN ; P2_U5153
g9034 nand P2_U4644 P2_U2432 ; P2_U5154
g9035 nand P2_U4451 P2_U2412 ; P2_U5155
g9036 nand P2_U5113 P2_U2411 ; P2_U5156
g9037 nand P2_U2401 P2_U5128 ; P2_U5157
g9038 nand P2_U5123 P2_INSTQUEUE_REG_7__2__SCAN_IN ; P2_U5158
g9039 nand P2_U4644 P2_U2428 ; P2_U5159
g9040 nand P2_U4451 P2_U2410 ; P2_U5160
g9041 nand P2_U5113 P2_U2409 ; P2_U5161
g9042 nand P2_U2400 P2_U5128 ; P2_U5162
g9043 nand P2_U5123 P2_INSTQUEUE_REG_7__1__SCAN_IN ; P2_U5163
g9044 nand P2_U4644 P2_U2431 ; P2_U5164
g9045 nand P2_U4451 P2_U2408 ; P2_U5165
g9046 nand P2_U5113 P2_U2407 ; P2_U5166
g9047 nand P2_U2399 P2_U5128 ; P2_U5167
g9048 nand P2_U5123 P2_INSTQUEUE_REG_7__0__SCAN_IN ; P2_U5168
g9049 not P2_U3440 ; P2_U5169
g9050 not P2_U3439 ; P2_U5170
g9051 not P2_U3249 ; P2_U5171
g9052 not P2_U3561 ; P2_U5172
g9053 not P2_U3441 ; P2_U5173
g9054 nand P2_U4633 P2_U2460 ; P2_U5174
g9055 nand P2_U2495 P2_U2362 ; P2_U5175
g9056 nand P2_U4445 P2_U5175 ; P2_U5176
g9057 nand P2_U5176 P2_U3249 ; P2_U5177
g9058 nand P2_U5173 P2_STATE2_REG_2__SCAN_IN ; P2_U5178
g9059 nand P2_U3439 P2_STATE2_REG_3__SCAN_IN ; P2_U5179
g9060 nand P2_U5177 P2_U3803 ; P2_U5180
g9061 nand P2_U2495 P2_U2398 ; P2_U5181
g9062 nand P2_U4445 P2_U5181 ; P2_U5182
g9063 nand P2_U5182 P2_U5171 ; P2_U5183
g9064 nand P2_U3441 P2_STATE2_REG_2__SCAN_IN ; P2_U5184
g9065 nand P2_U5184 P2_U5183 ; P2_U5185
g9066 nand P2_U5170 P2_U2425 ; P2_U5186
g9067 nand P2_U2494 P2_U2422 ; P2_U5187
g9068 nand P2_U5169 P2_U2421 ; P2_U5188
g9069 nand P2_U2406 P2_U5185 ; P2_U5189
g9070 nand P2_U5180 P2_INSTQUEUE_REG_6__7__SCAN_IN ; P2_U5190
g9071 nand P2_U5170 P2_U2426 ; P2_U5191
g9072 nand P2_U2494 P2_U2420 ; P2_U5192
g9073 nand P2_U5169 P2_U2419 ; P2_U5193
g9074 nand P2_U2405 P2_U5185 ; P2_U5194
g9075 nand P2_U5180 P2_INSTQUEUE_REG_6__6__SCAN_IN ; P2_U5195
g9076 nand P2_U5170 P2_U2429 ; P2_U5196
g9077 nand P2_U2494 P2_U2418 ; P2_U5197
g9078 nand P2_U5169 P2_U2417 ; P2_U5198
g9079 nand P2_U2404 P2_U5185 ; P2_U5199
g9080 nand P2_U5180 P2_INSTQUEUE_REG_6__5__SCAN_IN ; P2_U5200
g9081 nand P2_U5170 P2_U2424 ; P2_U5201
g9082 nand P2_U2494 P2_U2416 ; P2_U5202
g9083 nand P2_U5169 P2_U2415 ; P2_U5203
g9084 nand P2_U2403 P2_U5185 ; P2_U5204
g9085 nand P2_U5180 P2_INSTQUEUE_REG_6__4__SCAN_IN ; P2_U5205
g9086 nand P2_U5170 P2_U2423 ; P2_U5206
g9087 nand P2_U2494 P2_U2414 ; P2_U5207
g9088 nand P2_U5169 P2_U2413 ; P2_U5208
g9089 nand P2_U2402 P2_U5185 ; P2_U5209
g9090 nand P2_U5180 P2_INSTQUEUE_REG_6__3__SCAN_IN ; P2_U5210
g9091 nand P2_U5170 P2_U2432 ; P2_U5211
g9092 nand P2_U2494 P2_U2412 ; P2_U5212
g9093 nand P2_U5169 P2_U2411 ; P2_U5213
g9094 nand P2_U2401 P2_U5185 ; P2_U5214
g9095 nand P2_U5180 P2_INSTQUEUE_REG_6__2__SCAN_IN ; P2_U5215
g9096 nand P2_U5170 P2_U2428 ; P2_U5216
g9097 nand P2_U2494 P2_U2410 ; P2_U5217
g9098 nand P2_U5169 P2_U2409 ; P2_U5218
g9099 nand P2_U2400 P2_U5185 ; P2_U5219
g9100 nand P2_U5180 P2_INSTQUEUE_REG_6__1__SCAN_IN ; P2_U5220
g9101 nand P2_U5170 P2_U2431 ; P2_U5221
g9102 nand P2_U2494 P2_U2408 ; P2_U5222
g9103 nand P2_U5169 P2_U2407 ; P2_U5223
g9104 nand P2_U2399 P2_U5185 ; P2_U5224
g9105 nand P2_U5180 P2_INSTQUEUE_REG_6__0__SCAN_IN ; P2_U5225
g9106 not P2_U3451 ; P2_U5226
g9107 not P2_U3450 ; P2_U5227
g9108 nand P2_U2441 P2_U2445 ; P2_U5228
g9109 not P2_U3452 ; P2_U5229
g9110 not P2_U3560 ; P2_U5230
g9111 not P2_U3453 ; P2_U5231
g9112 nand P2_U4634 P2_U2460 ; P2_U5232
g9113 nand P2_U2497 P2_U2362 ; P2_U5233
g9114 nand P2_U4445 P2_U5233 ; P2_U5234
g9115 nand P2_U5229 P2_U5234 ; P2_U5235
g9116 nand P2_U5231 P2_STATE2_REG_2__SCAN_IN ; P2_U5236
g9117 nand P2_U3450 P2_STATE2_REG_3__SCAN_IN ; P2_U5237
g9118 nand P2_U5235 P2_U3812 ; P2_U5238
g9119 nand P2_U2497 P2_U2398 ; P2_U5239
g9120 nand P2_U4445 P2_U5239 ; P2_U5240
g9121 nand P2_U5240 P2_U3452 ; P2_U5241
g9122 nand P2_U3453 P2_STATE2_REG_2__SCAN_IN ; P2_U5242
g9123 nand P2_U5242 P2_U5241 ; P2_U5243
g9124 nand P2_U5227 P2_U2425 ; P2_U5244
g9125 nand P2_U2496 P2_U2422 ; P2_U5245
g9126 nand P2_U5226 P2_U2421 ; P2_U5246
g9127 nand P2_U2406 P2_U5243 ; P2_U5247
g9128 nand P2_U5238 P2_INSTQUEUE_REG_5__7__SCAN_IN ; P2_U5248
g9129 nand P2_U5227 P2_U2426 ; P2_U5249
g9130 nand P2_U2496 P2_U2420 ; P2_U5250
g9131 nand P2_U5226 P2_U2419 ; P2_U5251
g9132 nand P2_U2405 P2_U5243 ; P2_U5252
g9133 nand P2_U5238 P2_INSTQUEUE_REG_5__6__SCAN_IN ; P2_U5253
g9134 nand P2_U5227 P2_U2429 ; P2_U5254
g9135 nand P2_U2496 P2_U2418 ; P2_U5255
g9136 nand P2_U5226 P2_U2417 ; P2_U5256
g9137 nand P2_U2404 P2_U5243 ; P2_U5257
g9138 nand P2_U5238 P2_INSTQUEUE_REG_5__5__SCAN_IN ; P2_U5258
g9139 nand P2_U5227 P2_U2424 ; P2_U5259
g9140 nand P2_U2496 P2_U2416 ; P2_U5260
g9141 nand P2_U5226 P2_U2415 ; P2_U5261
g9142 nand P2_U2403 P2_U5243 ; P2_U5262
g9143 nand P2_U5238 P2_INSTQUEUE_REG_5__4__SCAN_IN ; P2_U5263
g9144 nand P2_U5227 P2_U2423 ; P2_U5264
g9145 nand P2_U2496 P2_U2414 ; P2_U5265
g9146 nand P2_U5226 P2_U2413 ; P2_U5266
g9147 nand P2_U2402 P2_U5243 ; P2_U5267
g9148 nand P2_U5238 P2_INSTQUEUE_REG_5__3__SCAN_IN ; P2_U5268
g9149 nand P2_U5227 P2_U2432 ; P2_U5269
g9150 nand P2_U2496 P2_U2412 ; P2_U5270
g9151 nand P2_U5226 P2_U2411 ; P2_U5271
g9152 nand P2_U2401 P2_U5243 ; P2_U5272
g9153 nand P2_U5238 P2_INSTQUEUE_REG_5__2__SCAN_IN ; P2_U5273
g9154 nand P2_U5227 P2_U2428 ; P2_U5274
g9155 nand P2_U2496 P2_U2410 ; P2_U5275
g9156 nand P2_U5226 P2_U2409 ; P2_U5276
g9157 nand P2_U2400 P2_U5243 ; P2_U5277
g9158 nand P2_U5238 P2_INSTQUEUE_REG_5__1__SCAN_IN ; P2_U5278
g9159 nand P2_U5227 P2_U2431 ; P2_U5279
g9160 nand P2_U2496 P2_U2408 ; P2_U5280
g9161 nand P2_U5226 P2_U2407 ; P2_U5281
g9162 nand P2_U2399 P2_U5243 ; P2_U5282
g9163 nand P2_U5238 P2_INSTQUEUE_REG_5__0__SCAN_IN ; P2_U5283
g9164 not P2_U3463 ; P2_U5284
g9165 not P2_U3462 ; P2_U5285
g9166 not P2_U3250 ; P2_U5286
g9167 not P2_U3559 ; P2_U5287
g9168 not P2_U3464 ; P2_U5288
g9169 nand P2_U2476 P2_U2460 ; P2_U5289
g9170 nand P2_U2499 P2_U2362 ; P2_U5290
g9171 nand P2_U4445 P2_U5290 ; P2_U5291
g9172 nand P2_U5291 P2_U3250 ; P2_U5292
g9173 nand P2_U5288 P2_STATE2_REG_2__SCAN_IN ; P2_U5293
g9174 nand P2_U3462 P2_STATE2_REG_3__SCAN_IN ; P2_U5294
g9175 nand P2_U5292 P2_U3821 ; P2_U5295
g9176 nand P2_U2499 P2_U2398 ; P2_U5296
g9177 nand P2_U4445 P2_U5296 ; P2_U5297
g9178 nand P2_U5297 P2_U5286 ; P2_U5298
g9179 nand P2_U3464 P2_STATE2_REG_2__SCAN_IN ; P2_U5299
g9180 nand P2_U5299 P2_U5298 ; P2_U5300
g9181 nand P2_U5285 P2_U2425 ; P2_U5301
g9182 nand P2_U2498 P2_U2422 ; P2_U5302
g9183 nand P2_U5284 P2_U2421 ; P2_U5303
g9184 nand P2_U2406 P2_U5300 ; P2_U5304
g9185 nand P2_U5295 P2_INSTQUEUE_REG_4__7__SCAN_IN ; P2_U5305
g9186 nand P2_U5285 P2_U2426 ; P2_U5306
g9187 nand P2_U2498 P2_U2420 ; P2_U5307
g9188 nand P2_U5284 P2_U2419 ; P2_U5308
g9189 nand P2_U2405 P2_U5300 ; P2_U5309
g9190 nand P2_U5295 P2_INSTQUEUE_REG_4__6__SCAN_IN ; P2_U5310
g9191 nand P2_U5285 P2_U2429 ; P2_U5311
g9192 nand P2_U2498 P2_U2418 ; P2_U5312
g9193 nand P2_U5284 P2_U2417 ; P2_U5313
g9194 nand P2_U2404 P2_U5300 ; P2_U5314
g9195 nand P2_U5295 P2_INSTQUEUE_REG_4__5__SCAN_IN ; P2_U5315
g9196 nand P2_U5285 P2_U2424 ; P2_U5316
g9197 nand P2_U2498 P2_U2416 ; P2_U5317
g9198 nand P2_U5284 P2_U2415 ; P2_U5318
g9199 nand P2_U2403 P2_U5300 ; P2_U5319
g9200 nand P2_U5295 P2_INSTQUEUE_REG_4__4__SCAN_IN ; P2_U5320
g9201 nand P2_U5285 P2_U2423 ; P2_U5321
g9202 nand P2_U2498 P2_U2414 ; P2_U5322
g9203 nand P2_U5284 P2_U2413 ; P2_U5323
g9204 nand P2_U2402 P2_U5300 ; P2_U5324
g9205 nand P2_U5295 P2_INSTQUEUE_REG_4__3__SCAN_IN ; P2_U5325
g9206 nand P2_U5285 P2_U2432 ; P2_U5326
g9207 nand P2_U2498 P2_U2412 ; P2_U5327
g9208 nand P2_U5284 P2_U2411 ; P2_U5328
g9209 nand P2_U2401 P2_U5300 ; P2_U5329
g9210 nand P2_U5295 P2_INSTQUEUE_REG_4__2__SCAN_IN ; P2_U5330
g9211 nand P2_U5285 P2_U2428 ; P2_U5331
g9212 nand P2_U2498 P2_U2410 ; P2_U5332
g9213 nand P2_U5284 P2_U2409 ; P2_U5333
g9214 nand P2_U2400 P2_U5300 ; P2_U5334
g9215 nand P2_U5295 P2_INSTQUEUE_REG_4__1__SCAN_IN ; P2_U5335
g9216 nand P2_U5285 P2_U2431 ; P2_U5336
g9217 nand P2_U2498 P2_U2408 ; P2_U5337
g9218 nand P2_U5284 P2_U2407 ; P2_U5338
g9219 nand P2_U2399 P2_U5300 ; P2_U5339
g9220 nand P2_U5295 P2_INSTQUEUE_REG_4__0__SCAN_IN ; P2_U5340
g9221 not P2_U3474 ; P2_U5341
g9222 not P2_U3473 ; P2_U5342
g9223 nand P2_U2443 P2_U2444 ; P2_U5343
g9224 not P2_U3475 ; P2_U5344
g9225 not P2_U3558 ; P2_U5345
g9226 not P2_U3476 ; P2_U5346
g9227 nand P2_U2501 P2_U4637 ; P2_U5347
g9228 nand P2_U2505 P2_U2362 ; P2_U5348
g9229 nand P2_U4445 P2_U5348 ; P2_U5349
g9230 nand P2_U5344 P2_U5349 ; P2_U5350
g9231 nand P2_U5346 P2_STATE2_REG_2__SCAN_IN ; P2_U5351
g9232 nand P2_U3473 P2_STATE2_REG_3__SCAN_IN ; P2_U5352
g9233 nand P2_U5350 P2_U3830 ; P2_U5353
g9234 nand P2_U2505 P2_U2398 ; P2_U5354
g9235 nand P2_U4445 P2_U5354 ; P2_U5355
g9236 nand P2_U5355 P2_U3475 ; P2_U5356
g9237 nand P2_U3476 P2_STATE2_REG_2__SCAN_IN ; P2_U5357
g9238 nand P2_U5357 P2_U5356 ; P2_U5358
g9239 nand P2_U5342 P2_U2425 ; P2_U5359
g9240 nand P2_U2502 P2_U2422 ; P2_U5360
g9241 nand P2_U5341 P2_U2421 ; P2_U5361
g9242 nand P2_U2406 P2_U5358 ; P2_U5362
g9243 nand P2_U5353 P2_INSTQUEUE_REG_3__7__SCAN_IN ; P2_U5363
g9244 nand P2_U5342 P2_U2426 ; P2_U5364
g9245 nand P2_U2502 P2_U2420 ; P2_U5365
g9246 nand P2_U5341 P2_U2419 ; P2_U5366
g9247 nand P2_U2405 P2_U5358 ; P2_U5367
g9248 nand P2_U5353 P2_INSTQUEUE_REG_3__6__SCAN_IN ; P2_U5368
g9249 nand P2_U5342 P2_U2429 ; P2_U5369
g9250 nand P2_U2502 P2_U2418 ; P2_U5370
g9251 nand P2_U5341 P2_U2417 ; P2_U5371
g9252 nand P2_U2404 P2_U5358 ; P2_U5372
g9253 nand P2_U5353 P2_INSTQUEUE_REG_3__5__SCAN_IN ; P2_U5373
g9254 nand P2_U5342 P2_U2424 ; P2_U5374
g9255 nand P2_U2502 P2_U2416 ; P2_U5375
g9256 nand P2_U5341 P2_U2415 ; P2_U5376
g9257 nand P2_U2403 P2_U5358 ; P2_U5377
g9258 nand P2_U5353 P2_INSTQUEUE_REG_3__4__SCAN_IN ; P2_U5378
g9259 nand P2_U5342 P2_U2423 ; P2_U5379
g9260 nand P2_U2502 P2_U2414 ; P2_U5380
g9261 nand P2_U5341 P2_U2413 ; P2_U5381
g9262 nand P2_U2402 P2_U5358 ; P2_U5382
g9263 nand P2_U5353 P2_INSTQUEUE_REG_3__3__SCAN_IN ; P2_U5383
g9264 nand P2_U5342 P2_U2432 ; P2_U5384
g9265 nand P2_U2502 P2_U2412 ; P2_U5385
g9266 nand P2_U5341 P2_U2411 ; P2_U5386
g9267 nand P2_U2401 P2_U5358 ; P2_U5387
g9268 nand P2_U5353 P2_INSTQUEUE_REG_3__2__SCAN_IN ; P2_U5388
g9269 nand P2_U5342 P2_U2428 ; P2_U5389
g9270 nand P2_U2502 P2_U2410 ; P2_U5390
g9271 nand P2_U5341 P2_U2409 ; P2_U5391
g9272 nand P2_U2400 P2_U5358 ; P2_U5392
g9273 nand P2_U5353 P2_INSTQUEUE_REG_3__1__SCAN_IN ; P2_U5393
g9274 nand P2_U5342 P2_U2431 ; P2_U5394
g9275 nand P2_U2502 P2_U2408 ; P2_U5395
g9276 nand P2_U5341 P2_U2407 ; P2_U5396
g9277 nand P2_U2399 P2_U5358 ; P2_U5397
g9278 nand P2_U5353 P2_INSTQUEUE_REG_3__0__SCAN_IN ; P2_U5398
g9279 not P2_U3486 ; P2_U5399
g9280 not P2_U3485 ; P2_U5400
g9281 not P2_U3251 ; P2_U5401
g9282 not P2_U3557 ; P2_U5402
g9283 not P2_U3487 ; P2_U5403
g9284 nand P2_U2501 P2_U4633 ; P2_U5404
g9285 nand P2_U2507 P2_U2362 ; P2_U5405
g9286 nand P2_U4445 P2_U5405 ; P2_U5406
g9287 nand P2_U5406 P2_U3251 ; P2_U5407
g9288 nand P2_U5403 P2_STATE2_REG_2__SCAN_IN ; P2_U5408
g9289 nand P2_U3485 P2_STATE2_REG_3__SCAN_IN ; P2_U5409
g9290 nand P2_U5407 P2_U3839 ; P2_U5410
g9291 nand P2_U2507 P2_U2398 ; P2_U5411
g9292 nand P2_U4445 P2_U5411 ; P2_U5412
g9293 nand P2_U5412 P2_U5401 ; P2_U5413
g9294 nand P2_U3487 P2_STATE2_REG_2__SCAN_IN ; P2_U5414
g9295 nand P2_U5414 P2_U5413 ; P2_U5415
g9296 nand P2_U5400 P2_U2425 ; P2_U5416
g9297 nand P2_U2506 P2_U2422 ; P2_U5417
g9298 nand P2_U5399 P2_U2421 ; P2_U5418
g9299 nand P2_U2406 P2_U5415 ; P2_U5419
g9300 nand P2_U5410 P2_INSTQUEUE_REG_2__7__SCAN_IN ; P2_U5420
g9301 nand P2_U5400 P2_U2426 ; P2_U5421
g9302 nand P2_U2506 P2_U2420 ; P2_U5422
g9303 nand P2_U5399 P2_U2419 ; P2_U5423
g9304 nand P2_U2405 P2_U5415 ; P2_U5424
g9305 nand P2_U5410 P2_INSTQUEUE_REG_2__6__SCAN_IN ; P2_U5425
g9306 nand P2_U5400 P2_U2429 ; P2_U5426
g9307 nand P2_U2506 P2_U2418 ; P2_U5427
g9308 nand P2_U5399 P2_U2417 ; P2_U5428
g9309 nand P2_U2404 P2_U5415 ; P2_U5429
g9310 nand P2_U5410 P2_INSTQUEUE_REG_2__5__SCAN_IN ; P2_U5430
g9311 nand P2_U5400 P2_U2424 ; P2_U5431
g9312 nand P2_U2506 P2_U2416 ; P2_U5432
g9313 nand P2_U5399 P2_U2415 ; P2_U5433
g9314 nand P2_U2403 P2_U5415 ; P2_U5434
g9315 nand P2_U5410 P2_INSTQUEUE_REG_2__4__SCAN_IN ; P2_U5435
g9316 nand P2_U5400 P2_U2423 ; P2_U5436
g9317 nand P2_U2506 P2_U2414 ; P2_U5437
g9318 nand P2_U5399 P2_U2413 ; P2_U5438
g9319 nand P2_U2402 P2_U5415 ; P2_U5439
g9320 nand P2_U5410 P2_INSTQUEUE_REG_2__3__SCAN_IN ; P2_U5440
g9321 nand P2_U5400 P2_U2432 ; P2_U5441
g9322 nand P2_U2506 P2_U2412 ; P2_U5442
g9323 nand P2_U5399 P2_U2411 ; P2_U5443
g9324 nand P2_U2401 P2_U5415 ; P2_U5444
g9325 nand P2_U5410 P2_INSTQUEUE_REG_2__2__SCAN_IN ; P2_U5445
g9326 nand P2_U5400 P2_U2428 ; P2_U5446
g9327 nand P2_U2506 P2_U2410 ; P2_U5447
g9328 nand P2_U5399 P2_U2409 ; P2_U5448
g9329 nand P2_U2400 P2_U5415 ; P2_U5449
g9330 nand P2_U5410 P2_INSTQUEUE_REG_2__1__SCAN_IN ; P2_U5450
g9331 nand P2_U5400 P2_U2431 ; P2_U5451
g9332 nand P2_U2506 P2_U2408 ; P2_U5452
g9333 nand P2_U5399 P2_U2407 ; P2_U5453
g9334 nand P2_U2399 P2_U5415 ; P2_U5454
g9335 nand P2_U5410 P2_INSTQUEUE_REG_2__0__SCAN_IN ; P2_U5455
g9336 not P2_U3497 ; P2_U5456
g9337 not P2_U3496 ; P2_U5457
g9338 nand P2_U2443 P2_U2445 ; P2_U5458
g9339 not P2_U3498 ; P2_U5459
g9340 not P2_U3556 ; P2_U5460
g9341 not P2_U3499 ; P2_U5461
g9342 nand P2_U2501 P2_U4634 ; P2_U5462
g9343 nand P2_U2509 P2_U2362 ; P2_U5463
g9344 nand P2_U4445 P2_U5463 ; P2_U5464
g9345 nand P2_U5459 P2_U5464 ; P2_U5465
g9346 nand P2_U5461 P2_STATE2_REG_2__SCAN_IN ; P2_U5466
g9347 nand P2_U3496 P2_STATE2_REG_3__SCAN_IN ; P2_U5467
g9348 nand P2_U5465 P2_U3848 ; P2_U5468
g9349 nand P2_U2509 P2_U2398 ; P2_U5469
g9350 nand P2_U4445 P2_U5469 ; P2_U5470
g9351 nand P2_U5470 P2_U3498 ; P2_U5471
g9352 nand P2_U3499 P2_STATE2_REG_2__SCAN_IN ; P2_U5472
g9353 nand P2_U5472 P2_U5471 ; P2_U5473
g9354 nand P2_U5457 P2_U2425 ; P2_U5474
g9355 nand P2_U2508 P2_U2422 ; P2_U5475
g9356 nand P2_U5456 P2_U2421 ; P2_U5476
g9357 nand P2_U2406 P2_U5473 ; P2_U5477
g9358 nand P2_U5468 P2_INSTQUEUE_REG_1__7__SCAN_IN ; P2_U5478
g9359 nand P2_U5457 P2_U2426 ; P2_U5479
g9360 nand P2_U2508 P2_U2420 ; P2_U5480
g9361 nand P2_U5456 P2_U2419 ; P2_U5481
g9362 nand P2_U2405 P2_U5473 ; P2_U5482
g9363 nand P2_U5468 P2_INSTQUEUE_REG_1__6__SCAN_IN ; P2_U5483
g9364 nand P2_U5457 P2_U2429 ; P2_U5484
g9365 nand P2_U2508 P2_U2418 ; P2_U5485
g9366 nand P2_U5456 P2_U2417 ; P2_U5486
g9367 nand P2_U2404 P2_U5473 ; P2_U5487
g9368 nand P2_U5468 P2_INSTQUEUE_REG_1__5__SCAN_IN ; P2_U5488
g9369 nand P2_U5457 P2_U2424 ; P2_U5489
g9370 nand P2_U2508 P2_U2416 ; P2_U5490
g9371 nand P2_U5456 P2_U2415 ; P2_U5491
g9372 nand P2_U2403 P2_U5473 ; P2_U5492
g9373 nand P2_U5468 P2_INSTQUEUE_REG_1__4__SCAN_IN ; P2_U5493
g9374 nand P2_U5457 P2_U2423 ; P2_U5494
g9375 nand P2_U2508 P2_U2414 ; P2_U5495
g9376 nand P2_U5456 P2_U2413 ; P2_U5496
g9377 nand P2_U2402 P2_U5473 ; P2_U5497
g9378 nand P2_U5468 P2_INSTQUEUE_REG_1__3__SCAN_IN ; P2_U5498
g9379 nand P2_U5457 P2_U2432 ; P2_U5499
g9380 nand P2_U2508 P2_U2412 ; P2_U5500
g9381 nand P2_U5456 P2_U2411 ; P2_U5501
g9382 nand P2_U2401 P2_U5473 ; P2_U5502
g9383 nand P2_U5468 P2_INSTQUEUE_REG_1__2__SCAN_IN ; P2_U5503
g9384 nand P2_U5457 P2_U2428 ; P2_U5504
g9385 nand P2_U2508 P2_U2410 ; P2_U5505
g9386 nand P2_U5456 P2_U2409 ; P2_U5506
g9387 nand P2_U2400 P2_U5473 ; P2_U5507
g9388 nand P2_U5468 P2_INSTQUEUE_REG_1__1__SCAN_IN ; P2_U5508
g9389 nand P2_U5457 P2_U2431 ; P2_U5509
g9390 nand P2_U2508 P2_U2408 ; P2_U5510
g9391 nand P2_U5456 P2_U2407 ; P2_U5511
g9392 nand P2_U2399 P2_U5473 ; P2_U5512
g9393 nand P2_U5468 P2_INSTQUEUE_REG_1__0__SCAN_IN ; P2_U5513
g9394 not P2_U3509 ; P2_U5514
g9395 not P2_U3508 ; P2_U5515
g9396 not P2_U3252 ; P2_U5516
g9397 not P2_U3555 ; P2_U5517
g9398 not P2_U3510 ; P2_U5518
g9399 nand P2_U2501 P2_U2476 ; P2_U5519
g9400 nand P2_U2511 P2_U2362 ; P2_U5520
g9401 nand P2_U4445 P2_U5520 ; P2_U5521
g9402 nand P2_U5521 P2_U3252 ; P2_U5522
g9403 nand P2_U5518 P2_STATE2_REG_2__SCAN_IN ; P2_U5523
g9404 nand P2_U3508 P2_STATE2_REG_3__SCAN_IN ; P2_U5524
g9405 nand P2_U5522 P2_U3857 ; P2_U5525
g9406 nand P2_U2511 P2_U2398 ; P2_U5526
g9407 nand P2_U4445 P2_U5526 ; P2_U5527
g9408 nand P2_U5527 P2_U5516 ; P2_U5528
g9409 nand P2_U3510 P2_STATE2_REG_2__SCAN_IN ; P2_U5529
g9410 nand P2_U5529 P2_U5528 ; P2_U5530
g9411 nand P2_U5515 P2_U2425 ; P2_U5531
g9412 nand P2_U2510 P2_U2422 ; P2_U5532
g9413 nand P2_U5514 P2_U2421 ; P2_U5533
g9414 nand P2_U2406 P2_U5530 ; P2_U5534
g9415 nand P2_U5525 P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U5535
g9416 nand P2_U5515 P2_U2426 ; P2_U5536
g9417 nand P2_U2510 P2_U2420 ; P2_U5537
g9418 nand P2_U5514 P2_U2419 ; P2_U5538
g9419 nand P2_U2405 P2_U5530 ; P2_U5539
g9420 nand P2_U5525 P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U5540
g9421 nand P2_U5515 P2_U2429 ; P2_U5541
g9422 nand P2_U2510 P2_U2418 ; P2_U5542
g9423 nand P2_U5514 P2_U2417 ; P2_U5543
g9424 nand P2_U2404 P2_U5530 ; P2_U5544
g9425 nand P2_U5525 P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U5545
g9426 nand P2_U5515 P2_U2424 ; P2_U5546
g9427 nand P2_U2510 P2_U2416 ; P2_U5547
g9428 nand P2_U5514 P2_U2415 ; P2_U5548
g9429 nand P2_U2403 P2_U5530 ; P2_U5549
g9430 nand P2_U5525 P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U5550
g9431 nand P2_U5515 P2_U2423 ; P2_U5551
g9432 nand P2_U2510 P2_U2414 ; P2_U5552
g9433 nand P2_U5514 P2_U2413 ; P2_U5553
g9434 nand P2_U2402 P2_U5530 ; P2_U5554
g9435 nand P2_U5525 P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U5555
g9436 nand P2_U5515 P2_U2432 ; P2_U5556
g9437 nand P2_U2510 P2_U2412 ; P2_U5557
g9438 nand P2_U5514 P2_U2411 ; P2_U5558
g9439 nand P2_U2401 P2_U5530 ; P2_U5559
g9440 nand P2_U5525 P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U5560
g9441 nand P2_U5515 P2_U2428 ; P2_U5561
g9442 nand P2_U2510 P2_U2410 ; P2_U5562
g9443 nand P2_U5514 P2_U2409 ; P2_U5563
g9444 nand P2_U2400 P2_U5530 ; P2_U5564
g9445 nand P2_U5525 P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U5565
g9446 nand P2_U5515 P2_U2431 ; P2_U5566
g9447 nand P2_U2510 P2_U2408 ; P2_U5567
g9448 nand P2_U5514 P2_U2407 ; P2_U5568
g9449 nand P2_U2399 P2_U5530 ; P2_U5569
g9450 nand P2_U5525 P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U5570
g9451 nand P2_U3279 P2_U7869 ; P2_U5571
g9452 not P2_U3574 ; P2_U5572
g9453 nand P2_U7863 P2_U2617 P2_U7861 ; P2_U5573
g9454 nand P2_U7895 P2_U3521 P2_U3255 P2_U3289 ; P2_U5574
g9455 nand P2_U2357 P2_U7871 ; P2_U5575
g9456 nand P2_U4417 P2_U3574 ; P2_U5576
g9457 nand P2_U4428 P2_U4424 ; P2_U5577
g9458 nand P2_U3524 P2_U5577 ; P2_U5578
g9459 nand P2_U5578 P2_U3265 P2_R2088_U6 ; P2_U5579
g9460 nand P2_U4436 P2_R2167_U6 ; P2_U5580
g9461 not P2_U4406 ; P2_U5581
g9462 nand P2_U2374 P2_U4406 ; P2_U5582
g9463 nand P2_U3284 P2_STATE2_REG_3__SCAN_IN ; P2_U5583
g9464 not P2_U4394 ; P2_U5584
g9465 nand P2_U4591 P2_U3276 ; P2_U5585
g9466 nand P2_U2617 P2_U3295 P2_U3878 ; P2_U5586
g9467 nand P2_U3295 P2_U3255 ; P2_U5587
g9468 nand P2_U7865 P2_U3278 ; P2_U5588
g9469 nand P2_U8075 P2_U8074 P2_U3879 ; P2_U5589
g9470 not P2_U3525 ; P2_U5590
g9471 nand P2_U7738 P2_U3278 ; P2_U5591
g9472 nand P2_U3521 P2_U5591 P2_U5573 P2_U5571 ; P2_U5592
g9473 nand P2_U4417 P2_U3574 ; P2_U5593
g9474 nand P2_U5592 P2_U2616 ; P2_U5594
g9475 nand P2_U3877 P2_U5594 ; P2_U5595
g9476 nand P2_U3295 P2_U7873 ; P2_U5596
g9477 nand P2_U3279 P2_U7871 ; P2_U5597
g9478 nand P2_U2617 P2_U3521 ; P2_U5598
g9479 nand P2_U4427 P2_U5598 ; P2_U5599
g9480 nand P2_U5597 P2_U3280 ; P2_U5600
g9481 nand P2_U2436 P2_U7884 ; P2_U5601
g9482 nand P2_U3527 P2_U3278 ; P2_U5602
g9483 nand P2_U2514 P2_U3288 ; P2_U5603
g9484 nand P2_U8077 P2_U8076 P2_U4470 ; P2_U5604
g9485 nand P2_U3296 P2_U3522 ; P2_U5605
g9486 nand P2_U3578 P2_U4437 ; P2_U5606
g9487 nand P2_U4395 P2_U5605 ; P2_U5607
g9488 nand P2_U3581 P2_U5606 ; P2_U5608
g9489 nand P2_R2147_U8 P2_U5604 ; P2_U5609
g9490 nand P2_R2099_U95 P2_U5603 ; P2_U5610
g9491 nand P2_U3884 P2_U5610 ; P2_U5611
g9492 nand P2_R2182_U76 P2_U4469 ; P2_U5612
g9493 nand P2_U4466 P2_U5611 ; P2_U5613
g9494 nand P2_U5613 P2_U5612 ; P2_U5614
g9495 nand P2_U4591 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U5615
g9496 not P2_U3530 ; P2_U5616
g9497 nand P2_R2147_U9 P2_U5604 ; P2_U5617
g9498 nand P2_R2099_U96 P2_U5603 ; P2_U5618
g9499 nand P2_U3885 P2_U5618 ; P2_U5619
g9500 nand P2_U3598 P2_U3597 P2_STATE2_REG_1__SCAN_IN ; P2_U5620
g9501 nand P2_R2182_U40 P2_U4469 ; P2_U5621
g9502 nand P2_U4466 P2_U5619 ; P2_U5622
g9503 nand P2_U5621 P2_U5622 P2_U5620 ; P2_U5623
g9504 nand P2_U2449 P2_U7861 P2_U4429 ; P2_U5624
g9505 nand P2_U7882 P2_U5624 ; P2_U5625
g9506 nand P2_U3887 P2_U8097 ; P2_U5626
g9507 nand P2_R2147_U4 P2_U5604 ; P2_U5627
g9508 nand P2_R2099_U5 P2_U5603 ; P2_U5628
g9509 nand P2_U3888 P2_U5628 ; P2_U5629
g9510 nand P2_U8090 P2_U3597 P2_STATE2_REG_1__SCAN_IN ; P2_U5630
g9511 nand P2_R2182_U68 P2_U4469 ; P2_U5631
g9512 nand P2_U4466 P2_U5629 ; P2_U5632
g9513 nand P2_U5631 P2_U5632 P2_U5630 ; P2_U5633
g9514 nand P2_U3889 P2_U8097 ; P2_U5634
g9515 nand P2_U5604 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U5635
g9516 nand P2_R2099_U94 P2_U5603 ; P2_U5636
g9517 nand P2_U3890 P2_U5636 ; P2_U5637
g9518 nand P2_R2182_U69 P2_U4469 ; P2_U5638
g9519 nand P2_U4466 P2_U5637 ; P2_U5639
g9520 nand P2_U8087 P2_STATE2_REG_1__SCAN_IN ; P2_U5640
g9521 nand P2_U5639 P2_U5638 P2_U5640 ; P2_U5641
g9522 nand P2_U2448 P2_R2243_U8 P2_STATE2_REG_0__SCAN_IN ; P2_U5642
g9523 not P2_U3533 ; P2_U5643
g9524 nand P2_U4445 P2_U3303 ; P2_U5644
g9525 nand P2_U4636 P2_U3579 ; P2_U5645
g9526 nand P2_U3426 P2_U5645 ; P2_U5646
g9527 nand P2_U3427 P2_U5646 ; P2_U5647
g9528 nand P2_U2398 P2_U5647 ; P2_U5648
g9529 nand P2_R2182_U76 P2_U5644 ; P2_U5649
g9530 nand P2_R2096_U75 P2_STATE2_REG_3__SCAN_IN ; P2_U5650
g9531 nand P2_U3891 P2_U5648 ; P2_U5651
g9532 nand P2_U2398 P2_U8109 ; P2_U5652
g9533 nand P2_R2182_U40 P2_U5644 ; P2_U5653
g9534 nand P2_R2096_U77 P2_STATE2_REG_3__SCAN_IN ; P2_U5654
g9535 nand P2_U3892 P2_U5652 ; P2_U5655
g9536 nand P2_U3338 P2_U3353 ; P2_U5656
g9537 nand P2_U2398 P2_U5656 ; P2_U5657
g9538 nand P2_R2182_U68 P2_U5644 ; P2_U5658
g9539 nand P2_R2096_U51 P2_STATE2_REG_3__SCAN_IN ; P2_U5659
g9540 nand P2_U3893 P2_U5657 ; P2_U5660
g9541 nand P2_U3313 P2_U3303 ; P2_U5661
g9542 nand P2_R2182_U69 P2_U5661 ; P2_U5662
g9543 nand P2_R2096_U68 P2_STATE2_REG_3__SCAN_IN ; P2_U5663
g9544 nand P2_U5662 P2_U5663 P2_U4464 ; P2_U5664
g9545 nand P2_U2616 P2_U3292 ; P2_U5665
g9546 nand P2_GTE_370_U6 P2_U4417 ; P2_U5666
g9547 nand P2_U5666 P2_U5665 ; P2_U5667
g9548 nand P2_U8122 P2_U8121 P2_U3265 P2_R2088_U6 ; P2_U5668
g9549 nand P2_U4420 P2_U5667 ; P2_U5669
g9550 nand P2_U2512 P2_U3894 P2_U4397 P2_U5669 ; P2_U5670
g9551 nand P2_U2374 P2_U5670 ; P2_U5671
g9552 nand P2_U4461 P2_U3284 ; P2_U5672
g9553 not P2_U3535 ; P2_U5673
g9554 nand P2_U4427 P2_U4420 ; P2_U5674
g9555 nand P2_U3895 P2_U2514 ; P2_U5675
g9556 nand P2_U4417 P2_U4424 ; P2_U5676
g9557 nand P2_U5676 P2_U4470 P2_U4437 P2_U3524 ; P2_U5677
g9558 nand P2_U4428 P2_U4424 ; P2_U5678
g9559 nand P2_U3296 P2_U5678 P2_U3523 ; P2_U5679
g9560 nand P2_U2390 P2_R2096_U68 ; P2_U5680
g9561 nand P2_U2389 P2_R2099_U94 ; P2_U5681
g9562 nand P2_R2027_U5 P2_U2388 ; P2_U5682
g9563 nand P2_ADD_394_U4 P2_U2386 ; P2_U5683
g9564 nand P2_R2278_U83 P2_U2385 ; P2_U5684
g9565 nand P2_ADD_371_1212_U68 P2_U2384 ; P2_U5685
g9566 nand P2_U2381 P2_REIP_REG_0__SCAN_IN ; P2_U5686
g9567 nand P2_U5673 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_U5687
g9568 nand P2_U2390 P2_R2096_U51 ; P2_U5688
g9569 nand P2_U2389 P2_R2099_U5 ; P2_U5689
g9570 nand P2_R2027_U85 P2_U2388 ; P2_U5690
g9571 nand P2_ADD_394_U85 P2_U2386 ; P2_U5691
g9572 nand P2_R2278_U6 P2_U2385 ; P2_U5692
g9573 nand P2_ADD_371_1212_U25 P2_U2384 ; P2_U5693
g9574 nand P2_U2381 P2_REIP_REG_1__SCAN_IN ; P2_U5694
g9575 nand P2_U5673 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_U5695
g9576 nand P2_U2390 P2_R2096_U77 ; P2_U5696
g9577 nand P2_U2389 P2_R2099_U96 ; P2_U5697
g9578 nand P2_R2027_U74 P2_U2388 ; P2_U5698
g9579 nand P2_ADD_394_U5 P2_U2386 ; P2_U5699
g9580 nand P2_R2278_U92 P2_U2385 ; P2_U5700
g9581 nand P2_ADD_371_1212_U79 P2_U2384 ; P2_U5701
g9582 nand P2_U2381 P2_REIP_REG_2__SCAN_IN ; P2_U5702
g9583 nand P2_U5673 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_U5703
g9584 nand P2_U2390 P2_R2096_U75 ; P2_U5704
g9585 nand P2_U2389 P2_R2099_U95 ; P2_U5705
g9586 nand P2_R2027_U71 P2_U2388 ; P2_U5706
g9587 nand P2_ADD_394_U95 P2_U2386 ; P2_U5707
g9588 nand P2_R2278_U90 P2_U2385 ; P2_U5708
g9589 nand P2_ADD_371_1212_U84 P2_U2384 ; P2_U5709
g9590 nand P2_U2381 P2_REIP_REG_3__SCAN_IN ; P2_U5710
g9591 nand P2_U5673 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_U5711
g9592 nand P2_R2096_U74 P2_U2390 ; P2_U5712
g9593 nand P2_R2099_U98 P2_U2389 ; P2_U5713
g9594 nand P2_R2027_U70 P2_U2388 ; P2_U5714
g9595 nand P2_ADD_394_U76 P2_U2386 ; P2_U5715
g9596 nand P2_R2278_U89 P2_U2385 ; P2_U5716
g9597 nand P2_ADD_371_1212_U80 P2_U2384 ; P2_U5717
g9598 nand P2_U2381 P2_REIP_REG_4__SCAN_IN ; P2_U5718
g9599 nand P2_U5673 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_U5719
g9600 nand P2_R2096_U73 P2_U2390 ; P2_U5720
g9601 nand P2_R2099_U71 P2_U2389 ; P2_U5721
g9602 nand P2_R2027_U69 P2_U2388 ; P2_U5722
g9603 nand P2_ADD_394_U79 P2_U2386 ; P2_U5723
g9604 nand P2_R2278_U88 P2_U2385 ; P2_U5724
g9605 nand P2_ADD_371_1212_U81 P2_U2384 ; P2_U5725
g9606 nand P2_U2381 P2_REIP_REG_5__SCAN_IN ; P2_U5726
g9607 nand P2_U5673 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_U5727
g9608 nand P2_R2096_U72 P2_U2390 ; P2_U5728
g9609 nand P2_R2099_U70 P2_U2389 ; P2_U5729
g9610 nand P2_R2027_U68 P2_U2388 ; P2_U5730
g9611 nand P2_ADD_394_U63 P2_U2386 ; P2_U5731
g9612 nand P2_R2278_U87 P2_U2385 ; P2_U5732
g9613 nand P2_ADD_371_1212_U78 P2_U2384 ; P2_U5733
g9614 nand P2_U2381 P2_REIP_REG_6__SCAN_IN ; P2_U5734
g9615 nand P2_U5673 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_U5735
g9616 nand P2_R2096_U71 P2_U2390 ; P2_U5736
g9617 nand P2_R2099_U69 P2_U2389 ; P2_U5737
g9618 nand P2_R2027_U67 P2_U2388 ; P2_U5738
g9619 nand P2_ADD_394_U89 P2_U2386 ; P2_U5739
g9620 nand P2_R2278_U86 P2_U2385 ; P2_U5740
g9621 nand P2_ADD_371_1212_U85 P2_U2384 ; P2_U5741
g9622 nand P2_U2381 P2_REIP_REG_7__SCAN_IN ; P2_U5742
g9623 nand P2_U5673 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_U5743
g9624 nand P2_R2096_U70 P2_U2390 ; P2_U5744
g9625 nand P2_R2099_U68 P2_U2389 ; P2_U5745
g9626 nand P2_R2027_U66 P2_U2388 ; P2_U5746
g9627 nand P2_ADD_394_U80 P2_U2386 ; P2_U5747
g9628 nand P2_R2278_U85 P2_U2385 ; P2_U5748
g9629 nand P2_ADD_371_1212_U82 P2_U2384 ; P2_U5749
g9630 nand P2_U2381 P2_REIP_REG_8__SCAN_IN ; P2_U5750
g9631 nand P2_U5673 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_U5751
g9632 nand P2_R2096_U69 P2_U2390 ; P2_U5752
g9633 nand P2_R2099_U67 P2_U2389 ; P2_U5753
g9634 nand P2_R2027_U65 P2_U2388 ; P2_U5754
g9635 nand P2_ADD_394_U70 P2_U2386 ; P2_U5755
g9636 nand P2_R2278_U84 P2_U2385 ; P2_U5756
g9637 nand P2_ADD_371_1212_U118 P2_U2384 ; P2_U5757
g9638 nand P2_U2381 P2_REIP_REG_9__SCAN_IN ; P2_U5758
g9639 nand P2_U5673 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_U5759
g9640 nand P2_R2096_U97 P2_U2390 ; P2_U5760
g9641 nand P2_R2099_U93 P2_U2389 ; P2_U5761
g9642 nand P2_R2027_U95 P2_U2388 ; P2_U5762
g9643 nand P2_ADD_394_U83 P2_U2386 ; P2_U5763
g9644 nand P2_R2278_U112 P2_U2385 ; P2_U5764
g9645 nand P2_ADD_371_1212_U13 P2_U2384 ; P2_U5765
g9646 nand P2_U2381 P2_REIP_REG_10__SCAN_IN ; P2_U5766
g9647 nand P2_U5673 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_U5767
g9648 nand P2_R2096_U96 P2_U2390 ; P2_U5768
g9649 nand P2_R2099_U92 P2_U2389 ; P2_U5769
g9650 nand P2_R2027_U94 P2_U2388 ; P2_U5770
g9651 nand P2_ADD_394_U73 P2_U2386 ; P2_U5771
g9652 nand P2_R2278_U111 P2_U2385 ; P2_U5772
g9653 nand P2_ADD_371_1212_U14 P2_U2384 ; P2_U5773
g9654 nand P2_U2381 P2_REIP_REG_11__SCAN_IN ; P2_U5774
g9655 nand P2_U5673 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_U5775
g9656 nand P2_R2096_U95 P2_U2390 ; P2_U5776
g9657 nand P2_R2099_U91 P2_U2389 ; P2_U5777
g9658 nand P2_R2027_U93 P2_U2388 ; P2_U5778
g9659 nand P2_ADD_394_U88 P2_U2386 ; P2_U5779
g9660 nand P2_R2278_U110 P2_U2385 ; P2_U5780
g9661 nand P2_ADD_371_1212_U76 P2_U2384 ; P2_U5781
g9662 nand P2_U2381 P2_REIP_REG_12__SCAN_IN ; P2_U5782
g9663 nand P2_U5673 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_U5783
g9664 nand P2_R2096_U94 P2_U2390 ; P2_U5784
g9665 nand P2_R2099_U90 P2_U2389 ; P2_U5785
g9666 nand P2_R2027_U92 P2_U2388 ; P2_U5786
g9667 nand P2_ADD_394_U69 P2_U2386 ; P2_U5787
g9668 nand P2_R2278_U109 P2_U2385 ; P2_U5788
g9669 nand P2_ADD_371_1212_U15 P2_U2384 ; P2_U5789
g9670 nand P2_U2381 P2_REIP_REG_13__SCAN_IN ; P2_U5790
g9671 nand P2_U5673 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_U5791
g9672 nand P2_R2096_U93 P2_U2390 ; P2_U5792
g9673 nand P2_R2099_U89 P2_U2389 ; P2_U5793
g9674 nand P2_R2027_U91 P2_U2388 ; P2_U5794
g9675 nand P2_ADD_394_U78 P2_U2386 ; P2_U5795
g9676 nand P2_R2278_U108 P2_U2385 ; P2_U5796
g9677 nand P2_ADD_371_1212_U16 P2_U2384 ; P2_U5797
g9678 nand P2_U2381 P2_REIP_REG_14__SCAN_IN ; P2_U5798
g9679 nand P2_U5673 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_U5799
g9680 nand P2_R2096_U92 P2_U2390 ; P2_U5800
g9681 nand P2_R2099_U88 P2_U2389 ; P2_U5801
g9682 nand P2_R2027_U90 P2_U2388 ; P2_U5802
g9683 nand P2_ADD_394_U75 P2_U2386 ; P2_U5803
g9684 nand P2_R2278_U107 P2_U2385 ; P2_U5804
g9685 nand P2_ADD_371_1212_U73 P2_U2384 ; P2_U5805
g9686 nand P2_U2381 P2_REIP_REG_15__SCAN_IN ; P2_U5806
g9687 nand P2_U5673 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_U5807
g9688 nand P2_R2096_U91 P2_U2390 ; P2_U5808
g9689 nand P2_R2099_U87 P2_U2389 ; P2_U5809
g9690 nand P2_R2027_U89 P2_U2388 ; P2_U5810
g9691 nand P2_ADD_394_U91 P2_U2386 ; P2_U5811
g9692 nand P2_R2278_U106 P2_U2385 ; P2_U5812
g9693 nand P2_ADD_371_1212_U17 P2_U2384 ; P2_U5813
g9694 nand P2_U2381 P2_REIP_REG_16__SCAN_IN ; P2_U5814
g9695 nand P2_U5673 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_U5815
g9696 nand P2_R2096_U90 P2_U2390 ; P2_U5816
g9697 nand P2_R2099_U86 P2_U2389 ; P2_U5817
g9698 nand P2_R2027_U88 P2_U2388 ; P2_U5818
g9699 nand P2_ADD_394_U67 P2_U2386 ; P2_U5819
g9700 nand P2_R2278_U105 P2_U2385 ; P2_U5820
g9701 nand P2_ADD_371_1212_U71 P2_U2384 ; P2_U5821
g9702 nand P2_U2381 P2_REIP_REG_17__SCAN_IN ; P2_U5822
g9703 nand P2_U5673 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_U5823
g9704 nand P2_R2096_U89 P2_U2390 ; P2_U5824
g9705 nand P2_R2099_U85 P2_U2389 ; P2_U5825
g9706 nand P2_R2027_U87 P2_U2388 ; P2_U5826
g9707 nand P2_ADD_394_U72 P2_U2386 ; P2_U5827
g9708 nand P2_R2278_U104 P2_U2385 ; P2_U5828
g9709 nand P2_ADD_371_1212_U72 P2_U2384 ; P2_U5829
g9710 nand P2_U2381 P2_REIP_REG_18__SCAN_IN ; P2_U5830
g9711 nand P2_U5673 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_U5831
g9712 nand P2_R2096_U88 P2_U2390 ; P2_U5832
g9713 nand P2_R2099_U84 P2_U2389 ; P2_U5833
g9714 nand P2_R2027_U86 P2_U2388 ; P2_U5834
g9715 nand P2_ADD_394_U82 P2_U2386 ; P2_U5835
g9716 nand P2_R2278_U103 P2_U2385 ; P2_U5836
g9717 nand P2_ADD_371_1212_U18 P2_U2384 ; P2_U5837
g9718 nand P2_U2381 P2_REIP_REG_19__SCAN_IN ; P2_U5838
g9719 nand P2_U5673 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_U5839
g9720 nand P2_R2096_U87 P2_U2390 ; P2_U5840
g9721 nand P2_R2099_U83 P2_U2389 ; P2_U5841
g9722 nand P2_R2027_U84 P2_U2388 ; P2_U5842
g9723 nand P2_ADD_394_U68 P2_U2386 ; P2_U5843
g9724 nand P2_R2278_U102 P2_U2385 ; P2_U5844
g9725 nand P2_ADD_371_1212_U19 P2_U2384 ; P2_U5845
g9726 nand P2_U2381 P2_REIP_REG_20__SCAN_IN ; P2_U5846
g9727 nand P2_U5673 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_U5847
g9728 nand P2_R2096_U86 P2_U2390 ; P2_U5848
g9729 nand P2_R2099_U82 P2_U2389 ; P2_U5849
g9730 nand P2_R2027_U83 P2_U2388 ; P2_U5850
g9731 nand P2_ADD_394_U87 P2_U2386 ; P2_U5851
g9732 nand P2_R2278_U101 P2_U2385 ; P2_U5852
g9733 nand P2_ADD_371_1212_U75 P2_U2384 ; P2_U5853
g9734 nand P2_U2381 P2_REIP_REG_21__SCAN_IN ; P2_U5854
g9735 nand P2_U5673 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_U5855
g9736 nand P2_R2096_U85 P2_U2390 ; P2_U5856
g9737 nand P2_R2099_U81 P2_U2389 ; P2_U5857
g9738 nand P2_R2027_U82 P2_U2388 ; P2_U5858
g9739 nand P2_ADD_394_U71 P2_U2386 ; P2_U5859
g9740 nand P2_R2278_U100 P2_U2385 ; P2_U5860
g9741 nand P2_ADD_371_1212_U20 P2_U2384 ; P2_U5861
g9742 nand P2_U2381 P2_REIP_REG_22__SCAN_IN ; P2_U5862
g9743 nand P2_U5673 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_U5863
g9744 nand P2_R2096_U84 P2_U2390 ; P2_U5864
g9745 nand P2_R2099_U80 P2_U2389 ; P2_U5865
g9746 nand P2_R2027_U81 P2_U2388 ; P2_U5866
g9747 nand P2_ADD_394_U81 P2_U2386 ; P2_U5867
g9748 nand P2_R2278_U99 P2_U2385 ; P2_U5868
g9749 nand P2_ADD_371_1212_U21 P2_U2384 ; P2_U5869
g9750 nand P2_U2381 P2_REIP_REG_23__SCAN_IN ; P2_U5870
g9751 nand P2_U5673 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_U5871
g9752 nand P2_R2096_U83 P2_U2390 ; P2_U5872
g9753 nand P2_R2099_U79 P2_U2389 ; P2_U5873
g9754 nand P2_R2027_U80 P2_U2388 ; P2_U5874
g9755 nand P2_ADD_394_U66 P2_U2386 ; P2_U5875
g9756 nand P2_R2278_U98 P2_U2385 ; P2_U5876
g9757 nand P2_ADD_371_1212_U70 P2_U2384 ; P2_U5877
g9758 nand P2_U2381 P2_REIP_REG_24__SCAN_IN ; P2_U5878
g9759 nand P2_U5673 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_U5879
g9760 nand P2_R2096_U82 P2_U2390 ; P2_U5880
g9761 nand P2_R2099_U78 P2_U2389 ; P2_U5881
g9762 nand P2_R2027_U79 P2_U2388 ; P2_U5882
g9763 nand P2_ADD_394_U90 P2_U2386 ; P2_U5883
g9764 nand P2_R2278_U97 P2_U2385 ; P2_U5884
g9765 nand P2_ADD_371_1212_U77 P2_U2384 ; P2_U5885
g9766 nand P2_U2381 P2_REIP_REG_25__SCAN_IN ; P2_U5886
g9767 nand P2_U5673 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_U5887
g9768 nand P2_R2096_U81 P2_U2390 ; P2_U5888
g9769 nand P2_R2099_U77 P2_U2389 ; P2_U5889
g9770 nand P2_R2027_U78 P2_U2388 ; P2_U5890
g9771 nand P2_ADD_394_U74 P2_U2386 ; P2_U5891
g9772 nand P2_R2278_U96 P2_U2385 ; P2_U5892
g9773 nand P2_ADD_371_1212_U22 P2_U2384 ; P2_U5893
g9774 nand P2_U2381 P2_REIP_REG_26__SCAN_IN ; P2_U5894
g9775 nand P2_U5673 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_U5895
g9776 nand P2_R2096_U80 P2_U2390 ; P2_U5896
g9777 nand P2_R2099_U76 P2_U2389 ; P2_U5897
g9778 nand P2_R2027_U77 P2_U2388 ; P2_U5898
g9779 nand P2_ADD_394_U77 P2_U2386 ; P2_U5899
g9780 nand P2_R2278_U95 P2_U2385 ; P2_U5900
g9781 nand P2_ADD_371_1212_U74 P2_U2384 ; P2_U5901
g9782 nand P2_U2381 P2_REIP_REG_27__SCAN_IN ; P2_U5902
g9783 nand P2_U5673 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_U5903
g9784 nand P2_R2096_U79 P2_U2390 ; P2_U5904
g9785 nand P2_R2099_U75 P2_U2389 ; P2_U5905
g9786 nand P2_R2027_U76 P2_U2388 ; P2_U5906
g9787 nand P2_ADD_394_U86 P2_U2386 ; P2_U5907
g9788 nand P2_R2278_U94 P2_U2385 ; P2_U5908
g9789 nand P2_ADD_371_1212_U23 P2_U2384 ; P2_U5909
g9790 nand P2_U2381 P2_REIP_REG_28__SCAN_IN ; P2_U5910
g9791 nand P2_U5673 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_U5911
g9792 nand P2_R2096_U78 P2_U2390 ; P2_U5912
g9793 nand P2_R2099_U74 P2_U2389 ; P2_U5913
g9794 nand P2_R2027_U75 P2_U2388 ; P2_U5914
g9795 nand P2_ADD_394_U65 P2_U2386 ; P2_U5915
g9796 nand P2_R2278_U93 P2_U2385 ; P2_U5916
g9797 nand P2_ADD_371_1212_U24 P2_U2384 ; P2_U5917
g9798 nand P2_U2381 P2_REIP_REG_29__SCAN_IN ; P2_U5918
g9799 nand P2_U5673 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_U5919
g9800 nand P2_R2096_U76 P2_U2390 ; P2_U5920
g9801 nand P2_R2099_U73 P2_U2389 ; P2_U5921
g9802 nand P2_R2027_U73 P2_U2388 ; P2_U5922
g9803 nand P2_ADD_394_U64 P2_U2386 ; P2_U5923
g9804 nand P2_R2278_U91 P2_U2385 ; P2_U5924
g9805 nand P2_ADD_371_1212_U69 P2_U2384 ; P2_U5925
g9806 nand P2_U2381 P2_REIP_REG_30__SCAN_IN ; P2_U5926
g9807 nand P2_U5673 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_U5927
g9808 nand P2_R2096_U50 P2_U2390 ; P2_U5928
g9809 nand P2_R2099_U72 P2_U2389 ; P2_U5929
g9810 nand P2_R2027_U72 P2_U2388 ; P2_U5930
g9811 nand P2_ADD_394_U84 P2_U2386 ; P2_U5931
g9812 nand P2_R2278_U5 P2_U2385 ; P2_U5932
g9813 nand P2_ADD_371_1212_U83 P2_U2384 ; P2_U5933
g9814 nand P2_U2381 P2_REIP_REG_31__SCAN_IN ; P2_U5934
g9815 nand P2_U5673 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_U5935
g9816 nand P2_U4420 P2_U2374 P2_U4613 ; P2_U5936
g9817 nand P2_U5661 P2_U3284 ; P2_U5937
g9818 not P2_U3537 ; P2_U5938
g9819 nand P2_U3302 P2_STATE2_REG_1__SCAN_IN ; P2_U5939
g9820 nand P2_U3540 P2_U5939 ; P2_U5940
g9821 nand P2_U2387 P2_PHYADDRPOINTER_REG_0__SCAN_IN ; P2_U5941
g9822 nand P2_U2373 P2_ADD_371_1212_U68 ; P2_U5942
g9823 nand P2_U2372 P2_R2099_U94 ; P2_U5943
g9824 nand P2_U2371 P2_REIP_REG_0__SCAN_IN ; P2_U5944
g9825 nand P2_U2370 P2_R2278_U83 ; P2_U5945
g9826 nand P2_U5938 P2_PHYADDRPOINTER_REG_0__SCAN_IN ; P2_U5946
g9827 nand P2_R2337_U4 P2_U2387 ; P2_U5947
g9828 nand P2_U2373 P2_ADD_371_1212_U25 ; P2_U5948
g9829 nand P2_U2372 P2_R2099_U5 ; P2_U5949
g9830 nand P2_U2371 P2_REIP_REG_1__SCAN_IN ; P2_U5950
g9831 nand P2_U2370 P2_R2278_U6 ; P2_U5951
g9832 nand P2_U5938 P2_PHYADDRPOINTER_REG_1__SCAN_IN ; P2_U5952
g9833 nand P2_R2337_U70 P2_U2387 ; P2_U5953
g9834 nand P2_U2373 P2_ADD_371_1212_U79 ; P2_U5954
g9835 nand P2_U2372 P2_R2099_U96 ; P2_U5955
g9836 nand P2_U2371 P2_REIP_REG_2__SCAN_IN ; P2_U5956
g9837 nand P2_U2370 P2_R2278_U92 ; P2_U5957
g9838 nand P2_U5938 P2_PHYADDRPOINTER_REG_2__SCAN_IN ; P2_U5958
g9839 nand P2_R2337_U67 P2_U2387 ; P2_U5959
g9840 nand P2_U2373 P2_ADD_371_1212_U84 ; P2_U5960
g9841 nand P2_U2372 P2_R2099_U95 ; P2_U5961
g9842 nand P2_U2371 P2_REIP_REG_3__SCAN_IN ; P2_U5962
g9843 nand P2_U2370 P2_R2278_U90 ; P2_U5963
g9844 nand P2_U5938 P2_PHYADDRPOINTER_REG_3__SCAN_IN ; P2_U5964
g9845 nand P2_R2337_U66 P2_U2387 ; P2_U5965
g9846 nand P2_U2373 P2_ADD_371_1212_U80 ; P2_U5966
g9847 nand P2_U2372 P2_R2099_U98 ; P2_U5967
g9848 nand P2_U2371 P2_REIP_REG_4__SCAN_IN ; P2_U5968
g9849 nand P2_U2370 P2_R2278_U89 ; P2_U5969
g9850 nand P2_U5938 P2_PHYADDRPOINTER_REG_4__SCAN_IN ; P2_U5970
g9851 nand P2_R2337_U65 P2_U2387 ; P2_U5971
g9852 nand P2_U2373 P2_ADD_371_1212_U81 ; P2_U5972
g9853 nand P2_U2372 P2_R2099_U71 ; P2_U5973
g9854 nand P2_U2371 P2_REIP_REG_5__SCAN_IN ; P2_U5974
g9855 nand P2_U2370 P2_R2278_U88 ; P2_U5975
g9856 nand P2_U5938 P2_PHYADDRPOINTER_REG_5__SCAN_IN ; P2_U5976
g9857 nand P2_R2337_U64 P2_U2387 ; P2_U5977
g9858 nand P2_U2373 P2_ADD_371_1212_U78 ; P2_U5978
g9859 nand P2_U2372 P2_R2099_U70 ; P2_U5979
g9860 nand P2_U2371 P2_REIP_REG_6__SCAN_IN ; P2_U5980
g9861 nand P2_U2370 P2_R2278_U87 ; P2_U5981
g9862 nand P2_U5938 P2_PHYADDRPOINTER_REG_6__SCAN_IN ; P2_U5982
g9863 nand P2_R2337_U63 P2_U2387 ; P2_U5983
g9864 nand P2_U2373 P2_ADD_371_1212_U85 ; P2_U5984
g9865 nand P2_U2372 P2_R2099_U69 ; P2_U5985
g9866 nand P2_U2371 P2_REIP_REG_7__SCAN_IN ; P2_U5986
g9867 nand P2_U2370 P2_R2278_U86 ; P2_U5987
g9868 nand P2_U5938 P2_PHYADDRPOINTER_REG_7__SCAN_IN ; P2_U5988
g9869 nand P2_R2337_U62 P2_U2387 ; P2_U5989
g9870 nand P2_U2373 P2_ADD_371_1212_U82 ; P2_U5990
g9871 nand P2_U2372 P2_R2099_U68 ; P2_U5991
g9872 nand P2_U2371 P2_REIP_REG_8__SCAN_IN ; P2_U5992
g9873 nand P2_U2370 P2_R2278_U85 ; P2_U5993
g9874 nand P2_U5938 P2_PHYADDRPOINTER_REG_8__SCAN_IN ; P2_U5994
g9875 nand P2_R2337_U61 P2_U2387 ; P2_U5995
g9876 nand P2_U2373 P2_ADD_371_1212_U118 ; P2_U5996
g9877 nand P2_U2372 P2_R2099_U67 ; P2_U5997
g9878 nand P2_U2371 P2_REIP_REG_9__SCAN_IN ; P2_U5998
g9879 nand P2_U2370 P2_R2278_U84 ; P2_U5999
g9880 nand P2_U5938 P2_PHYADDRPOINTER_REG_9__SCAN_IN ; P2_U6000
g9881 nand P2_R2337_U90 P2_U2387 ; P2_U6001
g9882 nand P2_U2373 P2_ADD_371_1212_U13 ; P2_U6002
g9883 nand P2_U2372 P2_R2099_U93 ; P2_U6003
g9884 nand P2_U2371 P2_REIP_REG_10__SCAN_IN ; P2_U6004
g9885 nand P2_U2370 P2_R2278_U112 ; P2_U6005
g9886 nand P2_U5938 P2_PHYADDRPOINTER_REG_10__SCAN_IN ; P2_U6006
g9887 nand P2_R2337_U89 P2_U2387 ; P2_U6007
g9888 nand P2_U2373 P2_ADD_371_1212_U14 ; P2_U6008
g9889 nand P2_U2372 P2_R2099_U92 ; P2_U6009
g9890 nand P2_U2371 P2_REIP_REG_11__SCAN_IN ; P2_U6010
g9891 nand P2_U2370 P2_R2278_U111 ; P2_U6011
g9892 nand P2_U5938 P2_PHYADDRPOINTER_REG_11__SCAN_IN ; P2_U6012
g9893 nand P2_R2337_U88 P2_U2387 ; P2_U6013
g9894 nand P2_U2373 P2_ADD_371_1212_U76 ; P2_U6014
g9895 nand P2_U2372 P2_R2099_U91 ; P2_U6015
g9896 nand P2_U2371 P2_REIP_REG_12__SCAN_IN ; P2_U6016
g9897 nand P2_U2370 P2_R2278_U110 ; P2_U6017
g9898 nand P2_U5938 P2_PHYADDRPOINTER_REG_12__SCAN_IN ; P2_U6018
g9899 nand P2_R2337_U87 P2_U2387 ; P2_U6019
g9900 nand P2_U2373 P2_ADD_371_1212_U15 ; P2_U6020
g9901 nand P2_U2372 P2_R2099_U90 ; P2_U6021
g9902 nand P2_U2371 P2_REIP_REG_13__SCAN_IN ; P2_U6022
g9903 nand P2_U2370 P2_R2278_U109 ; P2_U6023
g9904 nand P2_U5938 P2_PHYADDRPOINTER_REG_13__SCAN_IN ; P2_U6024
g9905 nand P2_R2337_U86 P2_U2387 ; P2_U6025
g9906 nand P2_U2373 P2_ADD_371_1212_U16 ; P2_U6026
g9907 nand P2_U2372 P2_R2099_U89 ; P2_U6027
g9908 nand P2_U2371 P2_REIP_REG_14__SCAN_IN ; P2_U6028
g9909 nand P2_U2370 P2_R2278_U108 ; P2_U6029
g9910 nand P2_U5938 P2_PHYADDRPOINTER_REG_14__SCAN_IN ; P2_U6030
g9911 nand P2_R2337_U85 P2_U2387 ; P2_U6031
g9912 nand P2_U2373 P2_ADD_371_1212_U73 ; P2_U6032
g9913 nand P2_U2372 P2_R2099_U88 ; P2_U6033
g9914 nand P2_U2371 P2_REIP_REG_15__SCAN_IN ; P2_U6034
g9915 nand P2_U2370 P2_R2278_U107 ; P2_U6035
g9916 nand P2_U5938 P2_PHYADDRPOINTER_REG_15__SCAN_IN ; P2_U6036
g9917 nand P2_R2337_U84 P2_U2387 ; P2_U6037
g9918 nand P2_U2373 P2_ADD_371_1212_U17 ; P2_U6038
g9919 nand P2_U2372 P2_R2099_U87 ; P2_U6039
g9920 nand P2_U2371 P2_REIP_REG_16__SCAN_IN ; P2_U6040
g9921 nand P2_U2370 P2_R2278_U106 ; P2_U6041
g9922 nand P2_U5938 P2_PHYADDRPOINTER_REG_16__SCAN_IN ; P2_U6042
g9923 nand P2_R2337_U83 P2_U2387 ; P2_U6043
g9924 nand P2_U2373 P2_ADD_371_1212_U71 ; P2_U6044
g9925 nand P2_U2372 P2_R2099_U86 ; P2_U6045
g9926 nand P2_U2371 P2_REIP_REG_17__SCAN_IN ; P2_U6046
g9927 nand P2_U2370 P2_R2278_U105 ; P2_U6047
g9928 nand P2_U5938 P2_PHYADDRPOINTER_REG_17__SCAN_IN ; P2_U6048
g9929 nand P2_R2337_U82 P2_U2387 ; P2_U6049
g9930 nand P2_U2373 P2_ADD_371_1212_U72 ; P2_U6050
g9931 nand P2_U2372 P2_R2099_U85 ; P2_U6051
g9932 nand P2_U2371 P2_REIP_REG_18__SCAN_IN ; P2_U6052
g9933 nand P2_U2370 P2_R2278_U104 ; P2_U6053
g9934 nand P2_U5938 P2_PHYADDRPOINTER_REG_18__SCAN_IN ; P2_U6054
g9935 nand P2_R2337_U81 P2_U2387 ; P2_U6055
g9936 nand P2_U2373 P2_ADD_371_1212_U18 ; P2_U6056
g9937 nand P2_U2372 P2_R2099_U84 ; P2_U6057
g9938 nand P2_U2371 P2_REIP_REG_19__SCAN_IN ; P2_U6058
g9939 nand P2_U2370 P2_R2278_U103 ; P2_U6059
g9940 nand P2_U5938 P2_PHYADDRPOINTER_REG_19__SCAN_IN ; P2_U6060
g9941 nand P2_R2337_U80 P2_U2387 ; P2_U6061
g9942 nand P2_U2373 P2_ADD_371_1212_U19 ; P2_U6062
g9943 nand P2_U2372 P2_R2099_U83 ; P2_U6063
g9944 nand P2_U2371 P2_REIP_REG_20__SCAN_IN ; P2_U6064
g9945 nand P2_U2370 P2_R2278_U102 ; P2_U6065
g9946 nand P2_U5938 P2_PHYADDRPOINTER_REG_20__SCAN_IN ; P2_U6066
g9947 nand P2_R2337_U79 P2_U2387 ; P2_U6067
g9948 nand P2_U2373 P2_ADD_371_1212_U75 ; P2_U6068
g9949 nand P2_U2372 P2_R2099_U82 ; P2_U6069
g9950 nand P2_U2371 P2_REIP_REG_21__SCAN_IN ; P2_U6070
g9951 nand P2_U2370 P2_R2278_U101 ; P2_U6071
g9952 nand P2_U5938 P2_PHYADDRPOINTER_REG_21__SCAN_IN ; P2_U6072
g9953 nand P2_R2337_U78 P2_U2387 ; P2_U6073
g9954 nand P2_U2373 P2_ADD_371_1212_U20 ; P2_U6074
g9955 nand P2_U2372 P2_R2099_U81 ; P2_U6075
g9956 nand P2_U2371 P2_REIP_REG_22__SCAN_IN ; P2_U6076
g9957 nand P2_U2370 P2_R2278_U100 ; P2_U6077
g9958 nand P2_U5938 P2_PHYADDRPOINTER_REG_22__SCAN_IN ; P2_U6078
g9959 nand P2_R2337_U77 P2_U2387 ; P2_U6079
g9960 nand P2_U2373 P2_ADD_371_1212_U21 ; P2_U6080
g9961 nand P2_U2372 P2_R2099_U80 ; P2_U6081
g9962 nand P2_U2371 P2_REIP_REG_23__SCAN_IN ; P2_U6082
g9963 nand P2_U2370 P2_R2278_U99 ; P2_U6083
g9964 nand P2_U5938 P2_PHYADDRPOINTER_REG_23__SCAN_IN ; P2_U6084
g9965 nand P2_R2337_U76 P2_U2387 ; P2_U6085
g9966 nand P2_U2373 P2_ADD_371_1212_U70 ; P2_U6086
g9967 nand P2_U2372 P2_R2099_U79 ; P2_U6087
g9968 nand P2_U2371 P2_REIP_REG_24__SCAN_IN ; P2_U6088
g9969 nand P2_U2370 P2_R2278_U98 ; P2_U6089
g9970 nand P2_U5938 P2_PHYADDRPOINTER_REG_24__SCAN_IN ; P2_U6090
g9971 nand P2_R2337_U75 P2_U2387 ; P2_U6091
g9972 nand P2_U2373 P2_ADD_371_1212_U77 ; P2_U6092
g9973 nand P2_U2372 P2_R2099_U78 ; P2_U6093
g9974 nand P2_U2371 P2_REIP_REG_25__SCAN_IN ; P2_U6094
g9975 nand P2_U2370 P2_R2278_U97 ; P2_U6095
g9976 nand P2_U5938 P2_PHYADDRPOINTER_REG_25__SCAN_IN ; P2_U6096
g9977 nand P2_R2337_U74 P2_U2387 ; P2_U6097
g9978 nand P2_U2373 P2_ADD_371_1212_U22 ; P2_U6098
g9979 nand P2_U2372 P2_R2099_U77 ; P2_U6099
g9980 nand P2_U2371 P2_REIP_REG_26__SCAN_IN ; P2_U6100
g9981 nand P2_U2370 P2_R2278_U96 ; P2_U6101
g9982 nand P2_U5938 P2_PHYADDRPOINTER_REG_26__SCAN_IN ; P2_U6102
g9983 nand P2_R2337_U73 P2_U2387 ; P2_U6103
g9984 nand P2_U2373 P2_ADD_371_1212_U74 ; P2_U6104
g9985 nand P2_U2372 P2_R2099_U76 ; P2_U6105
g9986 nand P2_U2371 P2_REIP_REG_27__SCAN_IN ; P2_U6106
g9987 nand P2_U2370 P2_R2278_U95 ; P2_U6107
g9988 nand P2_U5938 P2_PHYADDRPOINTER_REG_27__SCAN_IN ; P2_U6108
g9989 nand P2_R2337_U72 P2_U2387 ; P2_U6109
g9990 nand P2_U2373 P2_ADD_371_1212_U23 ; P2_U6110
g9991 nand P2_U2372 P2_R2099_U75 ; P2_U6111
g9992 nand P2_U2371 P2_REIP_REG_28__SCAN_IN ; P2_U6112
g9993 nand P2_U2370 P2_R2278_U94 ; P2_U6113
g9994 nand P2_U5938 P2_PHYADDRPOINTER_REG_28__SCAN_IN ; P2_U6114
g9995 nand P2_R2337_U71 P2_U2387 ; P2_U6115
g9996 nand P2_U2373 P2_ADD_371_1212_U24 ; P2_U6116
g9997 nand P2_U2372 P2_R2099_U74 ; P2_U6117
g9998 nand P2_U2371 P2_REIP_REG_29__SCAN_IN ; P2_U6118
g9999 nand P2_U2370 P2_R2278_U93 ; P2_U6119
g10000 nand P2_U5938 P2_PHYADDRPOINTER_REG_29__SCAN_IN ; P2_U6120
g10001 nand P2_R2337_U69 P2_U2387 ; P2_U6121
g10002 nand P2_U2373 P2_ADD_371_1212_U69 ; P2_U6122
g10003 nand P2_U2372 P2_R2099_U73 ; P2_U6123
g10004 nand P2_U2371 P2_REIP_REG_30__SCAN_IN ; P2_U6124
g10005 nand P2_U2370 P2_R2278_U91 ; P2_U6125
g10006 nand P2_U5938 P2_PHYADDRPOINTER_REG_30__SCAN_IN ; P2_U6126
g10007 nand P2_R2337_U68 P2_U2387 ; P2_U6127
g10008 nand P2_U2373 P2_ADD_371_1212_U83 ; P2_U6128
g10009 nand P2_U2372 P2_R2099_U72 ; P2_U6129
g10010 nand P2_U2371 P2_REIP_REG_31__SCAN_IN ; P2_U6130
g10011 nand P2_U2370 P2_R2278_U5 ; P2_U6131
g10012 nand P2_U5938 P2_PHYADDRPOINTER_REG_31__SCAN_IN ; P2_U6132
g10013 nand U211 P2_U2616 ; P2_U6133
g10014 nand P2_U2395 P2_EAX_REG_15__SCAN_IN ; P2_U6134
g10015 nand U308 P2_U2394 ; P2_U6135
g10016 nand P2_U3538 P2_LWORD_REG_15__SCAN_IN ; P2_U6136
g10017 nand P2_U2395 P2_EAX_REG_14__SCAN_IN ; P2_U6137
g10018 nand U309 P2_U2394 ; P2_U6138
g10019 nand P2_U3538 P2_LWORD_REG_14__SCAN_IN ; P2_U6139
g10020 nand P2_U2395 P2_EAX_REG_13__SCAN_IN ; P2_U6140
g10021 nand U310 P2_U2394 ; P2_U6141
g10022 nand P2_U3538 P2_LWORD_REG_13__SCAN_IN ; P2_U6142
g10023 nand P2_U2395 P2_EAX_REG_12__SCAN_IN ; P2_U6143
g10024 nand U311 P2_U2394 ; P2_U6144
g10025 nand P2_U3538 P2_LWORD_REG_12__SCAN_IN ; P2_U6145
g10026 nand P2_U2395 P2_EAX_REG_11__SCAN_IN ; P2_U6146
g10027 nand U312 P2_U2394 ; P2_U6147
g10028 nand P2_U3538 P2_LWORD_REG_11__SCAN_IN ; P2_U6148
g10029 nand P2_U2395 P2_EAX_REG_10__SCAN_IN ; P2_U6149
g10030 nand U313 P2_U2394 ; P2_U6150
g10031 nand P2_U3538 P2_LWORD_REG_10__SCAN_IN ; P2_U6151
g10032 nand P2_U2395 P2_EAX_REG_9__SCAN_IN ; P2_U6152
g10033 nand U283 P2_U2394 ; P2_U6153
g10034 nand P2_U3538 P2_LWORD_REG_9__SCAN_IN ; P2_U6154
g10035 nand P2_U2395 P2_EAX_REG_8__SCAN_IN ; P2_U6155
g10036 nand U284 P2_U2394 ; P2_U6156
g10037 nand P2_U3538 P2_LWORD_REG_8__SCAN_IN ; P2_U6157
g10038 nand P2_U2395 P2_EAX_REG_7__SCAN_IN ; P2_U6158
g10039 nand P2_U2394 U285 ; P2_U6159
g10040 nand P2_U3538 P2_LWORD_REG_7__SCAN_IN ; P2_U6160
g10041 nand P2_U2395 P2_EAX_REG_6__SCAN_IN ; P2_U6161
g10042 nand P2_U2394 U286 ; P2_U6162
g10043 nand P2_U3538 P2_LWORD_REG_6__SCAN_IN ; P2_U6163
g10044 nand P2_U2395 P2_EAX_REG_5__SCAN_IN ; P2_U6164
g10045 nand P2_U2394 U287 ; P2_U6165
g10046 nand P2_U3538 P2_LWORD_REG_5__SCAN_IN ; P2_U6166
g10047 nand P2_U2395 P2_EAX_REG_4__SCAN_IN ; P2_U6167
g10048 nand P2_U2394 U288 ; P2_U6168
g10049 nand P2_U3538 P2_LWORD_REG_4__SCAN_IN ; P2_U6169
g10050 nand P2_U2395 P2_EAX_REG_3__SCAN_IN ; P2_U6170
g10051 nand P2_U2394 U289 ; P2_U6171
g10052 nand P2_U3538 P2_LWORD_REG_3__SCAN_IN ; P2_U6172
g10053 nand P2_U2395 P2_EAX_REG_2__SCAN_IN ; P2_U6173
g10054 nand P2_U2394 U292 ; P2_U6174
g10055 nand P2_U3538 P2_LWORD_REG_2__SCAN_IN ; P2_U6175
g10056 nand P2_U2395 P2_EAX_REG_1__SCAN_IN ; P2_U6176
g10057 nand P2_U2394 U303 ; P2_U6177
g10058 nand P2_U3538 P2_LWORD_REG_1__SCAN_IN ; P2_U6178
g10059 nand P2_U2395 P2_EAX_REG_0__SCAN_IN ; P2_U6179
g10060 nand P2_U2394 U314 ; P2_U6180
g10061 nand P2_U3538 P2_LWORD_REG_0__SCAN_IN ; P2_U6181
g10062 nand P2_U2395 P2_EAX_REG_30__SCAN_IN ; P2_U6182
g10063 nand U309 P2_U2394 ; P2_U6183
g10064 nand P2_U3538 P2_UWORD_REG_14__SCAN_IN ; P2_U6184
g10065 nand P2_U2395 P2_EAX_REG_29__SCAN_IN ; P2_U6185
g10066 nand U310 P2_U2394 ; P2_U6186
g10067 nand P2_U3538 P2_UWORD_REG_13__SCAN_IN ; P2_U6187
g10068 nand P2_U2395 P2_EAX_REG_28__SCAN_IN ; P2_U6188
g10069 nand U311 P2_U2394 ; P2_U6189
g10070 nand P2_U3538 P2_UWORD_REG_12__SCAN_IN ; P2_U6190
g10071 nand P2_U2395 P2_EAX_REG_27__SCAN_IN ; P2_U6191
g10072 nand U312 P2_U2394 ; P2_U6192
g10073 nand P2_U3538 P2_UWORD_REG_11__SCAN_IN ; P2_U6193
g10074 nand P2_U2395 P2_EAX_REG_26__SCAN_IN ; P2_U6194
g10075 nand U313 P2_U2394 ; P2_U6195
g10076 nand P2_U3538 P2_UWORD_REG_10__SCAN_IN ; P2_U6196
g10077 nand P2_U2395 P2_EAX_REG_25__SCAN_IN ; P2_U6197
g10078 nand U283 P2_U2394 ; P2_U6198
g10079 nand P2_U3538 P2_UWORD_REG_9__SCAN_IN ; P2_U6199
g10080 nand P2_U2395 P2_EAX_REG_24__SCAN_IN ; P2_U6200
g10081 nand U284 P2_U2394 ; P2_U6201
g10082 nand P2_U3538 P2_UWORD_REG_8__SCAN_IN ; P2_U6202
g10083 nand P2_U2395 P2_EAX_REG_23__SCAN_IN ; P2_U6203
g10084 nand P2_U2394 U285 ; P2_U6204
g10085 nand P2_U3538 P2_UWORD_REG_7__SCAN_IN ; P2_U6205
g10086 nand P2_U2395 P2_EAX_REG_22__SCAN_IN ; P2_U6206
g10087 nand P2_U2394 U286 ; P2_U6207
g10088 nand P2_U3538 P2_UWORD_REG_6__SCAN_IN ; P2_U6208
g10089 nand P2_U2395 P2_EAX_REG_21__SCAN_IN ; P2_U6209
g10090 nand P2_U2394 U287 ; P2_U6210
g10091 nand P2_U3538 P2_UWORD_REG_5__SCAN_IN ; P2_U6211
g10092 nand P2_U2395 P2_EAX_REG_20__SCAN_IN ; P2_U6212
g10093 nand P2_U2394 U288 ; P2_U6213
g10094 nand P2_U3538 P2_UWORD_REG_4__SCAN_IN ; P2_U6214
g10095 nand P2_U2395 P2_EAX_REG_19__SCAN_IN ; P2_U6215
g10096 nand P2_U2394 U289 ; P2_U6216
g10097 nand P2_U3538 P2_UWORD_REG_3__SCAN_IN ; P2_U6217
g10098 nand P2_U2395 P2_EAX_REG_18__SCAN_IN ; P2_U6218
g10099 nand P2_U2394 U292 ; P2_U6219
g10100 nand P2_U3538 P2_UWORD_REG_2__SCAN_IN ; P2_U6220
g10101 nand P2_U2395 P2_EAX_REG_17__SCAN_IN ; P2_U6221
g10102 nand P2_U2394 U303 ; P2_U6222
g10103 nand P2_U3538 P2_UWORD_REG_1__SCAN_IN ; P2_U6223
g10104 nand P2_U2395 P2_EAX_REG_16__SCAN_IN ; P2_U6224
g10105 nand P2_U2394 U314 ; P2_U6225
g10106 nand P2_U3538 P2_UWORD_REG_0__SCAN_IN ; P2_U6226
g10107 nand P2_U4057 P2_U4421 P2_R2167_U6 ; P2_U6227
g10108 nand P2_U4058 P2_U2446 ; P2_U6228
g10109 nand P2_U6228 P2_U6227 ; P2_U6229
g10110 nand P2_U4411 P2_U6229 ; P2_U6230
g10111 nand P2_U4467 P2_STATE2_REG_1__SCAN_IN ; P2_U6231
g10112 not P2_U3541 ; P2_U6232
g10113 nand P2_U2430 P2_EAX_REG_0__SCAN_IN ; P2_U6233
g10114 nand P2_U2396 P2_LWORD_REG_0__SCAN_IN ; P2_U6234
g10115 nand P2_U6232 P2_DATAO_REG_0__SCAN_IN ; P2_U6235
g10116 nand P2_U2430 P2_EAX_REG_1__SCAN_IN ; P2_U6236
g10117 nand P2_U2396 P2_LWORD_REG_1__SCAN_IN ; P2_U6237
g10118 nand P2_U6232 P2_DATAO_REG_1__SCAN_IN ; P2_U6238
g10119 nand P2_U2430 P2_EAX_REG_2__SCAN_IN ; P2_U6239
g10120 nand P2_U2396 P2_LWORD_REG_2__SCAN_IN ; P2_U6240
g10121 nand P2_U6232 P2_DATAO_REG_2__SCAN_IN ; P2_U6241
g10122 nand P2_U2430 P2_EAX_REG_3__SCAN_IN ; P2_U6242
g10123 nand P2_U2396 P2_LWORD_REG_3__SCAN_IN ; P2_U6243
g10124 nand P2_U6232 P2_DATAO_REG_3__SCAN_IN ; P2_U6244
g10125 nand P2_U2430 P2_EAX_REG_4__SCAN_IN ; P2_U6245
g10126 nand P2_U2396 P2_LWORD_REG_4__SCAN_IN ; P2_U6246
g10127 nand P2_U6232 P2_DATAO_REG_4__SCAN_IN ; P2_U6247
g10128 nand P2_U2430 P2_EAX_REG_5__SCAN_IN ; P2_U6248
g10129 nand P2_U2396 P2_LWORD_REG_5__SCAN_IN ; P2_U6249
g10130 nand P2_U6232 P2_DATAO_REG_5__SCAN_IN ; P2_U6250
g10131 nand P2_U2430 P2_EAX_REG_6__SCAN_IN ; P2_U6251
g10132 nand P2_U2396 P2_LWORD_REG_6__SCAN_IN ; P2_U6252
g10133 nand P2_U6232 P2_DATAO_REG_6__SCAN_IN ; P2_U6253
g10134 nand P2_U2430 P2_EAX_REG_7__SCAN_IN ; P2_U6254
g10135 nand P2_U2396 P2_LWORD_REG_7__SCAN_IN ; P2_U6255
g10136 nand P2_U6232 P2_DATAO_REG_7__SCAN_IN ; P2_U6256
g10137 nand P2_U2430 P2_EAX_REG_8__SCAN_IN ; P2_U6257
g10138 nand P2_U2396 P2_LWORD_REG_8__SCAN_IN ; P2_U6258
g10139 nand P2_U6232 P2_DATAO_REG_8__SCAN_IN ; P2_U6259
g10140 nand P2_U2430 P2_EAX_REG_9__SCAN_IN ; P2_U6260
g10141 nand P2_U2396 P2_LWORD_REG_9__SCAN_IN ; P2_U6261
g10142 nand P2_U6232 P2_DATAO_REG_9__SCAN_IN ; P2_U6262
g10143 nand P2_U2430 P2_EAX_REG_10__SCAN_IN ; P2_U6263
g10144 nand P2_U2396 P2_LWORD_REG_10__SCAN_IN ; P2_U6264
g10145 nand P2_U6232 P2_DATAO_REG_10__SCAN_IN ; P2_U6265
g10146 nand P2_U2430 P2_EAX_REG_11__SCAN_IN ; P2_U6266
g10147 nand P2_U2396 P2_LWORD_REG_11__SCAN_IN ; P2_U6267
g10148 nand P2_U6232 P2_DATAO_REG_11__SCAN_IN ; P2_U6268
g10149 nand P2_U2430 P2_EAX_REG_12__SCAN_IN ; P2_U6269
g10150 nand P2_U2396 P2_LWORD_REG_12__SCAN_IN ; P2_U6270
g10151 nand P2_U6232 P2_DATAO_REG_12__SCAN_IN ; P2_U6271
g10152 nand P2_U2430 P2_EAX_REG_13__SCAN_IN ; P2_U6272
g10153 nand P2_U2396 P2_LWORD_REG_13__SCAN_IN ; P2_U6273
g10154 nand P2_U6232 P2_DATAO_REG_13__SCAN_IN ; P2_U6274
g10155 nand P2_U2430 P2_EAX_REG_14__SCAN_IN ; P2_U6275
g10156 nand P2_U2396 P2_LWORD_REG_14__SCAN_IN ; P2_U6276
g10157 nand P2_U6232 P2_DATAO_REG_14__SCAN_IN ; P2_U6277
g10158 nand P2_U2430 P2_EAX_REG_15__SCAN_IN ; P2_U6278
g10159 nand P2_U2396 P2_LWORD_REG_15__SCAN_IN ; P2_U6279
g10160 nand P2_U6232 P2_DATAO_REG_15__SCAN_IN ; P2_U6280
g10161 nand P2_U2435 P2_EAX_REG_16__SCAN_IN ; P2_U6281
g10162 nand P2_U2396 P2_UWORD_REG_0__SCAN_IN ; P2_U6282
g10163 nand P2_U6232 P2_DATAO_REG_16__SCAN_IN ; P2_U6283
g10164 nand P2_U2435 P2_EAX_REG_17__SCAN_IN ; P2_U6284
g10165 nand P2_U2396 P2_UWORD_REG_1__SCAN_IN ; P2_U6285
g10166 nand P2_U6232 P2_DATAO_REG_17__SCAN_IN ; P2_U6286
g10167 nand P2_U2435 P2_EAX_REG_18__SCAN_IN ; P2_U6287
g10168 nand P2_U2396 P2_UWORD_REG_2__SCAN_IN ; P2_U6288
g10169 nand P2_U6232 P2_DATAO_REG_18__SCAN_IN ; P2_U6289
g10170 nand P2_U2435 P2_EAX_REG_19__SCAN_IN ; P2_U6290
g10171 nand P2_U2396 P2_UWORD_REG_3__SCAN_IN ; P2_U6291
g10172 nand P2_U6232 P2_DATAO_REG_19__SCAN_IN ; P2_U6292
g10173 nand P2_U2435 P2_EAX_REG_20__SCAN_IN ; P2_U6293
g10174 nand P2_U2396 P2_UWORD_REG_4__SCAN_IN ; P2_U6294
g10175 nand P2_U6232 P2_DATAO_REG_20__SCAN_IN ; P2_U6295
g10176 nand P2_U2435 P2_EAX_REG_21__SCAN_IN ; P2_U6296
g10177 nand P2_U2396 P2_UWORD_REG_5__SCAN_IN ; P2_U6297
g10178 nand P2_U6232 P2_DATAO_REG_21__SCAN_IN ; P2_U6298
g10179 nand P2_U2435 P2_EAX_REG_22__SCAN_IN ; P2_U6299
g10180 nand P2_U2396 P2_UWORD_REG_6__SCAN_IN ; P2_U6300
g10181 nand P2_U6232 P2_DATAO_REG_22__SCAN_IN ; P2_U6301
g10182 nand P2_U2435 P2_EAX_REG_23__SCAN_IN ; P2_U6302
g10183 nand P2_U2396 P2_UWORD_REG_7__SCAN_IN ; P2_U6303
g10184 nand P2_U6232 P2_DATAO_REG_23__SCAN_IN ; P2_U6304
g10185 nand P2_U2435 P2_EAX_REG_24__SCAN_IN ; P2_U6305
g10186 nand P2_U2396 P2_UWORD_REG_8__SCAN_IN ; P2_U6306
g10187 nand P2_U6232 P2_DATAO_REG_24__SCAN_IN ; P2_U6307
g10188 nand P2_U2435 P2_EAX_REG_25__SCAN_IN ; P2_U6308
g10189 nand P2_U2396 P2_UWORD_REG_9__SCAN_IN ; P2_U6309
g10190 nand P2_U6232 P2_DATAO_REG_25__SCAN_IN ; P2_U6310
g10191 nand P2_U2435 P2_EAX_REG_26__SCAN_IN ; P2_U6311
g10192 nand P2_U2396 P2_UWORD_REG_10__SCAN_IN ; P2_U6312
g10193 nand P2_U6232 P2_DATAO_REG_26__SCAN_IN ; P2_U6313
g10194 nand P2_U2435 P2_EAX_REG_27__SCAN_IN ; P2_U6314
g10195 nand P2_U2396 P2_UWORD_REG_11__SCAN_IN ; P2_U6315
g10196 nand P2_U6232 P2_DATAO_REG_27__SCAN_IN ; P2_U6316
g10197 nand P2_U2435 P2_EAX_REG_28__SCAN_IN ; P2_U6317
g10198 nand P2_U2396 P2_UWORD_REG_12__SCAN_IN ; P2_U6318
g10199 nand P2_U6232 P2_DATAO_REG_28__SCAN_IN ; P2_U6319
g10200 nand P2_U2435 P2_EAX_REG_29__SCAN_IN ; P2_U6320
g10201 nand P2_U2396 P2_UWORD_REG_13__SCAN_IN ; P2_U6321
g10202 nand P2_U6232 P2_DATAO_REG_29__SCAN_IN ; P2_U6322
g10203 nand P2_U2435 P2_EAX_REG_30__SCAN_IN ; P2_U6323
g10204 nand P2_U2396 P2_UWORD_REG_14__SCAN_IN ; P2_U6324
g10205 nand P2_U6232 P2_DATAO_REG_30__SCAN_IN ; P2_U6325
g10206 nand P2_U2513 P2_U3254 ; P2_U6326
g10207 nand P2_U2433 U314 ; P2_U6327
g10208 nand P2_ADD_391_1196_U87 P2_U2397 ; P2_U6328
g10209 nand P2_U2380 P2_R2096_U68 ; P2_U6329
g10210 nand P2_U3542 P2_EAX_REG_0__SCAN_IN ; P2_U6330
g10211 nand P2_U2433 U303 ; P2_U6331
g10212 nand P2_ADD_391_1196_U12 P2_U2397 ; P2_U6332
g10213 nand P2_U2380 P2_R2096_U51 ; P2_U6333
g10214 nand P2_U3542 P2_EAX_REG_1__SCAN_IN ; P2_U6334
g10215 nand P2_U2433 U292 ; P2_U6335
g10216 nand P2_ADD_391_1196_U92 P2_U2397 ; P2_U6336
g10217 nand P2_U2380 P2_R2096_U77 ; P2_U6337
g10218 nand P2_U3542 P2_EAX_REG_2__SCAN_IN ; P2_U6338
g10219 nand P2_U2433 U289 ; P2_U6339
g10220 nand P2_ADD_391_1196_U91 P2_U2397 ; P2_U6340
g10221 nand P2_U2380 P2_R2096_U75 ; P2_U6341
g10222 nand P2_U3542 P2_EAX_REG_3__SCAN_IN ; P2_U6342
g10223 nand P2_U2433 U288 ; P2_U6343
g10224 nand P2_ADD_391_1196_U90 P2_U2397 ; P2_U6344
g10225 nand P2_U2380 P2_R2096_U74 ; P2_U6345
g10226 nand P2_U3542 P2_EAX_REG_4__SCAN_IN ; P2_U6346
g10227 nand P2_U2433 U287 ; P2_U6347
g10228 nand P2_ADD_391_1196_U9 P2_U2397 ; P2_U6348
g10229 nand P2_U2380 P2_R2096_U73 ; P2_U6349
g10230 nand P2_U3542 P2_EAX_REG_5__SCAN_IN ; P2_U6350
g10231 nand P2_U2433 U286 ; P2_U6351
g10232 nand P2_ADD_391_1196_U89 P2_U2397 ; P2_U6352
g10233 nand P2_U2380 P2_R2096_U72 ; P2_U6353
g10234 nand P2_U3542 P2_EAX_REG_6__SCAN_IN ; P2_U6354
g10235 nand P2_U2433 U285 ; P2_U6355
g10236 nand P2_ADD_391_1196_U10 P2_U2397 ; P2_U6356
g10237 nand P2_U2380 P2_R2096_U71 ; P2_U6357
g10238 nand P2_U3542 P2_EAX_REG_7__SCAN_IN ; P2_U6358
g10239 nand P2_U2433 U284 ; P2_U6359
g10240 nand P2_ADD_391_1196_U88 P2_U2397 ; P2_U6360
g10241 nand P2_U2380 P2_R2096_U70 ; P2_U6361
g10242 nand P2_U3542 P2_EAX_REG_8__SCAN_IN ; P2_U6362
g10243 nand P2_U2433 U283 ; P2_U6363
g10244 nand P2_ADD_391_1196_U11 P2_U2397 ; P2_U6364
g10245 nand P2_U2380 P2_R2096_U69 ; P2_U6365
g10246 nand P2_U3542 P2_EAX_REG_9__SCAN_IN ; P2_U6366
g10247 nand P2_U2433 U313 ; P2_U6367
g10248 nand P2_ADD_391_1196_U109 P2_U2397 ; P2_U6368
g10249 nand P2_U2380 P2_R2096_U97 ; P2_U6369
g10250 nand P2_U3542 P2_EAX_REG_10__SCAN_IN ; P2_U6370
g10251 nand P2_U2433 U312 ; P2_U6371
g10252 nand P2_ADD_391_1196_U5 P2_U2397 ; P2_U6372
g10253 nand P2_U2380 P2_R2096_U96 ; P2_U6373
g10254 nand P2_U3542 P2_EAX_REG_11__SCAN_IN ; P2_U6374
g10255 nand P2_U2433 U311 ; P2_U6375
g10256 nand P2_ADD_391_1196_U108 P2_U2397 ; P2_U6376
g10257 nand P2_U2380 P2_R2096_U95 ; P2_U6377
g10258 nand P2_U3542 P2_EAX_REG_12__SCAN_IN ; P2_U6378
g10259 nand P2_U2433 U310 ; P2_U6379
g10260 nand P2_ADD_391_1196_U6 P2_U2397 ; P2_U6380
g10261 nand P2_U2380 P2_R2096_U94 ; P2_U6381
g10262 nand P2_U3542 P2_EAX_REG_13__SCAN_IN ; P2_U6382
g10263 nand P2_U2433 U309 ; P2_U6383
g10264 nand P2_ADD_391_1196_U107 P2_U2397 ; P2_U6384
g10265 nand P2_U2380 P2_R2096_U93 ; P2_U6385
g10266 nand P2_U3542 P2_EAX_REG_14__SCAN_IN ; P2_U6386
g10267 nand P2_U2433 U308 ; P2_U6387
g10268 nand P2_ADD_391_1196_U7 P2_U2397 ; P2_U6388
g10269 nand P2_U2380 P2_R2096_U92 ; P2_U6389
g10270 nand P2_U3542 P2_EAX_REG_15__SCAN_IN ; P2_U6390
g10271 nand P2_U2434 U314 ; P2_U6391
g10272 nand P2_U2427 U307 ; P2_U6392
g10273 nand P2_ADD_391_1196_U106 P2_U2397 ; P2_U6393
g10274 nand P2_U2380 P2_R2096_U91 ; P2_U6394
g10275 nand P2_U3542 P2_EAX_REG_16__SCAN_IN ; P2_U6395
g10276 nand P2_U2434 U303 ; P2_U6396
g10277 nand P2_U2427 U306 ; P2_U6397
g10278 nand P2_ADD_391_1196_U105 P2_U2397 ; P2_U6398
g10279 nand P2_U2380 P2_R2096_U90 ; P2_U6399
g10280 nand P2_U3542 P2_EAX_REG_17__SCAN_IN ; P2_U6400
g10281 nand P2_U2434 U292 ; P2_U6401
g10282 nand P2_U2427 U305 ; P2_U6402
g10283 nand P2_ADD_391_1196_U104 P2_U2397 ; P2_U6403
g10284 nand P2_U2380 P2_R2096_U89 ; P2_U6404
g10285 nand P2_U3542 P2_EAX_REG_18__SCAN_IN ; P2_U6405
g10286 nand P2_U2434 U289 ; P2_U6406
g10287 nand P2_U2427 U304 ; P2_U6407
g10288 nand P2_ADD_391_1196_U103 P2_U2397 ; P2_U6408
g10289 nand P2_U2380 P2_R2096_U88 ; P2_U6409
g10290 nand P2_U3542 P2_EAX_REG_19__SCAN_IN ; P2_U6410
g10291 nand P2_U2434 U288 ; P2_U6411
g10292 nand P2_U2427 U302 ; P2_U6412
g10293 nand P2_ADD_391_1196_U102 P2_U2397 ; P2_U6413
g10294 nand P2_U2380 P2_R2096_U87 ; P2_U6414
g10295 nand P2_U3542 P2_EAX_REG_20__SCAN_IN ; P2_U6415
g10296 nand P2_U2434 U287 ; P2_U6416
g10297 nand P2_U2427 U301 ; P2_U6417
g10298 nand P2_ADD_391_1196_U101 P2_U2397 ; P2_U6418
g10299 nand P2_U2380 P2_R2096_U86 ; P2_U6419
g10300 nand P2_U3542 P2_EAX_REG_21__SCAN_IN ; P2_U6420
g10301 nand P2_U2434 U286 ; P2_U6421
g10302 nand P2_U2427 U300 ; P2_U6422
g10303 nand P2_ADD_391_1196_U100 P2_U2397 ; P2_U6423
g10304 nand P2_U2380 P2_R2096_U85 ; P2_U6424
g10305 nand P2_U3542 P2_EAX_REG_22__SCAN_IN ; P2_U6425
g10306 nand P2_U2434 U285 ; P2_U6426
g10307 nand P2_U2427 U299 ; P2_U6427
g10308 nand P2_ADD_391_1196_U99 P2_U2397 ; P2_U6428
g10309 nand P2_U2380 P2_R2096_U84 ; P2_U6429
g10310 nand P2_U3542 P2_EAX_REG_23__SCAN_IN ; P2_U6430
g10311 nand P2_U2434 U284 ; P2_U6431
g10312 nand P2_U2427 U298 ; P2_U6432
g10313 nand P2_ADD_391_1196_U98 P2_U2397 ; P2_U6433
g10314 nand P2_U2380 P2_R2096_U83 ; P2_U6434
g10315 nand P2_U3542 P2_EAX_REG_24__SCAN_IN ; P2_U6435
g10316 nand P2_U2434 U283 ; P2_U6436
g10317 nand P2_U2427 U297 ; P2_U6437
g10318 nand P2_ADD_391_1196_U97 P2_U2397 ; P2_U6438
g10319 nand P2_U2380 P2_R2096_U82 ; P2_U6439
g10320 nand P2_U3542 P2_EAX_REG_25__SCAN_IN ; P2_U6440
g10321 nand P2_U2434 U313 ; P2_U6441
g10322 nand P2_U2427 U296 ; P2_U6442
g10323 nand P2_ADD_391_1196_U96 P2_U2397 ; P2_U6443
g10324 nand P2_U2380 P2_R2096_U81 ; P2_U6444
g10325 nand P2_U3542 P2_EAX_REG_26__SCAN_IN ; P2_U6445
g10326 nand P2_U2434 U312 ; P2_U6446
g10327 nand P2_U2427 U295 ; P2_U6447
g10328 nand P2_ADD_391_1196_U95 P2_U2397 ; P2_U6448
g10329 nand P2_U2380 P2_R2096_U80 ; P2_U6449
g10330 nand P2_U3542 P2_EAX_REG_27__SCAN_IN ; P2_U6450
g10331 nand P2_U2434 U311 ; P2_U6451
g10332 nand P2_U2427 U294 ; P2_U6452
g10333 nand P2_ADD_391_1196_U94 P2_U2397 ; P2_U6453
g10334 nand P2_U2380 P2_R2096_U79 ; P2_U6454
g10335 nand P2_U3542 P2_EAX_REG_28__SCAN_IN ; P2_U6455
g10336 nand P2_U2434 U310 ; P2_U6456
g10337 nand P2_U2427 U293 ; P2_U6457
g10338 nand P2_ADD_391_1196_U93 P2_U2397 ; P2_U6458
g10339 nand P2_U2380 P2_R2096_U78 ; P2_U6459
g10340 nand P2_U3542 P2_EAX_REG_29__SCAN_IN ; P2_U6460
g10341 nand P2_U2434 U309 ; P2_U6461
g10342 nand P2_U2427 U291 ; P2_U6462
g10343 nand P2_ADD_391_1196_U8 P2_U2397 ; P2_U6463
g10344 nand P2_U2380 P2_R2096_U76 ; P2_U6464
g10345 nand P2_U3542 P2_EAX_REG_30__SCAN_IN ; P2_U6465
g10346 nand P2_U2427 U290 ; P2_U6466
g10347 nand P2_U2380 P2_R2096_U50 ; P2_U6467
g10348 nand P2_U3542 P2_EAX_REG_31__SCAN_IN ; P2_U6468
g10349 nand P2_U4435 P2_U3297 ; P2_U6469
g10350 nand P2_U3578 P2_U6469 ; P2_U6470
g10351 nand P2_U2393 P2_R2182_U69 ; P2_U6471
g10352 nand P2_U2379 P2_R2099_U94 ; P2_U6472
g10353 nand P2_U3543 P2_EBX_REG_0__SCAN_IN ; P2_U6473
g10354 nand P2_U2393 P2_R2182_U68 ; P2_U6474
g10355 nand P2_U2379 P2_R2099_U5 ; P2_U6475
g10356 nand P2_U3543 P2_EBX_REG_1__SCAN_IN ; P2_U6476
g10357 nand P2_U2393 P2_R2182_U40 ; P2_U6477
g10358 nand P2_U2379 P2_R2099_U96 ; P2_U6478
g10359 nand P2_U3543 P2_EBX_REG_2__SCAN_IN ; P2_U6479
g10360 nand P2_U2393 P2_R2182_U76 ; P2_U6480
g10361 nand P2_U2379 P2_R2099_U95 ; P2_U6481
g10362 nand P2_U3543 P2_EBX_REG_3__SCAN_IN ; P2_U6482
g10363 nand P2_R2182_U75 P2_U2393 ; P2_U6483
g10364 nand P2_U2379 P2_R2099_U98 ; P2_U6484
g10365 nand P2_U3543 P2_EBX_REG_4__SCAN_IN ; P2_U6485
g10366 nand P2_R2182_U74 P2_U2393 ; P2_U6486
g10367 nand P2_U2379 P2_R2099_U71 ; P2_U6487
g10368 nand P2_U3543 P2_EBX_REG_5__SCAN_IN ; P2_U6488
g10369 nand P2_R2182_U73 P2_U2393 ; P2_U6489
g10370 nand P2_U2379 P2_R2099_U70 ; P2_U6490
g10371 nand P2_U3543 P2_EBX_REG_6__SCAN_IN ; P2_U6491
g10372 nand P2_R2182_U72 P2_U2393 ; P2_U6492
g10373 nand P2_U2379 P2_R2099_U69 ; P2_U6493
g10374 nand P2_U3543 P2_EBX_REG_7__SCAN_IN ; P2_U6494
g10375 nand P2_R2182_U71 P2_U2393 ; P2_U6495
g10376 nand P2_U2379 P2_R2099_U68 ; P2_U6496
g10377 nand P2_U3543 P2_EBX_REG_8__SCAN_IN ; P2_U6497
g10378 nand P2_R2182_U70 P2_U2393 ; P2_U6498
g10379 nand P2_U2379 P2_R2099_U67 ; P2_U6499
g10380 nand P2_U3543 P2_EBX_REG_9__SCAN_IN ; P2_U6500
g10381 nand P2_R2182_U96 P2_U2393 ; P2_U6501
g10382 nand P2_U2379 P2_R2099_U93 ; P2_U6502
g10383 nand P2_U3543 P2_EBX_REG_10__SCAN_IN ; P2_U6503
g10384 nand P2_R2182_U95 P2_U2393 ; P2_U6504
g10385 nand P2_U2379 P2_R2099_U92 ; P2_U6505
g10386 nand P2_U3543 P2_EBX_REG_11__SCAN_IN ; P2_U6506
g10387 nand P2_R2182_U94 P2_U2393 ; P2_U6507
g10388 nand P2_U2379 P2_R2099_U91 ; P2_U6508
g10389 nand P2_U3543 P2_EBX_REG_12__SCAN_IN ; P2_U6509
g10390 nand P2_R2182_U93 P2_U2393 ; P2_U6510
g10391 nand P2_U2379 P2_R2099_U90 ; P2_U6511
g10392 nand P2_U3543 P2_EBX_REG_13__SCAN_IN ; P2_U6512
g10393 nand P2_R2182_U92 P2_U2393 ; P2_U6513
g10394 nand P2_U2379 P2_R2099_U89 ; P2_U6514
g10395 nand P2_U3543 P2_EBX_REG_14__SCAN_IN ; P2_U6515
g10396 nand P2_R2182_U91 P2_U2393 ; P2_U6516
g10397 nand P2_U2379 P2_R2099_U88 ; P2_U6517
g10398 nand P2_U3543 P2_EBX_REG_15__SCAN_IN ; P2_U6518
g10399 nand P2_R2182_U90 P2_U2393 ; P2_U6519
g10400 nand P2_U2379 P2_R2099_U87 ; P2_U6520
g10401 nand P2_U3543 P2_EBX_REG_16__SCAN_IN ; P2_U6521
g10402 nand P2_R2182_U89 P2_U2393 ; P2_U6522
g10403 nand P2_U2379 P2_R2099_U86 ; P2_U6523
g10404 nand P2_U3543 P2_EBX_REG_17__SCAN_IN ; P2_U6524
g10405 nand P2_R2182_U88 P2_U2393 ; P2_U6525
g10406 nand P2_U2379 P2_R2099_U85 ; P2_U6526
g10407 nand P2_U3543 P2_EBX_REG_18__SCAN_IN ; P2_U6527
g10408 nand P2_R2182_U87 P2_U2393 ; P2_U6528
g10409 nand P2_U2379 P2_R2099_U84 ; P2_U6529
g10410 nand P2_U3543 P2_EBX_REG_19__SCAN_IN ; P2_U6530
g10411 nand P2_R2182_U86 P2_U2393 ; P2_U6531
g10412 nand P2_U2379 P2_R2099_U83 ; P2_U6532
g10413 nand P2_U3543 P2_EBX_REG_20__SCAN_IN ; P2_U6533
g10414 nand P2_R2182_U85 P2_U2393 ; P2_U6534
g10415 nand P2_U2379 P2_R2099_U82 ; P2_U6535
g10416 nand P2_U3543 P2_EBX_REG_21__SCAN_IN ; P2_U6536
g10417 nand P2_R2182_U84 P2_U2393 ; P2_U6537
g10418 nand P2_U2379 P2_R2099_U81 ; P2_U6538
g10419 nand P2_U3543 P2_EBX_REG_22__SCAN_IN ; P2_U6539
g10420 nand P2_R2182_U83 P2_U2393 ; P2_U6540
g10421 nand P2_U2379 P2_R2099_U80 ; P2_U6541
g10422 nand P2_U3543 P2_EBX_REG_23__SCAN_IN ; P2_U6542
g10423 nand P2_R2182_U82 P2_U2393 ; P2_U6543
g10424 nand P2_U2379 P2_R2099_U79 ; P2_U6544
g10425 nand P2_U3543 P2_EBX_REG_24__SCAN_IN ; P2_U6545
g10426 nand P2_R2182_U81 P2_U2393 ; P2_U6546
g10427 nand P2_U2379 P2_R2099_U78 ; P2_U6547
g10428 nand P2_U3543 P2_EBX_REG_25__SCAN_IN ; P2_U6548
g10429 nand P2_R2182_U80 P2_U2393 ; P2_U6549
g10430 nand P2_U2379 P2_R2099_U77 ; P2_U6550
g10431 nand P2_U3543 P2_EBX_REG_26__SCAN_IN ; P2_U6551
g10432 nand P2_R2182_U79 P2_U2393 ; P2_U6552
g10433 nand P2_U2379 P2_R2099_U76 ; P2_U6553
g10434 nand P2_U3543 P2_EBX_REG_27__SCAN_IN ; P2_U6554
g10435 nand P2_R2182_U78 P2_U2393 ; P2_U6555
g10436 nand P2_U2379 P2_R2099_U75 ; P2_U6556
g10437 nand P2_U3543 P2_EBX_REG_28__SCAN_IN ; P2_U6557
g10438 nand P2_R2182_U77 P2_U2393 ; P2_U6558
g10439 nand P2_U2379 P2_R2099_U74 ; P2_U6559
g10440 nand P2_U3543 P2_EBX_REG_29__SCAN_IN ; P2_U6560
g10441 nand P2_R2182_U41 P2_U2393 ; P2_U6561
g10442 nand P2_U2379 P2_R2099_U73 ; P2_U6562
g10443 nand P2_U3543 P2_EBX_REG_30__SCAN_IN ; P2_U6563
g10444 nand P2_U2379 P2_R2099_U72 ; P2_U6564
g10445 nand P2_U3543 P2_EBX_REG_31__SCAN_IN ; P2_U6565
g10446 nand P2_R2088_U6 P2_U4603 ; P2_U6566
g10447 nand P2_U4433 P2_R2167_U6 ; P2_U6567
g10448 nand P2_U6567 P2_U6566 ; P2_U6568
g10449 nand P2_U4461 P2_U3284 ; P2_U6569
g10450 not P2_U3546 ; P2_U6570
g10451 not P2_U3545 ; P2_U6571
g10452 or U211 P2_STATEBS16_REG_SCAN_IN ; P2_U6572
g10453 nand P2_R2267_U21 P2_U2587 ; P2_U6573
g10454 nand P2_U2588 P2_R2096_U68 ; P2_U6574
g10455 nand P2_U7743 P2_EBX_REG_0__SCAN_IN ; P2_U6575
g10456 nand P2_U2437 P2_R2182_U69 ; P2_U6576
g10457 nand P2_U2392 P2_R2099_U94 ; P2_U6577
g10458 nand P2_U2383 P2_PHYADDRPOINTER_REG_0__SCAN_IN ; P2_U6578
g10459 nand P2_U2382 P2_U3683 ; P2_U6579
g10460 nand P2_U2378 P2_PHYADDRPOINTER_REG_0__SCAN_IN ; P2_U6580
g10461 nand P2_U6570 P2_REIP_REG_0__SCAN_IN ; P2_U6581
g10462 nand P2_R2267_U43 P2_U2587 ; P2_U6582
g10463 nand P2_U2588 P2_R2096_U51 ; P2_U6583
g10464 nand P2_U7743 P2_EBX_REG_1__SCAN_IN ; P2_U6584
g10465 nand P2_U2437 P2_R2182_U68 ; P2_U6585
g10466 nand P2_U2392 P2_R2099_U5 ; P2_U6586
g10467 nand P2_U2383 P2_R2337_U4 ; P2_U6587
g10468 nand P2_U2382 P2_R1957_U49 ; P2_U6588
g10469 nand P2_U2378 P2_PHYADDRPOINTER_REG_1__SCAN_IN ; P2_U6589
g10470 nand P2_U6570 P2_REIP_REG_1__SCAN_IN ; P2_U6590
g10471 nand P2_R2267_U65 P2_U2587 ; P2_U6591
g10472 nand P2_U2588 P2_R2096_U77 ; P2_U6592
g10473 nand P2_U7743 P2_EBX_REG_2__SCAN_IN ; P2_U6593
g10474 nand P2_U2437 P2_R2182_U40 ; P2_U6594
g10475 nand P2_U2392 P2_R2099_U96 ; P2_U6595
g10476 nand P2_U2383 P2_R2337_U70 ; P2_U6596
g10477 nand P2_R1957_U17 P2_U2382 ; P2_U6597
g10478 nand P2_U2378 P2_PHYADDRPOINTER_REG_2__SCAN_IN ; P2_U6598
g10479 nand P2_U6570 P2_REIP_REG_2__SCAN_IN ; P2_U6599
g10480 nand P2_R2267_U17 P2_U2587 ; P2_U6600
g10481 nand P2_U2588 P2_R2096_U75 ; P2_U6601
g10482 nand P2_U7743 P2_EBX_REG_3__SCAN_IN ; P2_U6602
g10483 nand P2_U2437 P2_R2182_U76 ; P2_U6603
g10484 nand P2_U2392 P2_R2099_U95 ; P2_U6604
g10485 nand P2_U2383 P2_R2337_U67 ; P2_U6605
g10486 nand P2_R1957_U59 P2_U2382 ; P2_U6606
g10487 nand P2_U2378 P2_PHYADDRPOINTER_REG_3__SCAN_IN ; P2_U6607
g10488 nand P2_U6570 P2_REIP_REG_3__SCAN_IN ; P2_U6608
g10489 nand P2_R2267_U60 P2_U2587 ; P2_U6609
g10490 nand P2_U2588 P2_R2096_U74 ; P2_U6610
g10491 nand P2_U7743 P2_EBX_REG_4__SCAN_IN ; P2_U6611
g10492 nand P2_U2437 P2_R2182_U75 ; P2_U6612
g10493 nand P2_U2392 P2_R2099_U98 ; P2_U6613
g10494 nand P2_U2383 P2_R2337_U66 ; P2_U6614
g10495 nand P2_R1957_U18 P2_U2382 ; P2_U6615
g10496 nand P2_U2378 P2_PHYADDRPOINTER_REG_4__SCAN_IN ; P2_U6616
g10497 nand P2_U6570 P2_REIP_REG_4__SCAN_IN ; P2_U6617
g10498 nand P2_R2267_U18 P2_U2587 ; P2_U6618
g10499 nand P2_U2588 P2_R2096_U73 ; P2_U6619
g10500 nand P2_U7743 P2_EBX_REG_5__SCAN_IN ; P2_U6620
g10501 nand P2_U2437 P2_R2182_U74 ; P2_U6621
g10502 nand P2_U2392 P2_R2099_U71 ; P2_U6622
g10503 nand P2_U2383 P2_R2337_U65 ; P2_U6623
g10504 nand P2_R1957_U57 P2_U2382 ; P2_U6624
g10505 nand P2_U2378 P2_PHYADDRPOINTER_REG_5__SCAN_IN ; P2_U6625
g10506 nand P2_U6570 P2_REIP_REG_5__SCAN_IN ; P2_U6626
g10507 nand P2_R2267_U58 P2_U2587 ; P2_U6627
g10508 nand P2_U2588 P2_R2096_U72 ; P2_U6628
g10509 nand P2_U7743 P2_EBX_REG_6__SCAN_IN ; P2_U6629
g10510 nand P2_U2392 P2_R2099_U70 ; P2_U6630
g10511 nand P2_U2383 P2_R2337_U64 ; P2_U6631
g10512 nand P2_R1957_U19 P2_U2382 ; P2_U6632
g10513 nand P2_U2378 P2_PHYADDRPOINTER_REG_6__SCAN_IN ; P2_U6633
g10514 nand P2_U6570 P2_REIP_REG_6__SCAN_IN ; P2_U6634
g10515 nand P2_R2267_U19 P2_U2587 ; P2_U6635
g10516 nand P2_U2588 P2_R2096_U71 ; P2_U6636
g10517 nand P2_U7743 P2_EBX_REG_7__SCAN_IN ; P2_U6637
g10518 nand P2_U2392 P2_R2099_U69 ; P2_U6638
g10519 nand P2_U2383 P2_R2337_U63 ; P2_U6639
g10520 nand P2_R1957_U55 P2_U2382 ; P2_U6640
g10521 nand P2_U2378 P2_PHYADDRPOINTER_REG_7__SCAN_IN ; P2_U6641
g10522 nand P2_U6570 P2_REIP_REG_7__SCAN_IN ; P2_U6642
g10523 nand P2_R2267_U56 P2_U2587 ; P2_U6643
g10524 nand P2_U2588 P2_R2096_U70 ; P2_U6644
g10525 nand P2_U7743 P2_EBX_REG_8__SCAN_IN ; P2_U6645
g10526 nand P2_U2392 P2_R2099_U68 ; P2_U6646
g10527 nand P2_U2383 P2_R2337_U62 ; P2_U6647
g10528 nand P2_R1957_U20 P2_U2382 ; P2_U6648
g10529 nand P2_U2378 P2_PHYADDRPOINTER_REG_8__SCAN_IN ; P2_U6649
g10530 nand P2_U6570 P2_REIP_REG_8__SCAN_IN ; P2_U6650
g10531 nand P2_R2267_U20 P2_U2587 ; P2_U6651
g10532 nand P2_U2588 P2_R2096_U69 ; P2_U6652
g10533 nand P2_U7743 P2_EBX_REG_9__SCAN_IN ; P2_U6653
g10534 nand P2_U2392 P2_R2099_U67 ; P2_U6654
g10535 nand P2_U2383 P2_R2337_U61 ; P2_U6655
g10536 nand P2_R1957_U53 P2_U2382 ; P2_U6656
g10537 nand P2_U2378 P2_PHYADDRPOINTER_REG_9__SCAN_IN ; P2_U6657
g10538 nand P2_U6570 P2_REIP_REG_9__SCAN_IN ; P2_U6658
g10539 nand P2_R2267_U87 P2_U2587 ; P2_U6659
g10540 nand P2_U2588 P2_R2096_U97 ; P2_U6660
g10541 nand P2_U7743 P2_EBX_REG_10__SCAN_IN ; P2_U6661
g10542 nand P2_U2392 P2_R2099_U93 ; P2_U6662
g10543 nand P2_U2383 P2_R2337_U90 ; P2_U6663
g10544 nand P2_R1957_U6 P2_U2382 ; P2_U6664
g10545 nand P2_U2378 P2_PHYADDRPOINTER_REG_10__SCAN_IN ; P2_U6665
g10546 nand P2_U6570 P2_REIP_REG_10__SCAN_IN ; P2_U6666
g10547 nand P2_R2267_U6 P2_U2587 ; P2_U6667
g10548 nand P2_U2588 P2_R2096_U96 ; P2_U6668
g10549 nand P2_U7743 P2_EBX_REG_11__SCAN_IN ; P2_U6669
g10550 nand P2_U2392 P2_R2099_U92 ; P2_U6670
g10551 nand P2_U2383 P2_R2337_U89 ; P2_U6671
g10552 nand P2_R1957_U82 P2_U2382 ; P2_U6672
g10553 nand P2_U2378 P2_PHYADDRPOINTER_REG_11__SCAN_IN ; P2_U6673
g10554 nand P2_U6570 P2_REIP_REG_11__SCAN_IN ; P2_U6674
g10555 nand P2_R2267_U85 P2_U2587 ; P2_U6675
g10556 nand P2_U2588 P2_R2096_U95 ; P2_U6676
g10557 nand P2_U7743 P2_EBX_REG_12__SCAN_IN ; P2_U6677
g10558 nand P2_U2392 P2_R2099_U91 ; P2_U6678
g10559 nand P2_U2383 P2_R2337_U88 ; P2_U6679
g10560 nand P2_R1957_U7 P2_U2382 ; P2_U6680
g10561 nand P2_U2378 P2_PHYADDRPOINTER_REG_12__SCAN_IN ; P2_U6681
g10562 nand P2_U6570 P2_REIP_REG_12__SCAN_IN ; P2_U6682
g10563 nand P2_R2267_U7 P2_U2587 ; P2_U6683
g10564 nand P2_U2588 P2_R2096_U94 ; P2_U6684
g10565 nand P2_U7743 P2_EBX_REG_13__SCAN_IN ; P2_U6685
g10566 nand P2_U2392 P2_R2099_U90 ; P2_U6686
g10567 nand P2_U2383 P2_R2337_U87 ; P2_U6687
g10568 nand P2_R1957_U80 P2_U2382 ; P2_U6688
g10569 nand P2_U2378 P2_PHYADDRPOINTER_REG_13__SCAN_IN ; P2_U6689
g10570 nand P2_U6570 P2_REIP_REG_13__SCAN_IN ; P2_U6690
g10571 nand P2_R2267_U83 P2_U2587 ; P2_U6691
g10572 nand P2_U2588 P2_R2096_U93 ; P2_U6692
g10573 nand P2_U7743 P2_EBX_REG_14__SCAN_IN ; P2_U6693
g10574 nand P2_U2392 P2_R2099_U89 ; P2_U6694
g10575 nand P2_U2383 P2_R2337_U86 ; P2_U6695
g10576 nand P2_R1957_U8 P2_U2382 ; P2_U6696
g10577 nand P2_U2378 P2_PHYADDRPOINTER_REG_14__SCAN_IN ; P2_U6697
g10578 nand P2_U6570 P2_REIP_REG_14__SCAN_IN ; P2_U6698
g10579 nand P2_R2267_U8 P2_U2587 ; P2_U6699
g10580 nand P2_U2588 P2_R2096_U92 ; P2_U6700
g10581 nand P2_U7743 P2_EBX_REG_15__SCAN_IN ; P2_U6701
g10582 nand P2_U2392 P2_R2099_U88 ; P2_U6702
g10583 nand P2_U2383 P2_R2337_U85 ; P2_U6703
g10584 nand P2_R1957_U78 P2_U2382 ; P2_U6704
g10585 nand P2_U2378 P2_PHYADDRPOINTER_REG_15__SCAN_IN ; P2_U6705
g10586 nand P2_U6570 P2_REIP_REG_15__SCAN_IN ; P2_U6706
g10587 nand P2_R2267_U81 P2_U2587 ; P2_U6707
g10588 nand P2_U2588 P2_R2096_U91 ; P2_U6708
g10589 nand P2_U7743 P2_EBX_REG_16__SCAN_IN ; P2_U6709
g10590 nand P2_U2392 P2_R2099_U87 ; P2_U6710
g10591 nand P2_U2383 P2_R2337_U84 ; P2_U6711
g10592 nand P2_R1957_U9 P2_U2382 ; P2_U6712
g10593 nand P2_U2378 P2_PHYADDRPOINTER_REG_16__SCAN_IN ; P2_U6713
g10594 nand P2_U6570 P2_REIP_REG_16__SCAN_IN ; P2_U6714
g10595 nand P2_R2267_U9 P2_U2587 ; P2_U6715
g10596 nand P2_U2588 P2_R2096_U90 ; P2_U6716
g10597 nand P2_U7743 P2_EBX_REG_17__SCAN_IN ; P2_U6717
g10598 nand P2_U2392 P2_R2099_U86 ; P2_U6718
g10599 nand P2_U2383 P2_R2337_U83 ; P2_U6719
g10600 nand P2_R1957_U76 P2_U2382 ; P2_U6720
g10601 nand P2_U2378 P2_PHYADDRPOINTER_REG_17__SCAN_IN ; P2_U6721
g10602 nand P2_U6570 P2_REIP_REG_17__SCAN_IN ; P2_U6722
g10603 nand P2_R2267_U79 P2_U2587 ; P2_U6723
g10604 nand P2_U2588 P2_R2096_U89 ; P2_U6724
g10605 nand P2_U7743 P2_EBX_REG_18__SCAN_IN ; P2_U6725
g10606 nand P2_U2392 P2_R2099_U85 ; P2_U6726
g10607 nand P2_U2383 P2_R2337_U82 ; P2_U6727
g10608 nand P2_R1957_U10 P2_U2382 ; P2_U6728
g10609 nand P2_U2378 P2_PHYADDRPOINTER_REG_18__SCAN_IN ; P2_U6729
g10610 nand P2_U6570 P2_REIP_REG_18__SCAN_IN ; P2_U6730
g10611 nand P2_R2267_U10 P2_U2587 ; P2_U6731
g10612 nand P2_U2588 P2_R2096_U88 ; P2_U6732
g10613 nand P2_U7743 P2_EBX_REG_19__SCAN_IN ; P2_U6733
g10614 nand P2_U2392 P2_R2099_U84 ; P2_U6734
g10615 nand P2_U2383 P2_R2337_U81 ; P2_U6735
g10616 nand P2_R1957_U74 P2_U2382 ; P2_U6736
g10617 nand P2_U2378 P2_PHYADDRPOINTER_REG_19__SCAN_IN ; P2_U6737
g10618 nand P2_U6570 P2_REIP_REG_19__SCAN_IN ; P2_U6738
g10619 nand P2_R2267_U75 P2_U2587 ; P2_U6739
g10620 nand P2_U2588 P2_R2096_U87 ; P2_U6740
g10621 nand P2_U7743 P2_EBX_REG_20__SCAN_IN ; P2_U6741
g10622 nand P2_U2392 P2_R2099_U83 ; P2_U6742
g10623 nand P2_U2383 P2_R2337_U80 ; P2_U6743
g10624 nand P2_R1957_U11 P2_U2382 ; P2_U6744
g10625 nand P2_U2378 P2_PHYADDRPOINTER_REG_20__SCAN_IN ; P2_U6745
g10626 nand P2_U6570 P2_REIP_REG_20__SCAN_IN ; P2_U6746
g10627 nand P2_R2267_U11 P2_U2587 ; P2_U6747
g10628 nand P2_U2588 P2_R2096_U86 ; P2_U6748
g10629 nand P2_U7743 P2_EBX_REG_21__SCAN_IN ; P2_U6749
g10630 nand P2_U2392 P2_R2099_U82 ; P2_U6750
g10631 nand P2_U2383 P2_R2337_U79 ; P2_U6751
g10632 nand P2_R1957_U70 P2_U2382 ; P2_U6752
g10633 nand P2_U2378 P2_PHYADDRPOINTER_REG_21__SCAN_IN ; P2_U6753
g10634 nand P2_U6570 P2_REIP_REG_21__SCAN_IN ; P2_U6754
g10635 nand P2_R2267_U73 P2_U2587 ; P2_U6755
g10636 nand P2_U2588 P2_R2096_U85 ; P2_U6756
g10637 nand P2_U7743 P2_EBX_REG_22__SCAN_IN ; P2_U6757
g10638 nand P2_U2392 P2_R2099_U81 ; P2_U6758
g10639 nand P2_U2383 P2_R2337_U78 ; P2_U6759
g10640 nand P2_R1957_U12 P2_U2382 ; P2_U6760
g10641 nand P2_U2378 P2_PHYADDRPOINTER_REG_22__SCAN_IN ; P2_U6761
g10642 nand P2_U6570 P2_REIP_REG_22__SCAN_IN ; P2_U6762
g10643 nand P2_R2267_U12 P2_U2587 ; P2_U6763
g10644 nand P2_U2588 P2_R2096_U84 ; P2_U6764
g10645 nand P2_U7743 P2_EBX_REG_23__SCAN_IN ; P2_U6765
g10646 nand P2_U2392 P2_R2099_U80 ; P2_U6766
g10647 nand P2_U2383 P2_R2337_U77 ; P2_U6767
g10648 nand P2_R1957_U68 P2_U2382 ; P2_U6768
g10649 nand P2_U2378 P2_PHYADDRPOINTER_REG_23__SCAN_IN ; P2_U6769
g10650 nand P2_U6570 P2_REIP_REG_23__SCAN_IN ; P2_U6770
g10651 nand P2_R2267_U71 P2_U2587 ; P2_U6771
g10652 nand P2_U2588 P2_R2096_U83 ; P2_U6772
g10653 nand P2_U7743 P2_EBX_REG_24__SCAN_IN ; P2_U6773
g10654 nand P2_U2392 P2_R2099_U79 ; P2_U6774
g10655 nand P2_U2383 P2_R2337_U76 ; P2_U6775
g10656 nand P2_R1957_U13 P2_U2382 ; P2_U6776
g10657 nand P2_U2378 P2_PHYADDRPOINTER_REG_24__SCAN_IN ; P2_U6777
g10658 nand P2_U6570 P2_REIP_REG_24__SCAN_IN ; P2_U6778
g10659 nand P2_R2267_U13 P2_U2587 ; P2_U6779
g10660 nand P2_U2588 P2_R2096_U82 ; P2_U6780
g10661 nand P2_U7743 P2_EBX_REG_25__SCAN_IN ; P2_U6781
g10662 nand P2_U2392 P2_R2099_U78 ; P2_U6782
g10663 nand P2_U2383 P2_R2337_U75 ; P2_U6783
g10664 nand P2_R1957_U66 P2_U2382 ; P2_U6784
g10665 nand P2_U2378 P2_PHYADDRPOINTER_REG_25__SCAN_IN ; P2_U6785
g10666 nand P2_U6570 P2_REIP_REG_25__SCAN_IN ; P2_U6786
g10667 nand P2_R2267_U69 P2_U2587 ; P2_U6787
g10668 nand P2_U2588 P2_R2096_U81 ; P2_U6788
g10669 nand P2_U7743 P2_EBX_REG_26__SCAN_IN ; P2_U6789
g10670 nand P2_U2392 P2_R2099_U77 ; P2_U6790
g10671 nand P2_U2383 P2_R2337_U74 ; P2_U6791
g10672 nand P2_R1957_U14 P2_U2382 ; P2_U6792
g10673 nand P2_U2378 P2_PHYADDRPOINTER_REG_26__SCAN_IN ; P2_U6793
g10674 nand P2_U6570 P2_REIP_REG_26__SCAN_IN ; P2_U6794
g10675 nand P2_R2267_U14 P2_U2587 ; P2_U6795
g10676 nand P2_U2588 P2_R2096_U80 ; P2_U6796
g10677 nand P2_U7743 P2_EBX_REG_27__SCAN_IN ; P2_U6797
g10678 nand P2_U2392 P2_R2099_U76 ; P2_U6798
g10679 nand P2_U2383 P2_R2337_U73 ; P2_U6799
g10680 nand P2_R1957_U64 P2_U2382 ; P2_U6800
g10681 nand P2_U2378 P2_PHYADDRPOINTER_REG_27__SCAN_IN ; P2_U6801
g10682 nand P2_U6570 P2_REIP_REG_27__SCAN_IN ; P2_U6802
g10683 nand P2_R2267_U67 P2_U2587 ; P2_U6803
g10684 nand P2_U2588 P2_R2096_U79 ; P2_U6804
g10685 nand P2_U7743 P2_EBX_REG_28__SCAN_IN ; P2_U6805
g10686 nand P2_U2392 P2_R2099_U75 ; P2_U6806
g10687 nand P2_U2383 P2_R2337_U72 ; P2_U6807
g10688 nand P2_R1957_U15 P2_U2382 ; P2_U6808
g10689 nand P2_U2378 P2_PHYADDRPOINTER_REG_28__SCAN_IN ; P2_U6809
g10690 nand P2_U6570 P2_REIP_REG_28__SCAN_IN ; P2_U6810
g10691 nand P2_R2267_U15 P2_U2587 ; P2_U6811
g10692 nand P2_U2588 P2_R2096_U78 ; P2_U6812
g10693 nand P2_U7743 P2_EBX_REG_29__SCAN_IN ; P2_U6813
g10694 nand P2_U2392 P2_R2099_U74 ; P2_U6814
g10695 nand P2_U2383 P2_R2337_U71 ; P2_U6815
g10696 nand P2_R1957_U16 P2_U2382 ; P2_U6816
g10697 nand P2_U2378 P2_PHYADDRPOINTER_REG_29__SCAN_IN ; P2_U6817
g10698 nand P2_U6570 P2_REIP_REG_29__SCAN_IN ; P2_U6818
g10699 nand P2_R2267_U16 P2_U2587 ; P2_U6819
g10700 nand P2_U2588 P2_R2096_U76 ; P2_U6820
g10701 nand P2_U7743 P2_EBX_REG_30__SCAN_IN ; P2_U6821
g10702 nand P2_U2392 P2_R2099_U73 ; P2_U6822
g10703 nand P2_U2383 P2_R2337_U69 ; P2_U6823
g10704 nand P2_R1957_U62 P2_U2382 ; P2_U6824
g10705 nand P2_U2378 P2_PHYADDRPOINTER_REG_30__SCAN_IN ; P2_U6825
g10706 nand P2_U6570 P2_REIP_REG_30__SCAN_IN ; P2_U6826
g10707 nand P2_R2267_U63 P2_U2587 ; P2_U6827
g10708 nand P2_U2588 P2_R2096_U50 ; P2_U6828
g10709 nand P2_U7743 P2_EBX_REG_31__SCAN_IN ; P2_U6829
g10710 nand P2_U2392 P2_R2099_U72 ; P2_U6830
g10711 nand P2_U2383 P2_R2337_U68 ; P2_U6831
g10712 nand P2_R1957_U50 P2_U2382 ; P2_U6832
g10713 nand P2_U2378 P2_PHYADDRPOINTER_REG_31__SCAN_IN ; P2_U6833
g10714 nand P2_U6570 P2_REIP_REG_31__SCAN_IN ; P2_U6834
g10715 nand P2_DATAWIDTH_REG_0__SCAN_IN P2_DATAWIDTH_REG_1__SCAN_IN ; P2_U6835
g10716 nand P2_U4477 P2_REIP_REG_0__SCAN_IN ; P2_U6836
g10717 nand P2_U3547 P2_BYTEENABLE_REG_1__SCAN_IN ; P2_U6837
g10718 not P2_U4400 ; P2_U6838
g10719 nand P2_U4426 P2_U4468 P2_U4399 ; P2_U6839
g10720 nand P2_U4400 P2_FLUSH_REG_SCAN_IN ; P2_U6840
g10721 nand P2_U4187 P2_U4467 ; P2_U6841
g10722 nand P2_U4466 P2_U3284 ; P2_U6842
g10723 not P2_U4402 ; P2_U6843
g10724 nand P2_U4411 P2_STATEBS16_REG_SCAN_IN ; P2_U6844
g10725 not P2_U2715 ; P2_U6845
g10726 nand P2_U2715 P2_U3536 ; P2_U6846
g10727 nand P2_U4411 P2_U3265 ; P2_U6847
g10728 nand P2_U4184 P2_U2356 ; P2_U6848
g10729 nand P2_U4418 P2_U6847 ; P2_U6849
g10730 nand U211 P2_U6846 ; P2_U6850
g10731 or P2_STATE2_REG_2__SCAN_IN P2_STATE2_REG_1__SCAN_IN ; P2_U6851
g10732 nand P2_U6851 P2_U6850 P2_U4186 ; P2_U6852
g10733 nand P2_U2374 P2_U2459 ; P2_U6853
g10734 nand P2_U6853 P2_CODEFETCH_REG_SCAN_IN ; P2_U6854
g10735 nand P2_U4461 P2_STATE2_REG_0__SCAN_IN ; P2_U6855
g10736 nand P2_STATE_REG_0__SCAN_IN P2_ADS_N_REG_SCAN_IN ; P2_U6856
g10737 not P2_U4403 ; P2_U6857
g10738 nand P2_U3286 P2_U3294 P2_STATE2_REG_2__SCAN_IN ; P2_U6858
g10739 nand P2_U4421 P2_U4468 P2_U4404 ; P2_U6859
g10740 nand P2_U4189 P2_U2446 ; P2_U6860
g10741 nand P2_U6859 P2_MEMORYFETCH_REG_SCAN_IN ; P2_U6861
g10742 nand P2_U2538 P2_INSTQUEUE_REG_8__7__SCAN_IN ; P2_U6862
g10743 nand P2_U2537 P2_INSTQUEUE_REG_9__7__SCAN_IN ; P2_U6863
g10744 nand P2_U2536 P2_INSTQUEUE_REG_10__7__SCAN_IN ; P2_U6864
g10745 nand P2_U2535 P2_INSTQUEUE_REG_11__7__SCAN_IN ; P2_U6865
g10746 nand P2_U2534 P2_INSTQUEUE_REG_12__7__SCAN_IN ; P2_U6866
g10747 nand P2_U2533 P2_INSTQUEUE_REG_13__7__SCAN_IN ; P2_U6867
g10748 nand P2_U2531 P2_INSTQUEUE_REG_14__7__SCAN_IN ; P2_U6868
g10749 nand P2_U2530 P2_INSTQUEUE_REG_15__7__SCAN_IN ; P2_U6869
g10750 nand P2_U2528 P2_INSTQUEUE_REG_7__7__SCAN_IN ; P2_U6870
g10751 nand P2_U2527 P2_INSTQUEUE_REG_6__7__SCAN_IN ; P2_U6871
g10752 nand P2_U2526 P2_INSTQUEUE_REG_5__7__SCAN_IN ; P2_U6872
g10753 nand P2_U2524 P2_INSTQUEUE_REG_4__7__SCAN_IN ; P2_U6873
g10754 nand P2_U2522 P2_INSTQUEUE_REG_3__7__SCAN_IN ; P2_U6874
g10755 nand P2_U2521 P2_INSTQUEUE_REG_2__7__SCAN_IN ; P2_U6875
g10756 nand P2_U2519 P2_INSTQUEUE_REG_1__7__SCAN_IN ; P2_U6876
g10757 nand P2_U2517 P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U6877
g10758 nand P2_U2562 P2_INSTQUEUE_REG_15__7__SCAN_IN ; P2_U6878
g10759 nand P2_U2561 P2_INSTQUEUE_REG_14__7__SCAN_IN ; P2_U6879
g10760 nand P2_U2560 P2_INSTQUEUE_REG_13__7__SCAN_IN ; P2_U6880
g10761 nand P2_U2559 P2_INSTQUEUE_REG_12__7__SCAN_IN ; P2_U6881
g10762 nand P2_U2558 P2_INSTQUEUE_REG_11__7__SCAN_IN ; P2_U6882
g10763 nand P2_U2557 P2_INSTQUEUE_REG_10__7__SCAN_IN ; P2_U6883
g10764 nand P2_U2555 P2_INSTQUEUE_REG_9__7__SCAN_IN ; P2_U6884
g10765 nand P2_U2554 P2_INSTQUEUE_REG_8__7__SCAN_IN ; P2_U6885
g10766 nand P2_U2552 P2_INSTQUEUE_REG_7__7__SCAN_IN ; P2_U6886
g10767 nand P2_U2551 P2_INSTQUEUE_REG_6__7__SCAN_IN ; P2_U6887
g10768 nand P2_U2550 P2_INSTQUEUE_REG_5__7__SCAN_IN ; P2_U6888
g10769 nand P2_U2548 P2_INSTQUEUE_REG_4__7__SCAN_IN ; P2_U6889
g10770 nand P2_U2546 P2_INSTQUEUE_REG_3__7__SCAN_IN ; P2_U6890
g10771 nand P2_U2545 P2_INSTQUEUE_REG_2__7__SCAN_IN ; P2_U6891
g10772 nand P2_U2543 P2_INSTQUEUE_REG_1__7__SCAN_IN ; P2_U6892
g10773 nand P2_U2541 P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U6893
g10774 nand P2_U2562 P2_INSTQUEUE_REG_15__6__SCAN_IN ; P2_U6894
g10775 nand P2_U2561 P2_INSTQUEUE_REG_14__6__SCAN_IN ; P2_U6895
g10776 nand P2_U2560 P2_INSTQUEUE_REG_13__6__SCAN_IN ; P2_U6896
g10777 nand P2_U2559 P2_INSTQUEUE_REG_12__6__SCAN_IN ; P2_U6897
g10778 nand P2_U2558 P2_INSTQUEUE_REG_11__6__SCAN_IN ; P2_U6898
g10779 nand P2_U2557 P2_INSTQUEUE_REG_10__6__SCAN_IN ; P2_U6899
g10780 nand P2_U2555 P2_INSTQUEUE_REG_9__6__SCAN_IN ; P2_U6900
g10781 nand P2_U2554 P2_INSTQUEUE_REG_8__6__SCAN_IN ; P2_U6901
g10782 nand P2_U2552 P2_INSTQUEUE_REG_7__6__SCAN_IN ; P2_U6902
g10783 nand P2_U2551 P2_INSTQUEUE_REG_6__6__SCAN_IN ; P2_U6903
g10784 nand P2_U2550 P2_INSTQUEUE_REG_5__6__SCAN_IN ; P2_U6904
g10785 nand P2_U2548 P2_INSTQUEUE_REG_4__6__SCAN_IN ; P2_U6905
g10786 nand P2_U2546 P2_INSTQUEUE_REG_3__6__SCAN_IN ; P2_U6906
g10787 nand P2_U2545 P2_INSTQUEUE_REG_2__6__SCAN_IN ; P2_U6907
g10788 nand P2_U2543 P2_INSTQUEUE_REG_1__6__SCAN_IN ; P2_U6908
g10789 nand P2_U2541 P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U6909
g10790 nand P2_U2562 P2_INSTQUEUE_REG_15__5__SCAN_IN ; P2_U6910
g10791 nand P2_U2561 P2_INSTQUEUE_REG_14__5__SCAN_IN ; P2_U6911
g10792 nand P2_U2560 P2_INSTQUEUE_REG_13__5__SCAN_IN ; P2_U6912
g10793 nand P2_U2559 P2_INSTQUEUE_REG_12__5__SCAN_IN ; P2_U6913
g10794 nand P2_U2558 P2_INSTQUEUE_REG_11__5__SCAN_IN ; P2_U6914
g10795 nand P2_U2557 P2_INSTQUEUE_REG_10__5__SCAN_IN ; P2_U6915
g10796 nand P2_U2555 P2_INSTQUEUE_REG_9__5__SCAN_IN ; P2_U6916
g10797 nand P2_U2554 P2_INSTQUEUE_REG_8__5__SCAN_IN ; P2_U6917
g10798 nand P2_U2552 P2_INSTQUEUE_REG_7__5__SCAN_IN ; P2_U6918
g10799 nand P2_U2551 P2_INSTQUEUE_REG_6__5__SCAN_IN ; P2_U6919
g10800 nand P2_U2550 P2_INSTQUEUE_REG_5__5__SCAN_IN ; P2_U6920
g10801 nand P2_U2548 P2_INSTQUEUE_REG_4__5__SCAN_IN ; P2_U6921
g10802 nand P2_U2546 P2_INSTQUEUE_REG_3__5__SCAN_IN ; P2_U6922
g10803 nand P2_U2545 P2_INSTQUEUE_REG_2__5__SCAN_IN ; P2_U6923
g10804 nand P2_U2543 P2_INSTQUEUE_REG_1__5__SCAN_IN ; P2_U6924
g10805 nand P2_U2541 P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U6925
g10806 nand P2_U2562 P2_INSTQUEUE_REG_15__4__SCAN_IN ; P2_U6926
g10807 nand P2_U2561 P2_INSTQUEUE_REG_14__4__SCAN_IN ; P2_U6927
g10808 nand P2_U2560 P2_INSTQUEUE_REG_13__4__SCAN_IN ; P2_U6928
g10809 nand P2_U2559 P2_INSTQUEUE_REG_12__4__SCAN_IN ; P2_U6929
g10810 nand P2_U2558 P2_INSTQUEUE_REG_11__4__SCAN_IN ; P2_U6930
g10811 nand P2_U2557 P2_INSTQUEUE_REG_10__4__SCAN_IN ; P2_U6931
g10812 nand P2_U2555 P2_INSTQUEUE_REG_9__4__SCAN_IN ; P2_U6932
g10813 nand P2_U2554 P2_INSTQUEUE_REG_8__4__SCAN_IN ; P2_U6933
g10814 nand P2_U2552 P2_INSTQUEUE_REG_7__4__SCAN_IN ; P2_U6934
g10815 nand P2_U2551 P2_INSTQUEUE_REG_6__4__SCAN_IN ; P2_U6935
g10816 nand P2_U2550 P2_INSTQUEUE_REG_5__4__SCAN_IN ; P2_U6936
g10817 nand P2_U2548 P2_INSTQUEUE_REG_4__4__SCAN_IN ; P2_U6937
g10818 nand P2_U2546 P2_INSTQUEUE_REG_3__4__SCAN_IN ; P2_U6938
g10819 nand P2_U2545 P2_INSTQUEUE_REG_2__4__SCAN_IN ; P2_U6939
g10820 nand P2_U2543 P2_INSTQUEUE_REG_1__4__SCAN_IN ; P2_U6940
g10821 nand P2_U2541 P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U6941
g10822 nand P2_U2562 P2_INSTQUEUE_REG_15__3__SCAN_IN ; P2_U6942
g10823 nand P2_U2561 P2_INSTQUEUE_REG_14__3__SCAN_IN ; P2_U6943
g10824 nand P2_U2560 P2_INSTQUEUE_REG_13__3__SCAN_IN ; P2_U6944
g10825 nand P2_U2559 P2_INSTQUEUE_REG_12__3__SCAN_IN ; P2_U6945
g10826 nand P2_U2558 P2_INSTQUEUE_REG_11__3__SCAN_IN ; P2_U6946
g10827 nand P2_U2557 P2_INSTQUEUE_REG_10__3__SCAN_IN ; P2_U6947
g10828 nand P2_U2555 P2_INSTQUEUE_REG_9__3__SCAN_IN ; P2_U6948
g10829 nand P2_U2554 P2_INSTQUEUE_REG_8__3__SCAN_IN ; P2_U6949
g10830 nand P2_U2552 P2_INSTQUEUE_REG_7__3__SCAN_IN ; P2_U6950
g10831 nand P2_U2551 P2_INSTQUEUE_REG_6__3__SCAN_IN ; P2_U6951
g10832 nand P2_U2550 P2_INSTQUEUE_REG_5__3__SCAN_IN ; P2_U6952
g10833 nand P2_U2548 P2_INSTQUEUE_REG_4__3__SCAN_IN ; P2_U6953
g10834 nand P2_U2546 P2_INSTQUEUE_REG_3__3__SCAN_IN ; P2_U6954
g10835 nand P2_U2545 P2_INSTQUEUE_REG_2__3__SCAN_IN ; P2_U6955
g10836 nand P2_U2543 P2_INSTQUEUE_REG_1__3__SCAN_IN ; P2_U6956
g10837 nand P2_U2541 P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U6957
g10838 nand P2_U2562 P2_INSTQUEUE_REG_15__2__SCAN_IN ; P2_U6958
g10839 nand P2_U2561 P2_INSTQUEUE_REG_14__2__SCAN_IN ; P2_U6959
g10840 nand P2_U2560 P2_INSTQUEUE_REG_13__2__SCAN_IN ; P2_U6960
g10841 nand P2_U2559 P2_INSTQUEUE_REG_12__2__SCAN_IN ; P2_U6961
g10842 nand P2_U2558 P2_INSTQUEUE_REG_11__2__SCAN_IN ; P2_U6962
g10843 nand P2_U2557 P2_INSTQUEUE_REG_10__2__SCAN_IN ; P2_U6963
g10844 nand P2_U2555 P2_INSTQUEUE_REG_9__2__SCAN_IN ; P2_U6964
g10845 nand P2_U2554 P2_INSTQUEUE_REG_8__2__SCAN_IN ; P2_U6965
g10846 nand P2_U2552 P2_INSTQUEUE_REG_7__2__SCAN_IN ; P2_U6966
g10847 nand P2_U2551 P2_INSTQUEUE_REG_6__2__SCAN_IN ; P2_U6967
g10848 nand P2_U2550 P2_INSTQUEUE_REG_5__2__SCAN_IN ; P2_U6968
g10849 nand P2_U2548 P2_INSTQUEUE_REG_4__2__SCAN_IN ; P2_U6969
g10850 nand P2_U2546 P2_INSTQUEUE_REG_3__2__SCAN_IN ; P2_U6970
g10851 nand P2_U2545 P2_INSTQUEUE_REG_2__2__SCAN_IN ; P2_U6971
g10852 nand P2_U2543 P2_INSTQUEUE_REG_1__2__SCAN_IN ; P2_U6972
g10853 nand P2_U2541 P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U6973
g10854 nand P2_U2562 P2_INSTQUEUE_REG_15__1__SCAN_IN ; P2_U6974
g10855 nand P2_U2561 P2_INSTQUEUE_REG_14__1__SCAN_IN ; P2_U6975
g10856 nand P2_U2560 P2_INSTQUEUE_REG_13__1__SCAN_IN ; P2_U6976
g10857 nand P2_U2559 P2_INSTQUEUE_REG_12__1__SCAN_IN ; P2_U6977
g10858 nand P2_U2558 P2_INSTQUEUE_REG_11__1__SCAN_IN ; P2_U6978
g10859 nand P2_U2557 P2_INSTQUEUE_REG_10__1__SCAN_IN ; P2_U6979
g10860 nand P2_U2555 P2_INSTQUEUE_REG_9__1__SCAN_IN ; P2_U6980
g10861 nand P2_U2554 P2_INSTQUEUE_REG_8__1__SCAN_IN ; P2_U6981
g10862 nand P2_U2552 P2_INSTQUEUE_REG_7__1__SCAN_IN ; P2_U6982
g10863 nand P2_U2551 P2_INSTQUEUE_REG_6__1__SCAN_IN ; P2_U6983
g10864 nand P2_U2550 P2_INSTQUEUE_REG_5__1__SCAN_IN ; P2_U6984
g10865 nand P2_U2548 P2_INSTQUEUE_REG_4__1__SCAN_IN ; P2_U6985
g10866 nand P2_U2546 P2_INSTQUEUE_REG_3__1__SCAN_IN ; P2_U6986
g10867 nand P2_U2545 P2_INSTQUEUE_REG_2__1__SCAN_IN ; P2_U6987
g10868 nand P2_U2543 P2_INSTQUEUE_REG_1__1__SCAN_IN ; P2_U6988
g10869 nand P2_U2541 P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U6989
g10870 nand P2_U2562 P2_INSTQUEUE_REG_15__0__SCAN_IN ; P2_U6990
g10871 nand P2_U2561 P2_INSTQUEUE_REG_14__0__SCAN_IN ; P2_U6991
g10872 nand P2_U2560 P2_INSTQUEUE_REG_13__0__SCAN_IN ; P2_U6992
g10873 nand P2_U2559 P2_INSTQUEUE_REG_12__0__SCAN_IN ; P2_U6993
g10874 nand P2_U2558 P2_INSTQUEUE_REG_11__0__SCAN_IN ; P2_U6994
g10875 nand P2_U2557 P2_INSTQUEUE_REG_10__0__SCAN_IN ; P2_U6995
g10876 nand P2_U2555 P2_INSTQUEUE_REG_9__0__SCAN_IN ; P2_U6996
g10877 nand P2_U2554 P2_INSTQUEUE_REG_8__0__SCAN_IN ; P2_U6997
g10878 nand P2_U2552 P2_INSTQUEUE_REG_7__0__SCAN_IN ; P2_U6998
g10879 nand P2_U2551 P2_INSTQUEUE_REG_6__0__SCAN_IN ; P2_U6999
g10880 nand P2_U2550 P2_INSTQUEUE_REG_5__0__SCAN_IN ; P2_U7000
g10881 nand P2_U2548 P2_INSTQUEUE_REG_4__0__SCAN_IN ; P2_U7001
g10882 nand P2_U2546 P2_INSTQUEUE_REG_3__0__SCAN_IN ; P2_U7002
g10883 nand P2_U2545 P2_INSTQUEUE_REG_2__0__SCAN_IN ; P2_U7003
g10884 nand P2_U2543 P2_INSTQUEUE_REG_1__0__SCAN_IN ; P2_U7004
g10885 nand P2_U2541 P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U7005
g10886 or P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U7006
g10887 not P2_U4405 ; P2_U7007
g10888 nand P2_U2586 P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U7008
g10889 nand P2_U2585 P2_INSTQUEUE_REG_1__7__SCAN_IN ; P2_U7009
g10890 nand P2_U2584 P2_INSTQUEUE_REG_2__7__SCAN_IN ; P2_U7010
g10891 nand P2_U2583 P2_INSTQUEUE_REG_3__7__SCAN_IN ; P2_U7011
g10892 nand P2_U2581 P2_INSTQUEUE_REG_4__7__SCAN_IN ; P2_U7012
g10893 nand P2_U2580 P2_INSTQUEUE_REG_5__7__SCAN_IN ; P2_U7013
g10894 nand P2_U2579 P2_INSTQUEUE_REG_6__7__SCAN_IN ; P2_U7014
g10895 nand P2_U2578 P2_INSTQUEUE_REG_7__7__SCAN_IN ; P2_U7015
g10896 nand P2_U2576 P2_INSTQUEUE_REG_8__7__SCAN_IN ; P2_U7016
g10897 nand P2_U2575 P2_INSTQUEUE_REG_9__7__SCAN_IN ; P2_U7017
g10898 nand P2_U2574 P2_INSTQUEUE_REG_10__7__SCAN_IN ; P2_U7018
g10899 nand P2_U2573 P2_INSTQUEUE_REG_11__7__SCAN_IN ; P2_U7019
g10900 nand P2_U2571 P2_INSTQUEUE_REG_12__7__SCAN_IN ; P2_U7020
g10901 nand P2_U2569 P2_INSTQUEUE_REG_13__7__SCAN_IN ; P2_U7021
g10902 nand P2_U2567 P2_INSTQUEUE_REG_14__7__SCAN_IN ; P2_U7022
g10903 nand P2_U2565 P2_INSTQUEUE_REG_15__7__SCAN_IN ; P2_U7023
g10904 nand P2_U2586 P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U7024
g10905 nand P2_U2585 P2_INSTQUEUE_REG_1__6__SCAN_IN ; P2_U7025
g10906 nand P2_U2584 P2_INSTQUEUE_REG_2__6__SCAN_IN ; P2_U7026
g10907 nand P2_U2583 P2_INSTQUEUE_REG_3__6__SCAN_IN ; P2_U7027
g10908 nand P2_U2581 P2_INSTQUEUE_REG_4__6__SCAN_IN ; P2_U7028
g10909 nand P2_U2580 P2_INSTQUEUE_REG_5__6__SCAN_IN ; P2_U7029
g10910 nand P2_U2579 P2_INSTQUEUE_REG_6__6__SCAN_IN ; P2_U7030
g10911 nand P2_U2578 P2_INSTQUEUE_REG_7__6__SCAN_IN ; P2_U7031
g10912 nand P2_U2576 P2_INSTQUEUE_REG_8__6__SCAN_IN ; P2_U7032
g10913 nand P2_U2575 P2_INSTQUEUE_REG_9__6__SCAN_IN ; P2_U7033
g10914 nand P2_U2574 P2_INSTQUEUE_REG_10__6__SCAN_IN ; P2_U7034
g10915 nand P2_U2573 P2_INSTQUEUE_REG_11__6__SCAN_IN ; P2_U7035
g10916 nand P2_U2571 P2_INSTQUEUE_REG_12__6__SCAN_IN ; P2_U7036
g10917 nand P2_U2569 P2_INSTQUEUE_REG_13__6__SCAN_IN ; P2_U7037
g10918 nand P2_U2567 P2_INSTQUEUE_REG_14__6__SCAN_IN ; P2_U7038
g10919 nand P2_U2565 P2_INSTQUEUE_REG_15__6__SCAN_IN ; P2_U7039
g10920 nand P2_U2586 P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U7040
g10921 nand P2_U2585 P2_INSTQUEUE_REG_1__5__SCAN_IN ; P2_U7041
g10922 nand P2_U2584 P2_INSTQUEUE_REG_2__5__SCAN_IN ; P2_U7042
g10923 nand P2_U2583 P2_INSTQUEUE_REG_3__5__SCAN_IN ; P2_U7043
g10924 nand P2_U2581 P2_INSTQUEUE_REG_4__5__SCAN_IN ; P2_U7044
g10925 nand P2_U2580 P2_INSTQUEUE_REG_5__5__SCAN_IN ; P2_U7045
g10926 nand P2_U2579 P2_INSTQUEUE_REG_6__5__SCAN_IN ; P2_U7046
g10927 nand P2_U2578 P2_INSTQUEUE_REG_7__5__SCAN_IN ; P2_U7047
g10928 nand P2_U2576 P2_INSTQUEUE_REG_8__5__SCAN_IN ; P2_U7048
g10929 nand P2_U2575 P2_INSTQUEUE_REG_9__5__SCAN_IN ; P2_U7049
g10930 nand P2_U2574 P2_INSTQUEUE_REG_10__5__SCAN_IN ; P2_U7050
g10931 nand P2_U2573 P2_INSTQUEUE_REG_11__5__SCAN_IN ; P2_U7051
g10932 nand P2_U2571 P2_INSTQUEUE_REG_12__5__SCAN_IN ; P2_U7052
g10933 nand P2_U2569 P2_INSTQUEUE_REG_13__5__SCAN_IN ; P2_U7053
g10934 nand P2_U2567 P2_INSTQUEUE_REG_14__5__SCAN_IN ; P2_U7054
g10935 nand P2_U2565 P2_INSTQUEUE_REG_15__5__SCAN_IN ; P2_U7055
g10936 nand P2_U2586 P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U7056
g10937 nand P2_U2585 P2_INSTQUEUE_REG_1__4__SCAN_IN ; P2_U7057
g10938 nand P2_U2584 P2_INSTQUEUE_REG_2__4__SCAN_IN ; P2_U7058
g10939 nand P2_U2583 P2_INSTQUEUE_REG_3__4__SCAN_IN ; P2_U7059
g10940 nand P2_U2581 P2_INSTQUEUE_REG_4__4__SCAN_IN ; P2_U7060
g10941 nand P2_U2580 P2_INSTQUEUE_REG_5__4__SCAN_IN ; P2_U7061
g10942 nand P2_U2579 P2_INSTQUEUE_REG_6__4__SCAN_IN ; P2_U7062
g10943 nand P2_U2578 P2_INSTQUEUE_REG_7__4__SCAN_IN ; P2_U7063
g10944 nand P2_U2576 P2_INSTQUEUE_REG_8__4__SCAN_IN ; P2_U7064
g10945 nand P2_U2575 P2_INSTQUEUE_REG_9__4__SCAN_IN ; P2_U7065
g10946 nand P2_U2574 P2_INSTQUEUE_REG_10__4__SCAN_IN ; P2_U7066
g10947 nand P2_U2573 P2_INSTQUEUE_REG_11__4__SCAN_IN ; P2_U7067
g10948 nand P2_U2571 P2_INSTQUEUE_REG_12__4__SCAN_IN ; P2_U7068
g10949 nand P2_U2569 P2_INSTQUEUE_REG_13__4__SCAN_IN ; P2_U7069
g10950 nand P2_U2567 P2_INSTQUEUE_REG_14__4__SCAN_IN ; P2_U7070
g10951 nand P2_U2565 P2_INSTQUEUE_REG_15__4__SCAN_IN ; P2_U7071
g10952 nand P2_U2586 P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U7072
g10953 nand P2_U2585 P2_INSTQUEUE_REG_1__3__SCAN_IN ; P2_U7073
g10954 nand P2_U2584 P2_INSTQUEUE_REG_2__3__SCAN_IN ; P2_U7074
g10955 nand P2_U2583 P2_INSTQUEUE_REG_3__3__SCAN_IN ; P2_U7075
g10956 nand P2_U2581 P2_INSTQUEUE_REG_4__3__SCAN_IN ; P2_U7076
g10957 nand P2_U2580 P2_INSTQUEUE_REG_5__3__SCAN_IN ; P2_U7077
g10958 nand P2_U2579 P2_INSTQUEUE_REG_6__3__SCAN_IN ; P2_U7078
g10959 nand P2_U2578 P2_INSTQUEUE_REG_7__3__SCAN_IN ; P2_U7079
g10960 nand P2_U2576 P2_INSTQUEUE_REG_8__3__SCAN_IN ; P2_U7080
g10961 nand P2_U2575 P2_INSTQUEUE_REG_9__3__SCAN_IN ; P2_U7081
g10962 nand P2_U2574 P2_INSTQUEUE_REG_10__3__SCAN_IN ; P2_U7082
g10963 nand P2_U2573 P2_INSTQUEUE_REG_11__3__SCAN_IN ; P2_U7083
g10964 nand P2_U2571 P2_INSTQUEUE_REG_12__3__SCAN_IN ; P2_U7084
g10965 nand P2_U2569 P2_INSTQUEUE_REG_13__3__SCAN_IN ; P2_U7085
g10966 nand P2_U2567 P2_INSTQUEUE_REG_14__3__SCAN_IN ; P2_U7086
g10967 nand P2_U2565 P2_INSTQUEUE_REG_15__3__SCAN_IN ; P2_U7087
g10968 nand P2_U2586 P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U7088
g10969 nand P2_U2585 P2_INSTQUEUE_REG_1__2__SCAN_IN ; P2_U7089
g10970 nand P2_U2584 P2_INSTQUEUE_REG_2__2__SCAN_IN ; P2_U7090
g10971 nand P2_U2583 P2_INSTQUEUE_REG_3__2__SCAN_IN ; P2_U7091
g10972 nand P2_U2581 P2_INSTQUEUE_REG_4__2__SCAN_IN ; P2_U7092
g10973 nand P2_U2580 P2_INSTQUEUE_REG_5__2__SCAN_IN ; P2_U7093
g10974 nand P2_U2579 P2_INSTQUEUE_REG_6__2__SCAN_IN ; P2_U7094
g10975 nand P2_U2578 P2_INSTQUEUE_REG_7__2__SCAN_IN ; P2_U7095
g10976 nand P2_U2576 P2_INSTQUEUE_REG_8__2__SCAN_IN ; P2_U7096
g10977 nand P2_U2575 P2_INSTQUEUE_REG_9__2__SCAN_IN ; P2_U7097
g10978 nand P2_U2574 P2_INSTQUEUE_REG_10__2__SCAN_IN ; P2_U7098
g10979 nand P2_U2573 P2_INSTQUEUE_REG_11__2__SCAN_IN ; P2_U7099
g10980 nand P2_U2571 P2_INSTQUEUE_REG_12__2__SCAN_IN ; P2_U7100
g10981 nand P2_U2569 P2_INSTQUEUE_REG_13__2__SCAN_IN ; P2_U7101
g10982 nand P2_U2567 P2_INSTQUEUE_REG_14__2__SCAN_IN ; P2_U7102
g10983 nand P2_U2565 P2_INSTQUEUE_REG_15__2__SCAN_IN ; P2_U7103
g10984 nand P2_U2586 P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U7104
g10985 nand P2_U2585 P2_INSTQUEUE_REG_1__1__SCAN_IN ; P2_U7105
g10986 nand P2_U2584 P2_INSTQUEUE_REG_2__1__SCAN_IN ; P2_U7106
g10987 nand P2_U2583 P2_INSTQUEUE_REG_3__1__SCAN_IN ; P2_U7107
g10988 nand P2_U2581 P2_INSTQUEUE_REG_4__1__SCAN_IN ; P2_U7108
g10989 nand P2_U2580 P2_INSTQUEUE_REG_5__1__SCAN_IN ; P2_U7109
g10990 nand P2_U2579 P2_INSTQUEUE_REG_6__1__SCAN_IN ; P2_U7110
g10991 nand P2_U2578 P2_INSTQUEUE_REG_7__1__SCAN_IN ; P2_U7111
g10992 nand P2_U2576 P2_INSTQUEUE_REG_8__1__SCAN_IN ; P2_U7112
g10993 nand P2_U2575 P2_INSTQUEUE_REG_9__1__SCAN_IN ; P2_U7113
g10994 nand P2_U2574 P2_INSTQUEUE_REG_10__1__SCAN_IN ; P2_U7114
g10995 nand P2_U2573 P2_INSTQUEUE_REG_11__1__SCAN_IN ; P2_U7115
g10996 nand P2_U2571 P2_INSTQUEUE_REG_12__1__SCAN_IN ; P2_U7116
g10997 nand P2_U2569 P2_INSTQUEUE_REG_13__1__SCAN_IN ; P2_U7117
g10998 nand P2_U2567 P2_INSTQUEUE_REG_14__1__SCAN_IN ; P2_U7118
g10999 nand P2_U2565 P2_INSTQUEUE_REG_15__1__SCAN_IN ; P2_U7119
g11000 nand P2_U2586 P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U7120
g11001 nand P2_U2585 P2_INSTQUEUE_REG_1__0__SCAN_IN ; P2_U7121
g11002 nand P2_U2584 P2_INSTQUEUE_REG_2__0__SCAN_IN ; P2_U7122
g11003 nand P2_U2583 P2_INSTQUEUE_REG_3__0__SCAN_IN ; P2_U7123
g11004 nand P2_U2581 P2_INSTQUEUE_REG_4__0__SCAN_IN ; P2_U7124
g11005 nand P2_U2580 P2_INSTQUEUE_REG_5__0__SCAN_IN ; P2_U7125
g11006 nand P2_U2579 P2_INSTQUEUE_REG_6__0__SCAN_IN ; P2_U7126
g11007 nand P2_U2578 P2_INSTQUEUE_REG_7__0__SCAN_IN ; P2_U7127
g11008 nand P2_U2576 P2_INSTQUEUE_REG_8__0__SCAN_IN ; P2_U7128
g11009 nand P2_U2575 P2_INSTQUEUE_REG_9__0__SCAN_IN ; P2_U7129
g11010 nand P2_U2574 P2_INSTQUEUE_REG_10__0__SCAN_IN ; P2_U7130
g11011 nand P2_U2573 P2_INSTQUEUE_REG_11__0__SCAN_IN ; P2_U7131
g11012 nand P2_U2571 P2_INSTQUEUE_REG_12__0__SCAN_IN ; P2_U7132
g11013 nand P2_U2569 P2_INSTQUEUE_REG_13__0__SCAN_IN ; P2_U7133
g11014 nand P2_U2567 P2_INSTQUEUE_REG_14__0__SCAN_IN ; P2_U7134
g11015 nand P2_U2565 P2_INSTQUEUE_REG_15__0__SCAN_IN ; P2_U7135
g11016 not P2_U3554 ; P2_U7136
g11017 nand P2_U7136 P2_U3300 ; P2_U7137
g11018 nand P2_U4467 P2_R2099_U95 ; P2_U7138
g11019 nand P2_U7137 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7139
g11020 nand P2_U4430 P2_U3428 ; P2_U7140
g11021 nand P2_ADD_402_1132_U23 P2_U2355 ; P2_U7141
g11022 nand P2_U2354 P2_U2606 ; P2_U7142
g11023 nand P2_U2605 P2_U2355 ; P2_U7143
g11024 nand P2_U2354 P2_U2605 ; P2_U7144
g11025 nand P2_U2604 P2_U2355 ; P2_U7145
g11026 nand P2_U2354 P2_U2604 ; P2_U7146
g11027 nand P2_U2603 P2_U2355 ; P2_U7147
g11028 nand P2_U2354 P2_U2603 ; P2_U7148
g11029 nand P2_U4467 P2_R2099_U96 ; P2_U7149
g11030 nand P2_U7137 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U7150
g11031 nand P2_U4430 P2_U3580 ; P2_U7151
g11032 nand P2_U2602 P2_U2355 ; P2_U7152
g11033 nand P2_U2354 P2_U2602 ; P2_U7153
g11034 nand P2_U2601 P2_U2355 ; P2_U7154
g11035 nand P2_U2354 P2_U2601 ; P2_U7155
g11036 nand P2_U2600 P2_U2355 ; P2_U7156
g11037 nand P2_U2354 P2_U2600 ; P2_U7157
g11038 nand P2_U2599 P2_U2355 ; P2_U7158
g11039 nand P2_U2354 P2_U2599 ; P2_U7159
g11040 nand P2_U4467 P2_R2099_U5 ; P2_U7160
g11041 nand P2_U7137 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U7161
g11042 nand P2_U4430 P2_U3243 ; P2_U7162
g11043 nand P2_U4467 P2_R2099_U94 ; P2_U7163
g11044 nand P2_U7137 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U7164
g11045 nand P2_U4430 P2_U3307 ; P2_U7165
g11046 nand P2_U2355 P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U7166
g11047 nand P2_U5517 P2_INSTQUEUE_REG_0__7__SCAN_IN ; P2_U7167
g11048 nand P2_U5460 P2_INSTQUEUE_REG_1__7__SCAN_IN ; P2_U7168
g11049 nand P2_U5402 P2_INSTQUEUE_REG_2__7__SCAN_IN ; P2_U7169
g11050 nand P2_U5345 P2_INSTQUEUE_REG_3__7__SCAN_IN ; P2_U7170
g11051 nand P2_U5287 P2_INSTQUEUE_REG_4__7__SCAN_IN ; P2_U7171
g11052 nand P2_U5230 P2_INSTQUEUE_REG_5__7__SCAN_IN ; P2_U7172
g11053 nand P2_U5172 P2_INSTQUEUE_REG_6__7__SCAN_IN ; P2_U7173
g11054 nand P2_U5116 P2_INSTQUEUE_REG_7__7__SCAN_IN ; P2_U7174
g11055 nand P2_U5059 P2_INSTQUEUE_REG_8__7__SCAN_IN ; P2_U7175
g11056 nand P2_U5002 P2_INSTQUEUE_REG_9__7__SCAN_IN ; P2_U7176
g11057 nand P2_U4944 P2_INSTQUEUE_REG_10__7__SCAN_IN ; P2_U7177
g11058 nand P2_U4887 P2_INSTQUEUE_REG_11__7__SCAN_IN ; P2_U7178
g11059 nand P2_U4829 P2_INSTQUEUE_REG_12__7__SCAN_IN ; P2_U7179
g11060 nand P2_U4772 P2_INSTQUEUE_REG_13__7__SCAN_IN ; P2_U7180
g11061 nand P2_U4713 P2_INSTQUEUE_REG_14__7__SCAN_IN ; P2_U7181
g11062 nand P2_U4653 P2_INSTQUEUE_REG_15__7__SCAN_IN ; P2_U7182
g11063 nand P2_U4280 P2_U4279 P2_U4278 P2_U4277 ; P2_U7183
g11064 nand P2_U5517 P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U7184
g11065 nand P2_U5460 P2_INSTQUEUE_REG_1__6__SCAN_IN ; P2_U7185
g11066 nand P2_U5402 P2_INSTQUEUE_REG_2__6__SCAN_IN ; P2_U7186
g11067 nand P2_U5345 P2_INSTQUEUE_REG_3__6__SCAN_IN ; P2_U7187
g11068 nand P2_U5287 P2_INSTQUEUE_REG_4__6__SCAN_IN ; P2_U7188
g11069 nand P2_U5230 P2_INSTQUEUE_REG_5__6__SCAN_IN ; P2_U7189
g11070 nand P2_U5172 P2_INSTQUEUE_REG_6__6__SCAN_IN ; P2_U7190
g11071 nand P2_U5116 P2_INSTQUEUE_REG_7__6__SCAN_IN ; P2_U7191
g11072 nand P2_U5059 P2_INSTQUEUE_REG_8__6__SCAN_IN ; P2_U7192
g11073 nand P2_U5002 P2_INSTQUEUE_REG_9__6__SCAN_IN ; P2_U7193
g11074 nand P2_U4944 P2_INSTQUEUE_REG_10__6__SCAN_IN ; P2_U7194
g11075 nand P2_U4887 P2_INSTQUEUE_REG_11__6__SCAN_IN ; P2_U7195
g11076 nand P2_U4829 P2_INSTQUEUE_REG_12__6__SCAN_IN ; P2_U7196
g11077 nand P2_U4772 P2_INSTQUEUE_REG_13__6__SCAN_IN ; P2_U7197
g11078 nand P2_U4713 P2_INSTQUEUE_REG_14__6__SCAN_IN ; P2_U7198
g11079 nand P2_U4653 P2_INSTQUEUE_REG_15__6__SCAN_IN ; P2_U7199
g11080 nand P2_U4284 P2_U4283 P2_U4282 P2_U4281 ; P2_U7200
g11081 nand P2_U2538 P2_INSTQUEUE_REG_8__6__SCAN_IN ; P2_U7201
g11082 nand P2_U2537 P2_INSTQUEUE_REG_9__6__SCAN_IN ; P2_U7202
g11083 nand P2_U2536 P2_INSTQUEUE_REG_10__6__SCAN_IN ; P2_U7203
g11084 nand P2_U2535 P2_INSTQUEUE_REG_11__6__SCAN_IN ; P2_U7204
g11085 nand P2_U2534 P2_INSTQUEUE_REG_12__6__SCAN_IN ; P2_U7205
g11086 nand P2_U2533 P2_INSTQUEUE_REG_13__6__SCAN_IN ; P2_U7206
g11087 nand P2_U2531 P2_INSTQUEUE_REG_14__6__SCAN_IN ; P2_U7207
g11088 nand P2_U2530 P2_INSTQUEUE_REG_15__6__SCAN_IN ; P2_U7208
g11089 nand P2_U2528 P2_INSTQUEUE_REG_7__6__SCAN_IN ; P2_U7209
g11090 nand P2_U2527 P2_INSTQUEUE_REG_6__6__SCAN_IN ; P2_U7210
g11091 nand P2_U2526 P2_INSTQUEUE_REG_5__6__SCAN_IN ; P2_U7211
g11092 nand P2_U2524 P2_INSTQUEUE_REG_4__6__SCAN_IN ; P2_U7212
g11093 nand P2_U2522 P2_INSTQUEUE_REG_3__6__SCAN_IN ; P2_U7213
g11094 nand P2_U2521 P2_INSTQUEUE_REG_2__6__SCAN_IN ; P2_U7214
g11095 nand P2_U2519 P2_INSTQUEUE_REG_1__6__SCAN_IN ; P2_U7215
g11096 nand P2_U2517 P2_INSTQUEUE_REG_0__6__SCAN_IN ; P2_U7216
g11097 nand P2_U4288 P2_U4287 P2_U4286 P2_U4285 ; P2_U7217
g11098 nand P2_U5517 P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U7218
g11099 nand P2_U5460 P2_INSTQUEUE_REG_1__5__SCAN_IN ; P2_U7219
g11100 nand P2_U5402 P2_INSTQUEUE_REG_2__5__SCAN_IN ; P2_U7220
g11101 nand P2_U5345 P2_INSTQUEUE_REG_3__5__SCAN_IN ; P2_U7221
g11102 nand P2_U5287 P2_INSTQUEUE_REG_4__5__SCAN_IN ; P2_U7222
g11103 nand P2_U5230 P2_INSTQUEUE_REG_5__5__SCAN_IN ; P2_U7223
g11104 nand P2_U5172 P2_INSTQUEUE_REG_6__5__SCAN_IN ; P2_U7224
g11105 nand P2_U5116 P2_INSTQUEUE_REG_7__5__SCAN_IN ; P2_U7225
g11106 nand P2_U5059 P2_INSTQUEUE_REG_8__5__SCAN_IN ; P2_U7226
g11107 nand P2_U5002 P2_INSTQUEUE_REG_9__5__SCAN_IN ; P2_U7227
g11108 nand P2_U4944 P2_INSTQUEUE_REG_10__5__SCAN_IN ; P2_U7228
g11109 nand P2_U4887 P2_INSTQUEUE_REG_11__5__SCAN_IN ; P2_U7229
g11110 nand P2_U4829 P2_INSTQUEUE_REG_12__5__SCAN_IN ; P2_U7230
g11111 nand P2_U4772 P2_INSTQUEUE_REG_13__5__SCAN_IN ; P2_U7231
g11112 nand P2_U4713 P2_INSTQUEUE_REG_14__5__SCAN_IN ; P2_U7232
g11113 nand P2_U4653 P2_INSTQUEUE_REG_15__5__SCAN_IN ; P2_U7233
g11114 nand P2_U4292 P2_U4291 P2_U4290 P2_U4289 ; P2_U7234
g11115 nand P2_U2538 P2_INSTQUEUE_REG_8__5__SCAN_IN ; P2_U7235
g11116 nand P2_U2537 P2_INSTQUEUE_REG_9__5__SCAN_IN ; P2_U7236
g11117 nand P2_U2536 P2_INSTQUEUE_REG_10__5__SCAN_IN ; P2_U7237
g11118 nand P2_U2535 P2_INSTQUEUE_REG_11__5__SCAN_IN ; P2_U7238
g11119 nand P2_U2534 P2_INSTQUEUE_REG_12__5__SCAN_IN ; P2_U7239
g11120 nand P2_U2533 P2_INSTQUEUE_REG_13__5__SCAN_IN ; P2_U7240
g11121 nand P2_U2531 P2_INSTQUEUE_REG_14__5__SCAN_IN ; P2_U7241
g11122 nand P2_U2530 P2_INSTQUEUE_REG_15__5__SCAN_IN ; P2_U7242
g11123 nand P2_U2528 P2_INSTQUEUE_REG_7__5__SCAN_IN ; P2_U7243
g11124 nand P2_U2527 P2_INSTQUEUE_REG_6__5__SCAN_IN ; P2_U7244
g11125 nand P2_U2526 P2_INSTQUEUE_REG_5__5__SCAN_IN ; P2_U7245
g11126 nand P2_U2524 P2_INSTQUEUE_REG_4__5__SCAN_IN ; P2_U7246
g11127 nand P2_U2522 P2_INSTQUEUE_REG_3__5__SCAN_IN ; P2_U7247
g11128 nand P2_U2521 P2_INSTQUEUE_REG_2__5__SCAN_IN ; P2_U7248
g11129 nand P2_U2519 P2_INSTQUEUE_REG_1__5__SCAN_IN ; P2_U7249
g11130 nand P2_U2517 P2_INSTQUEUE_REG_0__5__SCAN_IN ; P2_U7250
g11131 nand P2_U4296 P2_U4295 P2_U4294 P2_U4293 ; P2_U7251
g11132 nand P2_U5517 P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U7252
g11133 nand P2_U5460 P2_INSTQUEUE_REG_1__4__SCAN_IN ; P2_U7253
g11134 nand P2_U5402 P2_INSTQUEUE_REG_2__4__SCAN_IN ; P2_U7254
g11135 nand P2_U5345 P2_INSTQUEUE_REG_3__4__SCAN_IN ; P2_U7255
g11136 nand P2_U5287 P2_INSTQUEUE_REG_4__4__SCAN_IN ; P2_U7256
g11137 nand P2_U5230 P2_INSTQUEUE_REG_5__4__SCAN_IN ; P2_U7257
g11138 nand P2_U5172 P2_INSTQUEUE_REG_6__4__SCAN_IN ; P2_U7258
g11139 nand P2_U5116 P2_INSTQUEUE_REG_7__4__SCAN_IN ; P2_U7259
g11140 nand P2_U5059 P2_INSTQUEUE_REG_8__4__SCAN_IN ; P2_U7260
g11141 nand P2_U5002 P2_INSTQUEUE_REG_9__4__SCAN_IN ; P2_U7261
g11142 nand P2_U4944 P2_INSTQUEUE_REG_10__4__SCAN_IN ; P2_U7262
g11143 nand P2_U4887 P2_INSTQUEUE_REG_11__4__SCAN_IN ; P2_U7263
g11144 nand P2_U4829 P2_INSTQUEUE_REG_12__4__SCAN_IN ; P2_U7264
g11145 nand P2_U4772 P2_INSTQUEUE_REG_13__4__SCAN_IN ; P2_U7265
g11146 nand P2_U4713 P2_INSTQUEUE_REG_14__4__SCAN_IN ; P2_U7266
g11147 nand P2_U4653 P2_INSTQUEUE_REG_15__4__SCAN_IN ; P2_U7267
g11148 nand P2_U4300 P2_U4299 P2_U4298 P2_U4297 ; P2_U7268
g11149 nand P2_U2538 P2_INSTQUEUE_REG_8__4__SCAN_IN ; P2_U7269
g11150 nand P2_U2537 P2_INSTQUEUE_REG_9__4__SCAN_IN ; P2_U7270
g11151 nand P2_U2536 P2_INSTQUEUE_REG_10__4__SCAN_IN ; P2_U7271
g11152 nand P2_U2535 P2_INSTQUEUE_REG_11__4__SCAN_IN ; P2_U7272
g11153 nand P2_U2534 P2_INSTQUEUE_REG_12__4__SCAN_IN ; P2_U7273
g11154 nand P2_U2533 P2_INSTQUEUE_REG_13__4__SCAN_IN ; P2_U7274
g11155 nand P2_U2531 P2_INSTQUEUE_REG_14__4__SCAN_IN ; P2_U7275
g11156 nand P2_U2530 P2_INSTQUEUE_REG_15__4__SCAN_IN ; P2_U7276
g11157 nand P2_U2528 P2_INSTQUEUE_REG_7__4__SCAN_IN ; P2_U7277
g11158 nand P2_U2527 P2_INSTQUEUE_REG_6__4__SCAN_IN ; P2_U7278
g11159 nand P2_U2526 P2_INSTQUEUE_REG_5__4__SCAN_IN ; P2_U7279
g11160 nand P2_U2524 P2_INSTQUEUE_REG_4__4__SCAN_IN ; P2_U7280
g11161 nand P2_U2522 P2_INSTQUEUE_REG_3__4__SCAN_IN ; P2_U7281
g11162 nand P2_U2521 P2_INSTQUEUE_REG_2__4__SCAN_IN ; P2_U7282
g11163 nand P2_U2519 P2_INSTQUEUE_REG_1__4__SCAN_IN ; P2_U7283
g11164 nand P2_U2517 P2_INSTQUEUE_REG_0__4__SCAN_IN ; P2_U7284
g11165 nand P2_U4304 P2_U4303 P2_U4302 P2_U4301 ; P2_U7285
g11166 nand P2_U5517 P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U7286
g11167 nand P2_U5460 P2_INSTQUEUE_REG_1__3__SCAN_IN ; P2_U7287
g11168 nand P2_U5402 P2_INSTQUEUE_REG_2__3__SCAN_IN ; P2_U7288
g11169 nand P2_U5345 P2_INSTQUEUE_REG_3__3__SCAN_IN ; P2_U7289
g11170 nand P2_U5287 P2_INSTQUEUE_REG_4__3__SCAN_IN ; P2_U7290
g11171 nand P2_U5230 P2_INSTQUEUE_REG_5__3__SCAN_IN ; P2_U7291
g11172 nand P2_U5172 P2_INSTQUEUE_REG_6__3__SCAN_IN ; P2_U7292
g11173 nand P2_U5116 P2_INSTQUEUE_REG_7__3__SCAN_IN ; P2_U7293
g11174 nand P2_U5059 P2_INSTQUEUE_REG_8__3__SCAN_IN ; P2_U7294
g11175 nand P2_U5002 P2_INSTQUEUE_REG_9__3__SCAN_IN ; P2_U7295
g11176 nand P2_U4944 P2_INSTQUEUE_REG_10__3__SCAN_IN ; P2_U7296
g11177 nand P2_U4887 P2_INSTQUEUE_REG_11__3__SCAN_IN ; P2_U7297
g11178 nand P2_U4829 P2_INSTQUEUE_REG_12__3__SCAN_IN ; P2_U7298
g11179 nand P2_U4772 P2_INSTQUEUE_REG_13__3__SCAN_IN ; P2_U7299
g11180 nand P2_U4713 P2_INSTQUEUE_REG_14__3__SCAN_IN ; P2_U7300
g11181 nand P2_U4653 P2_INSTQUEUE_REG_15__3__SCAN_IN ; P2_U7301
g11182 nand P2_U4308 P2_U4307 P2_U4306 P2_U4305 ; P2_U7302
g11183 nand P2_U2538 P2_INSTQUEUE_REG_8__3__SCAN_IN ; P2_U7303
g11184 nand P2_U2537 P2_INSTQUEUE_REG_9__3__SCAN_IN ; P2_U7304
g11185 nand P2_U2536 P2_INSTQUEUE_REG_10__3__SCAN_IN ; P2_U7305
g11186 nand P2_U2535 P2_INSTQUEUE_REG_11__3__SCAN_IN ; P2_U7306
g11187 nand P2_U2534 P2_INSTQUEUE_REG_12__3__SCAN_IN ; P2_U7307
g11188 nand P2_U2533 P2_INSTQUEUE_REG_13__3__SCAN_IN ; P2_U7308
g11189 nand P2_U2531 P2_INSTQUEUE_REG_14__3__SCAN_IN ; P2_U7309
g11190 nand P2_U2530 P2_INSTQUEUE_REG_15__3__SCAN_IN ; P2_U7310
g11191 nand P2_U2528 P2_INSTQUEUE_REG_7__3__SCAN_IN ; P2_U7311
g11192 nand P2_U2527 P2_INSTQUEUE_REG_6__3__SCAN_IN ; P2_U7312
g11193 nand P2_U2526 P2_INSTQUEUE_REG_5__3__SCAN_IN ; P2_U7313
g11194 nand P2_U2524 P2_INSTQUEUE_REG_4__3__SCAN_IN ; P2_U7314
g11195 nand P2_U2522 P2_INSTQUEUE_REG_3__3__SCAN_IN ; P2_U7315
g11196 nand P2_U2521 P2_INSTQUEUE_REG_2__3__SCAN_IN ; P2_U7316
g11197 nand P2_U2519 P2_INSTQUEUE_REG_1__3__SCAN_IN ; P2_U7317
g11198 nand P2_U2517 P2_INSTQUEUE_REG_0__3__SCAN_IN ; P2_U7318
g11199 nand P2_U4312 P2_U4311 P2_U4310 P2_U4309 ; P2_U7319
g11200 nand P2_U5517 P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U7320
g11201 nand P2_U5460 P2_INSTQUEUE_REG_1__2__SCAN_IN ; P2_U7321
g11202 nand P2_U5402 P2_INSTQUEUE_REG_2__2__SCAN_IN ; P2_U7322
g11203 nand P2_U5345 P2_INSTQUEUE_REG_3__2__SCAN_IN ; P2_U7323
g11204 nand P2_U5287 P2_INSTQUEUE_REG_4__2__SCAN_IN ; P2_U7324
g11205 nand P2_U5230 P2_INSTQUEUE_REG_5__2__SCAN_IN ; P2_U7325
g11206 nand P2_U5172 P2_INSTQUEUE_REG_6__2__SCAN_IN ; P2_U7326
g11207 nand P2_U5116 P2_INSTQUEUE_REG_7__2__SCAN_IN ; P2_U7327
g11208 nand P2_U5059 P2_INSTQUEUE_REG_8__2__SCAN_IN ; P2_U7328
g11209 nand P2_U5002 P2_INSTQUEUE_REG_9__2__SCAN_IN ; P2_U7329
g11210 nand P2_U4944 P2_INSTQUEUE_REG_10__2__SCAN_IN ; P2_U7330
g11211 nand P2_U4887 P2_INSTQUEUE_REG_11__2__SCAN_IN ; P2_U7331
g11212 nand P2_U4829 P2_INSTQUEUE_REG_12__2__SCAN_IN ; P2_U7332
g11213 nand P2_U4772 P2_INSTQUEUE_REG_13__2__SCAN_IN ; P2_U7333
g11214 nand P2_U4713 P2_INSTQUEUE_REG_14__2__SCAN_IN ; P2_U7334
g11215 nand P2_U4653 P2_INSTQUEUE_REG_15__2__SCAN_IN ; P2_U7335
g11216 nand P2_U4316 P2_U4315 P2_U4314 P2_U4313 ; P2_U7336
g11217 nand P2_U2538 P2_INSTQUEUE_REG_8__2__SCAN_IN ; P2_U7337
g11218 nand P2_U2537 P2_INSTQUEUE_REG_9__2__SCAN_IN ; P2_U7338
g11219 nand P2_U2536 P2_INSTQUEUE_REG_10__2__SCAN_IN ; P2_U7339
g11220 nand P2_U2535 P2_INSTQUEUE_REG_11__2__SCAN_IN ; P2_U7340
g11221 nand P2_U2534 P2_INSTQUEUE_REG_12__2__SCAN_IN ; P2_U7341
g11222 nand P2_U2533 P2_INSTQUEUE_REG_13__2__SCAN_IN ; P2_U7342
g11223 nand P2_U2531 P2_INSTQUEUE_REG_14__2__SCAN_IN ; P2_U7343
g11224 nand P2_U2530 P2_INSTQUEUE_REG_15__2__SCAN_IN ; P2_U7344
g11225 nand P2_U2528 P2_INSTQUEUE_REG_7__2__SCAN_IN ; P2_U7345
g11226 nand P2_U2527 P2_INSTQUEUE_REG_6__2__SCAN_IN ; P2_U7346
g11227 nand P2_U2526 P2_INSTQUEUE_REG_5__2__SCAN_IN ; P2_U7347
g11228 nand P2_U2524 P2_INSTQUEUE_REG_4__2__SCAN_IN ; P2_U7348
g11229 nand P2_U2522 P2_INSTQUEUE_REG_3__2__SCAN_IN ; P2_U7349
g11230 nand P2_U2521 P2_INSTQUEUE_REG_2__2__SCAN_IN ; P2_U7350
g11231 nand P2_U2519 P2_INSTQUEUE_REG_1__2__SCAN_IN ; P2_U7351
g11232 nand P2_U2517 P2_INSTQUEUE_REG_0__2__SCAN_IN ; P2_U7352
g11233 nand P2_U4320 P2_U4319 P2_U4318 P2_U4317 ; P2_U7353
g11234 nand P2_U5517 P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U7354
g11235 nand P2_U5460 P2_INSTQUEUE_REG_1__1__SCAN_IN ; P2_U7355
g11236 nand P2_U5402 P2_INSTQUEUE_REG_2__1__SCAN_IN ; P2_U7356
g11237 nand P2_U5345 P2_INSTQUEUE_REG_3__1__SCAN_IN ; P2_U7357
g11238 nand P2_U5287 P2_INSTQUEUE_REG_4__1__SCAN_IN ; P2_U7358
g11239 nand P2_U5230 P2_INSTQUEUE_REG_5__1__SCAN_IN ; P2_U7359
g11240 nand P2_U5172 P2_INSTQUEUE_REG_6__1__SCAN_IN ; P2_U7360
g11241 nand P2_U5116 P2_INSTQUEUE_REG_7__1__SCAN_IN ; P2_U7361
g11242 nand P2_U5059 P2_INSTQUEUE_REG_8__1__SCAN_IN ; P2_U7362
g11243 nand P2_U5002 P2_INSTQUEUE_REG_9__1__SCAN_IN ; P2_U7363
g11244 nand P2_U4944 P2_INSTQUEUE_REG_10__1__SCAN_IN ; P2_U7364
g11245 nand P2_U4887 P2_INSTQUEUE_REG_11__1__SCAN_IN ; P2_U7365
g11246 nand P2_U4829 P2_INSTQUEUE_REG_12__1__SCAN_IN ; P2_U7366
g11247 nand P2_U4772 P2_INSTQUEUE_REG_13__1__SCAN_IN ; P2_U7367
g11248 nand P2_U4713 P2_INSTQUEUE_REG_14__1__SCAN_IN ; P2_U7368
g11249 nand P2_U4653 P2_INSTQUEUE_REG_15__1__SCAN_IN ; P2_U7369
g11250 nand P2_U4324 P2_U4323 P2_U4322 P2_U4321 ; P2_U7370
g11251 nand P2_U2538 P2_INSTQUEUE_REG_8__1__SCAN_IN ; P2_U7371
g11252 nand P2_U2537 P2_INSTQUEUE_REG_9__1__SCAN_IN ; P2_U7372
g11253 nand P2_U2536 P2_INSTQUEUE_REG_10__1__SCAN_IN ; P2_U7373
g11254 nand P2_U2535 P2_INSTQUEUE_REG_11__1__SCAN_IN ; P2_U7374
g11255 nand P2_U2534 P2_INSTQUEUE_REG_12__1__SCAN_IN ; P2_U7375
g11256 nand P2_U2533 P2_INSTQUEUE_REG_13__1__SCAN_IN ; P2_U7376
g11257 nand P2_U2531 P2_INSTQUEUE_REG_14__1__SCAN_IN ; P2_U7377
g11258 nand P2_U2530 P2_INSTQUEUE_REG_15__1__SCAN_IN ; P2_U7378
g11259 nand P2_U2528 P2_INSTQUEUE_REG_7__1__SCAN_IN ; P2_U7379
g11260 nand P2_U2527 P2_INSTQUEUE_REG_6__1__SCAN_IN ; P2_U7380
g11261 nand P2_U2526 P2_INSTQUEUE_REG_5__1__SCAN_IN ; P2_U7381
g11262 nand P2_U2524 P2_INSTQUEUE_REG_4__1__SCAN_IN ; P2_U7382
g11263 nand P2_U2522 P2_INSTQUEUE_REG_3__1__SCAN_IN ; P2_U7383
g11264 nand P2_U2521 P2_INSTQUEUE_REG_2__1__SCAN_IN ; P2_U7384
g11265 nand P2_U2519 P2_INSTQUEUE_REG_1__1__SCAN_IN ; P2_U7385
g11266 nand P2_U2517 P2_INSTQUEUE_REG_0__1__SCAN_IN ; P2_U7386
g11267 nand P2_U4328 P2_U4327 P2_U4326 P2_U4325 ; P2_U7387
g11268 nand P2_U5517 P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U7388
g11269 nand P2_U5460 P2_INSTQUEUE_REG_1__0__SCAN_IN ; P2_U7389
g11270 nand P2_U5402 P2_INSTQUEUE_REG_2__0__SCAN_IN ; P2_U7390
g11271 nand P2_U5345 P2_INSTQUEUE_REG_3__0__SCAN_IN ; P2_U7391
g11272 nand P2_U5287 P2_INSTQUEUE_REG_4__0__SCAN_IN ; P2_U7392
g11273 nand P2_U5230 P2_INSTQUEUE_REG_5__0__SCAN_IN ; P2_U7393
g11274 nand P2_U5172 P2_INSTQUEUE_REG_6__0__SCAN_IN ; P2_U7394
g11275 nand P2_U5116 P2_INSTQUEUE_REG_7__0__SCAN_IN ; P2_U7395
g11276 nand P2_U5059 P2_INSTQUEUE_REG_8__0__SCAN_IN ; P2_U7396
g11277 nand P2_U5002 P2_INSTQUEUE_REG_9__0__SCAN_IN ; P2_U7397
g11278 nand P2_U4944 P2_INSTQUEUE_REG_10__0__SCAN_IN ; P2_U7398
g11279 nand P2_U4887 P2_INSTQUEUE_REG_11__0__SCAN_IN ; P2_U7399
g11280 nand P2_U4829 P2_INSTQUEUE_REG_12__0__SCAN_IN ; P2_U7400
g11281 nand P2_U4772 P2_INSTQUEUE_REG_13__0__SCAN_IN ; P2_U7401
g11282 nand P2_U4713 P2_INSTQUEUE_REG_14__0__SCAN_IN ; P2_U7402
g11283 nand P2_U4653 P2_INSTQUEUE_REG_15__0__SCAN_IN ; P2_U7403
g11284 nand P2_U4332 P2_U4331 P2_U4330 P2_U4329 ; P2_U7404
g11285 nand P2_U2538 P2_INSTQUEUE_REG_8__0__SCAN_IN ; P2_U7405
g11286 nand P2_U2537 P2_INSTQUEUE_REG_9__0__SCAN_IN ; P2_U7406
g11287 nand P2_U2536 P2_INSTQUEUE_REG_10__0__SCAN_IN ; P2_U7407
g11288 nand P2_U2535 P2_INSTQUEUE_REG_11__0__SCAN_IN ; P2_U7408
g11289 nand P2_U2534 P2_INSTQUEUE_REG_12__0__SCAN_IN ; P2_U7409
g11290 nand P2_U2533 P2_INSTQUEUE_REG_13__0__SCAN_IN ; P2_U7410
g11291 nand P2_U2531 P2_INSTQUEUE_REG_14__0__SCAN_IN ; P2_U7411
g11292 nand P2_U2530 P2_INSTQUEUE_REG_15__0__SCAN_IN ; P2_U7412
g11293 nand P2_U2528 P2_INSTQUEUE_REG_7__0__SCAN_IN ; P2_U7413
g11294 nand P2_U2527 P2_INSTQUEUE_REG_6__0__SCAN_IN ; P2_U7414
g11295 nand P2_U2526 P2_INSTQUEUE_REG_5__0__SCAN_IN ; P2_U7415
g11296 nand P2_U2524 P2_INSTQUEUE_REG_4__0__SCAN_IN ; P2_U7416
g11297 nand P2_U2522 P2_INSTQUEUE_REG_3__0__SCAN_IN ; P2_U7417
g11298 nand P2_U2521 P2_INSTQUEUE_REG_2__0__SCAN_IN ; P2_U7418
g11299 nand P2_U2519 P2_INSTQUEUE_REG_1__0__SCAN_IN ; P2_U7419
g11300 nand P2_U2517 P2_INSTQUEUE_REG_0__0__SCAN_IN ; P2_U7420
g11301 nand P2_U4336 P2_U4335 P2_U4334 P2_U4333 ; P2_U7421
g11302 nand P2_U2352 P2_U7319 ; P2_U7422
g11303 nand P2_STATE2_REG_3__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U7423
g11304 nand P2_U2352 P2_U7353 ; P2_U7424
g11305 nand P2_STATE2_REG_3__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U7425
g11306 nand P2_U2439 P2_U3295 ; P2_U7426
g11307 nand P2_U2352 P2_U7387 ; P2_U7427
g11308 nand P2_STATE2_REG_3__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_U7428
g11309 nand P2_U2352 P2_U7421 ; P2_U7429
g11310 nand P2_STATE2_REG_3__SCAN_IN P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U7430
g11311 nand P2_U2439 P2_U3279 ; P2_U7431
g11312 nand P2_U4414 P2_U7431 P2_U4413 ; P2_U7432
g11313 nand P2_U7432 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_U7433
g11314 nand P2_U2353 P2_REIP_REG_9__SCAN_IN ; P2_U7434
g11315 nand P2_U4412 P2_EAX_REG_9__SCAN_IN ; P2_U7435
g11316 nand P2_U2352 P2_U2608 ; P2_U7436
g11317 nand P2_U7432 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_U7437
g11318 nand P2_U2353 P2_REIP_REG_8__SCAN_IN ; P2_U7438
g11319 nand P2_U4412 P2_EAX_REG_8__SCAN_IN ; P2_U7439
g11320 nand P2_U2352 P2_U2607 ; P2_U7440
g11321 nand P2_U7432 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_U7441
g11322 nand P2_U2353 P2_REIP_REG_7__SCAN_IN ; P2_U7442
g11323 nand P2_U4412 P2_EAX_REG_7__SCAN_IN ; P2_U7443
g11324 nand P2_U7432 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_U7444
g11325 nand P2_U2353 P2_REIP_REG_6__SCAN_IN ; P2_U7445
g11326 nand P2_U4412 P2_EAX_REG_6__SCAN_IN ; P2_U7446
g11327 nand P2_U7432 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_U7447
g11328 nand P2_U2353 P2_REIP_REG_5__SCAN_IN ; P2_U7448
g11329 nand P2_U4412 P2_EAX_REG_5__SCAN_IN ; P2_U7449
g11330 nand P2_U7432 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_U7450
g11331 nand P2_U2353 P2_REIP_REG_4__SCAN_IN ; P2_U7451
g11332 nand P2_U4412 P2_EAX_REG_4__SCAN_IN ; P2_U7452
g11333 nand P2_U7432 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_U7453
g11334 nand P2_U2353 P2_REIP_REG_31__SCAN_IN ; P2_U7454
g11335 nand P2_U4412 P2_EAX_REG_31__SCAN_IN ; P2_U7455
g11336 nand P2_U7432 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_U7456
g11337 nand P2_U2353 P2_REIP_REG_30__SCAN_IN ; P2_U7457
g11338 nand P2_U4412 P2_EAX_REG_30__SCAN_IN ; P2_U7458
g11339 nand P2_U7432 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_U7459
g11340 nand P2_U2353 P2_REIP_REG_3__SCAN_IN ; P2_U7460
g11341 nand P2_U4412 P2_EAX_REG_3__SCAN_IN ; P2_U7461
g11342 nand P2_U7432 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_U7462
g11343 nand P2_U2353 P2_REIP_REG_29__SCAN_IN ; P2_U7463
g11344 nand P2_U4412 P2_EAX_REG_29__SCAN_IN ; P2_U7464
g11345 nand P2_U7432 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_U7465
g11346 nand P2_U2353 P2_REIP_REG_28__SCAN_IN ; P2_U7466
g11347 nand P2_U4412 P2_EAX_REG_28__SCAN_IN ; P2_U7467
g11348 nand P2_U7432 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_U7468
g11349 nand P2_U2353 P2_REIP_REG_27__SCAN_IN ; P2_U7469
g11350 nand P2_U4412 P2_EAX_REG_27__SCAN_IN ; P2_U7470
g11351 nand P2_U7432 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_U7471
g11352 nand P2_U2353 P2_REIP_REG_26__SCAN_IN ; P2_U7472
g11353 nand P2_U4412 P2_EAX_REG_26__SCAN_IN ; P2_U7473
g11354 nand P2_U7432 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_U7474
g11355 nand P2_U2353 P2_REIP_REG_25__SCAN_IN ; P2_U7475
g11356 nand P2_U4412 P2_EAX_REG_25__SCAN_IN ; P2_U7476
g11357 nand P2_U7432 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_U7477
g11358 nand P2_U2353 P2_REIP_REG_24__SCAN_IN ; P2_U7478
g11359 nand P2_U4412 P2_EAX_REG_24__SCAN_IN ; P2_U7479
g11360 nand P2_U7432 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_U7480
g11361 nand P2_U2353 P2_REIP_REG_23__SCAN_IN ; P2_U7481
g11362 nand P2_U4412 P2_EAX_REG_23__SCAN_IN ; P2_U7482
g11363 nand P2_U7432 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_U7483
g11364 nand P2_U2353 P2_REIP_REG_22__SCAN_IN ; P2_U7484
g11365 nand P2_U4412 P2_EAX_REG_22__SCAN_IN ; P2_U7485
g11366 nand P2_U7432 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_U7486
g11367 nand P2_U2353 P2_REIP_REG_21__SCAN_IN ; P2_U7487
g11368 nand P2_U4412 P2_EAX_REG_21__SCAN_IN ; P2_U7488
g11369 nand P2_U7432 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_U7489
g11370 nand P2_U2353 P2_REIP_REG_20__SCAN_IN ; P2_U7490
g11371 nand P2_U4412 P2_EAX_REG_20__SCAN_IN ; P2_U7491
g11372 nand P2_U7432 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_U7492
g11373 nand P2_U2353 P2_REIP_REG_2__SCAN_IN ; P2_U7493
g11374 nand P2_U4412 P2_EAX_REG_2__SCAN_IN ; P2_U7494
g11375 nand P2_U7432 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_U7495
g11376 nand P2_U2353 P2_REIP_REG_19__SCAN_IN ; P2_U7496
g11377 nand P2_U4412 P2_EAX_REG_19__SCAN_IN ; P2_U7497
g11378 nand P2_U7432 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_U7498
g11379 nand P2_U2353 P2_REIP_REG_18__SCAN_IN ; P2_U7499
g11380 nand P2_U4412 P2_EAX_REG_18__SCAN_IN ; P2_U7500
g11381 nand P2_U7432 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_U7501
g11382 nand P2_U2353 P2_REIP_REG_17__SCAN_IN ; P2_U7502
g11383 nand P2_U4412 P2_EAX_REG_17__SCAN_IN ; P2_U7503
g11384 nand P2_U7432 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_U7504
g11385 nand P2_U2353 P2_REIP_REG_16__SCAN_IN ; P2_U7505
g11386 nand P2_U4412 P2_EAX_REG_16__SCAN_IN ; P2_U7506
g11387 nand P2_U7432 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_U7507
g11388 nand P2_U2353 P2_REIP_REG_15__SCAN_IN ; P2_U7508
g11389 nand P2_U4412 P2_EAX_REG_15__SCAN_IN ; P2_U7509
g11390 nand P2_U2352 P2_U2614 ; P2_U7510
g11391 nand P2_U7432 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_U7511
g11392 nand P2_U2353 P2_REIP_REG_14__SCAN_IN ; P2_U7512
g11393 nand P2_U4412 P2_EAX_REG_14__SCAN_IN ; P2_U7513
g11394 nand P2_U2352 P2_U2613 ; P2_U7514
g11395 nand P2_U7432 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_U7515
g11396 nand P2_U2353 P2_REIP_REG_13__SCAN_IN ; P2_U7516
g11397 nand P2_U4412 P2_EAX_REG_13__SCAN_IN ; P2_U7517
g11398 nand P2_U2352 P2_U2612 ; P2_U7518
g11399 nand P2_U7432 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_U7519
g11400 nand P2_U2353 P2_REIP_REG_12__SCAN_IN ; P2_U7520
g11401 nand P2_U4412 P2_EAX_REG_12__SCAN_IN ; P2_U7521
g11402 nand P2_U2352 P2_U2611 ; P2_U7522
g11403 nand P2_U7432 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_U7523
g11404 nand P2_U2353 P2_REIP_REG_11__SCAN_IN ; P2_U7524
g11405 nand P2_U4412 P2_EAX_REG_11__SCAN_IN ; P2_U7525
g11406 nand P2_U2352 P2_U2610 ; P2_U7526
g11407 nand P2_U7432 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_U7527
g11408 nand P2_U2353 P2_REIP_REG_10__SCAN_IN ; P2_U7528
g11409 nand P2_U4412 P2_EAX_REG_10__SCAN_IN ; P2_U7529
g11410 nand P2_U2352 P2_U2609 ; P2_U7530
g11411 nand P2_U7432 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_U7531
g11412 nand P2_U2353 P2_REIP_REG_1__SCAN_IN ; P2_U7532
g11413 nand P2_U4412 P2_EAX_REG_1__SCAN_IN ; P2_U7533
g11414 nand P2_U7432 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_U7534
g11415 nand P2_U2353 P2_REIP_REG_0__SCAN_IN ; P2_U7535
g11416 nand P2_U4412 P2_EAX_REG_0__SCAN_IN ; P2_U7536
g11417 nand P2_U7869 P2_EBX_REG_9__SCAN_IN ; P2_U7537
g11418 nand P2_U7869 P2_EBX_REG_8__SCAN_IN ; P2_U7538
g11419 nand P2_U7869 P2_EBX_REG_31__SCAN_IN ; P2_U7539
g11420 nand P2_U7869 P2_EBX_REG_30__SCAN_IN ; P2_U7540
g11421 nand P2_U7869 P2_EBX_REG_29__SCAN_IN ; P2_U7541
g11422 nand P2_U7869 P2_EBX_REG_28__SCAN_IN ; P2_U7542
g11423 nand P2_U7869 P2_EBX_REG_27__SCAN_IN ; P2_U7543
g11424 nand P2_U7869 P2_EBX_REG_26__SCAN_IN ; P2_U7544
g11425 nand P2_U7869 P2_EBX_REG_25__SCAN_IN ; P2_U7545
g11426 nand P2_U7869 P2_EBX_REG_24__SCAN_IN ; P2_U7546
g11427 nand P2_U7869 P2_EBX_REG_23__SCAN_IN ; P2_U7547
g11428 nand P2_U7869 P2_EBX_REG_22__SCAN_IN ; P2_U7548
g11429 nand P2_U7869 P2_EBX_REG_21__SCAN_IN ; P2_U7549
g11430 nand P2_U7869 P2_EBX_REG_20__SCAN_IN ; P2_U7550
g11431 nand P2_U7869 P2_EBX_REG_19__SCAN_IN ; P2_U7551
g11432 nand P2_U7869 P2_EBX_REG_18__SCAN_IN ; P2_U7552
g11433 nand P2_U7869 P2_EBX_REG_17__SCAN_IN ; P2_U7553
g11434 nand P2_U7869 P2_EBX_REG_16__SCAN_IN ; P2_U7554
g11435 nand P2_U7869 P2_EBX_REG_15__SCAN_IN ; P2_U7555
g11436 nand P2_U7869 P2_EBX_REG_14__SCAN_IN ; P2_U7556
g11437 nand P2_U7869 P2_EBX_REG_13__SCAN_IN ; P2_U7557
g11438 nand P2_U7869 P2_EBX_REG_12__SCAN_IN ; P2_U7558
g11439 nand P2_U7869 P2_EBX_REG_11__SCAN_IN ; P2_U7559
g11440 nand P2_U7869 P2_EBX_REG_10__SCAN_IN ; P2_U7560
g11441 nand P2_U4596 P2_U3294 ; P2_U7561
g11442 nand P2_U4428 P2_U7285 ; P2_U7562
g11443 nand P2_U7561 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U7563
g11444 nand P2_U4428 P2_U7319 ; P2_U7564
g11445 nand P2_U7561 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7565
g11446 nand P2_U4428 P2_U7353 ; P2_U7566
g11447 nand P2_U7561 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U7567
g11448 nand P2_U4428 P2_U7387 ; P2_U7568
g11449 nand P2_U7561 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U7569
g11450 nand P2_U4428 P2_U7421 ; P2_U7570
g11451 nand P2_U7561 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U7571
g11452 nand P2_U7561 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_U7572
g11453 nand P2_U7561 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U7573
g11454 nand P2_U7561 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U7574
g11455 nand P2_U7561 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_U7575
g11456 nand P2_U7561 P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U7576
g11457 nand P2_U4377 P2_U5572 ; P2_U7577
g11458 nand P2_U4432 P2_STATE2_REG_0__SCAN_IN ; P2_U7578
g11459 nand P2_U2617 P2_U2450 ; P2_U7579
g11460 nand P2_U4376 P2_U5592 ; P2_U7580
g11461 nand P2_U3525 P2_U6845 P2_U7867 ; P2_U7581
g11462 nand P2_U4471 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U7582
g11463 nand P2_U7890 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7583
g11464 nand P2_U7890 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U7584
g11465 nand P2_U3284 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U7585
g11466 nand P2_U4381 P2_U4424 ; P2_U7586
g11467 nand P2_U4471 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_U7587
g11468 nand P2_U7890 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U7588
g11469 nand P2_U2590 P2_U6845 ; P2_U7589
g11470 nand P2_U4471 P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U7590
g11471 nand P2_U2376 P2_U7871 P2_U4416 ; P2_U7591
g11472 nand P2_U7591 P2_U3285 P2_U4422 P2_U3539 ; P2_U7592
g11473 nand P2_U7592 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_U7593
g11474 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_9__SCAN_IN ; P2_U7594
g11475 nand P2_U4423 P2_REIP_REG_9__SCAN_IN ; P2_U7595
g11476 nand P2_U2358 P2_EBX_REG_9__SCAN_IN ; P2_U7596
g11477 nand P2_U7592 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_U7597
g11478 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_8__SCAN_IN ; P2_U7598
g11479 nand P2_U4423 P2_REIP_REG_8__SCAN_IN ; P2_U7599
g11480 nand P2_U2358 P2_EBX_REG_8__SCAN_IN ; P2_U7600
g11481 nand P2_U7592 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_U7601
g11482 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_7__SCAN_IN ; P2_U7602
g11483 nand P2_U4423 P2_REIP_REG_7__SCAN_IN ; P2_U7603
g11484 nand P2_U2358 P2_EBX_REG_7__SCAN_IN ; P2_U7604
g11485 nand P2_U7592 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_U7605
g11486 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_6__SCAN_IN ; P2_U7606
g11487 nand P2_U4423 P2_REIP_REG_6__SCAN_IN ; P2_U7607
g11488 nand P2_U2358 P2_EBX_REG_6__SCAN_IN ; P2_U7608
g11489 nand P2_U7592 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_U7609
g11490 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_5__SCAN_IN ; P2_U7610
g11491 nand P2_U4423 P2_REIP_REG_5__SCAN_IN ; P2_U7611
g11492 nand P2_U2358 P2_EBX_REG_5__SCAN_IN ; P2_U7612
g11493 nand P2_U7592 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_U7613
g11494 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_4__SCAN_IN ; P2_U7614
g11495 nand P2_U4423 P2_REIP_REG_4__SCAN_IN ; P2_U7615
g11496 nand P2_U2358 P2_EBX_REG_4__SCAN_IN ; P2_U7616
g11497 nand P2_U7592 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_U7617
g11498 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_31__SCAN_IN ; P2_U7618
g11499 nand P2_U4423 P2_REIP_REG_31__SCAN_IN ; P2_U7619
g11500 nand P2_U2358 P2_EBX_REG_31__SCAN_IN ; P2_U7620
g11501 nand P2_U7592 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_U7621
g11502 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_30__SCAN_IN ; P2_U7622
g11503 nand P2_U4423 P2_REIP_REG_30__SCAN_IN ; P2_U7623
g11504 nand P2_U2358 P2_EBX_REG_30__SCAN_IN ; P2_U7624
g11505 nand P2_U7592 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_U7625
g11506 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_3__SCAN_IN ; P2_U7626
g11507 nand P2_U4423 P2_REIP_REG_3__SCAN_IN ; P2_U7627
g11508 nand P2_U2358 P2_EBX_REG_3__SCAN_IN ; P2_U7628
g11509 nand P2_U7592 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_U7629
g11510 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_29__SCAN_IN ; P2_U7630
g11511 nand P2_U4423 P2_REIP_REG_29__SCAN_IN ; P2_U7631
g11512 nand P2_U2358 P2_EBX_REG_29__SCAN_IN ; P2_U7632
g11513 nand P2_U7592 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_U7633
g11514 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_28__SCAN_IN ; P2_U7634
g11515 nand P2_U4423 P2_REIP_REG_28__SCAN_IN ; P2_U7635
g11516 nand P2_U2358 P2_EBX_REG_28__SCAN_IN ; P2_U7636
g11517 nand P2_U7592 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_U7637
g11518 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_27__SCAN_IN ; P2_U7638
g11519 nand P2_U4423 P2_REIP_REG_27__SCAN_IN ; P2_U7639
g11520 nand P2_U2358 P2_EBX_REG_27__SCAN_IN ; P2_U7640
g11521 nand P2_U7592 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_U7641
g11522 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_26__SCAN_IN ; P2_U7642
g11523 nand P2_U4423 P2_REIP_REG_26__SCAN_IN ; P2_U7643
g11524 nand P2_U2358 P2_EBX_REG_26__SCAN_IN ; P2_U7644
g11525 nand P2_U7592 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_U7645
g11526 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_25__SCAN_IN ; P2_U7646
g11527 nand P2_U4423 P2_REIP_REG_25__SCAN_IN ; P2_U7647
g11528 nand P2_U2358 P2_EBX_REG_25__SCAN_IN ; P2_U7648
g11529 nand P2_U7592 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_U7649
g11530 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_24__SCAN_IN ; P2_U7650
g11531 nand P2_U4423 P2_REIP_REG_24__SCAN_IN ; P2_U7651
g11532 nand P2_U2358 P2_EBX_REG_24__SCAN_IN ; P2_U7652
g11533 nand P2_U7592 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_U7653
g11534 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_23__SCAN_IN ; P2_U7654
g11535 nand P2_U4423 P2_REIP_REG_23__SCAN_IN ; P2_U7655
g11536 nand P2_U2358 P2_EBX_REG_23__SCAN_IN ; P2_U7656
g11537 nand P2_U7592 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_U7657
g11538 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_22__SCAN_IN ; P2_U7658
g11539 nand P2_U4423 P2_REIP_REG_22__SCAN_IN ; P2_U7659
g11540 nand P2_U2358 P2_EBX_REG_22__SCAN_IN ; P2_U7660
g11541 nand P2_U7592 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_U7661
g11542 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_21__SCAN_IN ; P2_U7662
g11543 nand P2_U4423 P2_REIP_REG_21__SCAN_IN ; P2_U7663
g11544 nand P2_U2358 P2_EBX_REG_21__SCAN_IN ; P2_U7664
g11545 nand P2_U7592 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_U7665
g11546 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_20__SCAN_IN ; P2_U7666
g11547 nand P2_U4423 P2_REIP_REG_20__SCAN_IN ; P2_U7667
g11548 nand P2_U2358 P2_EBX_REG_20__SCAN_IN ; P2_U7668
g11549 nand P2_U7592 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_U7669
g11550 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_2__SCAN_IN ; P2_U7670
g11551 nand P2_U4423 P2_REIP_REG_2__SCAN_IN ; P2_U7671
g11552 nand P2_U2358 P2_EBX_REG_2__SCAN_IN ; P2_U7672
g11553 nand P2_U7592 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_U7673
g11554 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_19__SCAN_IN ; P2_U7674
g11555 nand P2_U4423 P2_REIP_REG_19__SCAN_IN ; P2_U7675
g11556 nand P2_U2358 P2_EBX_REG_19__SCAN_IN ; P2_U7676
g11557 nand P2_U7592 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_U7677
g11558 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_18__SCAN_IN ; P2_U7678
g11559 nand P2_U4423 P2_REIP_REG_18__SCAN_IN ; P2_U7679
g11560 nand P2_U2358 P2_EBX_REG_18__SCAN_IN ; P2_U7680
g11561 nand P2_U7592 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_U7681
g11562 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_17__SCAN_IN ; P2_U7682
g11563 nand P2_U4423 P2_REIP_REG_17__SCAN_IN ; P2_U7683
g11564 nand P2_U2358 P2_EBX_REG_17__SCAN_IN ; P2_U7684
g11565 nand P2_U7592 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_U7685
g11566 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_16__SCAN_IN ; P2_U7686
g11567 nand P2_U4423 P2_REIP_REG_16__SCAN_IN ; P2_U7687
g11568 nand P2_U2358 P2_EBX_REG_16__SCAN_IN ; P2_U7688
g11569 nand P2_U7592 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_U7689
g11570 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_15__SCAN_IN ; P2_U7690
g11571 nand P2_U4423 P2_REIP_REG_15__SCAN_IN ; P2_U7691
g11572 nand P2_U2358 P2_EBX_REG_15__SCAN_IN ; P2_U7692
g11573 nand P2_U7592 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_U7693
g11574 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_14__SCAN_IN ; P2_U7694
g11575 nand P2_U4423 P2_REIP_REG_14__SCAN_IN ; P2_U7695
g11576 nand P2_U2358 P2_EBX_REG_14__SCAN_IN ; P2_U7696
g11577 nand P2_U7592 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_U7697
g11578 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_13__SCAN_IN ; P2_U7698
g11579 nand P2_U4423 P2_REIP_REG_13__SCAN_IN ; P2_U7699
g11580 nand P2_U2358 P2_EBX_REG_13__SCAN_IN ; P2_U7700
g11581 nand P2_U7592 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_U7701
g11582 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_12__SCAN_IN ; P2_U7702
g11583 nand P2_U4423 P2_REIP_REG_12__SCAN_IN ; P2_U7703
g11584 nand P2_U2358 P2_EBX_REG_12__SCAN_IN ; P2_U7704
g11585 nand P2_U7592 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_U7705
g11586 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_11__SCAN_IN ; P2_U7706
g11587 nand P2_U4423 P2_REIP_REG_11__SCAN_IN ; P2_U7707
g11588 nand P2_U2358 P2_EBX_REG_11__SCAN_IN ; P2_U7708
g11589 nand P2_U7592 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_U7709
g11590 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_10__SCAN_IN ; P2_U7710
g11591 nand P2_U4423 P2_REIP_REG_10__SCAN_IN ; P2_U7711
g11592 nand P2_U2358 P2_EBX_REG_10__SCAN_IN ; P2_U7712
g11593 nand P2_U7592 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_U7713
g11594 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_1__SCAN_IN ; P2_U7714
g11595 nand P2_U4423 P2_REIP_REG_1__SCAN_IN ; P2_U7715
g11596 nand P2_U2358 P2_EBX_REG_1__SCAN_IN ; P2_U7716
g11597 nand P2_U4387 P2_U7885 ; P2_U7717
g11598 nand P2_U7739 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_U7718
g11599 nand P2_STATE2_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_0__SCAN_IN ; P2_U7719
g11600 nand P2_U4423 P2_REIP_REG_0__SCAN_IN ; P2_U7720
g11601 nand P2_U2358 P2_EBX_REG_0__SCAN_IN ; P2_U7721
g11602 nand P2_U7720 P2_U3575 ; P2_U7722
g11603 nand P2_U3550 P2_U3536 ; P2_U7723
g11604 nand P2_R2219_U28 P2_U7723 ; P2_U7724
g11605 nand P2_R2219_U30 P2_U7723 ; P2_U7725
g11606 nand P2_R2238_U19 P2_U2356 ; P2_U7726
g11607 nand P2_U3284 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U7727
g11608 nand P2_R2238_U20 P2_U2356 ; P2_U7728
g11609 nand P2_U3284 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7729
g11610 nand P2_R2238_U21 P2_U2356 ; P2_U7730
g11611 nand P2_U3284 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U7731
g11612 nand P2_R2238_U22 P2_U2356 ; P2_U7732
g11613 nand P2_U3284 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U7733
g11614 nand P2_R2238_U7 P2_U2356 ; P2_U7734
g11615 nand P2_U3284 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U7735
g11616 nand P2_U3295 P2_U7873 P2_U3525 ; P2_U7736
g11617 nand P2_U7590 P2_U7589 P2_U4422 P2_U3272 ; P2_U7737
g11618 nand P2_U7861 P2_U2617 ; P2_U7738
g11619 nand P2_U7591 P2_U3285 P2_U4422 P2_U3539 ; P2_U7739
g11620 nand P2_U3521 P2_U7744 P2_U5573 P2_U5571 ; P2_U7740
g11621 nand P2_U2391 P2_U3544 ; P2_U7741
g11622 nand P2_U2377 P2_U6572 ; P2_U7742
g11623 nand P2_U7741 P2_U4448 P2_U7742 ; P2_U7743
g11624 nand P2_U7745 P2_U3278 ; P2_U7744
g11625 nand P2_U7861 P2_U2617 ; P2_U7745
g11626 nand P2_U8003 P2_U8002 P2_U4592 ; P2_U7746
g11627 nand P2_U7971 P2_U7970 P2_U4592 ; P2_U7747
g11628 nand P2_U7955 P2_U7954 P2_U4592 ; P2_U7748
g11629 nand P2_U8035 P2_U8034 P2_U4592 ; P2_U7749
g11630 nand P2_U8019 P2_U8018 P2_U4592 ; P2_U7750
g11631 nand P2_U7987 P2_U7986 P2_U4592 ; P2_U7751
g11632 nand P2_U7939 P2_U7938 P2_U4592 ; P2_U7752
g11633 nand P2_U7923 P2_U7922 P2_U4592 ; P2_U7753
g11634 nand P2_U8154 P2_U8153 P2_U4592 ; P2_U7754
g11635 nand P2_U8170 P2_U8169 P2_U4592 ; P2_U7755
g11636 nand P2_U8186 P2_U8185 P2_U4592 ; P2_U7756
g11637 nand P2_U8202 P2_U8201 P2_U4592 ; P2_U7757
g11638 nand P2_U8218 P2_U8217 P2_U4592 ; P2_U7758
g11639 nand P2_U8234 P2_U8233 P2_U4592 ; P2_U7759
g11640 nand P2_U8250 P2_U8249 P2_U4592 ; P2_U7760
g11641 nand P2_U8266 P2_U8265 P2_U4592 ; P2_U7761
g11642 nand P2_U8005 P2_U8004 P2_U4593 ; P2_U7762
g11643 nand P2_U7973 P2_U7972 P2_U4593 ; P2_U7763
g11644 nand P2_U7957 P2_U7956 P2_U4593 ; P2_U7764
g11645 nand P2_U8037 P2_U8036 P2_U4593 ; P2_U7765
g11646 nand P2_U8021 P2_U8020 P2_U4593 ; P2_U7766
g11647 nand P2_U7989 P2_U7988 P2_U4593 ; P2_U7767
g11648 nand P2_U7941 P2_U7940 P2_U4593 ; P2_U7768
g11649 nand P2_U7925 P2_U7924 P2_U4593 ; P2_U7769
g11650 nand P2_U8156 P2_U8155 P2_U4593 ; P2_U7770
g11651 nand P2_U8172 P2_U8171 P2_U4593 ; P2_U7771
g11652 nand P2_U8188 P2_U8187 P2_U4593 ; P2_U7772
g11653 nand P2_U8204 P2_U8203 P2_U4593 ; P2_U7773
g11654 nand P2_U8220 P2_U8219 P2_U4593 ; P2_U7774
g11655 nand P2_U8236 P2_U8235 P2_U4593 ; P2_U7775
g11656 nand P2_U8252 P2_U8251 P2_U4593 ; P2_U7776
g11657 nand P2_U8268 P2_U8267 P2_U4593 ; P2_U7777
g11658 nand P2_U8007 P2_U8006 P2_U2456 ; P2_U7778
g11659 nand P2_U7975 P2_U7974 P2_U2456 ; P2_U7779
g11660 nand P2_U7959 P2_U7958 P2_U2456 ; P2_U7780
g11661 nand P2_U8039 P2_U8038 P2_U2456 ; P2_U7781
g11662 nand P2_U8023 P2_U8022 P2_U2456 ; P2_U7782
g11663 nand P2_U7991 P2_U7990 P2_U2456 ; P2_U7783
g11664 nand P2_U7943 P2_U7942 P2_U2456 ; P2_U7784
g11665 nand P2_U7927 P2_U7926 P2_U2456 ; P2_U7785
g11666 nand P2_U8158 P2_U8157 P2_U2456 ; P2_U7786
g11667 nand P2_U8174 P2_U8173 P2_U2456 ; P2_U7787
g11668 nand P2_U8190 P2_U8189 P2_U2456 ; P2_U7788
g11669 nand P2_U8206 P2_U8205 P2_U2456 ; P2_U7789
g11670 nand P2_U8222 P2_U8221 P2_U2456 ; P2_U7790
g11671 nand P2_U8238 P2_U8237 P2_U2456 ; P2_U7791
g11672 nand P2_U8254 P2_U8253 P2_U2456 ; P2_U7792
g11673 nand P2_U8270 P2_U8269 P2_U2456 ; P2_U7793
g11674 nand P2_U8009 P2_U8008 P2_U2454 ; P2_U7794
g11675 nand P2_U7977 P2_U7976 P2_U2454 ; P2_U7795
g11676 nand P2_U7961 P2_U7960 P2_U2454 ; P2_U7796
g11677 nand P2_U8041 P2_U8040 P2_U2454 ; P2_U7797
g11678 nand P2_U8025 P2_U8024 P2_U2454 ; P2_U7798
g11679 nand P2_U7993 P2_U7992 P2_U2454 ; P2_U7799
g11680 nand P2_U7945 P2_U7944 P2_U2454 ; P2_U7800
g11681 nand P2_U7929 P2_U7928 P2_U2454 ; P2_U7801
g11682 nand P2_U8160 P2_U8159 P2_U2454 ; P2_U7802
g11683 nand P2_U8176 P2_U8175 P2_U2454 ; P2_U7803
g11684 nand P2_U8192 P2_U8191 P2_U2454 ; P2_U7804
g11685 nand P2_U8208 P2_U8207 P2_U2454 ; P2_U7805
g11686 nand P2_U8224 P2_U8223 P2_U2454 ; P2_U7806
g11687 nand P2_U8240 P2_U8239 P2_U2454 ; P2_U7807
g11688 nand P2_U8256 P2_U8255 P2_U2454 ; P2_U7808
g11689 nand P2_U8272 P2_U8271 P2_U2454 ; P2_U7809
g11690 nand P2_U8011 P2_U8010 P2_U4590 ; P2_U7810
g11691 nand P2_U7979 P2_U7978 P2_U4590 ; P2_U7811
g11692 nand P2_U7963 P2_U7962 P2_U4590 ; P2_U7812
g11693 nand P2_U8043 P2_U8042 P2_U4590 ; P2_U7813
g11694 nand P2_U8027 P2_U8026 P2_U4590 ; P2_U7814
g11695 nand P2_U7995 P2_U7994 P2_U4590 ; P2_U7815
g11696 nand P2_U7947 P2_U7946 P2_U4590 ; P2_U7816
g11697 nand P2_U7931 P2_U7930 P2_U4590 ; P2_U7817
g11698 nand P2_U8162 P2_U8161 P2_U4590 ; P2_U7818
g11699 nand P2_U8178 P2_U8177 P2_U4590 ; P2_U7819
g11700 nand P2_U8194 P2_U8193 P2_U4590 ; P2_U7820
g11701 nand P2_U8210 P2_U8209 P2_U4590 ; P2_U7821
g11702 nand P2_U8226 P2_U8225 P2_U4590 ; P2_U7822
g11703 nand P2_U8242 P2_U8241 P2_U4590 ; P2_U7823
g11704 nand P2_U8258 P2_U8257 P2_U4590 ; P2_U7824
g11705 nand P2_U8274 P2_U8273 P2_U4590 ; P2_U7825
g11706 nand P2_U8013 P2_U8012 P2_U2453 ; P2_U7826
g11707 nand P2_U7981 P2_U7980 P2_U2453 ; P2_U7827
g11708 nand P2_U7965 P2_U7964 P2_U2453 ; P2_U7828
g11709 nand P2_U8045 P2_U8044 P2_U2453 ; P2_U7829
g11710 nand P2_U8029 P2_U8028 P2_U2453 ; P2_U7830
g11711 nand P2_U7997 P2_U7996 P2_U2453 ; P2_U7831
g11712 nand P2_U7949 P2_U7948 P2_U2453 ; P2_U7832
g11713 nand P2_U7933 P2_U7932 P2_U2453 ; P2_U7833
g11714 nand P2_U8164 P2_U8163 P2_U2453 ; P2_U7834
g11715 nand P2_U8180 P2_U8179 P2_U2453 ; P2_U7835
g11716 nand P2_U8196 P2_U8195 P2_U2453 ; P2_U7836
g11717 nand P2_U8212 P2_U8211 P2_U2453 ; P2_U7837
g11718 nand P2_U8228 P2_U8227 P2_U2453 ; P2_U7838
g11719 nand P2_U8244 P2_U8243 P2_U2453 ; P2_U7839
g11720 nand P2_U8260 P2_U8259 P2_U2453 ; P2_U7840
g11721 nand P2_U8276 P2_U8275 P2_U2453 ; P2_U7841
g11722 nand P2_U8015 P2_U8014 P2_U2452 ; P2_U7842
g11723 nand P2_U7983 P2_U7982 P2_U2452 ; P2_U7843
g11724 nand P2_U7967 P2_U7966 P2_U2452 ; P2_U7844
g11725 nand P2_U8047 P2_U8046 P2_U2452 ; P2_U7845
g11726 nand P2_U8031 P2_U8030 P2_U2452 ; P2_U7846
g11727 nand P2_U7999 P2_U7998 P2_U2452 ; P2_U7847
g11728 nand P2_U7951 P2_U7950 P2_U2452 ; P2_U7848
g11729 nand P2_U7935 P2_U7934 P2_U2452 ; P2_U7849
g11730 nand P2_U8166 P2_U8165 P2_U2452 ; P2_U7850
g11731 nand P2_U8182 P2_U8181 P2_U2452 ; P2_U7851
g11732 nand P2_U8198 P2_U8197 P2_U2452 ; P2_U7852
g11733 nand P2_U8214 P2_U8213 P2_U2452 ; P2_U7853
g11734 nand P2_U8230 P2_U8229 P2_U2452 ; P2_U7854
g11735 nand P2_U8246 P2_U8245 P2_U2452 ; P2_U7855
g11736 nand P2_U8262 P2_U8261 P2_U2452 ; P2_U7856
g11737 nand P2_U8278 P2_U8277 P2_U2452 ; P2_U7857
g11738 nand P2_U8017 P2_U8016 P2_U2455 ; P2_U7858
g11739 not P2_U3280 ; P2_U7859
g11740 nand P2_U7985 P2_U7984 P2_U2455 ; P2_U7860
g11741 not P2_U3279 ; P2_U7861
g11742 nand P2_U7969 P2_U7968 P2_U2455 ; P2_U7862
g11743 not P2_U3278 ; P2_U7863
g11744 nand P2_U8049 P2_U8048 P2_U2455 ; P2_U7864
g11745 not P2_U3521 ; P2_U7865
g11746 nand P2_U8033 P2_U8032 P2_U2455 ; P2_U7866
g11747 not P2_U3255 ; P2_U7867
g11748 nand P2_U8001 P2_U8000 P2_U2455 ; P2_U7868
g11749 not P2_U2617 ; P2_U7869
g11750 nand P2_U7953 P2_U7952 P2_U2455 ; P2_U7870
g11751 not P2_U3253 ; P2_U7871
g11752 nand P2_U7937 P2_U7936 P2_U2455 ; P2_U7872
g11753 not P2_U2616 ; P2_U7873
g11754 nand P2_U8168 P2_U8167 P2_U2455 ; P2_U7874
g11755 nand P2_U8184 P2_U8183 P2_U2455 ; P2_U7875
g11756 nand P2_U8200 P2_U8199 P2_U2455 ; P2_U7876
g11757 nand P2_U8216 P2_U8215 P2_U2455 ; P2_U7877
g11758 nand P2_U8232 P2_U8231 P2_U2455 ; P2_U7878
g11759 nand P2_U8248 P2_U8247 P2_U2455 ; P2_U7879
g11760 nand P2_U8264 P2_U8263 P2_U2455 ; P2_U7880
g11761 nand P2_U8280 P2_U8279 P2_U2455 ; P2_U7881
g11762 nand P2_U5590 P2_U4428 ; P2_U7882
g11763 nand P2_U5596 P2_U3525 ; P2_U7883
g11764 nand P2_U4596 P2_U7883 ; P2_U7884
g11765 nand P2_U8348 P2_U8347 P2_U3253 ; P2_U7885
g11766 nand P2_U7722 P2_U5589 ; P2_U7886
g11767 nand P2_U4459 P2_U5589 ; P2_U7887
g11768 nand P2_U4386 P2_U7887 P2_U2589 P2_U4385 P2_U4384 ; P2_U7888
g11769 nand P2_U4459 P2_U5589 ; P2_U7889
g11770 nand P2_U7889 P2_U4458 P2_U2589 P2_U4379 ; P2_U7890
g11771 nand P2_U4572 P2_U4569 P2_STATE_REG_1__SCAN_IN ; P2_U7891
g11772 nand P2_U3244 P2_STATE_REG_0__SCAN_IN P2_REQUESTPENDING_REG_SCAN_IN ; P2_U7892
g11773 nand P2_U4569 P2_STATE_REG_1__SCAN_IN ; P2_U7893
g11774 nand P2_U4600 P2_U4615 ; P2_U7894
g11775 nand P2_U7863 P2_U7871 ; P2_U7895
g11776 nand P2_U3255 P2_U5595 ; P2_U7896
g11777 nand P2_U4429 P2_U5589 ; P2_U7897
g11778 nand P2_DATAWIDTH_REG_0__SCAN_IN P2_REIP_REG_0__SCAN_IN ; P2_U7898
g11779 nand P2_U3259 P2_BE_N_REG_3__SCAN_IN ; P2_U7899
g11780 nand P2_U4439 P2_BYTEENABLE_REG_3__SCAN_IN ; P2_U7900
g11781 nand P2_U3259 P2_BE_N_REG_2__SCAN_IN ; P2_U7901
g11782 nand P2_U4439 P2_BYTEENABLE_REG_2__SCAN_IN ; P2_U7902
g11783 nand P2_U3259 P2_BE_N_REG_1__SCAN_IN ; P2_U7903
g11784 nand P2_U4439 P2_BYTEENABLE_REG_1__SCAN_IN ; P2_U7904
g11785 nand P2_U3259 P2_BE_N_REG_0__SCAN_IN ; P2_U7905
g11786 nand P2_U4439 P2_BYTEENABLE_REG_0__SCAN_IN ; P2_U7906
g11787 nand P2_U3268 P2_U3267 P2_STATE_REG_0__SCAN_IN ; P2_U7907
g11788 or NA P2_STATE_REG_0__SCAN_IN ; P2_U7908
g11789 nand P2_U3266 P2_STATE_REG_2__SCAN_IN ; P2_U7909
g11790 nand P2_U4568 P2_STATE_REG_0__SCAN_IN ; P2_U7910
g11791 nand P2_U4581 P2_U4572 P2_STATE_REG_1__SCAN_IN ; P2_U7911
g11792 nand P2_U4582 P2_U3258 ; P2_U7912
g11793 nand P2_U3267 P2_STATE_REG_2__SCAN_IN P2_STATE_REG_0__SCAN_IN ; P2_U7913
g11794 nand P2_U4584 P2_U3244 ; P2_U7914
g11795 or P2_STATE_REG_1__SCAN_IN P2_STATE_REG_0__SCAN_IN ; P2_U7915
g11796 nand P2_U4473 P2_STATE_REG_0__SCAN_IN ; P2_U7916
g11797 not P2_U3589 ; P2_U7917
g11798 nand P2_U7917 P2_DATAWIDTH_REG_0__SCAN_IN ; P2_U7918
g11799 nand P2_U3590 P2_U3589 ; P2_U7919
g11800 nand P2_U3589 P2_U4589 ; P2_U7920
g11801 nand P2_U7917 P2_DATAWIDTH_REG_1__SCAN_IN ; P2_U7921
g11802 nand P2_U3388 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7922
g11803 or P2_INSTQUEUE_REG_3__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7923
g11804 or P2_INSTQUEUE_REG_0__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7924
g11805 nand P2_U3422 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7925
g11806 or P2_INSTQUEUE_REG_1__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7926
g11807 nand P2_U3411 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7927
g11808 nand P2_U3374 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7928
g11809 or P2_INSTQUEUE_REG_4__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7929
g11810 nand P2_U3333 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7930
g11811 or P2_INSTQUEUE_REG_7__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7931
g11812 nand P2_U3363 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7932
g11813 or P2_INSTQUEUE_REG_5__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7933
g11814 nand P2_U3347 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7934
g11815 or P2_INSTQUEUE_REG_6__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7935
g11816 nand P2_U3399 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7936
g11817 or P2_INSTQUEUE_REG_2__1__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7937
g11818 nand P2_U3389 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7938
g11819 or P2_INSTQUEUE_REG_3__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7939
g11820 or P2_INSTQUEUE_REG_0__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7940
g11821 nand P2_U3423 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7941
g11822 or P2_INSTQUEUE_REG_1__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7942
g11823 nand P2_U3412 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7943
g11824 nand P2_U3375 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7944
g11825 or P2_INSTQUEUE_REG_4__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7945
g11826 nand P2_U3334 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7946
g11827 or P2_INSTQUEUE_REG_7__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7947
g11828 nand P2_U3364 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7948
g11829 or P2_INSTQUEUE_REG_5__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7949
g11830 nand P2_U3348 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7950
g11831 or P2_INSTQUEUE_REG_6__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7951
g11832 nand P2_U3400 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7952
g11833 or P2_INSTQUEUE_REG_2__0__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7953
g11834 nand P2_U3385 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7954
g11835 or P2_INSTQUEUE_REG_3__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7955
g11836 or P2_INSTQUEUE_REG_0__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7956
g11837 nand P2_U3419 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7957
g11838 or P2_INSTQUEUE_REG_1__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7958
g11839 nand P2_U3408 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7959
g11840 nand P2_U3371 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7960
g11841 or P2_INSTQUEUE_REG_4__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7961
g11842 nand P2_U3330 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7962
g11843 or P2_INSTQUEUE_REG_7__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7963
g11844 nand P2_U3360 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7964
g11845 or P2_INSTQUEUE_REG_5__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7965
g11846 nand P2_U3344 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7966
g11847 or P2_INSTQUEUE_REG_6__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7967
g11848 nand P2_U3396 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7968
g11849 or P2_INSTQUEUE_REG_2__4__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7969
g11850 nand P2_U3383 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7970
g11851 or P2_INSTQUEUE_REG_3__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7971
g11852 or P2_INSTQUEUE_REG_0__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7972
g11853 nand P2_U3417 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7973
g11854 or P2_INSTQUEUE_REG_1__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7974
g11855 nand P2_U3406 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7975
g11856 nand P2_U3369 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7976
g11857 or P2_INSTQUEUE_REG_4__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7977
g11858 nand P2_U3328 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7978
g11859 or P2_INSTQUEUE_REG_7__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7979
g11860 nand P2_U3358 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7980
g11861 or P2_INSTQUEUE_REG_5__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7981
g11862 nand P2_U3342 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7982
g11863 or P2_INSTQUEUE_REG_6__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7983
g11864 nand P2_U3394 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7984
g11865 or P2_INSTQUEUE_REG_2__6__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7985
g11866 nand P2_U3384 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7986
g11867 or P2_INSTQUEUE_REG_3__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7987
g11868 or P2_INSTQUEUE_REG_0__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7988
g11869 nand P2_U3418 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7989
g11870 or P2_INSTQUEUE_REG_1__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7990
g11871 nand P2_U3407 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7991
g11872 nand P2_U3370 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7992
g11873 or P2_INSTQUEUE_REG_4__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7993
g11874 nand P2_U3329 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7994
g11875 or P2_INSTQUEUE_REG_7__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7995
g11876 nand P2_U3359 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7996
g11877 or P2_INSTQUEUE_REG_5__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7997
g11878 nand P2_U3343 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7998
g11879 or P2_INSTQUEUE_REG_6__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U7999
g11880 nand P2_U3395 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8000
g11881 or P2_INSTQUEUE_REG_2__5__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8001
g11882 nand P2_U3387 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8002
g11883 or P2_INSTQUEUE_REG_3__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8003
g11884 or P2_INSTQUEUE_REG_0__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8004
g11885 nand P2_U3421 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8005
g11886 or P2_INSTQUEUE_REG_1__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8006
g11887 nand P2_U3410 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8007
g11888 nand P2_U3373 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8008
g11889 or P2_INSTQUEUE_REG_4__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8009
g11890 nand P2_U3332 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8010
g11891 or P2_INSTQUEUE_REG_7__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8011
g11892 nand P2_U3362 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8012
g11893 or P2_INSTQUEUE_REG_5__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8013
g11894 nand P2_U3346 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8014
g11895 or P2_INSTQUEUE_REG_6__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8015
g11896 nand P2_U3398 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8016
g11897 or P2_INSTQUEUE_REG_2__2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8017
g11898 nand P2_U3386 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8018
g11899 or P2_INSTQUEUE_REG_3__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8019
g11900 or P2_INSTQUEUE_REG_0__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8020
g11901 nand P2_U3420 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8021
g11902 or P2_INSTQUEUE_REG_1__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8022
g11903 nand P2_U3409 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8023
g11904 nand P2_U3372 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8024
g11905 or P2_INSTQUEUE_REG_4__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8025
g11906 nand P2_U3331 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8026
g11907 or P2_INSTQUEUE_REG_7__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8027
g11908 nand P2_U3361 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8028
g11909 or P2_INSTQUEUE_REG_5__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8029
g11910 nand P2_U3345 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8030
g11911 or P2_INSTQUEUE_REG_6__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8031
g11912 nand P2_U3397 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8032
g11913 or P2_INSTQUEUE_REG_2__3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8033
g11914 nand P2_U3382 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8034
g11915 or P2_INSTQUEUE_REG_3__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8035
g11916 or P2_INSTQUEUE_REG_0__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8036
g11917 nand P2_U3416 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8037
g11918 or P2_INSTQUEUE_REG_1__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8038
g11919 nand P2_U3405 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8039
g11920 nand P2_U3368 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8040
g11921 or P2_INSTQUEUE_REG_4__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8041
g11922 nand P2_U3327 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8042
g11923 or P2_INSTQUEUE_REG_7__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8043
g11924 nand P2_U3357 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8044
g11925 or P2_INSTQUEUE_REG_5__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8045
g11926 nand P2_U3341 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8046
g11927 or P2_INSTQUEUE_REG_6__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8047
g11928 nand P2_U3393 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8048
g11929 or P2_INSTQUEUE_REG_2__7__SCAN_IN P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8049
g11930 nand P2_R2167_U6 P2_U4435 ; P2_U8050
g11931 nand P2_U4604 P2_U3297 ; P2_U8051
g11932 nand P2_U7871 P2_U3293 ; P2_U8052
g11933 nand P2_U3253 P2_U3282 ; P2_U8053
g11934 nand P2_U4427 P2_U3297 ; P2_U8054
g11935 nand P2_U3289 P2_U3520 ; P2_U8055
g11936 or U211 P2_STATE2_REG_0__SCAN_IN ; P2_U8056
g11937 nand P2_U4617 P2_STATE2_REG_0__SCAN_IN ; P2_U8057
g11938 nand P2_U3299 P2_STATE2_REG_3__SCAN_IN ; P2_U8058
g11939 nand P2_U2448 P2_U4620 ; P2_U8059
g11940 nand P2_U4631 P2_STATE2_REG_0__SCAN_IN ; P2_U8060
g11941 nand P2_U4630 P2_U4619 P2_U3284 ; P2_U8061
g11942 nand P2_R2182_U40 P2_U3318 ; P2_U8062
g11943 nand P2_U4637 P2_U3316 ; P2_U8063
g11944 not P2_U3579 ; P2_U8064
g11945 nand P2_U3311 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U8065
g11946 nand P2_U4642 P2_U3310 ; P2_U8066
g11947 not P2_U3580 ; P2_U8067
g11948 nand P2_U7859 P2_U5574 ; P2_U8068
g11949 nand P2_U3280 P2_U5575 ; P2_U8069
g11950 nand P2_U4435 P2_U3297 ; P2_U8070
g11951 nand P2_U4433 P2_U2359 P2_R2167_U6 ; P2_U8071
g11952 nand P2_U3594 P2_U4394 ; P2_U8072
g11953 nand P2_U5584 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U8073
g11954 nand P2_U3280 P2_U5586 ; P2_U8074
g11955 nand P2_U2617 P2_U3279 P2_U7859 ; P2_U8075
g11956 nand P2_U4424 P2_U3253 ; P2_U8076
g11957 nand P2_U4475 P2_U7871 ; P2_U8077
g11958 nand P2_U5585 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8078
g11959 nand P2_U4591 P2_U3276 P2_U3273 ; P2_U8079
g11960 nand P2_U3277 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8080
g11961 nand P2_U4590 P2_U3273 ; P2_U8081
g11962 not P2_U3581 ; P2_U8082
g11963 nand P2_U5584 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8083
g11964 nand P2_U5614 P2_U4394 ; P2_U8084
g11965 nand P2_U3528 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_U8085
g11966 nand P2_U3647 P2_U3683 ; P2_U8086
g11967 not P2_U3597 ; P2_U8087
g11968 nand P2_U3528 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_U8088
g11969 nand P2_R1957_U49 P2_U3647 ; P2_U8089
g11970 not P2_U3598 ; P2_U8090
g11971 nand P2_U5616 P2_U5605 ; P2_U8091
g11972 nand P2_U3530 P2_U5606 ; P2_U8092
g11973 nand P2_U5584 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U8093
g11974 nand P2_U5623 P2_U4394 ; P2_U8094
g11975 nand P2_U3886 P2_U4597 P2_U3255 ; P2_U8095
g11976 nand P2_U7869 P2_U5625 P2_U7867 ; P2_U8096
g11977 nand P2_U8096 P2_U8095 ; P2_U8097
g11978 nand P2_U3271 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U8098
g11979 nand P2_U3272 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U8099
g11980 not P2_U3582 ; P2_U8100
g11981 nand P2_U5584 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U8101
g11982 nand P2_U5633 P2_U4394 ; P2_U8102
g11983 nand P2_U5584 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U8103
g11984 nand P2_U5641 P2_U4394 ; P2_U8104
g11985 nand P2_U5643 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_U8105
g11986 nand P2_U5651 P2_U3533 ; P2_U8106
g11987 nand P2_U8064 P2_U4636 ; P2_U8107
g11988 nand P2_U3579 P2_U3319 ; P2_U8108
g11989 nand P2_U8108 P2_U8107 ; P2_U8109
g11990 nand P2_U5643 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_U8110
g11991 nand P2_U5655 P2_U3533 ; P2_U8111
g11992 nand P2_U5643 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_U8112
g11993 nand P2_U5660 P2_U3533 ; P2_U8113
g11994 nand P2_U5643 P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_U8114
g11995 nand P2_U5664 P2_U3533 ; P2_U8115
g11996 nand P2_U2359 P2_U3280 P2_U2616 ; P2_U8116
g11997 nand P2_U2438 P2_U7873 ; P2_U8117
g11998 nand P2_U8117 P2_U8116 ; P2_U8118
g11999 nand P2_U3253 P2_U3278 P2_U3297 ; P2_U8119
g12000 nand P2_U8118 P2_R2167_U6 ; P2_U8120
g12001 nand P2_U7859 P2_U7873 ; P2_U8121
g12002 nand P2_U2616 P2_U3282 ; P2_U8122
g12003 nand P2_U3547 P2_BYTEENABLE_REG_3__SCAN_IN ; P2_U8123
g12004 nand P2_U3606 P2_U4438 ; P2_U8124
g12005 nand P2_U3547 P2_BYTEENABLE_REG_2__SCAN_IN ; P2_U8125
g12006 nand P2_U3607 P2_U4438 ; P2_U8126
g12007 nand P2_U3547 P2_BYTEENABLE_REG_0__SCAN_IN ; P2_U8127
g12008 nand P2_U4438 P2_REIP_REG_0__SCAN_IN ; P2_U8128
g12009 nand P2_U4439 P2_U3552 ; P2_U8129
g12010 nand P2_U3259 P2_W_R_N_REG_SCAN_IN ; P2_U8130
g12011 nand P2_U3287 P2_U7873 ; P2_U8131
g12012 nand P2_R2243_U8 P2_U2616 ; P2_U8132
g12013 nand P2_U6838 P2_U3257 ; P2_U8133
g12014 nand P2_U4400 P2_MORE_REG_SCAN_IN ; P2_U8134
g12015 nand P2_U7917 P2_STATEBS16_REG_SCAN_IN ; P2_U8135
g12016 nand BS16 P2_U3589 ; P2_U8136
g12017 nand P2_U6843 P2_REQUESTPENDING_REG_SCAN_IN ; P2_U8137
g12018 nand P2_U6852 P2_U4402 ; P2_U8138
g12019 nand P2_U4439 P2_U3551 ; P2_U8139
g12020 nand P2_U3259 P2_D_C_N_REG_SCAN_IN ; P2_U8140
g12021 nand P2_U3259 P2_M_IO_N_REG_SCAN_IN ; P2_U8141
g12022 nand P2_U4439 P2_MEMORYFETCH_REG_SCAN_IN ; P2_U8142
g12023 nand P2_U6857 P2_READREQUEST_REG_SCAN_IN ; P2_U8143
g12024 nand P2_U6858 P2_U4403 ; P2_U8144
g12025 nand P2_U7873 P2_U3520 ; P2_U8145
g12026 nand P2_U2616 P2_U3297 ; P2_U8146
g12027 nand P2_U4405 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8147
g12028 nand P2_U7007 P2_U3273 ; P2_U8148
g12029 not P2_U3583 ; P2_U8149
g12030 nand P2_U3273 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U8150
g12031 nand P2_U3276 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8151
g12032 not P2_U3584 ; P2_U8152
g12033 nand P2_U3584 P2_U3327 ; P2_U8153
g12034 nand P2_U8152 P2_U3431 ; P2_U8154
g12035 nand P2_U3584 P2_U3368 ; P2_U8155
g12036 nand P2_U8152 P2_U3465 ; P2_U8156
g12037 nand P2_U3584 P2_U3357 ; P2_U8157
g12038 nand P2_U8152 P2_U3454 ; P2_U8158
g12039 nand P2_U3584 P2_U3416 ; P2_U8159
g12040 nand P2_U8152 P2_U3511 ; P2_U8160
g12041 nand P2_U3584 P2_U3382 ; P2_U8161
g12042 nand P2_U8152 P2_U3477 ; P2_U8162
g12043 nand P2_U3584 P2_U3405 ; P2_U8163
g12044 nand P2_U8152 P2_U3500 ; P2_U8164
g12045 nand P2_U3584 P2_U3393 ; P2_U8165
g12046 nand P2_U8152 P2_U3488 ; P2_U8166
g12047 nand P2_U3584 P2_U3341 ; P2_U8167
g12048 nand P2_U8152 P2_U3442 ; P2_U8168
g12049 nand P2_U3584 P2_U3328 ; P2_U8169
g12050 nand P2_U8152 P2_U3432 ; P2_U8170
g12051 nand P2_U3584 P2_U3369 ; P2_U8171
g12052 nand P2_U8152 P2_U3466 ; P2_U8172
g12053 nand P2_U3584 P2_U3358 ; P2_U8173
g12054 nand P2_U8152 P2_U3455 ; P2_U8174
g12055 nand P2_U3584 P2_U3417 ; P2_U8175
g12056 nand P2_U8152 P2_U3512 ; P2_U8176
g12057 nand P2_U3584 P2_U3383 ; P2_U8177
g12058 nand P2_U8152 P2_U3478 ; P2_U8178
g12059 nand P2_U3584 P2_U3406 ; P2_U8179
g12060 nand P2_U8152 P2_U3501 ; P2_U8180
g12061 nand P2_U3584 P2_U3394 ; P2_U8181
g12062 nand P2_U8152 P2_U3489 ; P2_U8182
g12063 nand P2_U3584 P2_U3342 ; P2_U8183
g12064 nand P2_U8152 P2_U3443 ; P2_U8184
g12065 nand P2_U3584 P2_U3329 ; P2_U8185
g12066 nand P2_U8152 P2_U3433 ; P2_U8186
g12067 nand P2_U3584 P2_U3370 ; P2_U8187
g12068 nand P2_U8152 P2_U3467 ; P2_U8188
g12069 nand P2_U3584 P2_U3359 ; P2_U8189
g12070 nand P2_U8152 P2_U3456 ; P2_U8190
g12071 nand P2_U3584 P2_U3418 ; P2_U8191
g12072 nand P2_U8152 P2_U3513 ; P2_U8192
g12073 nand P2_U3584 P2_U3384 ; P2_U8193
g12074 nand P2_U8152 P2_U3479 ; P2_U8194
g12075 nand P2_U3584 P2_U3407 ; P2_U8195
g12076 nand P2_U8152 P2_U3502 ; P2_U8196
g12077 nand P2_U3584 P2_U3395 ; P2_U8197
g12078 nand P2_U8152 P2_U3490 ; P2_U8198
g12079 nand P2_U3584 P2_U3343 ; P2_U8199
g12080 nand P2_U8152 P2_U3444 ; P2_U8200
g12081 nand P2_U3584 P2_U3330 ; P2_U8201
g12082 nand P2_U8152 P2_U3434 ; P2_U8202
g12083 nand P2_U3584 P2_U3371 ; P2_U8203
g12084 nand P2_U8152 P2_U3468 ; P2_U8204
g12085 nand P2_U3584 P2_U3360 ; P2_U8205
g12086 nand P2_U8152 P2_U3457 ; P2_U8206
g12087 nand P2_U3584 P2_U3419 ; P2_U8207
g12088 nand P2_U8152 P2_U3514 ; P2_U8208
g12089 nand P2_U3584 P2_U3385 ; P2_U8209
g12090 nand P2_U8152 P2_U3480 ; P2_U8210
g12091 nand P2_U3584 P2_U3408 ; P2_U8211
g12092 nand P2_U8152 P2_U3503 ; P2_U8212
g12093 nand P2_U3584 P2_U3396 ; P2_U8213
g12094 nand P2_U8152 P2_U3491 ; P2_U8214
g12095 nand P2_U3584 P2_U3344 ; P2_U8215
g12096 nand P2_U8152 P2_U3445 ; P2_U8216
g12097 nand P2_U3584 P2_U3331 ; P2_U8217
g12098 nand P2_U8152 P2_U3435 ; P2_U8218
g12099 nand P2_U3584 P2_U3372 ; P2_U8219
g12100 nand P2_U8152 P2_U3469 ; P2_U8220
g12101 nand P2_U3584 P2_U3361 ; P2_U8221
g12102 nand P2_U8152 P2_U3458 ; P2_U8222
g12103 nand P2_U3584 P2_U3420 ; P2_U8223
g12104 nand P2_U8152 P2_U3515 ; P2_U8224
g12105 nand P2_U3584 P2_U3386 ; P2_U8225
g12106 nand P2_U8152 P2_U3481 ; P2_U8226
g12107 nand P2_U3584 P2_U3409 ; P2_U8227
g12108 nand P2_U8152 P2_U3504 ; P2_U8228
g12109 nand P2_U3584 P2_U3397 ; P2_U8229
g12110 nand P2_U8152 P2_U3492 ; P2_U8230
g12111 nand P2_U3584 P2_U3345 ; P2_U8231
g12112 nand P2_U8152 P2_U3446 ; P2_U8232
g12113 nand P2_U3584 P2_U3332 ; P2_U8233
g12114 nand P2_U8152 P2_U3436 ; P2_U8234
g12115 nand P2_U3584 P2_U3373 ; P2_U8235
g12116 nand P2_U8152 P2_U3470 ; P2_U8236
g12117 nand P2_U3584 P2_U3362 ; P2_U8237
g12118 nand P2_U8152 P2_U3459 ; P2_U8238
g12119 nand P2_U3584 P2_U3421 ; P2_U8239
g12120 nand P2_U8152 P2_U3516 ; P2_U8240
g12121 nand P2_U3584 P2_U3387 ; P2_U8241
g12122 nand P2_U8152 P2_U3482 ; P2_U8242
g12123 nand P2_U3584 P2_U3410 ; P2_U8243
g12124 nand P2_U8152 P2_U3505 ; P2_U8244
g12125 nand P2_U3584 P2_U3398 ; P2_U8245
g12126 nand P2_U8152 P2_U3493 ; P2_U8246
g12127 nand P2_U3584 P2_U3346 ; P2_U8247
g12128 nand P2_U8152 P2_U3447 ; P2_U8248
g12129 nand P2_U3584 P2_U3333 ; P2_U8249
g12130 nand P2_U8152 P2_U3437 ; P2_U8250
g12131 nand P2_U3584 P2_U3374 ; P2_U8251
g12132 nand P2_U8152 P2_U3471 ; P2_U8252
g12133 nand P2_U3584 P2_U3363 ; P2_U8253
g12134 nand P2_U8152 P2_U3460 ; P2_U8254
g12135 nand P2_U3584 P2_U3422 ; P2_U8255
g12136 nand P2_U8152 P2_U3517 ; P2_U8256
g12137 nand P2_U3584 P2_U3388 ; P2_U8257
g12138 nand P2_U8152 P2_U3483 ; P2_U8258
g12139 nand P2_U3584 P2_U3411 ; P2_U8259
g12140 nand P2_U8152 P2_U3506 ; P2_U8260
g12141 nand P2_U3584 P2_U3399 ; P2_U8261
g12142 nand P2_U8152 P2_U3494 ; P2_U8262
g12143 nand P2_U3584 P2_U3347 ; P2_U8263
g12144 nand P2_U8152 P2_U3448 ; P2_U8264
g12145 nand P2_U3584 P2_U3334 ; P2_U8265
g12146 nand P2_U8152 P2_U3438 ; P2_U8266
g12147 nand P2_U3584 P2_U3375 ; P2_U8267
g12148 nand P2_U8152 P2_U3472 ; P2_U8268
g12149 nand P2_U3584 P2_U3364 ; P2_U8269
g12150 nand P2_U8152 P2_U3461 ; P2_U8270
g12151 nand P2_U3584 P2_U3423 ; P2_U8271
g12152 nand P2_U8152 P2_U3518 ; P2_U8272
g12153 nand P2_U3584 P2_U3389 ; P2_U8273
g12154 nand P2_U8152 P2_U3484 ; P2_U8274
g12155 nand P2_U3584 P2_U3412 ; P2_U8275
g12156 nand P2_U8152 P2_U3507 ; P2_U8276
g12157 nand P2_U3584 P2_U3400 ; P2_U8277
g12158 nand P2_U8152 P2_U3495 ; P2_U8278
g12159 nand P2_U3584 P2_U3348 ; P2_U8279
g12160 nand P2_U8152 P2_U3449 ; P2_U8280
g12161 nand P2_U3519 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U8281
g12162 nand P2_U3598 P2_U3597 P2_FLUSH_REG_SCAN_IN ; P2_U8282
g12163 nand P2_U3519 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U8283
g12164 nand P2_U3597 P2_U8090 P2_FLUSH_REG_SCAN_IN ; P2_U8284
g12165 nand P2_U3519 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U8285
g12166 nand P2_U8087 P2_FLUSH_REG_SCAN_IN ; P2_U8286
g12167 nand P2_U3616 P2_U4406 ; P2_U8287
g12168 nand P2_U5581 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_U8288
g12169 nand P2_U5581 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_U8289
g12170 nand P2_U5611 P2_U4406 ; P2_U8290
g12171 nand P2_U5581 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_U8291
g12172 nand P2_U5619 P2_U4406 ; P2_U8292
g12173 nand P2_U5581 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_U8293
g12174 nand P2_U5629 P2_U4406 ; P2_U8294
g12175 nand P2_U5581 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_U8295
g12176 nand P2_U5637 P2_U4406 ; P2_U8296
g12177 nand P2_U3242 P2_U7873 ; P2_U8297
g12178 nand P2_U2616 P2_U7183 ; P2_U8298
g12179 nand P2_U7217 P2_U7873 ; P2_U8299
g12180 nand P2_U2616 P2_U7200 ; P2_U8300
g12181 nand P2_U7251 P2_U7873 ; P2_U8301
g12182 nand P2_U2616 P2_U7234 ; P2_U8302
g12183 nand P2_U7285 P2_U7873 ; P2_U8303
g12184 nand P2_U2616 P2_U7268 ; P2_U8304
g12185 nand P2_U7319 P2_U7873 ; P2_U8305
g12186 nand P2_U2616 P2_U7302 ; P2_U8306
g12187 nand P2_U7353 P2_U7873 ; P2_U8307
g12188 nand P2_U2616 P2_U7336 ; P2_U8308
g12189 nand P2_U7387 P2_U7873 ; P2_U8309
g12190 nand P2_U2616 P2_U7370 ; P2_U8310
g12191 nand P2_U7421 P2_U7873 ; P2_U8311
g12192 nand P2_U2616 P2_U7404 ; P2_U8312
g12193 nand P2_R2256_U5 P2_U3572 ; P2_U8313
g12194 nand P2_U3242 P2_R2267_U56 ; P2_U8314
g12195 nand P2_R2256_U17 P2_U3572 ; P2_U8315
g12196 nand P2_U3242 P2_R2267_U19 ; P2_U8316
g12197 nand P2_R2256_U18 P2_U3572 ; P2_U8317
g12198 nand P2_U3242 P2_R2267_U58 ; P2_U8318
g12199 nand P2_R2256_U19 P2_U3572 ; P2_U8319
g12200 nand P2_U3242 P2_R2267_U18 ; P2_U8320
g12201 nand P2_R2256_U20 P2_U3572 ; P2_U8321
g12202 nand P2_U3242 P2_R2267_U60 ; P2_U8322
g12203 nand P2_R2256_U26 P2_U3572 ; P2_U8323
g12204 nand P2_U3242 P2_R2267_U17 ; P2_U8324
g12205 nand P2_R2256_U22 P2_U3572 ; P2_U8325
g12206 nand P2_U3242 P2_R2267_U65 ; P2_U8326
g12207 nand P2_R2256_U4 P2_U3572 ; P2_U8327
g12208 nand P2_U3242 P2_R2267_U43 ; P2_U8328
g12209 nand P2_R2256_U21 P2_U3572 ; P2_U8329
g12210 nand P2_U3242 P2_R2267_U21 ; P2_U8330
g12211 nand P2_R2219_U24 P2_U2617 ; P2_U8331
g12212 nand P2_U7869 P2_EBX_REG_7__SCAN_IN ; P2_U8332
g12213 nand P2_R2219_U25 P2_U2617 ; P2_U8333
g12214 nand P2_U7869 P2_EBX_REG_6__SCAN_IN ; P2_U8334
g12215 nand P2_R2219_U26 P2_U2617 ; P2_U8335
g12216 nand P2_U7869 P2_EBX_REG_5__SCAN_IN ; P2_U8336
g12217 nand P2_R2219_U27 P2_U2617 ; P2_U8337
g12218 nand P2_U7869 P2_EBX_REG_4__SCAN_IN ; P2_U8338
g12219 nand P2_R2219_U28 P2_U2617 ; P2_U8339
g12220 nand P2_U7869 P2_EBX_REG_3__SCAN_IN ; P2_U8340
g12221 nand P2_R2219_U29 P2_U2617 ; P2_U8341
g12222 nand P2_U7869 P2_EBX_REG_2__SCAN_IN ; P2_U8342
g12223 nand P2_R2219_U30 P2_U2617 ; P2_U8343
g12224 nand P2_U7869 P2_EBX_REG_1__SCAN_IN ; P2_U8344
g12225 nand P2_R2219_U8 P2_U2617 ; P2_U8345
g12226 nand P2_U7869 P2_EBX_REG_0__SCAN_IN ; P2_U8346
g12227 nand P2_U3255 P2_U7740 ; P2_U8347
g12228 nand P2_U7867 P2_U3525 ; P2_U8348
g12229 nand P2_R2337_U68 P2_U3284 ; P2_U8349
g12230 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_U8350
g12231 nand P2_R2238_U6 P2_U3283 ; P2_U8351
g12232 nand P2_SUB_450_U6 P2_U4417 ; P2_U8352
g12233 nand P2_R2238_U19 P2_U3283 ; P2_U8353
g12234 nand P2_SUB_450_U17 P2_U4417 ; P2_U8354
g12235 nand P2_R2238_U20 P2_U3283 ; P2_U8355
g12236 nand P2_SUB_450_U18 P2_U4417 ; P2_U8356
g12237 nand P2_R2238_U21 P2_U3283 ; P2_U8357
g12238 nand P2_SUB_450_U19 P2_U4417 ; P2_U8358
g12239 nand P2_R2238_U22 P2_U3283 ; P2_U8359
g12240 nand P2_SUB_450_U20 P2_U4417 ; P2_U8360
g12241 nand P2_R2337_U61 P2_U3284 ; P2_U8361
g12242 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_U8362
g12243 nand P2_R2337_U62 P2_U3284 ; P2_U8363
g12244 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_U8364
g12245 nand P2_R2337_U63 P2_U3284 ; P2_U8365
g12246 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_U8366
g12247 nand P2_R2337_U64 P2_U3284 ; P2_U8367
g12248 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_U8368
g12249 nand P2_R2337_U65 P2_U3284 ; P2_U8369
g12250 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_U8370
g12251 nand P2_R2337_U66 P2_U3284 ; P2_U8371
g12252 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_U8372
g12253 nand P2_R2337_U69 P2_U3284 ; P2_U8373
g12254 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_U8374
g12255 nand P2_R2337_U67 P2_U3284 ; P2_U8375
g12256 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_U8376
g12257 nand P2_R2337_U71 P2_U3284 ; P2_U8377
g12258 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_U8378
g12259 nand P2_R2337_U72 P2_U3284 ; P2_U8379
g12260 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_U8380
g12261 nand P2_R2337_U73 P2_U3284 ; P2_U8381
g12262 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_U8382
g12263 nand P2_R2337_U74 P2_U3284 ; P2_U8383
g12264 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_U8384
g12265 nand P2_R2337_U75 P2_U3284 ; P2_U8385
g12266 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_U8386
g12267 nand P2_R2337_U76 P2_U3284 ; P2_U8387
g12268 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_U8388
g12269 nand P2_R2337_U77 P2_U3284 ; P2_U8389
g12270 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_U8390
g12271 nand P2_R2337_U78 P2_U3284 ; P2_U8391
g12272 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_U8392
g12273 nand P2_R2337_U79 P2_U3284 ; P2_U8393
g12274 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_U8394
g12275 nand P2_R2337_U80 P2_U3284 ; P2_U8395
g12276 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_U8396
g12277 nand P2_R2337_U70 P2_U3284 ; P2_U8397
g12278 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_U8398
g12279 nand P2_R2337_U81 P2_U3284 ; P2_U8399
g12280 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_U8400
g12281 nand P2_R2337_U82 P2_U3284 ; P2_U8401
g12282 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_U8402
g12283 nand P2_R2337_U83 P2_U3284 ; P2_U8403
g12284 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_U8404
g12285 nand P2_R2337_U84 P2_U3284 ; P2_U8405
g12286 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_U8406
g12287 nand P2_R2337_U85 P2_U3284 ; P2_U8407
g12288 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_U8408
g12289 nand P2_R2337_U86 P2_U3284 ; P2_U8409
g12290 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_U8410
g12291 nand P2_R2337_U87 P2_U3284 ; P2_U8411
g12292 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_U8412
g12293 nand P2_R2337_U88 P2_U3284 ; P2_U8413
g12294 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_U8414
g12295 nand P2_R2337_U89 P2_U3284 ; P2_U8415
g12296 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_U8416
g12297 nand P2_R2337_U90 P2_U3284 ; P2_U8417
g12298 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_U8418
g12299 nand P2_R2337_U4 P2_U3284 ; P2_U8419
g12300 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_U8420
g12301 nand P2_U3284 P2_PHYADDRPOINTER_REG_0__SCAN_IN ; P2_U8421
g12302 nand P2_STATE2_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_U8422
g12303 nand P2_R2238_U6 P2_U3269 ; P2_U8423
g12304 nand P2_U2615 P2_STATE2_REG_1__SCAN_IN ; P2_U8424
g12305 nand P2_R2238_U19 P2_U3269 ; P2_U8425
g12306 nand P2_U2615 P2_STATE2_REG_1__SCAN_IN ; P2_U8426
g12307 nand P2_R2238_U20 P2_U3269 ; P2_U8427
g12308 nand P2_SUB_589_U8 P2_STATE2_REG_1__SCAN_IN ; P2_U8428
g12309 nand P2_R2238_U21 P2_U3269 ; P2_U8429
g12310 nand P2_SUB_589_U9 P2_STATE2_REG_1__SCAN_IN ; P2_U8430
g12311 nand P2_R2238_U22 P2_U3269 ; P2_U8431
g12312 nand P2_SUB_589_U6 P2_STATE2_REG_1__SCAN_IN ; P2_U8432
g12313 nand P2_R2238_U7 P2_U3269 ; P2_U8433
g12314 nand P2_SUB_589_U7 P2_STATE2_REG_1__SCAN_IN ; P2_U8434
g12315 nor P1_STATE2_REG_2__SCAN_IN P1_STATEBS16_REG_SCAN_IN ; P1_U2352
g12316 and P1_U4231 P1_STATE2_REG_2__SCAN_IN ; P1_U2353
g12317 and P1_U4265 P1_U4477 ; P1_U2354
g12318 and P1_U3234 P1_U2450 ; P1_U2355
g12319 and P1_R2238_U6 P1_U4192 ; P1_U2356
g12320 and P1_U5959 P1_U3865 P1_R2167_U17 ; P1_U2357
g12321 and P1_U2388 P1_U4224 ; P1_U2358
g12322 and P1_U3431 P1_STATE2_REG_2__SCAN_IN ; P1_U2359
g12323 and P1_U3414 P1_STATE2_REG_2__SCAN_IN ; P1_U2360
g12324 and P1_U4224 P1_STATE2_REG_3__SCAN_IN ; P1_U2361
g12325 and P1_U2359 P1_U4208 ; P1_U2362
g12326 and P1_U2359 P1_U4210 ; P1_U2363
g12327 and P1_U3864 P1_U3416 ; P1_U2364
g12328 and P1_U4261 P1_U3416 ; P1_U2365
g12329 and P1_U3431 P1_U3430 P1_STATE2_REG_1__SCAN_IN ; P1_U2366
g12330 and P1_U3431 P1_R2337_U69 P1_STATE2_REG_1__SCAN_IN ; P1_U2367
g12331 and P1_U4235 P1_STATE2_REG_0__SCAN_IN ; P1_U2368
g12332 and P1_U2362 P1_U4497 ; P1_U2369
g12333 and P1_U3414 P1_U3263 ; P1_U2370
g12334 and P1_U4222 P1_U4449 ; P1_U2371
g12335 and P1_U3416 P1_STATE2_REG_0__SCAN_IN ; P1_U2372
g12336 and P1_U3431 P1_STATE2_REG_3__SCAN_IN ; P1_U2373
g12337 and P1_U2360 P1_U4214 ; P1_U2374
g12338 and P1_U2360 P1_U4216 ; P1_U2375
g12339 and P1_U5798 P1_U3416 ; P1_U2376
g12340 and P1_U3762 P1_U3414 ; P1_U2377
g12341 and P1_U2360 P1_U5569 ; P1_U2378
g12342 and P1_U2363 P1_U3280 ; P1_U2379
g12343 and P1_U2360 P1_U7608 ; P1_U2380
g12344 and P1_U2357 P1_U3271 ; P1_U2381
g12345 and P1_U2357 P1_U4477 ; P1_U2382
g12346 and P1_U4222 P1_U3391 ; P1_U2383
g12347 and P1_U3417 P1_STATE2_REG_0__SCAN_IN ; P1_U2384
g12348 and P1_U3417 P1_U3294 ; P1_U2385
g12349 and P1_U4223 P1_U3423 ; P1_U2386
g12350 and P1_U3884 P1_U4223 ; P1_U2387
g12351 and P1_U4209 P1_STATEBS16_REG_SCAN_IN ; P1_U2388
g12352 and P1_U2452 P1_U7494 ; P1_U2389
g12353 and U346 P1_U4224 ; P1_U2390
g12354 and U335 P1_U4224 ; P1_U2391
g12355 and U324 P1_U4224 ; P1_U2392
g12356 and U321 P1_U4224 ; P1_U2393
g12357 and U320 P1_U4224 ; P1_U2394
g12358 and U319 P1_U4224 ; P1_U2395
g12359 and U318 P1_U4224 ; P1_U2396
g12360 and U317 P1_U4224 ; P1_U2397
g12361 and U330 P1_U2358 ; P1_U2398
g12362 and U339 P1_U2358 ; P1_U2399
g12363 and U329 P1_U2358 ; P1_U2400
g12364 and U338 P1_U2358 ; P1_U2401
g12365 and U328 P1_U2358 ; P1_U2402
g12366 and U337 P1_U2358 ; P1_U2403
g12367 and U327 P1_U2358 ; P1_U2404
g12368 and U336 P1_U2358 ; P1_U2405
g12369 and U326 P1_U2358 ; P1_U2406
g12370 and U334 P1_U2358 ; P1_U2407
g12371 and U325 P1_U2358 ; P1_U2408
g12372 and U333 P1_U2358 ; P1_U2409
g12373 and U323 P1_U2358 ; P1_U2410
g12374 and U332 P1_U2358 ; P1_U2411
g12375 and U322 P1_U2358 ; P1_U2412
g12376 and U331 P1_U2358 ; P1_U2413
g12377 and P1_U2361 P1_U3271 ; P1_U2414
g12378 and P1_U2361 P1_U3391 ; P1_U2415
g12379 and P1_U2361 P1_U3277 ; P1_U2416
g12380 and P1_U2361 P1_U3284 ; P1_U2417
g12381 and P1_U2361 P1_U3283 ; P1_U2418
g12382 and P1_U2361 P1_U3278 ; P1_U2419
g12383 and P1_U2361 P1_U4173 ; P1_U2420
g12384 and P1_U2361 P1_U4171 ; P1_U2421
g12385 and P1_U4223 P1_U5461 ; P1_U2422
g12386 and P1_U4223 P1_U4231 ; P1_U2423
g12387 and P1_U2384 P1_U3284 ; P1_U2424
g12388 and P1_U2368 P1_U2448 ; P1_U2425
g12389 and P1_U3889 P1_U3431 ; P1_U2426
g12390 nor P1_STATE2_REG_3__SCAN_IN P1_STATE2_REG_1__SCAN_IN ; P1_U2427
g12391 and P1_STATE2_REG_2__SCAN_IN P1_STATE2_REG_1__SCAN_IN ; P1_U2428
g12392 and P1_U6366 P1_U3431 ; P1_U2429
g12393 and P1_U3387 P1_STATE2_REG_1__SCAN_IN ; P1_U2430
g12394 and P1_U4199 P1_U7494 ; P1_U2431
g12395 and P1_U3455 P1_U3360 ; P1_U2432
g12396 and P1_U4540 P1_U3455 ; P1_U2433
g12397 and P1_U7696 P1_U3360 ; P1_U2434
g12398 and P1_U4540 P1_U7696 ; P1_U2435
g12399 and P1_U3235 P1_U3301 ; P1_U2436
g12400 and P1_U4543 P1_U3301 ; P1_U2437
g12401 and P1_R2182_U42 P1_R2182_U25 ; P1_U2438
g12402 and P1_R2182_U42 P1_U3316 ; P1_U2439
g12403 and P1_R2182_U25 P1_U3317 ; P1_U2440
g12404 nor P1_R2182_U42 P1_R2182_U25 ; P1_U2441
g12405 and P1_R2182_U33 P1_R2182_U34 ; P1_U2442
g12406 and P1_R2182_U33 P1_U3318 ; P1_U2443
g12407 and P1_R2182_U34 P1_U3319 ; P1_U2444
g12408 nor P1_R2182_U33 P1_R2182_U34 ; P1_U2445
g12409 and P1_U3471 P1_STATE2_REG_1__SCAN_IN ; P1_U2446
g12410 and P1_U3577 P1_U2452 ; P1_U2447
g12411 and P1_R2167_U17 P1_U3284 ; P1_U2448
g12412 and P1_U4494 P1_U3271 ; P1_U2449
g12413 and P1_U4400 P1_STATE2_REG_0__SCAN_IN ; P1_U2450
g12414 and P1_U4251 P1_STATE2_REG_0__SCAN_IN ; P1_U2451
g12415 and P1_U4400 P1_U3277 P1_U3391 P1_U4173 ; P1_U2452
g12416 and P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2453
g12417 and P1_U3266 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U2454
g12418 and P1_U3266 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U2455
g12419 and P1_U3265 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2456
g12420 and P1_U3265 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2457
g12421 and P1_U3507 P1_U4378 ; P1_U2458
g12422 and P1_U3264 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2459
g12423 and P1_U3264 P1_U3266 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U2460
g12424 and P1_U3506 P1_U3505 ; P1_U2461
g12425 and P1_U3264 P1_U3265 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2462
g12426 and P1_U3504 P1_U3503 ; P1_U2463
g12427 and P1_U4380 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U2464
g12428 and P1_U3502 P1_U3501 ; P1_U2465
g12429 and P1_U3500 P1_U3499 ; P1_U2466
g12430 and P1_U3270 P1_U4378 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U2467
g12431 and P1_U3498 P1_U3497 ; P1_U2468
g12432 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U2469
g12433 and P1_U3266 P1_U2469 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U2470
g12434 and P1_U3265 P1_U2469 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2471
g12435 and P1_U4380 P1_U3270 ; P1_U2472
g12436 and P1_U7680 P1_U7679 P1_U3406 ; P1_U2473
g12437 and P1_R2144_U49 P1_U3312 ; P1_U2474
g12438 and P1_U3454 P1_U3358 ; P1_U2475
g12439 and P1_R2144_U8 P1_R2144_U49 ; P1_U2476
g12440 and P1_U4528 P1_U2476 ; P1_U2477
g12441 and P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U2478
g12442 and P1_U3303 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U2479
g12443 and P1_U3315 P1_U4548 ; P1_U2480
g12444 and P1_U4524 P1_U2476 ; P1_U2481
g12445 and P1_U3327 P1_U4606 ; P1_U2482
g12446 and P1_U4525 P1_U2476 ; P1_U2483
g12447 and P1_U3334 P1_U4665 ; P1_U2484
g12448 and P1_U4526 P1_R2144_U43 ; P1_U2485
g12449 nor P1_R2144_U43 P1_R2144_U50 ; P1_U2486
g12450 and P1_U2486 P1_U2476 ; P1_U2487
g12451 nor P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_U2488
g12452 and P1_U3338 P1_U4722 ; P1_U2489
g12453 and P1_U7693 P1_U3358 ; P1_U2490
g12454 and P1_U4529 P1_U4528 ; P1_U2491
g12455 and P1_U3343 P1_U4780 ; P1_U2492
g12456 and P1_U4529 P1_U4524 ; P1_U2493
g12457 and P1_U3347 P1_U4837 ; P1_U2494
g12458 and P1_U4529 P1_U4525 ; P1_U2495
g12459 and P1_U3350 P1_U4895 ; P1_U2496
g12460 and P1_U4529 P1_U2486 ; P1_U2497
g12461 and P1_U3354 P1_U4952 ; P1_U2498
g12462 and P1_U4531 P1_U3454 ; P1_U2499
g12463 and P1_U3359 P1_U3357 ; P1_U2500
g12464 and P1_U4524 P1_U2474 ; P1_U2501
g12465 and P1_U3364 P1_U5065 ; P1_U2502
g12466 and P1_U4525 P1_U2474 ; P1_U2503
g12467 and P1_U3367 P1_U5123 ; P1_U2504
g12468 and P1_U2486 P1_U2474 ; P1_U2505
g12469 and P1_U3371 P1_U5180 ; P1_U2506
g12470 and P1_U4531 P1_U7693 ; P1_U2507
g12471 nor P1_R2144_U49 P1_R2144_U8 ; P1_U2508
g12472 and P1_U2508 P1_U4528 ; P1_U2509
g12473 nor P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U2510
g12474 and P1_U3374 P1_U5238 ; P1_U2511
g12475 and P1_U2508 P1_U4524 ; P1_U2512
g12476 and P1_U3378 P1_U5295 ; P1_U2513
g12477 and P1_U2508 P1_U4525 ; P1_U2514
g12478 and P1_U3381 P1_U5353 ; P1_U2515
g12479 and P1_U2508 P1_U2486 ; P1_U2516
g12480 and P1_U3385 P1_U5410 ; P1_U2517
g12481 and P1_U7700 P1_U7699 P1_U5468 ; P1_U2518
g12482 and P1_U3744 P1_U5499 ; P1_U2519
g12483 and P1_U4219 P1_U3446 ; P1_U2520
g12484 and P1_U3402 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2521
g12485 and P1_U5483 P1_U5511 ; P1_U2522
g12486 and P1_U2522 P1_U2521 ; P1_U2523
g12487 and P1_U3266 P1_U3402 ; P1_U2524
g12488 and P1_U2522 P1_U2524 ; P1_U2525
g12489 and P1_U5519 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U2526
g12490 and P1_U2522 P1_U2526 ; P1_U2527
g12491 and P1_U5519 P1_U3266 ; P1_U2528
g12492 and P1_U2522 P1_U2528 ; P1_U2529
g12493 and P1_U5483 P1_U3401 ; P1_U2530
g12494 and P1_U2530 P1_U2521 ; P1_U2531
g12495 and P1_U2530 P1_U2524 ; P1_U2532
g12496 and P1_U2530 P1_U2526 ; P1_U2533
g12497 and P1_U2530 P1_U2528 ; P1_U2534
g12498 and P1_U5511 P1_U3438 ; P1_U2535
g12499 and P1_U2535 P1_U2521 ; P1_U2536
g12500 and P1_U2535 P1_U2524 ; P1_U2537
g12501 and P1_U2535 P1_U2526 ; P1_U2538
g12502 and P1_U2535 P1_U2528 ; P1_U2539
g12503 and P1_U3438 P1_U3401 ; P1_U2540
g12504 and P1_U2521 P1_U2540 ; P1_U2541
g12505 and P1_U2524 P1_U2540 ; P1_U2542
g12506 and P1_U2526 P1_U2540 ; P1_U2543
g12507 and P1_U2528 P1_U2540 ; P1_U2544
g12508 and P1_U5480 P1_U7720 ; P1_U2545
g12509 and P1_U2545 P1_U2454 ; P1_U2546
g12510 and P1_U2545 P1_U3498 ; P1_U2547
g12511 and P1_U2545 P1_U4378 ; P1_U2548
g12512 and P1_U2545 P1_U2456 ; P1_U2549
g12513 and P1_U5480 P1_U3456 ; P1_U2550
g12514 and P1_U2550 P1_U2454 ; P1_U2551
g12515 and P1_U2550 P1_U3498 ; P1_U2552
g12516 and P1_U2550 P1_U4378 ; P1_U2553
g12517 and P1_U2550 P1_U2456 ; P1_U2554
g12518 and P1_U7720 P1_U3442 ; P1_U2555
g12519 and P1_U2555 P1_U2454 ; P1_U2556
g12520 and P1_U2555 P1_U3498 ; P1_U2557
g12521 and P1_U2555 P1_U4378 ; P1_U2558
g12522 and P1_U2555 P1_U2456 ; P1_U2559
g12523 and P1_U3456 P1_U3442 ; P1_U2560
g12524 and P1_U2560 P1_U2454 ; P1_U2561
g12525 and P1_U2560 P1_U3498 ; P1_U2562
g12526 and P1_U2560 P1_U4378 ; P1_U2563
g12527 and P1_U2560 P1_U2456 ; P1_U2564
g12528 and P1_U7065 P1_U4379 ; P1_U2565
g12529 and P1_U7065 P1_U2460 ; P1_U2566
g12530 and P1_U7065 P1_U2462 ; P1_U2567
g12531 and P1_U7065 P1_U4380 ; P1_U2568
g12532 and P1_U7065 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U2569
g12533 and P1_U2569 P1_U3498 ; P1_U2570
g12534 and P1_U2569 P1_U2454 ; P1_U2571
g12535 and P1_U2569 P1_U2456 ; P1_U2572
g12536 and P1_U2569 P1_U4378 ; P1_U2573
g12537 and P1_U4379 P1_U3445 ; P1_U2574
g12538 and P1_U2460 P1_U3445 ; P1_U2575
g12539 and P1_U2462 P1_U3445 ; P1_U2576
g12540 and P1_U4380 P1_U3445 ; P1_U2577
g12541 and P1_U3445 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U2578
g12542 and P1_U2578 P1_U3498 ; P1_U2579
g12543 and P1_U2578 P1_U2454 ; P1_U2580
g12544 and P1_U2578 P1_U2456 ; P1_U2581
g12545 and P1_U2578 P1_U4378 ; P1_U2582
g12546 and P1_U7790 P1_U4184 ; P1_U2583
g12547 and P1_U2583 P1_U2524 ; P1_U2584
g12548 and P1_U2583 P1_U2521 ; P1_U2585
g12549 and P1_U2583 P1_U2528 ; P1_U2586
g12550 and P1_U2583 P1_U2526 ; P1_U2587
g12551 and P1_U7790 P1_U3452 ; P1_U2588
g12552 and P1_U2588 P1_U2524 ; P1_U2589
g12553 and P1_U2588 P1_U2521 ; P1_U2590
g12554 and P1_U2588 P1_U2528 ; P1_U2591
g12555 and P1_U2588 P1_U2526 ; P1_U2592
g12556 and P1_U4184 P1_U3457 ; P1_U2593
g12557 and P1_U2593 P1_U2524 ; P1_U2594
g12558 and P1_U2593 P1_U2521 ; P1_U2595
g12559 and P1_U2593 P1_U2528 ; P1_U2596
g12560 and P1_U2593 P1_U2526 ; P1_U2597
g12561 and P1_U3457 P1_U3452 ; P1_U2598
g12562 and P1_U2598 P1_U2524 ; P1_U2599
g12563 and P1_U2598 P1_U2521 ; P1_U2600
g12564 and P1_U2598 P1_U2528 ; P1_U2601
g12565 and P1_U2598 P1_U2526 ; P1_U2602
g12566 and P1_U3389 P1_STATE2_REG_0__SCAN_IN ; P1_U2603
g12567 and P1_U2379 P1_EBX_REG_31__SCAN_IN ; P1_U2604
g12568 and P1_U3533 P1_U2607 P1_U3532 P1_U3531 P1_U3530 ; P1_U2605
g12569 and P1_U7504 P1_U3427 ; P1_U2606
g12570 and P1_U7672 P1_U7671 ; P1_U2607
g12571 and P1_U7787 P1_U7786 ; P1_U2608
g12572 nand P1_U6853 P1_U6854 P1_U6855 ; P1_U2609
g12573 nand P1_U6856 P1_U4026 ; P1_U2610
g12574 nand P1_U6841 P1_U6842 P1_U6843 ; P1_U2611
g12575 nand P1_U6844 P1_U6845 P1_U6846 ; P1_U2612
g12576 nand P1_U6847 P1_U6848 P1_U6849 ; P1_U2613
g12577 nand P1_U6756 P1_U4005 ; P1_U2614
g12578 nand P1_U6753 P1_U4004 ; P1_U2615
g12579 nand P1_U6850 P1_U6851 P1_U6852 ; P1_U2616
g12580 nand P1_U6750 P1_U4003 ; P1_U2617
g12581 nand P1_U6747 P1_U4002 ; P1_U2618
g12582 and P1_R2144_U145 P1_U6746 ; P1_U2620
g12583 and P1_R2144_U145 P1_U6746 ; P1_U2621
g12584 and P1_R2144_U145 P1_U6746 ; P1_U2622
g12585 and P1_R2144_U145 P1_U6746 ; P1_U2623
g12586 and P1_R2144_U145 P1_U6746 ; P1_U2624
g12587 and P1_R2144_U145 P1_U6746 ; P1_U2625
g12588 and P1_R2144_U145 P1_U6746 ; P1_U2626
g12589 and P1_R2144_U145 P1_U6746 ; P1_U2627
g12590 and P1_R2144_U145 P1_U6746 ; P1_U2628
g12591 and P1_R2144_U145 P1_U6746 ; P1_U2629
g12592 and P1_R2144_U145 P1_U6746 ; P1_U2630
g12593 and P1_R2144_U145 P1_U6746 ; P1_U2631
g12594 and P1_R2144_U145 P1_U6746 ; P1_U2632
g12595 and P1_R2144_U145 P1_U6746 ; P1_U2633
g12596 and P1_R2144_U11 P1_U6746 ; P1_U2634
g12597 and P1_R2144_U37 P1_U6746 ; P1_U2635
g12598 and P1_R2144_U38 P1_U6746 ; P1_U2636
g12599 and P1_R2144_U39 P1_U6746 ; P1_U2637
g12600 and P1_R2144_U40 P1_U6746 ; P1_U2638
g12601 and P1_R2144_U41 P1_U6746 ; P1_U2639
g12602 and P1_R2144_U42 P1_U6746 ; P1_U2640
g12603 and P1_R2144_U30 P1_U6746 ; P1_U2641
g12604 and P1_R2144_U80 P1_U6746 ; P1_U2642
g12605 and P1_R2144_U10 P1_U6746 ; P1_U2643
g12606 and P1_R2144_U9 P1_U6746 ; P1_U2644
g12607 and P1_R2144_U45 P1_U6746 ; P1_U2645
g12608 and P1_R2144_U47 P1_U6746 ; P1_U2646
g12609 and P1_R2144_U8 P1_U6746 ; P1_U2647
g12610 nand P1_U3440 P1_U6869 ; P1_U2648
g12611 and P1_R2144_U50 P1_U6746 ; P1_U2649
g12612 and P1_U6870 P1_STATE2_REG_2__SCAN_IN ; P1_U2650
g12613 nand P1_U6769 P1_U6768 P1_U6770 ; P1_U2651
g12614 nand P1_U6771 P1_U4009 ; P1_U2652
g12615 nand P1_U6780 P1_U4011 ; P1_U2653
g12616 nand P1_U6784 P1_U4012 ; P1_U2654
g12617 nand P1_U6788 P1_U4013 ; P1_U2655
g12618 nand P1_U6792 P1_U4014 ; P1_U2656
g12619 nand P1_U6796 P1_U4015 ; P1_U2657
g12620 nand P1_U6800 P1_U4016 ; P1_U2658
g12621 nand P1_U6804 P1_U4017 ; P1_U2659
g12622 nand P1_U6808 P1_U4018 ; P1_U2660
g12623 nand P1_U6812 P1_U4019 ; P1_U2661
g12624 nand P1_U6816 P1_U4020 ; P1_U2662
g12625 nand P1_U6825 P1_U4022 ; P1_U2663
g12626 nand P1_U6829 P1_U4023 ; P1_U2664
g12627 nand P1_U6833 P1_U4024 ; P1_U2665
g12628 nand P1_U6837 P1_U4025 ; P1_U2666
g12629 nand P1_U6759 P1_U4006 ; P1_U2667
g12630 nand P1_U6767 P1_U6766 P1_U4008 P1_U6763 ; P1_U2668
g12631 nand P1_U6779 P1_U6778 P1_U4010 P1_U6775 ; P1_U2669
g12632 nand P1_U6824 P1_U6823 P1_U4021 P1_U6820 ; P1_U2670
g12633 nand P1_U6863 P1_U6862 P1_U4027 P1_U6859 ; P1_U2671
g12634 nand P1_U6866 P1_U6864 P1_U6865 P1_U6868 P1_U6867 ; P1_U2672
g12635 nand P1_U7458 P1_U7457 ; P1_U2673
g12636 nand P1_U7460 P1_U7459 ; P1_U2674
g12637 nand P1_U4168 P1_U7463 ; P1_U2675
g12638 nand P1_U4169 P1_U7466 ; P1_U2676
g12639 nand P1_U7794 P1_U7793 P1_U7467 ; P1_U2677
g12640 nand P1_U7456 P1_U3284 ; P1_U2678
g12641 nand P1_U7405 P1_U7404 ; P1_U2679
g12642 nand P1_U7407 P1_U7406 ; P1_U2680
g12643 nand P1_U7411 P1_U7410 ; P1_U2681
g12644 nand P1_U7413 P1_U7412 ; P1_U2682
g12645 nand P1_U7415 P1_U7414 ; P1_U2683
g12646 nand P1_U7417 P1_U7416 ; P1_U2684
g12647 nand P1_U7419 P1_U7418 ; P1_U2685
g12648 nand P1_U7421 P1_U7420 ; P1_U2686
g12649 nand P1_U7423 P1_U7422 ; P1_U2687
g12650 nand P1_U7425 P1_U7424 ; P1_U2688
g12651 nand P1_U7427 P1_U7426 ; P1_U2689
g12652 nand P1_U7429 P1_U7428 ; P1_U2690
g12653 nand P1_U7433 P1_U7432 ; P1_U2691
g12654 nand P1_U7435 P1_U7434 ; P1_U2692
g12655 nand P1_U7437 P1_U7436 ; P1_U2693
g12656 nand P1_U7439 P1_U7438 ; P1_U2694
g12657 nand P1_U7441 P1_U7440 ; P1_U2695
g12658 nand P1_U7443 P1_U7442 ; P1_U2696
g12659 nand P1_U7445 P1_U7444 ; P1_U2697
g12660 nand P1_U7447 P1_U7446 ; P1_U2698
g12661 nand P1_U7449 P1_U7448 ; P1_U2699
g12662 nand P1_U7451 P1_U7450 ; P1_U2700
g12663 nand P1_U7393 P1_U7392 ; P1_U2701
g12664 nand P1_U7395 P1_U7394 ; P1_U2702
g12665 nand P1_U7397 P1_U7396 ; P1_U2703
g12666 nand P1_U7399 P1_U7398 ; P1_U2704
g12667 nand P1_U7401 P1_U7400 ; P1_U2705
g12668 nand P1_U7403 P1_U7402 ; P1_U2706
g12669 nand P1_U7409 P1_U7408 ; P1_U2707
g12670 nand P1_U7431 P1_U7430 ; P1_U2708
g12671 nand P1_U7453 P1_U7452 ; P1_U2709
g12672 nand P1_U7455 P1_U7454 ; P1_U2710
g12673 nand P1_U7377 P1_U7376 ; P1_U2711
g12674 nand P1_U7379 P1_U7378 ; P1_U2712
g12675 nand P1_U4165 P1_U4239 ; P1_U2713
g12676 nand P1_U7386 P1_U7385 P1_U4166 P1_U3434 ; P1_U2714
g12677 nand P1_U4239 P1_U4167 ; P1_U2715
g12678 nand P1_U7365 P1_U7364 ; P1_U2716
g12679 nand P1_U7367 P1_U7366 ; P1_U2717
g12680 nand P1_U4161 P1_U7368 ; P1_U2718
g12681 nand P1_U4162 P1_U7370 ; P1_U2719
g12682 nand P1_U4163 P1_U7372 ; P1_U2720
g12683 nand P1_U4164 P1_U7374 ; P1_U2721
g12684 nand P1_U4159 P1_U4192 ; P1_U2722
g12685 and P1_U7236 P1_U7083 ; P1_U2723
g12686 and P1_U7253 P1_U7083 ; P1_U2724
g12687 and P1_U7270 P1_U7083 ; P1_U2725
g12688 and P1_U7620 P1_U7083 ; P1_U2726
g12689 and P1_U7302 P1_U7083 ; P1_U2727
g12690 and P1_U7319 P1_U7083 ; P1_U2728
g12691 and P1_U7336 P1_U7083 ; P1_U2729
g12692 and P1_U7353 P1_U7083 ; P1_U2730
g12693 nand P1_U2606 P1_U7354 ; P1_U2731
g12694 and P1_U7083 P1_U7082 ; P1_U2732
g12695 and P1_U7114 P1_U7083 ; P1_U2733
g12696 and P1_U7131 P1_U7083 ; P1_U2734
g12697 and P1_U7618 P1_U7083 ; P1_U2735
g12698 and P1_U7163 P1_U7083 ; P1_U2736
g12699 and P1_U7180 P1_U7083 ; P1_U2737
g12700 and P1_U7197 P1_U7083 ; P1_U2738
g12701 and P1_U7214 P1_U7083 ; P1_U2739
g12702 and P1_U7063 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_U2740
g12703 nand P1_U4078 P1_U7096 ; P1_U2741
g12704 and P1_U7492 P1_U7491 ; P1_U2742
g12705 and P1_U7506 P1_U7470 ; P1_U2743
g12706 and P1_U7479 P1_U7478 ; P1_U2744
g12707 nand P1_U7048 P1_U7047 ; P1_U2745
g12708 nand P1_U7050 P1_U7049 ; P1_U2746
g12709 nand P1_U7052 P1_U7051 ; P1_U2747
g12710 nand P1_U7616 P1_U7053 ; P1_U2748
g12711 nand P1_U7055 P1_U7054 ; P1_U2749
g12712 nand P1_U7057 P1_U7056 ; P1_U2750
g12713 nand P1_U4061 P1_U7058 ; P1_U2751
g12714 nand P1_U4062 P1_U7060 P1_U7061 ; P1_U2752
g12715 and P1_U6957 P1_U6909 ; P1_U2753
g12716 and P1_U6974 P1_U6909 ; P1_U2754
g12717 and P1_U6991 P1_U6909 ; P1_U2755
g12718 and P1_U7615 P1_U6909 ; P1_U2756
g12719 and P1_U7023 P1_U6909 ; P1_U2757
g12720 and P1_U7040 P1_U6909 ; P1_U2758
g12721 and P1_U6909 P1_U6908 ; P1_U2759
g12722 and P1_U6926 P1_U6909 ; P1_U2760
g12723 nand P1_U6928 P1_U6927 ; P1_U2761
g12724 nand P1_U6930 P1_U6929 ; P1_U2762
g12725 nand P1_U6932 P1_U6931 ; P1_U2763
g12726 nand P1_U6934 P1_U6933 ; P1_U2764
g12727 nand P1_U6936 P1_U6935 P1_U6937 ; P1_U2765
g12728 nand P1_U6939 P1_U6938 P1_U6940 ; P1_U2766
g12729 nand P1_U7043 P1_U7041 P1_U7042 ; P1_U2767
g12730 nand P1_U7046 P1_U7044 P1_U7045 ; P1_U2768
g12731 and P1_R2144_U145 P1_U4159 ; P1_U2769
g12732 and P1_U4159 P1_R2144_U145 ; P1_U2770
g12733 and P1_U4159 P1_R2144_U145 ; P1_U2771
g12734 and P1_U4159 P1_R2144_U145 ; P1_U2772
g12735 and P1_U4159 P1_R2144_U145 ; P1_U2773
g12736 and P1_U4159 P1_R2144_U145 ; P1_U2774
g12737 and P1_U4159 P1_R2144_U145 ; P1_U2775
g12738 and P1_U4159 P1_R2144_U145 ; P1_U2776
g12739 and P1_U4159 P1_R2144_U145 ; P1_U2777
g12740 and P1_U4159 P1_R2144_U145 ; P1_U2778
g12741 and P1_U4159 P1_R2144_U145 ; P1_U2779
g12742 and P1_U4159 P1_R2144_U145 ; P1_U2780
g12743 and P1_U4159 P1_R2144_U145 ; P1_U2781
g12744 and P1_U4159 P1_R2144_U145 ; P1_U2782
g12745 and P1_U4159 P1_R2144_U145 ; P1_U2783
g12746 and P1_U4159 P1_R2144_U11 ; P1_U2784
g12747 and P1_U4159 P1_R2144_U37 ; P1_U2785
g12748 and P1_U4159 P1_R2144_U38 ; P1_U2786
g12749 and P1_U4159 P1_R2144_U39 ; P1_U2787
g12750 and P1_U4159 P1_R2144_U40 ; P1_U2788
g12751 and P1_U4159 P1_R2144_U41 ; P1_U2789
g12752 and P1_U4159 P1_R2144_U42 ; P1_U2790
g12753 and P1_U4159 P1_R2144_U30 ; P1_U2791
g12754 nand P1_U6872 P1_U6871 ; P1_U2792
g12755 nand P1_U6874 P1_U6873 ; P1_U2793
g12756 nand P1_U6876 P1_U6875 ; P1_U2794
g12757 nand P1_U6878 P1_U6877 ; P1_U2795
g12758 nand P1_U6880 P1_U6879 ; P1_U2796
g12759 nand P1_U6882 P1_U6881 ; P1_U2797
g12760 nand P1_U6884 P1_U6885 P1_U6883 ; P1_U2798
g12761 nand P1_U4028 P1_U6887 P1_U6886 ; P1_U2799
g12762 nand P1_U6890 P1_U6891 P1_U6889 ; P1_U2800
g12763 nand P1_U6617 P1_U3432 P1_U7498 ; P1_U2801
g12764 nand P1_U7650 P1_U6613 ; P1_U2802
g12765 nand P1_U6612 P1_U6611 ; P1_U2803
g12766 nand P1_U7769 P1_U7768 P1_U4243 ; P1_U2804
g12767 nand P1_U7765 P1_U7764 P1_U4243 ; P1_U2805
g12768 nand P1_U6601 P1_U4248 ; P1_U2806
g12769 nand P1_U7757 P1_U7756 P1_U4240 ; P1_U2807
g12770 nand P1_U7747 P1_U7746 P1_U4240 ; P1_U2808
g12771 nand P1_U6593 P1_U3948 P1_U3949 P1_U6591 P1_U6595 ; P1_U2809
g12772 nand P1_U6586 P1_U3946 P1_U3947 P1_U6584 P1_U6588 ; P1_U2810
g12773 nand P1_U6579 P1_U3944 P1_U3945 P1_U6577 P1_U6581 ; P1_U2811
g12774 nand P1_U6572 P1_U3942 P1_U3943 P1_U6570 P1_U6574 ; P1_U2812
g12775 nand P1_U6565 P1_U3940 P1_U3941 P1_U6563 P1_U6567 ; P1_U2813
g12776 nand P1_U6558 P1_U3938 P1_U3939 P1_U6556 P1_U6560 ; P1_U2814
g12777 nand P1_U6551 P1_U3936 P1_U3937 P1_U6549 P1_U6553 ; P1_U2815
g12778 nand P1_U6544 P1_U3934 P1_U3935 P1_U6542 P1_U6546 ; P1_U2816
g12779 nand P1_U6537 P1_U3932 P1_U3933 P1_U6535 P1_U6539 ; P1_U2817
g12780 nand P1_U6530 P1_U3930 P1_U3931 P1_U6528 P1_U6532 ; P1_U2818
g12781 nand P1_U6523 P1_U3928 P1_U3929 P1_U6521 P1_U6525 ; P1_U2819
g12782 nand P1_U6516 P1_U3926 P1_U3927 P1_U6514 P1_U6518 ; P1_U2820
g12783 nand P1_U3924 P1_U6509 P1_U3925 P1_U6507 P1_U6511 ; P1_U2821
g12784 nand P1_U3922 P1_U6502 P1_U3923 P1_U6500 P1_U6504 ; P1_U2822
g12785 nand P1_U3920 P1_U6495 P1_U3921 P1_U6493 P1_U6497 ; P1_U2823
g12786 nand P1_U6488 P1_U6487 P1_U3919 P1_U3918 P1_U6490 ; P1_U2824
g12787 nand P1_U6481 P1_U6480 P1_U3917 P1_U3916 P1_U6483 ; P1_U2825
g12788 nand P1_U3915 P1_U6474 P1_U3914 P1_U6473 P1_U6476 ; P1_U2826
g12789 nand P1_U3913 P1_U6467 P1_U3912 P1_U6466 P1_U6469 ; P1_U2827
g12790 nand P1_U3911 P1_U6460 P1_U3910 P1_U6459 P1_U6462 ; P1_U2828
g12791 nand P1_U3909 P1_U6453 P1_U3908 P1_U6452 P1_U6455 ; P1_U2829
g12792 nand P1_U3907 P1_U6446 P1_U3906 P1_U6445 P1_U6448 ; P1_U2830
g12793 nand P1_U3905 P1_U6439 P1_U3904 P1_U6438 P1_U6441 ; P1_U2831
g12794 nand P1_U3903 P1_U6432 P1_U3902 P1_U6431 P1_U6434 ; P1_U2832
g12795 nand P1_U3901 P1_U6425 P1_U3900 P1_U6424 P1_U6427 ; P1_U2833
g12796 nand P1_U3899 P1_U6418 P1_U3898 P1_U6417 P1_U6420 ; P1_U2834
g12797 nand P1_U3896 P1_U6409 P1_U6410 P1_U3897 ; P1_U2835
g12798 nand P1_U3894 P1_U6401 P1_U3895 P1_U6403 P1_U6402 ; P1_U2836
g12799 nand P1_U6393 P1_U6392 P1_U6394 P1_U3893 ; P1_U2837
g12800 nand P1_U6385 P1_U6384 P1_U6386 P1_U3892 ; P1_U2838
g12801 nand P1_U6377 P1_U6376 P1_U6378 P1_U3891 ; P1_U2839
g12802 nand P1_U6369 P1_U6368 P1_U6370 P1_U3890 ; P1_U2840
g12803 nand P1_U6359 P1_U6358 ; P1_U2841
g12804 nand P1_U6356 P1_U6357 P1_U6355 ; P1_U2842
g12805 nand P1_U6353 P1_U6354 P1_U6352 ; P1_U2843
g12806 nand P1_U6350 P1_U6351 P1_U6349 ; P1_U2844
g12807 nand P1_U6347 P1_U6348 P1_U6346 ; P1_U2845
g12808 nand P1_U6344 P1_U6345 P1_U6343 ; P1_U2846
g12809 nand P1_U6341 P1_U6342 P1_U6340 ; P1_U2847
g12810 nand P1_U6338 P1_U6339 P1_U6337 ; P1_U2848
g12811 nand P1_U6335 P1_U6336 P1_U6334 ; P1_U2849
g12812 nand P1_U6332 P1_U6333 P1_U6331 ; P1_U2850
g12813 nand P1_U6329 P1_U6330 P1_U6328 ; P1_U2851
g12814 nand P1_U6326 P1_U6327 P1_U6325 ; P1_U2852
g12815 nand P1_U6323 P1_U6324 P1_U6322 ; P1_U2853
g12816 nand P1_U6320 P1_U6321 P1_U6319 ; P1_U2854
g12817 nand P1_U6317 P1_U6318 P1_U6316 ; P1_U2855
g12818 nand P1_U6314 P1_U6315 P1_U6313 ; P1_U2856
g12819 nand P1_U6311 P1_U6312 P1_U6310 ; P1_U2857
g12820 nand P1_U6308 P1_U6309 P1_U6307 ; P1_U2858
g12821 nand P1_U6305 P1_U6306 P1_U6304 ; P1_U2859
g12822 nand P1_U6302 P1_U6303 P1_U6301 ; P1_U2860
g12823 nand P1_U6299 P1_U6300 P1_U6298 ; P1_U2861
g12824 nand P1_U6296 P1_U6297 P1_U6295 ; P1_U2862
g12825 nand P1_U6293 P1_U6294 P1_U6292 ; P1_U2863
g12826 nand P1_U6290 P1_U6291 P1_U6289 ; P1_U2864
g12827 nand P1_U6287 P1_U6288 P1_U6286 ; P1_U2865
g12828 nand P1_U6284 P1_U6285 P1_U6283 ; P1_U2866
g12829 nand P1_U6281 P1_U6282 P1_U6280 ; P1_U2867
g12830 nand P1_U6278 P1_U6279 P1_U6277 ; P1_U2868
g12831 nand P1_U6275 P1_U6276 P1_U6274 ; P1_U2869
g12832 nand P1_U6272 P1_U6273 P1_U6271 ; P1_U2870
g12833 nand P1_U6269 P1_U6270 P1_U6268 ; P1_U2871
g12834 nand P1_U6266 P1_U6265 P1_U6267 ; P1_U2872
g12835 nand P1_U4176 P1_U6262 ; P1_U2873
g12836 nand P1_U6259 P1_U6258 P1_U6261 P1_U6260 ; P1_U2874
g12837 nand P1_U6255 P1_U6254 P1_U6257 P1_U6256 ; P1_U2875
g12838 nand P1_U6251 P1_U6250 P1_U6253 P1_U6252 ; P1_U2876
g12839 nand P1_U6247 P1_U6246 P1_U6249 P1_U6248 ; P1_U2877
g12840 nand P1_U6243 P1_U6242 P1_U6245 P1_U6244 ; P1_U2878
g12841 nand P1_U6239 P1_U6238 P1_U6241 P1_U6240 ; P1_U2879
g12842 nand P1_U6235 P1_U6234 P1_U6237 P1_U6236 ; P1_U2880
g12843 nand P1_U6231 P1_U6230 P1_U6233 P1_U6232 ; P1_U2881
g12844 nand P1_U6227 P1_U6226 P1_U6229 P1_U6228 ; P1_U2882
g12845 nand P1_U6223 P1_U6222 P1_U6225 P1_U6224 ; P1_U2883
g12846 nand P1_U6219 P1_U6218 P1_U6221 P1_U6220 ; P1_U2884
g12847 nand P1_U6215 P1_U6214 P1_U6217 P1_U6216 ; P1_U2885
g12848 nand P1_U6211 P1_U6210 P1_U6213 P1_U6212 ; P1_U2886
g12849 nand P1_U6207 P1_U6206 P1_U6209 P1_U6208 ; P1_U2887
g12850 nand P1_U6203 P1_U6202 P1_U6205 P1_U6204 ; P1_U2888
g12851 nand P1_U6201 P1_U6199 P1_U6200 ; P1_U2889
g12852 nand P1_U6198 P1_U6196 P1_U6197 ; P1_U2890
g12853 nand P1_U6195 P1_U6193 P1_U6194 ; P1_U2891
g12854 nand P1_U6192 P1_U6190 P1_U6191 ; P1_U2892
g12855 nand P1_U6189 P1_U6187 P1_U6188 ; P1_U2893
g12856 nand P1_U6186 P1_U6184 P1_U6185 ; P1_U2894
g12857 nand P1_U6183 P1_U6181 P1_U6182 ; P1_U2895
g12858 nand P1_U6180 P1_U6178 P1_U6179 ; P1_U2896
g12859 nand P1_U6177 P1_U6175 P1_U6176 ; P1_U2897
g12860 nand P1_U6174 P1_U6172 P1_U6173 ; P1_U2898
g12861 nand P1_U6171 P1_U6169 P1_U6170 ; P1_U2899
g12862 nand P1_U6168 P1_U6166 P1_U6167 ; P1_U2900
g12863 nand P1_U6165 P1_U6163 P1_U6164 ; P1_U2901
g12864 nand P1_U6162 P1_U6160 P1_U6161 ; P1_U2902
g12865 nand P1_U6158 P1_U6157 P1_U6159 ; P1_U2903
g12866 nand P1_U6155 P1_U6154 P1_U6156 ; P1_U2904
g12867 and P1_U6055 P1_DATAO_REG_31__SCAN_IN ; P1_U2905
g12868 nand P1_U3882 P1_U6146 ; P1_U2906
g12869 nand P1_U3881 P1_U6143 ; P1_U2907
g12870 nand P1_U3880 P1_U6140 ; P1_U2908
g12871 nand P1_U3879 P1_U6137 ; P1_U2909
g12872 nand P1_U3878 P1_U6134 ; P1_U2910
g12873 nand P1_U3877 P1_U6131 ; P1_U2911
g12874 nand P1_U3876 P1_U6128 ; P1_U2912
g12875 nand P1_U3875 P1_U6125 ; P1_U2913
g12876 nand P1_U3874 P1_U6122 ; P1_U2914
g12877 nand P1_U3873 P1_U6119 ; P1_U2915
g12878 nand P1_U3872 P1_U6116 ; P1_U2916
g12879 nand P1_U3871 P1_U6113 ; P1_U2917
g12880 nand P1_U3870 P1_U6110 ; P1_U2918
g12881 nand P1_U3869 P1_U6107 ; P1_U2919
g12882 nand P1_U3868 P1_U6104 ; P1_U2920
g12883 nand P1_U6102 P1_U6101 P1_U6103 ; P1_U2921
g12884 nand P1_U6099 P1_U6098 P1_U6100 ; P1_U2922
g12885 nand P1_U6096 P1_U6095 P1_U6097 ; P1_U2923
g12886 nand P1_U6093 P1_U6092 P1_U6094 ; P1_U2924
g12887 nand P1_U6090 P1_U6089 P1_U6091 ; P1_U2925
g12888 nand P1_U6087 P1_U6086 P1_U6088 ; P1_U2926
g12889 nand P1_U6084 P1_U6083 P1_U6085 ; P1_U2927
g12890 nand P1_U6081 P1_U6080 P1_U6082 ; P1_U2928
g12891 nand P1_U6078 P1_U6077 P1_U6079 ; P1_U2929
g12892 nand P1_U6075 P1_U6074 P1_U6076 ; P1_U2930
g12893 nand P1_U6072 P1_U6071 P1_U6073 ; P1_U2931
g12894 nand P1_U6069 P1_U6068 P1_U6070 ; P1_U2932
g12895 nand P1_U6066 P1_U6065 P1_U6067 ; P1_U2933
g12896 nand P1_U6063 P1_U6062 P1_U6064 ; P1_U2934
g12897 nand P1_U6060 P1_U6059 P1_U6061 ; P1_U2935
g12898 nand P1_U6057 P1_U6056 P1_U6058 ; P1_U2936
g12899 nand P1_U7540 P1_U7542 ; P1_U2937
g12900 nand P1_U7539 P1_U7544 ; P1_U2938
g12901 nand P1_U7538 P1_U7546 ; P1_U2939
g12902 nand P1_U7537 P1_U7548 ; P1_U2940
g12903 nand P1_U7536 P1_U7550 ; P1_U2941
g12904 nand P1_U7535 P1_U7552 ; P1_U2942
g12905 nand P1_U7534 P1_U7554 ; P1_U2943
g12906 nand P1_U7533 P1_U7556 ; P1_U2944
g12907 nand P1_U7532 P1_U7558 ; P1_U2945
g12908 nand P1_U7531 P1_U7560 ; P1_U2946
g12909 nand P1_U7530 P1_U7562 ; P1_U2947
g12910 nand P1_U7529 P1_U7564 ; P1_U2948
g12911 nand P1_U7528 P1_U7566 ; P1_U2949
g12912 nand P1_U7527 P1_U7568 ; P1_U2950
g12913 nand P1_U7526 P1_U7570 ; P1_U2951
g12914 nand P1_U7525 P1_U7572 ; P1_U2952
g12915 nand P1_U7524 P1_U7574 ; P1_U2953
g12916 nand P1_U7523 P1_U7576 ; P1_U2954
g12917 nand P1_U7522 P1_U7578 ; P1_U2955
g12918 nand P1_U7521 P1_U7580 ; P1_U2956
g12919 nand P1_U7520 P1_U7582 ; P1_U2957
g12920 nand P1_U7519 P1_U7584 ; P1_U2958
g12921 nand P1_U7518 P1_U7586 ; P1_U2959
g12922 nand P1_U7517 P1_U7588 ; P1_U2960
g12923 nand P1_U7516 P1_U7590 ; P1_U2961
g12924 nand P1_U7515 P1_U7592 ; P1_U2962
g12925 nand P1_U7514 P1_U7594 ; P1_U2963
g12926 nand P1_U7513 P1_U7596 ; P1_U2964
g12927 nand P1_U7512 P1_U7598 ; P1_U2965
g12928 nand P1_U7511 P1_U7600 ; P1_U2966
g12929 nand P1_U7510 P1_U7602 ; P1_U2967
g12930 nand P1_U5956 P1_U5954 P1_U5958 P1_U5955 P1_U5957 ; P1_U2968
g12931 nand P1_U5951 P1_U5949 P1_U5953 P1_U5950 P1_U5952 ; P1_U2969
g12932 nand P1_U5946 P1_U5944 P1_U5948 P1_U5945 P1_U5947 ; P1_U2970
g12933 nand P1_U5941 P1_U5939 P1_U5943 P1_U5940 P1_U5942 ; P1_U2971
g12934 nand P1_U5936 P1_U5934 P1_U5938 P1_U5935 P1_U5937 ; P1_U2972
g12935 nand P1_U5931 P1_U5929 P1_U5933 P1_U5930 P1_U5932 ; P1_U2973
g12936 nand P1_U5926 P1_U5924 P1_U5928 P1_U5925 P1_U5927 ; P1_U2974
g12937 nand P1_U5921 P1_U5919 P1_U5923 P1_U5920 P1_U5922 ; P1_U2975
g12938 nand P1_U5916 P1_U5914 P1_U5918 P1_U5915 P1_U5917 ; P1_U2976
g12939 nand P1_U5911 P1_U5909 P1_U5913 P1_U5910 P1_U5912 ; P1_U2977
g12940 nand P1_U5906 P1_U5904 P1_U5908 P1_U5905 P1_U5907 ; P1_U2978
g12941 nand P1_U5901 P1_U5899 P1_U5903 P1_U5900 P1_U5902 ; P1_U2979
g12942 nand P1_U5896 P1_U5894 P1_U5898 P1_U5895 P1_U5897 ; P1_U2980
g12943 nand P1_U5891 P1_U5889 P1_U5893 P1_U5890 P1_U5892 ; P1_U2981
g12944 nand P1_U5886 P1_U5884 P1_U5888 P1_U5885 P1_U5887 ; P1_U2982
g12945 nand P1_U5881 P1_U5879 P1_U5883 P1_U5880 P1_U5882 ; P1_U2983
g12946 nand P1_U5876 P1_U5874 P1_U5878 P1_U5875 P1_U5877 ; P1_U2984
g12947 nand P1_U5871 P1_U5869 P1_U5873 P1_U5870 P1_U5872 ; P1_U2985
g12948 nand P1_U5866 P1_U5864 P1_U5868 P1_U5865 P1_U5867 ; P1_U2986
g12949 nand P1_U5861 P1_U5859 P1_U5863 P1_U5860 P1_U5862 ; P1_U2987
g12950 nand P1_U5856 P1_U5854 P1_U5858 P1_U5855 P1_U5857 ; P1_U2988
g12951 nand P1_U5851 P1_U5849 P1_U5853 P1_U5850 P1_U5852 ; P1_U2989
g12952 nand P1_U5846 P1_U5844 P1_U5848 P1_U5845 P1_U5847 ; P1_U2990
g12953 nand P1_U5841 P1_U5839 P1_U5843 P1_U5840 P1_U5842 ; P1_U2991
g12954 nand P1_U5836 P1_U5834 P1_U5835 P1_U5838 P1_U5837 ; P1_U2992
g12955 nand P1_U5831 P1_U5829 P1_U5830 P1_U5833 P1_U5832 ; P1_U2993
g12956 nand P1_U5826 P1_U5824 P1_U5825 P1_U5828 P1_U5827 ; P1_U2994
g12957 nand P1_U5821 P1_U5819 P1_U5820 P1_U5823 P1_U5822 ; P1_U2995
g12958 nand P1_U5816 P1_U5814 P1_U5815 P1_U5818 P1_U5817 ; P1_U2996
g12959 nand P1_U5811 P1_U5809 P1_U5810 P1_U5813 P1_U5812 ; P1_U2997
g12960 nand P1_U5805 P1_U5804 P1_U5806 P1_U5808 P1_U5807 ; P1_U2998
g12961 nand P1_U5800 P1_U5799 P1_U5801 P1_U5803 P1_U5802 ; P1_U2999
g12962 nand P1_U3861 P1_U3859 P1_U5787 P1_U5789 ; P1_U3000
g12963 nand P1_U3858 P1_U3856 P1_U5780 P1_U5782 ; P1_U3001
g12964 nand P1_U3855 P1_U3853 P1_U5773 P1_U5775 ; P1_U3002
g12965 nand P1_U3852 P1_U3850 P1_U5766 P1_U5768 ; P1_U3003
g12966 nand P1_U3849 P1_U3847 P1_U5759 P1_U5761 ; P1_U3004
g12967 nand P1_U3846 P1_U3844 P1_U5752 P1_U5754 ; P1_U3005
g12968 nand P1_U3843 P1_U3841 P1_U5745 P1_U5747 ; P1_U3006
g12969 nand P1_U3840 P1_U3838 P1_U5738 P1_U5740 ; P1_U3007
g12970 nand P1_U3837 P1_U3835 P1_U5731 P1_U5733 ; P1_U3008
g12971 nand P1_U3834 P1_U3832 P1_U5724 P1_U5726 ; P1_U3009
g12972 nand P1_U3831 P1_U3829 P1_U5717 P1_U5719 ; P1_U3010
g12973 nand P1_U3828 P1_U3826 P1_U5710 P1_U5712 ; P1_U3011
g12974 nand P1_U3825 P1_U3823 P1_U5703 P1_U5705 ; P1_U3012
g12975 nand P1_U3822 P1_U3820 P1_U5696 P1_U5698 ; P1_U3013
g12976 nand P1_U3819 P1_U3817 P1_U5689 P1_U5691 ; P1_U3014
g12977 nand P1_U3816 P1_U3814 P1_U5682 P1_U5684 ; P1_U3015
g12978 nand P1_U3813 P1_U3811 P1_U5675 P1_U5677 ; P1_U3016
g12979 nand P1_U3810 P1_U3808 P1_U5668 P1_U5670 ; P1_U3017
g12980 nand P1_U3807 P1_U3805 P1_U5661 P1_U5663 ; P1_U3018
g12981 nand P1_U3802 P1_U3804 P1_U5656 ; P1_U3019
g12982 nand P1_U3799 P1_U3801 P1_U5649 ; P1_U3020
g12983 nand P1_U3796 P1_U3798 P1_U5642 ; P1_U3021
g12984 nand P1_U3793 P1_U3795 P1_U5635 ; P1_U3022
g12985 nand P1_U3790 P1_U3792 P1_U5628 ; P1_U3023
g12986 nand P1_U3787 P1_U3789 P1_U5621 ; P1_U3024
g12987 nand P1_U3784 P1_U3786 P1_U5614 ; P1_U3025
g12988 nand P1_U3781 P1_U3783 P1_U5607 ; P1_U3026
g12989 nand P1_U3778 P1_U3780 P1_U5600 ; P1_U3027
g12990 nand P1_U3775 P1_U3776 ; P1_U3028
g12991 nand P1_U3772 P1_U3771 P1_U3774 ; P1_U3029
g12992 nand P1_U3768 P1_U3767 P1_U3770 ; P1_U3030
g12993 nand P1_U3764 P1_U3763 P1_U3766 ; P1_U3031
g12994 and P1_U5537 P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_U3032
g12995 nand P1_U5460 P1_U5459 P1_U3730 ; P1_U3033
g12996 nand P1_U5455 P1_U5454 P1_U3729 ; P1_U3034
g12997 nand P1_U5450 P1_U5449 P1_U3728 ; P1_U3035
g12998 nand P1_U5445 P1_U5444 P1_U3727 ; P1_U3036
g12999 nand P1_U7612 P1_U5440 P1_U3726 ; P1_U3037
g13000 nand P1_U5436 P1_U5435 P1_U3725 ; P1_U3038
g13001 nand P1_U5431 P1_U5430 P1_U3724 ; P1_U3039
g13002 nand P1_U5426 P1_U5425 P1_U3723 ; P1_U3040
g13003 nand P1_U5404 P1_U5403 P1_U3721 ; P1_U3041
g13004 nand P1_U5399 P1_U5398 P1_U3720 ; P1_U3042
g13005 nand P1_U5394 P1_U5393 P1_U3719 ; P1_U3043
g13006 nand P1_U5389 P1_U5388 P1_U3718 ; P1_U3044
g13007 nand P1_U5384 P1_U5383 P1_U3717 ; P1_U3045
g13008 nand P1_U5379 P1_U5378 P1_U3716 ; P1_U3046
g13009 nand P1_U5374 P1_U5373 P1_U3715 ; P1_U3047
g13010 nand P1_U5369 P1_U5368 P1_U3714 ; P1_U3048
g13011 nand P1_U5346 P1_U5345 P1_U3712 ; P1_U3049
g13012 nand P1_U5341 P1_U5340 P1_U3711 ; P1_U3050
g13013 nand P1_U5336 P1_U5335 P1_U3710 ; P1_U3051
g13014 nand P1_U5331 P1_U5330 P1_U3709 ; P1_U3052
g13015 nand P1_U5326 P1_U5325 P1_U3708 ; P1_U3053
g13016 nand P1_U5321 P1_U5320 P1_U3707 ; P1_U3054
g13017 nand P1_U5316 P1_U5315 P1_U3706 ; P1_U3055
g13018 nand P1_U5311 P1_U5310 P1_U3705 ; P1_U3056
g13019 nand P1_U5289 P1_U5288 P1_U3703 ; P1_U3057
g13020 nand P1_U5284 P1_U5283 P1_U3702 ; P1_U3058
g13021 nand P1_U5279 P1_U5278 P1_U3701 ; P1_U3059
g13022 nand P1_U5274 P1_U5273 P1_U3700 ; P1_U3060
g13023 nand P1_U5269 P1_U5268 P1_U3699 ; P1_U3061
g13024 nand P1_U5264 P1_U5263 P1_U3698 ; P1_U3062
g13025 nand P1_U5259 P1_U5258 P1_U3697 ; P1_U3063
g13026 nand P1_U5254 P1_U5253 P1_U3696 ; P1_U3064
g13027 nand P1_U5231 P1_U5230 P1_U3694 ; P1_U3065
g13028 nand P1_U5226 P1_U5225 P1_U3693 ; P1_U3066
g13029 nand P1_U5221 P1_U5220 P1_U3692 ; P1_U3067
g13030 nand P1_U5216 P1_U5215 P1_U3691 ; P1_U3068
g13031 nand P1_U5211 P1_U5210 P1_U3690 ; P1_U3069
g13032 nand P1_U5206 P1_U5205 P1_U3689 ; P1_U3070
g13033 nand P1_U5201 P1_U5200 P1_U3688 ; P1_U3071
g13034 nand P1_U5196 P1_U5195 P1_U3687 ; P1_U3072
g13035 nand P1_U5174 P1_U5173 P1_U3685 ; P1_U3073
g13036 nand P1_U5169 P1_U5168 P1_U3684 ; P1_U3074
g13037 nand P1_U5164 P1_U5163 P1_U3683 ; P1_U3075
g13038 nand P1_U5159 P1_U5158 P1_U3682 ; P1_U3076
g13039 nand P1_U5154 P1_U5153 P1_U3681 ; P1_U3077
g13040 nand P1_U5149 P1_U5148 P1_U3680 ; P1_U3078
g13041 nand P1_U5144 P1_U5143 P1_U3679 ; P1_U3079
g13042 nand P1_U5139 P1_U5138 P1_U3678 ; P1_U3080
g13043 nand P1_U5116 P1_U5115 P1_U3676 ; P1_U3081
g13044 nand P1_U5111 P1_U5110 P1_U3675 ; P1_U3082
g13045 nand P1_U5106 P1_U5105 P1_U3674 ; P1_U3083
g13046 nand P1_U5101 P1_U5100 P1_U3673 ; P1_U3084
g13047 nand P1_U5096 P1_U5095 P1_U3672 ; P1_U3085
g13048 nand P1_U5091 P1_U5090 P1_U3671 ; P1_U3086
g13049 nand P1_U5086 P1_U5085 P1_U3670 ; P1_U3087
g13050 nand P1_U5081 P1_U5080 P1_U3669 ; P1_U3088
g13051 nand P1_U5059 P1_U5058 P1_U3667 ; P1_U3089
g13052 nand P1_U5054 P1_U5053 P1_U3666 ; P1_U3090
g13053 nand P1_U5049 P1_U5048 P1_U3665 ; P1_U3091
g13054 nand P1_U5044 P1_U5043 P1_U3664 ; P1_U3092
g13055 nand P1_U5039 P1_U5038 P1_U3663 ; P1_U3093
g13056 nand P1_U5034 P1_U5033 P1_U3662 ; P1_U3094
g13057 nand P1_U5029 P1_U5028 P1_U3661 ; P1_U3095
g13058 nand P1_U5024 P1_U5023 P1_U3660 ; P1_U3096
g13059 nand P1_U5003 P1_U5002 P1_U3658 ; P1_U3097
g13060 nand P1_U4998 P1_U4997 P1_U3657 ; P1_U3098
g13061 nand P1_U4993 P1_U4992 P1_U3656 ; P1_U3099
g13062 nand P1_U4988 P1_U4987 P1_U3655 ; P1_U3100
g13063 nand P1_U4983 P1_U4982 P1_U3654 ; P1_U3101
g13064 nand P1_U4978 P1_U4977 P1_U3653 ; P1_U3102
g13065 nand P1_U4973 P1_U4972 P1_U3652 ; P1_U3103
g13066 nand P1_U4968 P1_U4967 P1_U3651 ; P1_U3104
g13067 nand P1_U4946 P1_U4945 P1_U3649 ; P1_U3105
g13068 nand P1_U4941 P1_U4940 P1_U3648 ; P1_U3106
g13069 nand P1_U4936 P1_U4935 P1_U3647 ; P1_U3107
g13070 nand P1_U4931 P1_U4930 P1_U3646 ; P1_U3108
g13071 nand P1_U4926 P1_U4925 P1_U3645 ; P1_U3109
g13072 nand P1_U4921 P1_U4920 P1_U3644 ; P1_U3110
g13073 nand P1_U4916 P1_U4915 P1_U3643 ; P1_U3111
g13074 nand P1_U4911 P1_U4910 P1_U3642 ; P1_U3112
g13075 nand P1_U4888 P1_U4887 P1_U3640 ; P1_U3113
g13076 nand P1_U4883 P1_U4882 P1_U3639 ; P1_U3114
g13077 nand P1_U4878 P1_U4877 P1_U3638 ; P1_U3115
g13078 nand P1_U4873 P1_U4872 P1_U3637 ; P1_U3116
g13079 nand P1_U4868 P1_U4867 P1_U3636 ; P1_U3117
g13080 nand P1_U4863 P1_U4862 P1_U3635 ; P1_U3118
g13081 nand P1_U4858 P1_U4857 P1_U3634 ; P1_U3119
g13082 nand P1_U4853 P1_U4852 P1_U3633 ; P1_U3120
g13083 nand P1_U4831 P1_U4830 P1_U3631 ; P1_U3121
g13084 nand P1_U4826 P1_U4825 P1_U3630 ; P1_U3122
g13085 nand P1_U4821 P1_U4820 P1_U3629 ; P1_U3123
g13086 nand P1_U4816 P1_U4815 P1_U3628 ; P1_U3124
g13087 nand P1_U4811 P1_U4810 P1_U3627 ; P1_U3125
g13088 nand P1_U4806 P1_U4805 P1_U3626 ; P1_U3126
g13089 nand P1_U4801 P1_U4800 P1_U3625 ; P1_U3127
g13090 nand P1_U4796 P1_U4795 P1_U3624 ; P1_U3128
g13091 nand P1_U4773 P1_U4772 P1_U3622 ; P1_U3129
g13092 nand P1_U4768 P1_U4767 P1_U3621 ; P1_U3130
g13093 nand P1_U4763 P1_U4762 P1_U3620 ; P1_U3131
g13094 nand P1_U4758 P1_U4757 P1_U3619 ; P1_U3132
g13095 nand P1_U4753 P1_U4752 P1_U3618 ; P1_U3133
g13096 nand P1_U4748 P1_U4747 P1_U3617 ; P1_U3134
g13097 nand P1_U4743 P1_U4742 P1_U3616 ; P1_U3135
g13098 nand P1_U4738 P1_U4737 P1_U3615 ; P1_U3136
g13099 nand P1_U4716 P1_U4715 P1_U3613 ; P1_U3137
g13100 nand P1_U4711 P1_U4710 P1_U3612 ; P1_U3138
g13101 nand P1_U4706 P1_U4705 P1_U3611 ; P1_U3139
g13102 nand P1_U4701 P1_U4700 P1_U3610 ; P1_U3140
g13103 nand P1_U4696 P1_U4695 P1_U3609 ; P1_U3141
g13104 nand P1_U4691 P1_U4690 P1_U3608 ; P1_U3142
g13105 nand P1_U4686 P1_U4685 P1_U3607 ; P1_U3143
g13106 nand P1_U4681 P1_U4680 P1_U3606 ; P1_U3144
g13107 nand P1_U4657 P1_U4656 P1_U3604 ; P1_U3145
g13108 nand P1_U4652 P1_U4651 P1_U3603 ; P1_U3146
g13109 nand P1_U4647 P1_U4646 P1_U3602 ; P1_U3147
g13110 nand P1_U4642 P1_U4641 P1_U3601 ; P1_U3148
g13111 nand P1_U4637 P1_U4636 P1_U3600 ; P1_U3149
g13112 nand P1_U4632 P1_U4631 P1_U3599 ; P1_U3150
g13113 nand P1_U4627 P1_U4626 P1_U3598 ; P1_U3151
g13114 nand P1_U4622 P1_U4621 P1_U3597 ; P1_U3152
g13115 nand P1_U4599 P1_U4598 P1_U3595 ; P1_U3153
g13116 nand P1_U4594 P1_U4593 P1_U3594 ; P1_U3154
g13117 nand P1_U4589 P1_U4588 P1_U3593 ; P1_U3155
g13118 nand P1_U4584 P1_U4583 P1_U3592 ; P1_U3156
g13119 nand P1_U4579 P1_U4578 P1_U3591 ; P1_U3157
g13120 nand P1_U4574 P1_U4573 P1_U3590 ; P1_U3158
g13121 nand P1_U4569 P1_U4568 P1_U3589 ; P1_U3159
g13122 nand P1_U4564 P1_U4563 P1_U3588 ; P1_U3160
g13123 nand P1_U7690 P1_U7689 P1_U3586 ; P1_U3161
g13124 nand P1_U4520 P1_U4519 P1_U4518 P1_U4244 ; P1_U3162
g13125 nand P1_U3582 P1_U4516 ; P1_U3163
g13126 and P1_U7650 P1_DATAWIDTH_REG_31__SCAN_IN ; P1_U3164
g13127 and P1_U7650 P1_DATAWIDTH_REG_30__SCAN_IN ; P1_U3165
g13128 and P1_U7650 P1_DATAWIDTH_REG_29__SCAN_IN ; P1_U3166
g13129 and P1_U7650 P1_DATAWIDTH_REG_28__SCAN_IN ; P1_U3167
g13130 and P1_U7650 P1_DATAWIDTH_REG_27__SCAN_IN ; P1_U3168
g13131 and P1_U7650 P1_DATAWIDTH_REG_26__SCAN_IN ; P1_U3169
g13132 and P1_U7650 P1_DATAWIDTH_REG_25__SCAN_IN ; P1_U3170
g13133 and P1_U7650 P1_DATAWIDTH_REG_24__SCAN_IN ; P1_U3171
g13134 and P1_U7650 P1_DATAWIDTH_REG_23__SCAN_IN ; P1_U3172
g13135 and P1_U7650 P1_DATAWIDTH_REG_22__SCAN_IN ; P1_U3173
g13136 and P1_U7650 P1_DATAWIDTH_REG_21__SCAN_IN ; P1_U3174
g13137 and P1_U7650 P1_DATAWIDTH_REG_20__SCAN_IN ; P1_U3175
g13138 and P1_U7650 P1_DATAWIDTH_REG_19__SCAN_IN ; P1_U3176
g13139 and P1_U7650 P1_DATAWIDTH_REG_18__SCAN_IN ; P1_U3177
g13140 and P1_U7650 P1_DATAWIDTH_REG_17__SCAN_IN ; P1_U3178
g13141 and P1_U7650 P1_DATAWIDTH_REG_16__SCAN_IN ; P1_U3179
g13142 and P1_U7650 P1_DATAWIDTH_REG_15__SCAN_IN ; P1_U3180
g13143 and P1_U7650 P1_DATAWIDTH_REG_14__SCAN_IN ; P1_U3181
g13144 and P1_U7650 P1_DATAWIDTH_REG_13__SCAN_IN ; P1_U3182
g13145 and P1_U7650 P1_DATAWIDTH_REG_12__SCAN_IN ; P1_U3183
g13146 and P1_U7650 P1_DATAWIDTH_REG_11__SCAN_IN ; P1_U3184
g13147 and P1_U7650 P1_DATAWIDTH_REG_10__SCAN_IN ; P1_U3185
g13148 and P1_U7650 P1_DATAWIDTH_REG_9__SCAN_IN ; P1_U3186
g13149 and P1_U7650 P1_DATAWIDTH_REG_8__SCAN_IN ; P1_U3187
g13150 and P1_U7650 P1_DATAWIDTH_REG_7__SCAN_IN ; P1_U3188
g13151 and P1_U7650 P1_DATAWIDTH_REG_6__SCAN_IN ; P1_U3189
g13152 and P1_U7650 P1_DATAWIDTH_REG_5__SCAN_IN ; P1_U3190
g13153 and P1_U7650 P1_DATAWIDTH_REG_4__SCAN_IN ; P1_U3191
g13154 and P1_U7650 P1_DATAWIDTH_REG_3__SCAN_IN ; P1_U3192
g13155 and P1_U7650 P1_DATAWIDTH_REG_2__SCAN_IN ; P1_U3193
g13156 nand P1_U7647 P1_U7646 P1_U4375 ; P1_U3194
g13157 nand P1_U7645 P1_U7644 P1_U3495 ; P1_U3195
g13158 nand P1_U3494 P1_U4369 ; P1_U3196
g13159 nand P1_U4355 P1_U4354 P1_U4356 ; P1_U3197
g13160 nand P1_U4352 P1_U4351 P1_U4353 ; P1_U3198
g13161 nand P1_U4349 P1_U4348 P1_U4350 ; P1_U3199
g13162 nand P1_U4346 P1_U4345 P1_U4347 ; P1_U3200
g13163 nand P1_U4343 P1_U4342 P1_U4344 ; P1_U3201
g13164 nand P1_U4340 P1_U4339 P1_U4341 ; P1_U3202
g13165 nand P1_U4337 P1_U4336 P1_U4338 ; P1_U3203
g13166 nand P1_U4334 P1_U4333 P1_U4335 ; P1_U3204
g13167 nand P1_U4331 P1_U4330 P1_U4332 ; P1_U3205
g13168 nand P1_U4328 P1_U4327 P1_U4329 ; P1_U3206
g13169 nand P1_U4325 P1_U4324 P1_U4326 ; P1_U3207
g13170 nand P1_U4322 P1_U4321 P1_U4323 ; P1_U3208
g13171 nand P1_U4319 P1_U4318 P1_U4320 ; P1_U3209
g13172 nand P1_U4316 P1_U4315 P1_U4317 ; P1_U3210
g13173 nand P1_U4313 P1_U4312 P1_U4314 ; P1_U3211
g13174 nand P1_U4310 P1_U4309 P1_U4311 ; P1_U3212
g13175 nand P1_U4307 P1_U4306 P1_U4308 ; P1_U3213
g13176 nand P1_U4304 P1_U4303 P1_U4305 ; P1_U3214
g13177 nand P1_U4301 P1_U4300 P1_U4302 ; P1_U3215
g13178 nand P1_U4298 P1_U4297 P1_U4299 ; P1_U3216
g13179 nand P1_U4295 P1_U4294 P1_U4296 ; P1_U3217
g13180 nand P1_U4292 P1_U4291 P1_U4293 ; P1_U3218
g13181 nand P1_U4289 P1_U4288 P1_U4290 ; P1_U3219
g13182 nand P1_U4286 P1_U4285 P1_U4287 ; P1_U3220
g13183 nand P1_U4283 P1_U4282 P1_U4284 ; P1_U3221
g13184 nand P1_U4280 P1_U4279 P1_U4281 ; P1_U3222
g13185 nand P1_U4277 P1_U4276 P1_U4278 ; P1_U3223
g13186 nand P1_U4274 P1_U4273 P1_U4275 ; P1_U3224
g13187 nand P1_U4271 P1_U4270 P1_U4272 ; P1_U3225
g13188 nand P1_U4268 P1_U4267 P1_U4269 ; P1_U3226
g13189 nand P1_U4001 P1_U4000 P1_U3999 P1_U3998 ; P1_U3227
g13190 nand P1_U3997 P1_U3996 P1_U3995 P1_U3994 ; P1_U3228
g13191 nand P1_U3993 P1_U3992 P1_U3991 P1_U3990 ; P1_U3229
g13192 nand P1_U3989 P1_U3988 P1_U3987 P1_U3986 ; P1_U3230
g13193 nand P1_U3985 P1_U3984 P1_U3983 P1_U3982 ; P1_U3231
g13194 nand P1_U3981 P1_U3980 P1_U3979 P1_U3978 ; P1_U3232
g13195 nand P1_U3977 P1_U3976 P1_U3975 P1_U3974 ; P1_U3233
g13196 nand P1_U3973 P1_U3972 P1_U3971 P1_U3970 ; P1_U3234
g13197 nand P1_U3329 P1_U3323 ; P1_U3235
g13198 nand P1_U2432 P1_U3235 ; P1_U3236
g13199 nand P1_U2432 P1_U4543 ; P1_U3237
g13200 nand P1_U2434 P1_U3235 ; P1_U3238
g13201 nand P1_U2434 P1_U4543 ; P1_U3239
g13202 nand P1_U2433 P1_U3235 ; P1_U3240
g13203 nand P1_U2433 P1_U4543 ; P1_U3241
g13204 nand P1_U2435 P1_U3235 ; P1_U3242
g13205 nand P1_U2435 P1_U4543 ; P1_U3243
g13206 nand P1_U3391 P1_U3394 P1_U5463 ; P1_U3244
g13207 nand P1_U7086 P1_U5464 ; P1_U3245
g13208 nand P1_U7792 P1_U7791 P1_U4158 P1_U4156 ; P1_U3246
g13209 not P1_REQUESTPENDING_REG_SCAN_IN ; P1_U3247
g13210 not P1_STATE_REG_1__SCAN_IN ; P1_U3248
g13211 nand P1_U3258 P1_STATE_REG_1__SCAN_IN ; P1_U3249
g13212 nand P1_U4221 P1_U3251 ; P1_U3250
g13213 not P1_STATE_REG_2__SCAN_IN ; P1_U3251
g13214 nand P1_U4221 P1_STATE_REG_2__SCAN_IN ; P1_U3252
g13215 not P1_REIP_REG_1__SCAN_IN ; P1_U3253
g13216 nand P1_U3251 P1_STATE_REG_1__SCAN_IN ; P1_U3254
g13217 or P1_STATE_REG_2__SCAN_IN P1_STATE_REG_1__SCAN_IN ; P1_U3255
g13218 not HOLD ; P1_U3256
g13219 not U210 ; P1_U3257
g13220 not P1_STATE_REG_0__SCAN_IN ; P1_U3258
g13221 nand P1_U3260 P1_STATE_REG_0__SCAN_IN ; P1_U3259
g13222 nand P1_U3256 P1_REQUESTPENDING_REG_SCAN_IN ; P1_U3260
g13223 or HOLD P1_REQUESTPENDING_REG_SCAN_IN ; P1_U3261
g13224 not P1_STATE2_REG_1__SCAN_IN ; P1_U3262
g13225 not P1_STATE2_REG_2__SCAN_IN ; P1_U3263
g13226 not P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3264
g13227 not P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3265
g13228 not P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3266
g13229 nand P1_U3270 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3267
g13230 or P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3268
g13231 or P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3269
g13232 not P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3270
g13233 nand P1_U3567 P1_U3566 P1_U3565 P1_U3564 ; P1_U3271
g13234 nand P1_U4496 P1_U3258 ; P1_U3272
g13235 not P1_R2167_U17 ; P1_U3273
g13236 nand P1_U3270 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3274
g13237 nand P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3275
g13238 nand P1_U3519 P1_U3518 P1_U3517 P1_U3516 ; P1_U3276
g13239 nand P1_U3539 P1_U4170 P1_U3538 P1_U3537 P1_U3536 ; P1_U3277
g13240 nand P1_U3557 P1_U3556 P1_U3555 P1_U3554 ; P1_U3278
g13241 nand P1_U3559 P1_U3558 ; P1_U3279
g13242 or U210 P1_STATEBS16_REG_SCAN_IN ; P1_U3280
g13243 nand P1_R2167_U17 P1_U4497 ; P1_U3281
g13244 nand P1_U4477 P1_U3284 ; P1_U3282
g13245 nand P1_U3511 P1_U3510 P1_U3509 P1_U3508 ; P1_U3283
g13246 nand P1_U3563 P1_U3562 P1_U3561 P1_U3560 ; P1_U3284
g13247 nand P1_U2473 P1_U4501 ; P1_U3285
g13248 nand P1_U2389 P1_U3283 ; P1_U3286
g13249 nand P1_U4494 P1_U4477 ; P1_U3287
g13250 nand P1_U4249 P1_U2447 ; P1_U3288
g13251 nand P1_U4460 P1_U3391 P1_U4173 P1_U3278 ; P1_U3289
g13252 nand P1_U3271 P1_U3283 ; P1_U3290
g13253 nand P1_U4190 P1_U3284 ; P1_U3291
g13254 nand P1_U4256 P1_U2431 ; P1_U3292
g13255 nand P1_U4178 P1_U4509 P1_U7626 P1_U4225 P1_LT_563_U6 ; P1_U3293
g13256 not P1_STATE2_REG_0__SCAN_IN ; P1_U3294
g13257 nand P1_U7604 P1_STATE2_REG_0__SCAN_IN ; P1_U3295
g13258 not P1_STATE2_REG_3__SCAN_IN ; P1_U3296
g13259 nand P1_U3262 P1_STATE2_REG_2__SCAN_IN ; P1_U3297
g13260 or P1_STATE2_REG_2__SCAN_IN P1_STATE2_REG_1__SCAN_IN ; P1_U3298
g13261 nand P1_R2167_U17 P1_STATE2_REG_3__SCAN_IN ; P1_U3299
g13262 nand P1_U4547 P1_U3294 ; P1_U3300
g13263 not P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_U3301
g13264 not P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_U3302
g13265 not P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_U3303
g13266 not P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U3304
g13267 nand P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_U3305
g13268 nand P1_U4533 P1_U2478 ; P1_U3306
g13269 or P1_STATE2_REG_3__SCAN_IN P1_STATE2_REG_2__SCAN_IN ; P1_U3307
g13270 not P1_STATEBS16_REG_SCAN_IN ; P1_U3308
g13271 not P1_R2144_U43 ; P1_U3309
g13272 not P1_R2144_U50 ; P1_U3310
g13273 not P1_R2144_U49 ; P1_U3311
g13274 not P1_R2144_U8 ; P1_U3312
g13275 nand P1_R2144_U50 P1_R2144_U43 ; P1_U3313
g13276 nand P1_U3332 P1_U3309 ; P1_U3314
g13277 nand P1_U4527 P1_U2475 ; P1_U3315
g13278 not P1_R2182_U25 ; P1_U3316
g13279 not P1_R2182_U42 ; P1_U3317
g13280 not P1_R2182_U34 ; P1_U3318
g13281 not P1_R2182_U33 ; P1_U3319
g13282 nand P1_U4209 P1_U3308 ; P1_U3320
g13283 nand P1_U3306 P1_U4535 ; P1_U3321
g13284 nand P1_U3306 P1_U4544 ; P1_U3322
g13285 nand P1_U3301 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_U3323
g13286 nand P1_U4542 P1_U2478 ; P1_U3324
g13287 nand P1_R2144_U50 P1_U3309 ; P1_U3325
g13288 nand P1_R2144_U43 P1_U3332 ; P1_U3326
g13289 nand P1_U4600 P1_U2475 ; P1_U3327
g13290 nand P1_U3324 P1_U4603 ; P1_U3328
g13291 nand P1_U3302 P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_U3329
g13292 nand P1_U4541 P1_U2478 ; P1_U3330
g13293 nand P1_R2144_U43 P1_U3310 ; P1_U3331
g13294 nand P1_U3325 P1_U3331 ; P1_U3332
g13295 nand P1_U4526 P1_U3309 ; P1_U3333
g13296 nand P1_U4658 P1_U2475 ; P1_U3334
g13297 nand P1_U3330 P1_U4661 ; P1_U3335
g13298 nand P1_U3330 P1_U4663 ; P1_U3336
g13299 nand P1_U2488 P1_U2478 ; P1_U3337
g13300 nand P1_U2485 P1_U2475 ; P1_U3338
g13301 nand P1_U3337 P1_U4719 ; P1_U3339
g13302 nand P1_U3304 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_U3340
g13303 nand P1_U4538 P1_U4533 ; P1_U3341
g13304 nand P1_R2144_U8 P1_U3311 ; P1_U3342
g13305 nand P1_U2490 P1_U4527 ; P1_U3343
g13306 nand P1_U3341 P1_U4776 ; P1_U3344
g13307 nand P1_U3341 P1_U4778 ; P1_U3345
g13308 nand P1_U4538 P1_U4542 ; P1_U3346
g13309 nand P1_U2490 P1_U4600 ; P1_U3347
g13310 nand P1_U3346 P1_U4834 ; P1_U3348
g13311 nand P1_U4538 P1_U4541 ; P1_U3349
g13312 nand P1_U2490 P1_U4658 ; P1_U3350
g13313 nand P1_U3349 P1_U4891 ; P1_U3351
g13314 nand P1_U3349 P1_U4893 ; P1_U3352
g13315 nand P1_U4538 P1_U2488 ; P1_U3353
g13316 nand P1_U2490 P1_U2485 ; P1_U3354
g13317 nand P1_U3353 P1_U4949 ; P1_U3355
g13318 nand P1_U2479 P1_U4533 ; P1_U3356
g13319 nand P1_U2474 P1_U4528 ; P1_U3357
g13320 nand P1_U3342 P1_U4530 P1_U3357 ; P1_U3358
g13321 nand P1_U2499 P1_U4527 ; P1_U3359
g13322 nand P1_U3340 P1_U4539 P1_U3356 ; P1_U3360
g13323 nand P1_U3356 P1_U5005 ; P1_U3361
g13324 nand P1_U3356 P1_U5007 ; P1_U3362
g13325 nand P1_U4542 P1_U2479 ; P1_U3363
g13326 nand P1_U2499 P1_U4600 ; P1_U3364
g13327 nand P1_U3363 P1_U5062 ; P1_U3365
g13328 nand P1_U4541 P1_U2479 ; P1_U3366
g13329 nand P1_U2499 P1_U4658 ; P1_U3367
g13330 nand P1_U3366 P1_U5119 ; P1_U3368
g13331 nand P1_U3366 P1_U5121 ; P1_U3369
g13332 nand P1_U2488 P1_U2479 ; P1_U3370
g13333 nand P1_U2499 P1_U2485 ; P1_U3371
g13334 nand P1_U3370 P1_U5177 ; P1_U3372
g13335 nand P1_U2510 P1_U4533 ; P1_U3373
g13336 nand P1_U2507 P1_U4527 ; P1_U3374
g13337 nand P1_U3373 P1_U5234 ; P1_U3375
g13338 nand P1_U3373 P1_U5236 ; P1_U3376
g13339 nand P1_U2510 P1_U4542 ; P1_U3377
g13340 nand P1_U2507 P1_U4600 ; P1_U3378
g13341 nand P1_U3377 P1_U5292 ; P1_U3379
g13342 nand P1_U2510 P1_U4541 ; P1_U3380
g13343 nand P1_U2507 P1_U4658 ; P1_U3381
g13344 nand P1_U3380 P1_U5349 ; P1_U3382
g13345 nand P1_U3380 P1_U5351 ; P1_U3383
g13346 nand P1_U2510 P1_U2488 ; P1_U3384
g13347 nand P1_U2507 P1_U2485 ; P1_U3385
g13348 nand P1_U3384 P1_U5407 ; P1_U3386
g13349 not P1_FLUSH_REG_SCAN_IN ; P1_U3387
g13350 not P1_GTE_485_U6 ; P1_U3388
g13351 nand P1_U3284 P1_U3278 ; P1_U3389
g13352 nand P1_U3284 P1_U3271 ; P1_U3390
g13353 nand P1_U3515 P1_U3514 P1_U3513 P1_U3512 ; P1_U3391
g13354 nand P1_U5490 P1_U5489 P1_U7628 ; P1_U3392
g13355 nand P1_U4399 P1_U3284 ; P1_U3393
g13356 nand P1_U2605 P1_U3277 ; P1_U3394
g13357 nand P1_U4399 P1_U7494 P1_U4494 ; P1_U3395
g13358 nand P1_U3741 P1_U4247 ; P1_U3396
g13359 nand P1_U7494 P1_U4477 P1_U2605 P1_U4494 P1_U4399 ; P1_U3397
g13360 nand P1_U2605 P1_U4460 P1_U4171 P1_U4449 P1_U4400 ; P1_U3398
g13361 nand P1_U4199 P1_U4477 P1_U4234 ; P1_U3399
g13362 nand P1_U2449 P1_U2447 ; P1_U3400
g13363 nand P1_U3444 P1_U5510 ; P1_U3401
g13364 nand P1_U3269 P1_U3275 ; P1_U3402
g13365 not P1_LT_589_U6 ; P1_U3403
g13366 nand P1_U4242 P1_U3300 P1_U5536 ; P1_U3404
g13367 nand P1_U3278 P1_U3284 P1_STATE2_REG_0__SCAN_IN ; P1_U3405
g13368 nand P1_U3271 P1_U3273 ; P1_U3406
g13369 nand P1_U3277 P1_U3391 ; P1_U3407
g13370 nand P1_U2427 P1_U3294 ; P1_U3408
g13371 nand P1_U4460 P1_U3391 ; P1_U3409
g13372 nand P1_U4253 P1_U3278 ; P1_U3410
g13373 nand P1_U4190 P1_U2452 ; P1_U3411
g13374 nand P1_U3271 P1_STATE2_REG_2__SCAN_IN ; P1_U3412
g13375 not P1_REIP_REG_0__SCAN_IN ; P1_U3413
g13376 nand P1_U3756 P1_U5562 ; P1_U3414
g13377 nand P1_U4400 P1_U4173 ; P1_U3415
g13378 nand P1_U3863 P1_U4248 ; P1_U3416
g13379 nand P1_U6054 P1_U6053 ; P1_U3417
g13380 nand P1_U4494 P1_STATE2_REG_0__SCAN_IN ; P1_U3418
g13381 nand P1_U4399 P1_U7494 ; P1_U3419
g13382 nand P1_U4206 P1_U4477 ; P1_U3420
g13383 nand P1_U4194 P1_U2431 ; P1_U3421
g13384 nand P1_U4210 P1_STATE2_REG_0__SCAN_IN ; P1_U3422
g13385 nand P1_U4503 P1_U3391 ; P1_U3423
g13386 nand P1_U4235 P1_U6153 ; P1_U3424
g13387 nand P1_U4216 P1_STATE2_REG_0__SCAN_IN ; P1_U3425
g13388 nand P1_U4235 P1_U6264 ; P1_U3426
g13389 nand P1_U4249 P1_U3886 P1_U2452 P1_STATE2_REG_0__SCAN_IN ; P1_U3427
g13390 nand P1_U3866 P1_U2447 ; P1_U3428
g13391 not P1_EBX_REG_31__SCAN_IN ; P1_U3429
g13392 not P1_R2337_U69 ; P1_U3430
g13393 nand P1_U4228 P1_U3887 ; P1_U3431
g13394 nand P1_U4209 P1_U3262 ; P1_U3432
g13395 nand P1_U3962 P1_U3958 P1_U3955 P1_U3952 ; P1_U3433
g13396 nand P1_U4206 P1_U3271 ; P1_U3434
g13397 not P1_CODEFETCH_REG_SCAN_IN ; P1_U3435
g13398 not P1_READREQUEST_REG_SCAN_IN ; P1_U3436
g13399 nand P1_U2447 P1_U4498 ; P1_U3437
g13400 nand P1_U3267 P1_U5482 ; P1_U3438
g13401 nand P1_U4449 P1_STATE2_REG_2__SCAN_IN ; P1_U3439
g13402 nand P1_U3263 P1_STATEBS16_REG_SCAN_IN ; P1_U3440
g13403 not P1_U3234 ; P1_U3441
g13404 nand P1_U5479 P1_U5478 ; P1_U3442
g13405 nand P1_U2450 P1_U3441 ; P1_U3443
g13406 nand P1_U3264 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3444
g13407 nand P1_U3274 P1_U7064 ; P1_U3445
g13408 nand P1_U4197 P1_U4234 ; P1_U3446
g13409 nand P1_U4231 P1_U4400 P1_U4250 ; P1_U3447
g13410 nand P1_U4231 P1_U3278 P1_U4250 ; P1_U3448
g13411 nand P1_U4477 P1_U4496 ; P1_U3449
g13412 nand P1_U4074 P1_U7093 P1_U4075 P1_U4077 ; P1_U3450
g13413 nand P1_U4254 P1_U4266 ; P1_U3451
g13414 nand P1_U4183 P1_U3268 ; P1_U3452
g13415 nand P1_U2605 P1_STATE2_REG_0__SCAN_IN ; P1_U3453
g13416 nand P1_U7692 P1_U7691 ; P1_U3454
g13417 nand P1_U7695 P1_U7694 ; P1_U3455
g13418 nand P1_U7719 P1_U7718 ; P1_U3456
g13419 nand P1_U7789 P1_U7788 ; P1_U3457
g13420 nand P1_U7634 P1_U7633 ; P1_U3458
g13421 nand P1_U7636 P1_U7635 ; P1_U3459
g13422 nand P1_U7638 P1_U7637 ; P1_U3460
g13423 nand P1_U7640 P1_U7639 ; P1_U3461
g13424 nand P1_U7649 P1_U7648 ; P1_U3462
g13425 and P1_U3255 P1_U4179 ; P1_U3463
g13426 nand P1_U7652 P1_U7651 ; P1_U3464
g13427 nand P1_U7654 P1_U7653 ; P1_U3465
g13428 nand P1_U7686 P1_U7685 ; P1_U3466
g13429 and P1_U2427 P1_U4215 P1_R2182_U24 ; P1_U3467
g13430 nand P1_U7702 P1_U7701 ; P1_U3468
g13431 nand P1_U7709 P1_U7708 ; P1_U3469
g13432 nand P1_U7711 P1_U7710 ; P1_U3470
g13433 nand P1_U7714 P1_U7713 ; P1_U3471
g13434 nand P1_U7722 P1_U7721 ; P1_U3472
g13435 nand P1_U7724 P1_U7723 ; P1_U3473
g13436 nand P1_U7728 P1_U7727 ; P1_U3474
g13437 nand P1_U7730 P1_U7729 ; P1_U3475
g13438 nand P1_U7735 P1_U7734 ; P1_U3476
g13439 nand P1_U7737 P1_U7736 ; P1_U3477
g13440 nand P1_U7739 P1_U7738 ; P1_U3478
g13441 and P1_R2358_U22 P1_U4449 ; P1_U3479
g13442 nor P1_DATAWIDTH_REG_1__SCAN_IN P1_REIP_REG_1__SCAN_IN ; P1_U3480
g13443 nand P1_U7755 P1_U7754 ; P1_U3481
g13444 nand P1_U7759 P1_U7758 ; P1_U3482
g13445 nand P1_U7761 P1_U7760 ; P1_U3483
g13446 nand P1_U7763 P1_U7762 ; P1_U3484
g13447 nand P1_U7767 P1_U7766 ; P1_U3485
g13448 nand P1_U7771 P1_U7770 ; P1_U3486
g13449 nand P1_U7773 P1_U7772 ; P1_U3487
g13450 and P1_R2182_U24 P1_U4215 ; P1_U3488
g13451 nand P1_U7775 P1_U7774 ; P1_U3489
g13452 nand P1_U7777 P1_U7776 ; P1_U3490
g13453 nand P1_U7779 P1_U7778 ; P1_U3491
g13454 nand P1_U7781 P1_U7780 ; P1_U3492
g13455 nand P1_U7783 P1_U7782 ; P1_U3493
g13456 and P1_U4368 P1_U3252 ; P1_U3494
g13457 and P1_U4370 P1_U3250 ; P1_U3495
g13458 and P1_STATE_REG_0__SCAN_IN P1_REQUESTPENDING_REG_SCAN_IN ; P1_U3496
g13459 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3497
g13460 and P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3498
g13461 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3499
g13462 and P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3500
g13463 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3501
g13464 and P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3502
g13465 nor P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3503
g13466 and P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3504
g13467 nor P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3505
g13468 and P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3506
g13469 and P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3507
g13470 and P1_U4386 P1_U4385 P1_U4384 P1_U4383 ; P1_U3508
g13471 and P1_U4390 P1_U4389 P1_U4388 P1_U4387 ; P1_U3509
g13472 and P1_U4394 P1_U4393 P1_U4392 P1_U4391 ; P1_U3510
g13473 and P1_U4398 P1_U4397 P1_U4396 P1_U4395 ; P1_U3511
g13474 and P1_U4436 P1_U4435 P1_U4434 P1_U4433 ; P1_U3512
g13475 and P1_U4440 P1_U4439 P1_U4438 P1_U4437 ; P1_U3513
g13476 and P1_U4444 P1_U4443 P1_U4442 P1_U4441 ; P1_U3514
g13477 and P1_U4448 P1_U4447 P1_U4446 P1_U4445 ; P1_U3515
g13478 and P1_U4419 P1_U4418 P1_U4417 P1_U4416 ; P1_U3516
g13479 and P1_U4423 P1_U4422 P1_U4421 P1_U4420 ; P1_U3517
g13480 and P1_U4427 P1_U4426 P1_U4425 P1_U4424 ; P1_U3518
g13481 and P1_U4431 P1_U4430 P1_U4429 P1_U4428 ; P1_U3519
g13482 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3520
g13483 and P1_INSTQUEUE_REG_5__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3521
g13484 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3522
g13485 and P1_INSTQUEUE_REG_6__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3523
g13486 and P1_INSTQUEUE_REG_8__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3524
g13487 nor P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3525
g13488 and P1_INSTQUEUE_REG_10__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3526
g13489 and P1_INSTQUEUE_REG_12__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3527
g13490 nor P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3528
g13491 and P1_INSTQUEUE_REG_9__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3529
g13492 and P1_U4404 P1_U4403 P1_U4402 P1_U4401 ; P1_U3530
g13493 and P1_U4408 P1_U4407 P1_U4406 P1_U4405 ; P1_U3531
g13494 and P1_U4412 P1_U4411 P1_U4410 P1_U4409 ; P1_U3532
g13495 and P1_U4414 P1_U4413 ; P1_U3533
g13496 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3534
g13497 and P1_INSTQUEUE_REG_3__6__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3535
g13498 and P1_U4453 P1_U4452 P1_U4451 P1_U4450 ; P1_U3536
g13499 and P1_U4455 P1_U4454 P1_U4456 ; P1_U3537
g13500 and P1_U4458 P1_U4457 P1_U4459 ; P1_U3538
g13501 and P1_U7678 P1_U7677 P1_U7676 P1_U7675 ; P1_U3539
g13502 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3540
g13503 and P1_INSTQUEUE_REG_1__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3541
g13504 nor P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3542
g13505 and P1_INSTQUEUE_REG_4__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3543
g13506 nor P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3544
g13507 and P1_INSTQUEUE_REG_12__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3545
g13508 and P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3546
g13509 and P1_INSTQUEUE_REG_13__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3547
g13510 nor P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U3548
g13511 and P1_INSTQUEUE_REG_6__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U3549
g13512 and P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3550
g13513 and P1_INSTQUEUE_REG_14__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3551
g13514 nor P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U3552
g13515 and P1_INSTQUEUE_REG_9__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U3553
g13516 and P1_U7658 P1_U7657 P1_U7656 P1_U7655 ; P1_U3554
g13517 and P1_U7662 P1_U7661 P1_U7660 P1_U7659 ; P1_U3555
g13518 and P1_U7666 P1_U7665 P1_U7664 P1_U7663 ; P1_U3556
g13519 and P1_U7670 P1_U7669 P1_U7668 P1_U7667 ; P1_U3557
g13520 and P1_U3391 P1_U3283 P1_U7494 ; P1_U3558
g13521 and P1_U4460 P1_U2605 P1_U4400 ; P1_U3559
g13522 and P1_U4481 P1_U4480 P1_U4479 P1_U4478 ; P1_U3560
g13523 and P1_U4485 P1_U4484 P1_U4483 P1_U4482 ; P1_U3561
g13524 and P1_U4489 P1_U4488 P1_U4487 P1_U4486 ; P1_U3562
g13525 and P1_U4493 P1_U4492 P1_U4491 P1_U4490 ; P1_U3563
g13526 and P1_U4464 P1_U4463 P1_U4462 P1_U4461 ; P1_U3564
g13527 and P1_U4468 P1_U4467 P1_U4466 P1_U4465 ; P1_U3565
g13528 and P1_U4472 P1_U4471 P1_U4470 P1_U4469 ; P1_U3566
g13529 and P1_U4476 P1_U4475 P1_U4474 P1_U4473 ; P1_U3567
g13530 and P1_U4377 P1_U4208 ; P1_U3568
g13531 and P1_U4419 P1_U4418 P1_U4417 P1_U4416 ; P1_U3569
g13532 and P1_U4423 P1_U4422 P1_U4421 P1_U4420 ; P1_U3570
g13533 and P1_U4427 P1_U4426 P1_U4425 P1_U4424 ; P1_U3571
g13534 and P1_U4431 P1_U4430 P1_U4429 P1_U4428 ; P1_U3572
g13535 and P1_U4404 P1_U4403 P1_U4402 P1_U4401 ; P1_U3573
g13536 and P1_U4408 P1_U4407 P1_U4406 P1_U4405 ; P1_U3574
g13537 and P1_U4412 P1_U4411 P1_U4410 P1_U4409 ; P1_U3575
g13538 and P1_U4414 P1_U4413 ; P1_U3576
g13539 and P1_U4399 P1_U4171 ; P1_U3577
g13540 and P1_U4249 P1_U3283 ; P1_U3578
g13541 and P1_U3284 P1_U3283 P1_U4400 P1_U7494 ; P1_U3579
g13542 and P1_U4217 P1_U3400 ; P1_U3580
g13543 and P1_U7603 P1_STATE2_REG_2__SCAN_IN ; P1_U3581
g13544 and P1_U4515 P1_U3297 ; P1_U3582
g13545 and P1_U2427 P1_U3257 ; P1_U3583
g13546 and P1_STATE2_REG_3__SCAN_IN P1_STATE2_REG_0__SCAN_IN ; P1_U3584
g13547 and P1_U4246 P1_U4241 ; P1_U3585
g13548 and P1_U3585 P1_U4523 ; P1_U3586
g13549 and P1_U4552 P1_U4553 P1_U4224 ; P1_U3587
g13550 and P1_U4561 P1_U4560 P1_U4562 ; P1_U3588
g13551 and P1_U4566 P1_U4565 P1_U4567 ; P1_U3589
g13552 and P1_U4571 P1_U4570 P1_U4572 ; P1_U3590
g13553 and P1_U4576 P1_U4575 P1_U4577 ; P1_U3591
g13554 and P1_U4581 P1_U4580 P1_U4582 ; P1_U3592
g13555 and P1_U4586 P1_U4585 P1_U4587 ; P1_U3593
g13556 and P1_U4591 P1_U4590 P1_U4592 ; P1_U3594
g13557 and P1_U4596 P1_U4595 P1_U4597 ; P1_U3595
g13558 and P1_U4610 P1_U4611 P1_U4224 ; P1_U3596
g13559 and P1_U4619 P1_U4618 P1_U4620 ; P1_U3597
g13560 and P1_U4624 P1_U4623 P1_U4625 ; P1_U3598
g13561 and P1_U4629 P1_U4628 P1_U4630 ; P1_U3599
g13562 and P1_U4634 P1_U4633 P1_U4635 ; P1_U3600
g13563 and P1_U4639 P1_U4638 P1_U4640 ; P1_U3601
g13564 and P1_U4644 P1_U4643 P1_U4645 ; P1_U3602
g13565 and P1_U4649 P1_U4648 P1_U4650 ; P1_U3603
g13566 and P1_U4654 P1_U4653 P1_U4655 ; P1_U3604
g13567 and P1_U4669 P1_U4670 P1_U4224 ; P1_U3605
g13568 and P1_U4678 P1_U4677 P1_U4679 ; P1_U3606
g13569 and P1_U4683 P1_U4682 P1_U4684 ; P1_U3607
g13570 and P1_U4688 P1_U4687 P1_U4689 ; P1_U3608
g13571 and P1_U4693 P1_U4692 P1_U4694 ; P1_U3609
g13572 and P1_U4698 P1_U4697 P1_U4699 ; P1_U3610
g13573 and P1_U4703 P1_U4702 P1_U4704 ; P1_U3611
g13574 and P1_U4708 P1_U4707 P1_U4709 ; P1_U3612
g13575 and P1_U4713 P1_U4712 P1_U4714 ; P1_U3613
g13576 and P1_U4726 P1_U4727 P1_U4224 ; P1_U3614
g13577 and P1_U4735 P1_U4734 P1_U4736 ; P1_U3615
g13578 and P1_U4740 P1_U4739 P1_U4741 ; P1_U3616
g13579 and P1_U4745 P1_U4744 P1_U4746 ; P1_U3617
g13580 and P1_U4750 P1_U4749 P1_U4751 ; P1_U3618
g13581 and P1_U4755 P1_U4754 P1_U4756 ; P1_U3619
g13582 and P1_U4760 P1_U4759 P1_U4761 ; P1_U3620
g13583 and P1_U4765 P1_U4764 P1_U4766 ; P1_U3621
g13584 and P1_U4770 P1_U4769 P1_U4771 ; P1_U3622
g13585 and P1_U4784 P1_U4785 P1_U4224 ; P1_U3623
g13586 and P1_U4793 P1_U4792 P1_U4794 ; P1_U3624
g13587 and P1_U4798 P1_U4797 P1_U4799 ; P1_U3625
g13588 and P1_U4803 P1_U4802 P1_U4804 ; P1_U3626
g13589 and P1_U4808 P1_U4807 P1_U4809 ; P1_U3627
g13590 and P1_U4813 P1_U4812 P1_U4814 ; P1_U3628
g13591 and P1_U4818 P1_U4817 P1_U4819 ; P1_U3629
g13592 and P1_U4823 P1_U4822 P1_U4824 ; P1_U3630
g13593 and P1_U4828 P1_U4827 P1_U4829 ; P1_U3631
g13594 and P1_U4841 P1_U4842 P1_U4224 ; P1_U3632
g13595 and P1_U4850 P1_U4849 P1_U4851 ; P1_U3633
g13596 and P1_U4855 P1_U4854 P1_U4856 ; P1_U3634
g13597 and P1_U4860 P1_U4859 P1_U4861 ; P1_U3635
g13598 and P1_U4865 P1_U4864 P1_U4866 ; P1_U3636
g13599 and P1_U4870 P1_U4869 P1_U4871 ; P1_U3637
g13600 and P1_U4875 P1_U4874 P1_U4876 ; P1_U3638
g13601 and P1_U4880 P1_U4879 P1_U4881 ; P1_U3639
g13602 and P1_U4885 P1_U4884 P1_U4886 ; P1_U3640
g13603 and P1_U4899 P1_U4900 P1_U4224 ; P1_U3641
g13604 and P1_U4908 P1_U4907 P1_U4909 ; P1_U3642
g13605 and P1_U4913 P1_U4912 P1_U4914 ; P1_U3643
g13606 and P1_U4918 P1_U4917 P1_U4919 ; P1_U3644
g13607 and P1_U4923 P1_U4922 P1_U4924 ; P1_U3645
g13608 and P1_U4928 P1_U4927 P1_U4929 ; P1_U3646
g13609 and P1_U4933 P1_U4932 P1_U4934 ; P1_U3647
g13610 and P1_U4938 P1_U4937 P1_U4939 ; P1_U3648
g13611 and P1_U4943 P1_U4942 P1_U4944 ; P1_U3649
g13612 and P1_U4956 P1_U4957 P1_U4224 ; P1_U3650
g13613 and P1_U4965 P1_U4964 P1_U4966 ; P1_U3651
g13614 and P1_U4970 P1_U4969 P1_U4971 ; P1_U3652
g13615 and P1_U4975 P1_U4974 P1_U4976 ; P1_U3653
g13616 and P1_U4980 P1_U4979 P1_U4981 ; P1_U3654
g13617 and P1_U4985 P1_U4984 P1_U4986 ; P1_U3655
g13618 and P1_U4990 P1_U4989 P1_U4991 ; P1_U3656
g13619 and P1_U4995 P1_U4994 P1_U4996 ; P1_U3657
g13620 and P1_U5000 P1_U4999 P1_U5001 ; P1_U3658
g13621 and P1_U5012 P1_U5013 P1_U4224 ; P1_U3659
g13622 and P1_U5021 P1_U5020 P1_U5022 ; P1_U3660
g13623 and P1_U5026 P1_U5025 P1_U5027 ; P1_U3661
g13624 and P1_U5031 P1_U5030 P1_U5032 ; P1_U3662
g13625 and P1_U5036 P1_U5035 P1_U5037 ; P1_U3663
g13626 and P1_U5041 P1_U5040 P1_U5042 ; P1_U3664
g13627 and P1_U5046 P1_U5045 P1_U5047 ; P1_U3665
g13628 and P1_U5051 P1_U5050 P1_U5052 ; P1_U3666
g13629 and P1_U5056 P1_U5055 P1_U5057 ; P1_U3667
g13630 and P1_U5069 P1_U5070 P1_U4224 ; P1_U3668
g13631 and P1_U5078 P1_U5077 P1_U5079 ; P1_U3669
g13632 and P1_U5083 P1_U5082 P1_U5084 ; P1_U3670
g13633 and P1_U5088 P1_U5087 P1_U5089 ; P1_U3671
g13634 and P1_U5093 P1_U5092 P1_U5094 ; P1_U3672
g13635 and P1_U5098 P1_U5097 P1_U5099 ; P1_U3673
g13636 and P1_U5103 P1_U5102 P1_U5104 ; P1_U3674
g13637 and P1_U5108 P1_U5107 P1_U5109 ; P1_U3675
g13638 and P1_U5113 P1_U5112 P1_U5114 ; P1_U3676
g13639 and P1_U5127 P1_U5128 P1_U4224 ; P1_U3677
g13640 and P1_U5136 P1_U5135 P1_U5137 ; P1_U3678
g13641 and P1_U5141 P1_U5140 P1_U5142 ; P1_U3679
g13642 and P1_U5146 P1_U5145 P1_U5147 ; P1_U3680
g13643 and P1_U5151 P1_U5150 P1_U5152 ; P1_U3681
g13644 and P1_U5156 P1_U5155 P1_U5157 ; P1_U3682
g13645 and P1_U5161 P1_U5160 P1_U5162 ; P1_U3683
g13646 and P1_U5166 P1_U5165 P1_U5167 ; P1_U3684
g13647 and P1_U5171 P1_U5170 P1_U5172 ; P1_U3685
g13648 and P1_U5184 P1_U5185 P1_U4224 ; P1_U3686
g13649 and P1_U5193 P1_U5192 P1_U5194 ; P1_U3687
g13650 and P1_U5198 P1_U5197 P1_U5199 ; P1_U3688
g13651 and P1_U5203 P1_U5202 P1_U5204 ; P1_U3689
g13652 and P1_U5208 P1_U5207 P1_U5209 ; P1_U3690
g13653 and P1_U5213 P1_U5212 P1_U5214 ; P1_U3691
g13654 and P1_U5218 P1_U5217 P1_U5219 ; P1_U3692
g13655 and P1_U5223 P1_U5222 P1_U5224 ; P1_U3693
g13656 and P1_U5228 P1_U5227 P1_U5229 ; P1_U3694
g13657 and P1_U5242 P1_U5243 P1_U4224 ; P1_U3695
g13658 and P1_U5251 P1_U5250 P1_U5252 ; P1_U3696
g13659 and P1_U5256 P1_U5255 P1_U5257 ; P1_U3697
g13660 and P1_U5261 P1_U5260 P1_U5262 ; P1_U3698
g13661 and P1_U5266 P1_U5265 P1_U5267 ; P1_U3699
g13662 and P1_U5271 P1_U5270 P1_U5272 ; P1_U3700
g13663 and P1_U5276 P1_U5275 P1_U5277 ; P1_U3701
g13664 and P1_U5281 P1_U5280 P1_U5282 ; P1_U3702
g13665 and P1_U5286 P1_U5285 P1_U5287 ; P1_U3703
g13666 and P1_U5299 P1_U5300 P1_U4224 ; P1_U3704
g13667 and P1_U5308 P1_U5307 P1_U5309 ; P1_U3705
g13668 and P1_U5313 P1_U5312 P1_U5314 ; P1_U3706
g13669 and P1_U5318 P1_U5317 P1_U5319 ; P1_U3707
g13670 and P1_U5323 P1_U5322 P1_U5324 ; P1_U3708
g13671 and P1_U5328 P1_U5327 P1_U5329 ; P1_U3709
g13672 and P1_U5333 P1_U5332 P1_U5334 ; P1_U3710
g13673 and P1_U5338 P1_U5337 P1_U5339 ; P1_U3711
g13674 and P1_U5343 P1_U5342 P1_U5344 ; P1_U3712
g13675 and P1_U5357 P1_U5358 P1_U4224 ; P1_U3713
g13676 and P1_U5366 P1_U5365 P1_U5367 ; P1_U3714
g13677 and P1_U5371 P1_U5370 P1_U5372 ; P1_U3715
g13678 and P1_U5376 P1_U5375 P1_U5377 ; P1_U3716
g13679 and P1_U5381 P1_U5380 P1_U5382 ; P1_U3717
g13680 and P1_U5386 P1_U5385 P1_U5387 ; P1_U3718
g13681 and P1_U5391 P1_U5390 P1_U5392 ; P1_U3719
g13682 and P1_U5396 P1_U5395 P1_U5397 ; P1_U3720
g13683 and P1_U5401 P1_U5400 P1_U5402 ; P1_U3721
g13684 and P1_U5414 P1_U5415 P1_U4224 ; P1_U3722
g13685 and P1_U5423 P1_U5422 P1_U5424 ; P1_U3723
g13686 and P1_U5428 P1_U5427 P1_U5429 ; P1_U3724
g13687 and P1_U5433 P1_U5432 P1_U5434 ; P1_U3725
g13688 and P1_U5438 P1_U5437 P1_U5439 ; P1_U3726
g13689 and P1_U5442 P1_U5441 P1_U5443 ; P1_U3727
g13690 and P1_U5447 P1_U5446 P1_U5448 ; P1_U3728
g13691 and P1_U5452 P1_U5451 P1_U5453 ; P1_U3729
g13692 and P1_U5457 P1_U5456 P1_U5458 ; P1_U3730
g13693 and P1_STATE2_REG_0__SCAN_IN P1_FLUSH_REG_SCAN_IN ; P1_U3731
g13694 and P1_U4494 P1_U4399 ; P1_U3732
g13695 and P1_U4497 P1_U3257 ; P1_U3733
g13696 and P1_U4210 P1_U3257 ; P1_U3734
g13697 and P1_U7496 P1_U4217 ; P1_U3735
g13698 and P1_U5471 P1_U5472 ; P1_U3736
g13699 and P1_U3736 P1_U5470 ; P1_U3737
g13700 and P1_U3737 P1_U2518 ; P1_U3738
g13701 and P1_U5475 P1_U4242 ; P1_U3739
g13702 and P1_U5486 P1_U5485 ; P1_U3740
g13703 and P1_U4449 P1_U4400 ; P1_U3741
g13704 and P1_U5496 P1_U3393 ; P1_U3742
g13705 and P1_U5498 P1_U5497 ; P1_U3743
g13706 and P1_U5500 P1_U7627 P1_U3742 P1_U3743 ; P1_U3744
g13707 and P1_U4263 P1_U3397 ; P1_U3745
g13708 and P1_U3411 P1_U3288 P1_U3745 P1_U2520 P1_U3279 ; P1_U3746
g13709 and P1_U3748 P1_U5502 ; P1_U3747
g13710 and P1_U5505 P1_U5504 ; P1_U3748
g13711 and P1_U7717 P1_U7716 P1_U5513 ; P1_U3749
g13712 and P1_U5524 P1_U5522 ; P1_U3750
g13713 and P1_U5543 P1_U5544 ; P1_U3751
g13714 and P1_U5547 P1_U5548 ; P1_U3752
g13715 and P1_U5552 P1_U5553 ; P1_U3753
g13716 and P1_U5558 P1_U3257 ; P1_U3754
g13717 and P1_U3284 P1_U3407 ; P1_U3755
g13718 and P1_U5563 P1_U5561 ; P1_U3756
g13719 and P1_U3398 P1_U3399 P1_U5567 ; P1_U3757
g13720 and P1_U2520 P1_U5568 P1_U3757 ; P1_U3758
g13721 and P1_U4186 P1_U3284 ; P1_U3759
g13722 and P1_U3288 P1_U4217 P1_U3448 ; P1_U3760
g13723 and P1_U5566 P1_U7507 ; P1_U3761
g13724 and P1_U7508 P1_STATE2_REG_2__SCAN_IN ; P1_U3762
g13725 and P1_U5571 P1_U5570 ; P1_U3763
g13726 and P1_U5573 P1_U5572 ; P1_U3764
g13727 and P1_U5575 P1_U5576 ; P1_U3765
g13728 and P1_U3765 P1_U5574 ; P1_U3766
g13729 and P1_U5578 P1_U5577 ; P1_U3767
g13730 and P1_U5580 P1_U5579 ; P1_U3768
g13731 and P1_U5582 P1_U5583 ; P1_U3769
g13732 and P1_U3769 P1_U5581 ; P1_U3770
g13733 and P1_U5585 P1_U5584 ; P1_U3771
g13734 and P1_U5587 P1_U5586 ; P1_U3772
g13735 and P1_U5589 P1_U5590 ; P1_U3773
g13736 and P1_U3773 P1_U5588 ; P1_U3774
g13737 and P1_U5592 P1_U5591 P1_U5594 ; P1_U3775
g13738 and P1_U3777 P1_U5595 P1_U5593 ; P1_U3776
g13739 and P1_U5596 P1_U5597 ; P1_U3777
g13740 and P1_U5599 P1_U5598 P1_U5601 ; P1_U3778
g13741 and P1_U5603 P1_U5604 ; P1_U3779
g13742 and P1_U3779 P1_U5602 ; P1_U3780
g13743 and P1_U5606 P1_U5605 P1_U5608 ; P1_U3781
g13744 and P1_U5610 P1_U5611 ; P1_U3782
g13745 and P1_U3782 P1_U5609 ; P1_U3783
g13746 and P1_U5613 P1_U5612 P1_U5615 ; P1_U3784
g13747 and P1_U5617 P1_U5618 ; P1_U3785
g13748 and P1_U3785 P1_U5616 ; P1_U3786
g13749 and P1_U5620 P1_U5619 P1_U5622 ; P1_U3787
g13750 and P1_U5624 P1_U5625 ; P1_U3788
g13751 and P1_U3788 P1_U5623 ; P1_U3789
g13752 and P1_U5627 P1_U5626 P1_U5629 ; P1_U3790
g13753 and P1_U5631 P1_U5632 ; P1_U3791
g13754 and P1_U3791 P1_U5630 ; P1_U3792
g13755 and P1_U5634 P1_U5633 P1_U5636 ; P1_U3793
g13756 and P1_U5638 P1_U5639 ; P1_U3794
g13757 and P1_U3794 P1_U5637 ; P1_U3795
g13758 and P1_U5641 P1_U5640 P1_U5643 ; P1_U3796
g13759 and P1_U5645 P1_U5646 ; P1_U3797
g13760 and P1_U3797 P1_U5644 ; P1_U3798
g13761 and P1_U5648 P1_U5647 P1_U5650 ; P1_U3799
g13762 and P1_U5652 P1_U5653 ; P1_U3800
g13763 and P1_U3800 P1_U5651 ; P1_U3801
g13764 and P1_U5655 P1_U5654 P1_U5657 ; P1_U3802
g13765 and P1_U5659 P1_U5660 ; P1_U3803
g13766 and P1_U3803 P1_U5658 ; P1_U3804
g13767 and P1_U5662 P1_U5664 ; P1_U3805
g13768 and P1_U5666 P1_U5667 ; P1_U3806
g13769 and P1_U3806 P1_U5665 ; P1_U3807
g13770 and P1_U5669 P1_U5671 ; P1_U3808
g13771 and P1_U5673 P1_U5674 ; P1_U3809
g13772 and P1_U3809 P1_U5672 ; P1_U3810
g13773 and P1_U5676 P1_U5678 ; P1_U3811
g13774 and P1_U5680 P1_U5681 ; P1_U3812
g13775 and P1_U3812 P1_U5679 ; P1_U3813
g13776 and P1_U5683 P1_U5685 ; P1_U3814
g13777 and P1_U5687 P1_U5688 ; P1_U3815
g13778 and P1_U3815 P1_U5686 ; P1_U3816
g13779 and P1_U5690 P1_U5692 ; P1_U3817
g13780 and P1_U5694 P1_U5695 ; P1_U3818
g13781 and P1_U3818 P1_U5693 ; P1_U3819
g13782 and P1_U5697 P1_U5699 ; P1_U3820
g13783 and P1_U5701 P1_U5702 ; P1_U3821
g13784 and P1_U3821 P1_U5700 ; P1_U3822
g13785 and P1_U5704 P1_U5706 ; P1_U3823
g13786 and P1_U5708 P1_U5709 ; P1_U3824
g13787 and P1_U3824 P1_U5707 ; P1_U3825
g13788 and P1_U5711 P1_U5713 ; P1_U3826
g13789 and P1_U5715 P1_U5716 ; P1_U3827
g13790 and P1_U3827 P1_U5714 ; P1_U3828
g13791 and P1_U5718 P1_U5720 ; P1_U3829
g13792 and P1_U5722 P1_U5723 ; P1_U3830
g13793 and P1_U3830 P1_U5721 ; P1_U3831
g13794 and P1_U5725 P1_U5727 ; P1_U3832
g13795 and P1_U5729 P1_U5730 ; P1_U3833
g13796 and P1_U3833 P1_U5728 ; P1_U3834
g13797 and P1_U5732 P1_U5734 ; P1_U3835
g13798 and P1_U5736 P1_U5737 ; P1_U3836
g13799 and P1_U3836 P1_U5735 ; P1_U3837
g13800 and P1_U5739 P1_U5741 ; P1_U3838
g13801 and P1_U5743 P1_U5744 ; P1_U3839
g13802 and P1_U3839 P1_U5742 ; P1_U3840
g13803 and P1_U5746 P1_U5748 ; P1_U3841
g13804 and P1_U5750 P1_U5751 ; P1_U3842
g13805 and P1_U3842 P1_U5749 ; P1_U3843
g13806 and P1_U5753 P1_U5755 ; P1_U3844
g13807 and P1_U5757 P1_U5758 ; P1_U3845
g13808 and P1_U3845 P1_U5756 ; P1_U3846
g13809 and P1_U5760 P1_U5762 ; P1_U3847
g13810 and P1_U5764 P1_U5765 ; P1_U3848
g13811 and P1_U3848 P1_U5763 ; P1_U3849
g13812 and P1_U5767 P1_U5769 ; P1_U3850
g13813 and P1_U5771 P1_U5772 ; P1_U3851
g13814 and P1_U3851 P1_U5770 ; P1_U3852
g13815 and P1_U5774 P1_U5776 ; P1_U3853
g13816 and P1_U5778 P1_U5779 ; P1_U3854
g13817 and P1_U3854 P1_U5777 ; P1_U3855
g13818 and P1_U5781 P1_U5783 ; P1_U3856
g13819 and P1_U5785 P1_U5786 ; P1_U3857
g13820 and P1_U3857 P1_U5784 ; P1_U3858
g13821 and P1_U5788 P1_U5790 ; P1_U3859
g13822 and P1_U5792 P1_U5793 ; P1_U3860
g13823 and P1_U3860 P1_U5791 ; P1_U3861
g13824 and P1_U3283 P1_U3262 P1_U7494 ; P1_U3862
g13825 and P1_U5794 P1_U3408 ; P1_U3863
g13826 and P1_STATE2_REG_1__SCAN_IN P1_STATEBS16_REG_SCAN_IN ; P1_U3864
g13827 and P1_U2368 P1_U3284 ; P1_U3865
g13828 and P1_U2449 P1_STATE2_REG_0__SCAN_IN ; P1_U3866
g13829 and P1_U4208 P1_U2368 ; P1_U3867
g13830 and P1_U6105 P1_U6106 ; P1_U3868
g13831 and P1_U6108 P1_U6109 ; P1_U3869
g13832 and P1_U6111 P1_U6112 ; P1_U3870
g13833 and P1_U6114 P1_U6115 ; P1_U3871
g13834 and P1_U6117 P1_U6118 ; P1_U3872
g13835 and P1_U6120 P1_U6121 ; P1_U3873
g13836 and P1_U6123 P1_U6124 ; P1_U3874
g13837 and P1_U6126 P1_U6127 ; P1_U3875
g13838 and P1_U6129 P1_U6130 ; P1_U3876
g13839 and P1_U6132 P1_U6133 ; P1_U3877
g13840 and P1_U6135 P1_U6136 ; P1_U3878
g13841 and P1_U6138 P1_U6139 ; P1_U3879
g13842 and P1_U6141 P1_U6142 ; P1_U3880
g13843 and P1_U6144 P1_U6145 ; P1_U3881
g13844 and P1_U6147 P1_U6148 ; P1_U3882
g13845 and P1_U6151 P1_U6150 ; P1_U3883
g13846 and P1_U2605 P1_U3391 ; P1_U3884
g13847 and P1_U3271 P1_U7494 P1_STATE2_REG_0__SCAN_IN ; P1_U3885
g13848 and P1_U4399 P1_U4171 ; P1_U3886
g13849 and P1_U4241 P1_U4244 P1_U6362 ; P1_U3887
g13850 nor U210 P1_STATEBS16_REG_SCAN_IN ; P1_U3888
g13851 and P1_U4494 P1_U4186 ; P1_U3889
g13852 and P1_U6373 P1_U6372 P1_U6375 P1_U6374 P1_U6371 ; P1_U3890
g13853 and P1_U6381 P1_U6380 P1_U6383 P1_U6382 P1_U6379 ; P1_U3891
g13854 and P1_U6389 P1_U6388 P1_U6391 P1_U6390 P1_U6387 ; P1_U3892
g13855 and P1_U6397 P1_U6396 P1_U6399 P1_U6398 P1_U6395 ; P1_U3893
g13856 and P1_U6400 P1_U4227 ; P1_U3894
g13857 and P1_U6405 P1_U6404 P1_U6407 P1_U6406 ; P1_U3895
g13858 and P1_U6408 P1_U4227 ; P1_U3896
g13859 and P1_U6413 P1_U6412 P1_U6415 P1_U6414 P1_U6411 ; P1_U3897
g13860 and P1_U6416 P1_U4227 ; P1_U3898
g13861 and P1_U6422 P1_U6419 P1_U6421 ; P1_U3899
g13862 and P1_U6423 P1_U4227 ; P1_U3900
g13863 and P1_U6429 P1_U6426 P1_U6428 ; P1_U3901
g13864 and P1_U6430 P1_U4227 ; P1_U3902
g13865 and P1_U6436 P1_U6433 P1_U6435 ; P1_U3903
g13866 and P1_U6437 P1_U4227 ; P1_U3904
g13867 and P1_U6443 P1_U6440 P1_U6442 ; P1_U3905
g13868 and P1_U6444 P1_U4227 ; P1_U3906
g13869 and P1_U6450 P1_U6447 P1_U6449 ; P1_U3907
g13870 and P1_U6451 P1_U4227 ; P1_U3908
g13871 and P1_U6457 P1_U6454 P1_U6456 ; P1_U3909
g13872 and P1_U6458 P1_U4227 ; P1_U3910
g13873 and P1_U6464 P1_U6461 P1_U6463 ; P1_U3911
g13874 and P1_U6465 P1_U4227 ; P1_U3912
g13875 and P1_U6471 P1_U6468 P1_U6470 ; P1_U3913
g13876 and P1_U6472 P1_U4227 ; P1_U3914
g13877 and P1_U6478 P1_U6475 P1_U6477 ; P1_U3915
g13878 and P1_U6479 P1_U4227 ; P1_U3916
g13879 and P1_U6485 P1_U6482 P1_U6484 ; P1_U3917
g13880 and P1_U6486 P1_U4227 ; P1_U3918
g13881 and P1_U6492 P1_U6489 P1_U6491 ; P1_U3919
g13882 and P1_U4227 P1_U6494 ; P1_U3920
g13883 and P1_U6499 P1_U6496 P1_U6498 ; P1_U3921
g13884 and P1_U4227 P1_U6501 ; P1_U3922
g13885 and P1_U6506 P1_U6503 P1_U6505 ; P1_U3923
g13886 and P1_U4227 P1_U6508 ; P1_U3924
g13887 and P1_U6513 P1_U6510 P1_U6512 ; P1_U3925
g13888 and P1_U6517 P1_U6515 ; P1_U3926
g13889 and P1_U6519 P1_U6520 ; P1_U3927
g13890 and P1_U6524 P1_U6522 ; P1_U3928
g13891 and P1_U6526 P1_U6527 ; P1_U3929
g13892 and P1_U6531 P1_U6529 ; P1_U3930
g13893 and P1_U6533 P1_U6534 ; P1_U3931
g13894 and P1_U6538 P1_U6536 ; P1_U3932
g13895 and P1_U6540 P1_U6541 ; P1_U3933
g13896 and P1_U6545 P1_U6543 ; P1_U3934
g13897 and P1_U6547 P1_U6548 ; P1_U3935
g13898 and P1_U6552 P1_U6550 ; P1_U3936
g13899 and P1_U6554 P1_U6555 ; P1_U3937
g13900 and P1_U6559 P1_U6557 ; P1_U3938
g13901 and P1_U6561 P1_U6562 ; P1_U3939
g13902 and P1_U6566 P1_U6564 ; P1_U3940
g13903 and P1_U6568 P1_U6569 ; P1_U3941
g13904 and P1_U6573 P1_U6571 ; P1_U3942
g13905 and P1_U6575 P1_U6576 ; P1_U3943
g13906 and P1_U6580 P1_U6578 ; P1_U3944
g13907 and P1_U6582 P1_U6583 ; P1_U3945
g13908 and P1_U6587 P1_U6585 ; P1_U3946
g13909 and P1_U6589 P1_U6590 ; P1_U3947
g13910 and P1_U6594 P1_U6592 ; P1_U3948
g13911 and P1_U6596 P1_U6597 ; P1_U3949
g13912 nor P1_DATAWIDTH_REG_2__SCAN_IN P1_DATAWIDTH_REG_3__SCAN_IN P1_DATAWIDTH_REG_4__SCAN_IN P1_DATAWIDTH_REG_5__SCAN_IN ; P1_U3950
g13913 nor P1_DATAWIDTH_REG_6__SCAN_IN P1_DATAWIDTH_REG_7__SCAN_IN P1_DATAWIDTH_REG_8__SCAN_IN P1_DATAWIDTH_REG_9__SCAN_IN ; P1_U3951
g13914 and P1_U3951 P1_U3950 ; P1_U3952
g13915 nor P1_DATAWIDTH_REG_10__SCAN_IN P1_DATAWIDTH_REG_11__SCAN_IN P1_DATAWIDTH_REG_12__SCAN_IN P1_DATAWIDTH_REG_13__SCAN_IN ; P1_U3953
g13916 nor P1_DATAWIDTH_REG_14__SCAN_IN P1_DATAWIDTH_REG_15__SCAN_IN P1_DATAWIDTH_REG_16__SCAN_IN P1_DATAWIDTH_REG_17__SCAN_IN ; P1_U3954
g13917 and P1_U3954 P1_U3953 ; P1_U3955
g13918 nor P1_DATAWIDTH_REG_18__SCAN_IN P1_DATAWIDTH_REG_19__SCAN_IN P1_DATAWIDTH_REG_20__SCAN_IN P1_DATAWIDTH_REG_21__SCAN_IN ; P1_U3956
g13919 nor P1_DATAWIDTH_REG_22__SCAN_IN P1_DATAWIDTH_REG_23__SCAN_IN P1_DATAWIDTH_REG_24__SCAN_IN P1_DATAWIDTH_REG_25__SCAN_IN ; P1_U3957
g13920 and P1_U3957 P1_U3956 ; P1_U3958
g13921 nor P1_DATAWIDTH_REG_26__SCAN_IN P1_DATAWIDTH_REG_27__SCAN_IN ; P1_U3959
g13922 nor P1_DATAWIDTH_REG_28__SCAN_IN P1_DATAWIDTH_REG_29__SCAN_IN ; P1_U3960
g13923 nor P1_DATAWIDTH_REG_30__SCAN_IN P1_DATAWIDTH_REG_31__SCAN_IN ; P1_U3961
g13924 and P1_U3961 P1_U6598 P1_U3960 P1_U3959 ; P1_U3962
g13925 nor P1_DATAWIDTH_REG_0__SCAN_IN P1_DATAWIDTH_REG_1__SCAN_IN P1_REIP_REG_0__SCAN_IN ; P1_U3963
g13926 and P1_U3257 P1_STATE2_REG_2__SCAN_IN ; P1_U3964
g13927 and P1_U6608 P1_U3298 ; P1_U3965
g13928 nor U210 P1_STATE2_REG_0__SCAN_IN ; P1_U3966
g13929 and P1_U3307 P1_U3408 P1_U6602 ; P1_U3967
g13930 and P1_U3287 P1_STATE2_REG_2__SCAN_IN ; P1_U3968
g13931 and P1_U4235 P1_U4206 ; P1_U3969
g13932 and P1_U6621 P1_U6620 P1_U6619 P1_U6618 ; P1_U3970
g13933 and P1_U6625 P1_U6624 P1_U6623 P1_U6622 ; P1_U3971
g13934 and P1_U6629 P1_U6628 P1_U6627 P1_U6626 ; P1_U3972
g13935 and P1_U6633 P1_U6632 P1_U6631 P1_U6630 ; P1_U3973
g13936 and P1_U6637 P1_U6636 P1_U6635 P1_U6634 ; P1_U3974
g13937 and P1_U6641 P1_U6640 P1_U6639 P1_U6638 ; P1_U3975
g13938 and P1_U6645 P1_U6644 P1_U6643 P1_U6642 ; P1_U3976
g13939 and P1_U6649 P1_U6648 P1_U6647 P1_U6646 ; P1_U3977
g13940 and P1_U6653 P1_U6652 P1_U6651 P1_U6650 ; P1_U3978
g13941 and P1_U6657 P1_U6656 P1_U6655 P1_U6654 ; P1_U3979
g13942 and P1_U6661 P1_U6660 P1_U6659 P1_U6658 ; P1_U3980
g13943 and P1_U6665 P1_U6664 P1_U6663 P1_U6662 ; P1_U3981
g13944 and P1_U6669 P1_U6668 P1_U6667 P1_U6666 ; P1_U3982
g13945 and P1_U6673 P1_U6672 P1_U6671 P1_U6670 ; P1_U3983
g13946 and P1_U6677 P1_U6676 P1_U6675 P1_U6674 ; P1_U3984
g13947 and P1_U7613 P1_U6680 P1_U6679 P1_U6678 ; P1_U3985
g13948 and P1_U6684 P1_U6683 P1_U6682 P1_U6681 ; P1_U3986
g13949 and P1_U6688 P1_U6687 P1_U6686 P1_U6685 ; P1_U3987
g13950 and P1_U6692 P1_U6691 P1_U6690 P1_U6689 ; P1_U3988
g13951 and P1_U6696 P1_U6695 P1_U6694 P1_U6693 ; P1_U3989
g13952 and P1_U6700 P1_U6699 P1_U6698 P1_U6697 ; P1_U3990
g13953 and P1_U6704 P1_U6703 P1_U6702 P1_U6701 ; P1_U3991
g13954 and P1_U6708 P1_U6707 P1_U6706 P1_U6705 ; P1_U3992
g13955 and P1_U6712 P1_U6711 P1_U6710 P1_U6709 ; P1_U3993
g13956 and P1_U6716 P1_U6715 P1_U6714 P1_U6713 ; P1_U3994
g13957 and P1_U6720 P1_U6719 P1_U6718 P1_U6717 ; P1_U3995
g13958 and P1_U6724 P1_U6723 P1_U6722 P1_U6721 ; P1_U3996
g13959 and P1_U6728 P1_U6727 P1_U6726 P1_U6725 ; P1_U3997
g13960 and P1_U6732 P1_U6731 P1_U6730 P1_U6729 ; P1_U3998
g13961 and P1_U6736 P1_U6735 P1_U6734 P1_U6733 ; P1_U3999
g13962 and P1_U6740 P1_U6739 P1_U6738 P1_U6737 ; P1_U4000
g13963 and P1_U6744 P1_U6743 P1_U6742 P1_U6741 ; P1_U4001
g13964 and P1_U6749 P1_U6748 ; P1_U4002
g13965 and P1_U6752 P1_U6751 ; P1_U4003
g13966 and P1_U6755 P1_U6754 ; P1_U4004
g13967 and P1_U6758 P1_U6757 ; P1_U4005
g13968 and P1_U6760 P1_U4007 ; P1_U4006
g13969 and P1_U6762 P1_U6761 ; P1_U4007
g13970 and P1_U6764 P1_U6765 ; P1_U4008
g13971 and P1_U6772 P1_U6773 P1_U6774 ; P1_U4009
g13972 and P1_U6776 P1_U6777 ; P1_U4010
g13973 and P1_U6781 P1_U6782 P1_U6783 ; P1_U4011
g13974 and P1_U6785 P1_U6786 P1_U6787 ; P1_U4012
g13975 and P1_U6789 P1_U6790 P1_U6791 ; P1_U4013
g13976 and P1_U6793 P1_U6794 P1_U6795 ; P1_U4014
g13977 and P1_U6797 P1_U6798 P1_U6799 ; P1_U4015
g13978 and P1_U6801 P1_U6802 P1_U6803 ; P1_U4016
g13979 and P1_U6805 P1_U6806 P1_U6807 ; P1_U4017
g13980 and P1_U6809 P1_U6810 P1_U6811 ; P1_U4018
g13981 and P1_U6813 P1_U6814 P1_U6815 ; P1_U4019
g13982 and P1_U6817 P1_U6818 P1_U6819 ; P1_U4020
g13983 and P1_U6821 P1_U6822 ; P1_U4021
g13984 and P1_U6826 P1_U6827 P1_U6828 ; P1_U4022
g13985 and P1_U6830 P1_U6831 P1_U6832 ; P1_U4023
g13986 and P1_U6834 P1_U6835 P1_U6836 ; P1_U4024
g13987 and P1_U6838 P1_U6839 P1_U6840 ; P1_U4025
g13988 and P1_U6858 P1_U6857 ; P1_U4026
g13989 and P1_U6860 P1_U6861 ; P1_U4027
g13990 and P1_U7494 P1_U6888 P1_U3283 ; P1_U4028
g13991 and P1_U6895 P1_U6894 P1_U6893 P1_U6892 ; P1_U4029
g13992 and P1_U6899 P1_U6898 P1_U6897 P1_U6896 ; P1_U4030
g13993 and P1_U6903 P1_U6902 P1_U6901 P1_U6900 ; P1_U4031
g13994 and P1_U6907 P1_U6906 P1_U6905 P1_U6904 ; P1_U4032
g13995 and P1_U6913 P1_U6912 P1_U6911 P1_U6910 ; P1_U4033
g13996 and P1_U6917 P1_U6916 P1_U6915 P1_U6914 ; P1_U4034
g13997 and P1_U6921 P1_U6920 P1_U6919 P1_U6918 ; P1_U4035
g13998 and P1_U6925 P1_U6924 P1_U6923 P1_U6922 ; P1_U4036
g13999 and P1_U6944 P1_U6943 P1_U6942 P1_U6941 ; P1_U4037
g14000 and P1_U6948 P1_U6947 P1_U6946 P1_U6945 ; P1_U4038
g14001 and P1_U6952 P1_U6951 P1_U6950 P1_U6949 ; P1_U4039
g14002 and P1_U6956 P1_U6955 P1_U6954 P1_U6953 ; P1_U4040
g14003 and P1_U6961 P1_U6960 P1_U6959 P1_U6958 ; P1_U4041
g14004 and P1_U6965 P1_U6964 P1_U6963 P1_U6962 ; P1_U4042
g14005 and P1_U6969 P1_U6968 P1_U6967 P1_U6966 ; P1_U4043
g14006 and P1_U6973 P1_U6972 P1_U6971 P1_U6970 ; P1_U4044
g14007 and P1_U6978 P1_U6977 P1_U6976 P1_U6975 ; P1_U4045
g14008 and P1_U6982 P1_U6981 P1_U6980 P1_U6979 ; P1_U4046
g14009 and P1_U6986 P1_U6985 P1_U6984 P1_U6983 ; P1_U4047
g14010 and P1_U6990 P1_U6989 P1_U6988 P1_U6987 ; P1_U4048
g14011 and P1_U6995 P1_U6994 P1_U6993 P1_U6992 ; P1_U4049
g14012 and P1_U6999 P1_U6998 P1_U6997 P1_U6996 ; P1_U4050
g14013 and P1_U7003 P1_U7002 P1_U7001 P1_U7000 ; P1_U4051
g14014 and P1_U7614 P1_U7006 P1_U7005 P1_U7004 ; P1_U4052
g14015 and P1_U7010 P1_U7009 P1_U7008 P1_U7007 ; P1_U4053
g14016 and P1_U7014 P1_U7013 P1_U7012 P1_U7011 ; P1_U4054
g14017 and P1_U7018 P1_U7017 P1_U7016 P1_U7015 ; P1_U4055
g14018 and P1_U7022 P1_U7021 P1_U7020 P1_U7019 ; P1_U4056
g14019 and P1_U7027 P1_U7026 P1_U7025 P1_U7024 ; P1_U4057
g14020 and P1_U7031 P1_U7030 P1_U7029 P1_U7028 ; P1_U4058
g14021 and P1_U7035 P1_U7034 P1_U7033 P1_U7032 ; P1_U4059
g14022 and P1_U7039 P1_U7038 P1_U7037 P1_U7036 ; P1_U4060
g14023 and P1_U7059 P1_U3443 ; P1_U4061
g14024 and P1_U7062 P1_STATE2_REG_0__SCAN_IN ; P1_U4062
g14025 and P1_U7069 P1_U7068 P1_U7067 P1_U7066 ; P1_U4063
g14026 and P1_U7073 P1_U7072 P1_U7071 P1_U7070 ; P1_U4064
g14027 and P1_U7077 P1_U7076 P1_U7075 P1_U7074 ; P1_U4065
g14028 and P1_U7081 P1_U7080 P1_U7079 P1_U7078 ; P1_U4066
g14029 and P1_U4256 P1_STATE2_REG_0__SCAN_IN ; P1_U4067
g14030 and P1_U4405 P1_U4404 P1_U4403 P1_U4401 ; P1_U4068
g14031 and P1_U4407 P1_U4406 P1_U4408 ; P1_U4069
g14032 and P1_U4412 P1_U4411 P1_U4410 P1_U4409 ; P1_U4070
g14033 and P1_U4414 P1_U4413 ; P1_U4071
g14034 and P1_U4400 P1_U3391 ; P1_U4072
g14035 and P1_U3284 P1_STATE2_REG_0__SCAN_IN ; P1_U4073
g14036 and P1_U7090 P1_U7089 ; P1_U4074
g14037 and P1_U7472 P1_U3434 P1_U7473 ; P1_U4075
g14038 and P1_U7475 P1_U7476 P1_U7474 ; P1_U4076
g14039 and P1_U2606 P1_U7477 P1_U4076 ; P1_U4077
g14040 and P1_U7097 P1_U7095 ; P1_U4078
g14041 and P1_U7101 P1_U7100 P1_U7099 P1_U7098 ; P1_U4079
g14042 and P1_U7105 P1_U7104 P1_U7103 P1_U7102 ; P1_U4080
g14043 and P1_U7109 P1_U7108 P1_U7107 P1_U7106 ; P1_U4081
g14044 and P1_U7113 P1_U7112 P1_U7111 P1_U7110 ; P1_U4082
g14045 and P1_U7118 P1_U7117 P1_U7116 P1_U7115 ; P1_U4083
g14046 and P1_U7122 P1_U7121 P1_U7120 P1_U7119 ; P1_U4084
g14047 and P1_U7126 P1_U7125 P1_U7124 P1_U7123 ; P1_U4085
g14048 and P1_U7130 P1_U7129 P1_U7128 P1_U7127 ; P1_U4086
g14049 and P1_U7135 P1_U7134 P1_U7133 P1_U7132 ; P1_U4087
g14050 and P1_U7139 P1_U7138 P1_U7137 P1_U7136 ; P1_U4088
g14051 and P1_U7143 P1_U7142 P1_U7141 P1_U7140 ; P1_U4089
g14052 and P1_U7145 P1_U7144 ; P1_U4090
g14053 and P1_U7617 P1_U7146 P1_U4090 ; P1_U4091
g14054 and P1_U7150 P1_U7149 P1_U7148 P1_U7147 ; P1_U4092
g14055 and P1_U7154 P1_U7153 P1_U7152 P1_U7151 ; P1_U4093
g14056 and P1_U7158 P1_U7157 P1_U7156 P1_U7155 ; P1_U4094
g14057 and P1_U7162 P1_U7161 P1_U7160 P1_U7159 ; P1_U4095
g14058 and P1_U7167 P1_U7166 P1_U7165 P1_U7164 ; P1_U4096
g14059 and P1_U7171 P1_U7170 P1_U7169 P1_U7168 ; P1_U4097
g14060 and P1_U7175 P1_U7174 P1_U7173 P1_U7172 ; P1_U4098
g14061 and P1_U7179 P1_U7178 P1_U7177 P1_U7176 ; P1_U4099
g14062 and P1_U7184 P1_U7183 P1_U7182 P1_U7181 ; P1_U4100
g14063 and P1_U7188 P1_U7187 P1_U7186 P1_U7185 ; P1_U4101
g14064 and P1_U7192 P1_U7191 P1_U7190 P1_U7189 ; P1_U4102
g14065 and P1_U7196 P1_U7195 P1_U7194 P1_U7193 ; P1_U4103
g14066 and P1_U7201 P1_U7200 P1_U7199 P1_U7198 ; P1_U4104
g14067 and P1_U7205 P1_U7204 P1_U7203 P1_U7202 ; P1_U4105
g14068 and P1_U7209 P1_U7208 P1_U7207 P1_U7206 ; P1_U4106
g14069 and P1_U7213 P1_U7212 P1_U7211 P1_U7210 ; P1_U4107
g14070 and P1_U7215 P1_U3264 ; P1_U4108
g14071 and P1_U7216 P1_U7215 ; P1_U4109
g14072 and P1_U7217 P1_U3265 ; P1_U4110
g14073 and P1_U7089 P1_U3427 ; P1_U4111
g14074 and P1_U7218 P1_U7217 ; P1_U4112
g14075 and P1_U4112 P1_U7472 P1_U7473 ; P1_U4113
g14076 and P1_U7090 P1_U3434 P1_U4111 P1_U4113 ; P1_U4114
g14077 and P1_U7486 P1_U7480 P1_U7476 P1_U7474 ; P1_U4115
g14078 and P1_U7505 P1_U7489 P1_U7488 P1_U7487 ; P1_U4116
g14079 and P1_U7090 P1_U7089 ; P1_U4117
g14080 and P1_U7472 P1_U3434 P1_U7473 ; P1_U4118
g14081 and P1_U7475 P1_U7476 P1_U7474 ; P1_U4119
g14082 and P1_U2608 P1_U7477 P1_U2606 P1_U4119 ; P1_U4120
g14083 and P1_U7223 P1_U7222 P1_U7221 P1_U7220 ; P1_U4121
g14084 and P1_U7227 P1_U7226 P1_U7225 P1_U7224 ; P1_U4122
g14085 and P1_U7231 P1_U7230 P1_U7229 P1_U7228 ; P1_U4123
g14086 and P1_U7235 P1_U7234 P1_U7233 P1_U7232 ; P1_U4124
g14087 and P1_U7240 P1_U7239 P1_U7238 P1_U7237 ; P1_U4125
g14088 and P1_U7244 P1_U7243 P1_U7242 P1_U7241 ; P1_U4126
g14089 and P1_U7248 P1_U7247 P1_U7246 P1_U7245 ; P1_U4127
g14090 and P1_U7252 P1_U7251 P1_U7250 P1_U7249 ; P1_U4128
g14091 and P1_U7257 P1_U7256 P1_U7255 P1_U7254 ; P1_U4129
g14092 and P1_U7261 P1_U7260 P1_U7259 P1_U7258 ; P1_U4130
g14093 and P1_U7265 P1_U7264 P1_U7263 P1_U7262 ; P1_U4131
g14094 and P1_U7269 P1_U7268 P1_U7267 P1_U7266 ; P1_U4132
g14095 and P1_U7274 P1_U7273 P1_U7272 P1_U7271 ; P1_U4133
g14096 and P1_U7278 P1_U7277 P1_U7276 P1_U7275 ; P1_U4134
g14097 and P1_U7282 P1_U7281 P1_U7280 P1_U7279 ; P1_U4135
g14098 and P1_U7619 P1_U7285 P1_U7284 P1_U7283 ; P1_U4136
g14099 and P1_U7289 P1_U7288 P1_U7287 P1_U7286 ; P1_U4137
g14100 and P1_U7293 P1_U7292 P1_U7291 P1_U7290 ; P1_U4138
g14101 and P1_U7297 P1_U7296 P1_U7295 P1_U7294 ; P1_U4139
g14102 and P1_U7301 P1_U7300 P1_U7299 P1_U7298 ; P1_U4140
g14103 and P1_U7306 P1_U7305 P1_U7304 P1_U7303 ; P1_U4141
g14104 and P1_U7310 P1_U7309 P1_U7308 P1_U7307 ; P1_U4142
g14105 and P1_U7314 P1_U7313 P1_U7312 P1_U7311 ; P1_U4143
g14106 and P1_U7318 P1_U7317 P1_U7316 P1_U7315 ; P1_U4144
g14107 and P1_U7323 P1_U7322 P1_U7321 P1_U7320 ; P1_U4145
g14108 and P1_U7327 P1_U7326 P1_U7325 P1_U7324 ; P1_U4146
g14109 and P1_U7331 P1_U7330 P1_U7329 P1_U7328 ; P1_U4147
g14110 and P1_U7335 P1_U7334 P1_U7333 P1_U7332 ; P1_U4148
g14111 and P1_U7340 P1_U7339 P1_U7338 P1_U7337 ; P1_U4149
g14112 and P1_U7344 P1_U7343 P1_U7342 P1_U7341 ; P1_U4150
g14113 and P1_U7348 P1_U7347 P1_U7346 P1_U7345 ; P1_U4151
g14114 and P1_U7352 P1_U7351 P1_U7350 P1_U7349 ; P1_U4152
g14115 and P1_U3284 P1_U3419 ; P1_U4153
g14116 and P1_U3283 P1_U3391 ; P1_U4154
g14117 and P1_U7357 P1_U7358 P1_U4263 ; P1_U4155
g14118 and P1_U4155 P1_U7359 ; P1_U4156
g14119 and P1_U2427 P1_STATE2_REG_0__SCAN_IN ; P1_U4157
g14120 and P1_U4157 P1_U7360 ; P1_U4158
g14121 and P1_U3271 P1_U4173 ; P1_U4159
g14122 and P1_U4173 P1_STATE2_REG_0__SCAN_IN ; P1_U4160
g14123 and P1_U7369 P1_STATE2_REG_0__SCAN_IN ; P1_U4161
g14124 and P1_U7371 P1_U2603 ; P1_U4162
g14125 and P1_U7373 P1_STATE2_REG_0__SCAN_IN ; P1_U4163
g14126 and P1_U7375 P1_U2603 ; P1_U4164
g14127 and P1_U7382 P1_U7383 ; P1_U4165
g14128 and P1_U3453 P1_U7384 ; P1_U4166
g14129 and P1_U7389 P1_U7388 P1_U7387 ; P1_U4167
g14130 and P1_U7462 P1_U7461 ; P1_U4168
g14131 and P1_U7465 P1_U7464 ; P1_U4169
g14132 and P1_U7674 P1_U7673 ; P1_U4170
g14133 nand P1_U3572 P1_U3571 P1_U3570 P1_U3569 ; P1_U4171
g14134 nand P1_U3739 P1_U5474 ; P1_U4172
g14135 nand P1_U3576 P1_U2607 P1_U3575 P1_U3574 P1_U3573 ; P1_U4173
g14136 not P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_U4174
g14137 and P1_U7726 P1_U7725 ; P1_U4175
g14138 and P1_U7745 P1_U7744 ; P1_U4176
g14139 nand P1_U2368 P1_U3285 ; P1_U4177
g14140 nand P1_U4508 P1_U3391 ; P1_U4178
g14141 not BS16 ; P1_U4179
g14142 nand P1_U3967 P1_U4228 ; P1_U4180
g14143 nand P1_U4228 P1_U3432 ; P1_U4181
g14144 nand P1_U7698 P1_U7697 P1_U3738 ; P1_U4182
g14145 nand P1_U3269 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U4183
g14146 not P1_U3452 ; P1_U4184
g14147 nand HOLD P1_U3257 ; P1_U4185
g14148 not P1_U3412 ; P1_U4186
g14149 not P1_U3440 ; P1_U4187
g14150 not P1_U3439 ; P1_U4188
g14151 not P1_U3393 ; P1_U4189
g14152 not P1_U3290 ; P1_U4190
g14153 not P1_U3449 ; P1_U4191
g14154 not P1_U3405 ; P1_U4192
g14155 not P1_U3434 ; P1_U4193
g14156 not P1_U3420 ; P1_U4194
g14157 nand P1_U4265 P1_U3271 ; P1_U4195
g14158 nand P1_U4460 P1_U2605 ; P1_U4196
g14159 not P1_U3396 ; P1_U4197
g14160 not P1_U3425 ; P1_U4198
g14161 not P1_U3289 ; P1_U4199
g14162 not P1_U3421 ; P1_U4200
g14163 not P1_U3422 ; P1_U4201
g14164 not P1_U3428 ; P1_U4202
g14165 not P1_U3408 ; P1_U4203
g14166 not P1_U3427 ; P1_U4204
g14167 nand P1_U3885 P1_U4189 P1_U4197 ; P1_U4205
g14168 not P1_U3418 ; P1_U4206
g14169 not P1_U3443 ; P1_U4207
g14170 not P1_U3282 ; P1_U4208
g14171 not P1_U3307 ; P1_U4209
g14172 not P1_U3390 ; P1_U4210
g14173 not P1_U3446 ; P1_U4211
g14174 not P1_U3447 ; P1_U4212
g14175 not P1_U3448 ; P1_U4213
g14176 not P1_U3400 ; P1_U4214
g14177 not P1_U3288 ; P1_U4215
g14178 not P1_U3292 ; P1_U4216
g14179 nand P1_U3578 P1_U2431 ; P1_U4217
g14180 not P1_U3399 ; P1_U4218
g14181 nand P1_U4449 P1_U3271 ; P1_U4219
g14182 not P1_U3433 ; P1_U4220
g14183 not P1_U3249 ; P1_U4221
g14184 not P1_U3426 ; P1_U4222
g14185 not P1_U3424 ; P1_U4223
g14186 not P1_U3300 ; P1_U4224
g14187 not P1_LT_563_1260_U6 ; P1_U4225
g14188 not P1_U3320 ; P1_U4226
g14189 nand P1_U4255 P1_U3431 ; P1_U4227
g14190 nand P1_U4235 P1_U7500 ; P1_U4228
g14191 nand P1_U2362 P1_U3272 ; P1_U4229
g14192 nand P1_U2363 P1_U4377 ; P1_U4230
g14193 not P1_U3407 ; P1_U4231
g14194 not P1_U3252 ; P1_U4232
g14195 not P1_U3250 ; P1_U4233
g14196 not P1_U3395 ; P1_U4234
g14197 not P1_U3297 ; P1_U4235
g14198 not P1_U3398 ; P1_U4236
g14199 not P1_U4178 ; P1_U4237
g14200 not P1_U3357 ; P1_U4238
g14201 nand P1_U4477 P1_U7381 ; P1_U4239
g14202 nand P1_U3963 P1_U4220 ; P1_U4240
g14203 nand P1_U3584 P1_U4261 ; P1_U4241
g14204 nand P1_U3731 P1_U2428 ; P1_U4242
g14205 nand P1_U4364 P1_U3258 ; P1_U4243
g14206 nand P1_U3294 P1_U2352 P1_STATE2_REG_1__SCAN_IN ; P1_U4244
g14207 nand P1_U2428 P1_U3403 ; P1_U4245
g14208 nand P1_U3263 U210 P1_STATE2_REG_0__SCAN_IN ; P1_U4246
g14209 not P1_U3394 ; P1_U4247
g14210 nand P1_U2451 P1_U2353 P1_U3862 P1_U2448 ; P1_U4248
g14211 not P1_U3287 ; P1_U4249
g14212 not P1_U3397 ; P1_U4250
g14213 not P1_U3415 ; P1_U4251
g14214 not P1_U3299 ; P1_U4252
g14215 not P1_U3409 ; P1_U4253
g14216 not P1_U3419 ; P1_U4254
g14217 not P1_U3432 ; P1_U4255
g14218 not P1_U3291 ; P1_U4256
g14219 not P1_U3389 ; P1_U4257
g14220 not P1_U3254 ; P1_U4258
g14221 not P1_U3281 ; P1_U4259
g14222 not P1_U3406 ; P1_U4260
g14223 not P1_U3298 ; P1_U4261
g14224 not P1_U3286 ; P1_U4262
g14225 nand P1_U4236 P1_U4399 ; P1_U4263
g14226 not P1_U3411 ; P1_U4264
g14227 not P1_U3453 ; P1_U4265
g14228 not P1_U3410 ; P1_U4266
g14229 nand P1_U4233 P1_REIP_REG_31__SCAN_IN ; P1_U4267
g14230 nand P1_U4232 P1_REIP_REG_30__SCAN_IN ; P1_U4268
g14231 nand P1_U3249 P1_ADDRESS_REG_29__SCAN_IN ; P1_U4269
g14232 nand P1_U4233 P1_REIP_REG_30__SCAN_IN ; P1_U4270
g14233 nand P1_U4232 P1_REIP_REG_29__SCAN_IN ; P1_U4271
g14234 nand P1_U3249 P1_ADDRESS_REG_28__SCAN_IN ; P1_U4272
g14235 nand P1_U4233 P1_REIP_REG_29__SCAN_IN ; P1_U4273
g14236 nand P1_U4232 P1_REIP_REG_28__SCAN_IN ; P1_U4274
g14237 nand P1_U3249 P1_ADDRESS_REG_27__SCAN_IN ; P1_U4275
g14238 nand P1_U4233 P1_REIP_REG_28__SCAN_IN ; P1_U4276
g14239 nand P1_U4232 P1_REIP_REG_27__SCAN_IN ; P1_U4277
g14240 nand P1_U3249 P1_ADDRESS_REG_26__SCAN_IN ; P1_U4278
g14241 nand P1_U4233 P1_REIP_REG_27__SCAN_IN ; P1_U4279
g14242 nand P1_U4232 P1_REIP_REG_26__SCAN_IN ; P1_U4280
g14243 nand P1_U3249 P1_ADDRESS_REG_25__SCAN_IN ; P1_U4281
g14244 nand P1_U4233 P1_REIP_REG_26__SCAN_IN ; P1_U4282
g14245 nand P1_U4232 P1_REIP_REG_25__SCAN_IN ; P1_U4283
g14246 nand P1_U3249 P1_ADDRESS_REG_24__SCAN_IN ; P1_U4284
g14247 nand P1_U4233 P1_REIP_REG_25__SCAN_IN ; P1_U4285
g14248 nand P1_U4232 P1_REIP_REG_24__SCAN_IN ; P1_U4286
g14249 nand P1_U3249 P1_ADDRESS_REG_23__SCAN_IN ; P1_U4287
g14250 nand P1_U4233 P1_REIP_REG_24__SCAN_IN ; P1_U4288
g14251 nand P1_U4232 P1_REIP_REG_23__SCAN_IN ; P1_U4289
g14252 nand P1_U3249 P1_ADDRESS_REG_22__SCAN_IN ; P1_U4290
g14253 nand P1_U4233 P1_REIP_REG_23__SCAN_IN ; P1_U4291
g14254 nand P1_U4232 P1_REIP_REG_22__SCAN_IN ; P1_U4292
g14255 nand P1_U3249 P1_ADDRESS_REG_21__SCAN_IN ; P1_U4293
g14256 nand P1_U4233 P1_REIP_REG_22__SCAN_IN ; P1_U4294
g14257 nand P1_U4232 P1_REIP_REG_21__SCAN_IN ; P1_U4295
g14258 nand P1_U3249 P1_ADDRESS_REG_20__SCAN_IN ; P1_U4296
g14259 nand P1_U4233 P1_REIP_REG_21__SCAN_IN ; P1_U4297
g14260 nand P1_U4232 P1_REIP_REG_20__SCAN_IN ; P1_U4298
g14261 nand P1_U3249 P1_ADDRESS_REG_19__SCAN_IN ; P1_U4299
g14262 nand P1_U4233 P1_REIP_REG_20__SCAN_IN ; P1_U4300
g14263 nand P1_U4232 P1_REIP_REG_19__SCAN_IN ; P1_U4301
g14264 nand P1_U3249 P1_ADDRESS_REG_18__SCAN_IN ; P1_U4302
g14265 nand P1_U4233 P1_REIP_REG_19__SCAN_IN ; P1_U4303
g14266 nand P1_U4232 P1_REIP_REG_18__SCAN_IN ; P1_U4304
g14267 nand P1_U3249 P1_ADDRESS_REG_17__SCAN_IN ; P1_U4305
g14268 nand P1_U4233 P1_REIP_REG_18__SCAN_IN ; P1_U4306
g14269 nand P1_U4232 P1_REIP_REG_17__SCAN_IN ; P1_U4307
g14270 nand P1_U3249 P1_ADDRESS_REG_16__SCAN_IN ; P1_U4308
g14271 nand P1_U4233 P1_REIP_REG_17__SCAN_IN ; P1_U4309
g14272 nand P1_U4232 P1_REIP_REG_16__SCAN_IN ; P1_U4310
g14273 nand P1_U3249 P1_ADDRESS_REG_15__SCAN_IN ; P1_U4311
g14274 nand P1_U4233 P1_REIP_REG_16__SCAN_IN ; P1_U4312
g14275 nand P1_U4232 P1_REIP_REG_15__SCAN_IN ; P1_U4313
g14276 nand P1_U3249 P1_ADDRESS_REG_14__SCAN_IN ; P1_U4314
g14277 nand P1_U4233 P1_REIP_REG_15__SCAN_IN ; P1_U4315
g14278 nand P1_U4232 P1_REIP_REG_14__SCAN_IN ; P1_U4316
g14279 nand P1_U3249 P1_ADDRESS_REG_13__SCAN_IN ; P1_U4317
g14280 nand P1_U4233 P1_REIP_REG_14__SCAN_IN ; P1_U4318
g14281 nand P1_U4232 P1_REIP_REG_13__SCAN_IN ; P1_U4319
g14282 nand P1_U3249 P1_ADDRESS_REG_12__SCAN_IN ; P1_U4320
g14283 nand P1_U4233 P1_REIP_REG_13__SCAN_IN ; P1_U4321
g14284 nand P1_U4232 P1_REIP_REG_12__SCAN_IN ; P1_U4322
g14285 nand P1_U3249 P1_ADDRESS_REG_11__SCAN_IN ; P1_U4323
g14286 nand P1_U4233 P1_REIP_REG_12__SCAN_IN ; P1_U4324
g14287 nand P1_U4232 P1_REIP_REG_11__SCAN_IN ; P1_U4325
g14288 nand P1_U3249 P1_ADDRESS_REG_10__SCAN_IN ; P1_U4326
g14289 nand P1_U4233 P1_REIP_REG_11__SCAN_IN ; P1_U4327
g14290 nand P1_U4232 P1_REIP_REG_10__SCAN_IN ; P1_U4328
g14291 nand P1_U3249 P1_ADDRESS_REG_9__SCAN_IN ; P1_U4329
g14292 nand P1_U4233 P1_REIP_REG_10__SCAN_IN ; P1_U4330
g14293 nand P1_U4232 P1_REIP_REG_9__SCAN_IN ; P1_U4331
g14294 nand P1_U3249 P1_ADDRESS_REG_8__SCAN_IN ; P1_U4332
g14295 nand P1_U4233 P1_REIP_REG_9__SCAN_IN ; P1_U4333
g14296 nand P1_U4232 P1_REIP_REG_8__SCAN_IN ; P1_U4334
g14297 nand P1_U3249 P1_ADDRESS_REG_7__SCAN_IN ; P1_U4335
g14298 nand P1_U4233 P1_REIP_REG_8__SCAN_IN ; P1_U4336
g14299 nand P1_U4232 P1_REIP_REG_7__SCAN_IN ; P1_U4337
g14300 nand P1_U3249 P1_ADDRESS_REG_6__SCAN_IN ; P1_U4338
g14301 nand P1_U4233 P1_REIP_REG_7__SCAN_IN ; P1_U4339
g14302 nand P1_U4232 P1_REIP_REG_6__SCAN_IN ; P1_U4340
g14303 nand P1_U3249 P1_ADDRESS_REG_5__SCAN_IN ; P1_U4341
g14304 nand P1_U4233 P1_REIP_REG_6__SCAN_IN ; P1_U4342
g14305 nand P1_U4232 P1_REIP_REG_5__SCAN_IN ; P1_U4343
g14306 nand P1_U3249 P1_ADDRESS_REG_4__SCAN_IN ; P1_U4344
g14307 nand P1_U4233 P1_REIP_REG_5__SCAN_IN ; P1_U4345
g14308 nand P1_U4232 P1_REIP_REG_4__SCAN_IN ; P1_U4346
g14309 nand P1_U3249 P1_ADDRESS_REG_3__SCAN_IN ; P1_U4347
g14310 nand P1_U4233 P1_REIP_REG_4__SCAN_IN ; P1_U4348
g14311 nand P1_U4232 P1_REIP_REG_3__SCAN_IN ; P1_U4349
g14312 nand P1_U3249 P1_ADDRESS_REG_2__SCAN_IN ; P1_U4350
g14313 nand P1_U4233 P1_REIP_REG_3__SCAN_IN ; P1_U4351
g14314 nand P1_U4232 P1_REIP_REG_2__SCAN_IN ; P1_U4352
g14315 nand P1_U3249 P1_ADDRESS_REG_1__SCAN_IN ; P1_U4353
g14316 nand P1_U4233 P1_REIP_REG_2__SCAN_IN ; P1_U4354
g14317 nand P1_U4232 P1_REIP_REG_1__SCAN_IN ; P1_U4355
g14318 nand P1_U3249 P1_ADDRESS_REG_0__SCAN_IN ; P1_U4356
g14319 not P1_U3260 ; P1_U4357
g14320 nand P1_U4357 P1_U3257 ; P1_U4358
g14321 nand NA P1_U4258 ; P1_U4359
g14322 not P1_U3261 ; P1_U4360
g14323 nand P1_U4360 P1_U3257 ; P1_U4361
g14324 or NA P1_STATE_REG_0__SCAN_IN ; P1_U4362
g14325 nand P1_U7622 P1_U4362 P1_U7623 ; P1_U4363
g14326 not P1_U3255 ; P1_U4364
g14327 nand HOLD P1_U3247 P1_U4364 ; P1_U4365
g14328 nand P1_U3261 U210 P1_STATE_REG_1__SCAN_IN ; P1_U4366
g14329 nand P1_U4366 P1_U4365 ; P1_U4367
g14330 nand P1_U4359 P1_U4367 P1_STATE_REG_0__SCAN_IN ; P1_U4368
g14331 nand P1_U4363 P1_STATE_REG_2__SCAN_IN ; P1_U4369
g14332 nand U210 P1_U4221 ; P1_U4370
g14333 nand P1_U3496 P1_U7625 ; P1_U4371
g14334 nand P1_U3260 P1_STATE_REG_2__SCAN_IN ; P1_U4372
g14335 nand NA P1_U3258 ; P1_U4373
g14336 nand P1_U4373 P1_U4372 ; P1_U4374
g14337 nand P1_U4374 P1_U3248 ; P1_U4375
g14338 nand P1_U4179 P1_U3255 ; P1_U4376
g14339 not P1_U3280 ; P1_U4377
g14340 not P1_U3269 ; P1_U4378
g14341 not P1_U3444 ; P1_U4379
g14342 not P1_U3268 ; P1_U4380
g14343 not P1_U3274 ; P1_U4381
g14344 not P1_U3267 ; P1_U4382
g14345 nand P1_U4382 P1_INSTQUEUE_REG_7__3__SCAN_IN ; P1_U4383
g14346 nand P1_U2472 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U4384
g14347 nand P1_U2471 P1_INSTQUEUE_REG_1__3__SCAN_IN ; P1_U4385
g14348 nand P1_U2470 P1_INSTQUEUE_REG_2__3__SCAN_IN ; P1_U4386
g14349 nand P1_U2468 P1_INSTQUEUE_REG_3__3__SCAN_IN ; P1_U4387
g14350 nand P1_U2467 P1_INSTQUEUE_REG_4__3__SCAN_IN ; P1_U4388
g14351 nand P1_U2466 P1_INSTQUEUE_REG_5__3__SCAN_IN ; P1_U4389
g14352 nand P1_U2465 P1_INSTQUEUE_REG_6__3__SCAN_IN ; P1_U4390
g14353 nand P1_U2464 P1_INSTQUEUE_REG_8__3__SCAN_IN ; P1_U4391
g14354 nand P1_U2463 P1_INSTQUEUE_REG_9__3__SCAN_IN ; P1_U4392
g14355 nand P1_U2461 P1_INSTQUEUE_REG_10__3__SCAN_IN ; P1_U4393
g14356 nand P1_U2459 P1_INSTQUEUE_REG_11__3__SCAN_IN ; P1_U4394
g14357 nand P1_U2458 P1_INSTQUEUE_REG_12__3__SCAN_IN ; P1_U4395
g14358 nand P1_U2457 P1_INSTQUEUE_REG_13__3__SCAN_IN ; P1_U4396
g14359 nand P1_U2455 P1_INSTQUEUE_REG_14__3__SCAN_IN ; P1_U4397
g14360 nand P1_U2453 P1_INSTQUEUE_REG_15__3__SCAN_IN ; P1_U4398
g14361 not P1_U3283 ; P1_U4399
g14362 not P1_U3278 ; P1_U4400
g14363 nand P1_U3270 P1_INSTQUEUE_REG_7__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U4401
g14364 nand P1_U3270 P1_U4380 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U4402
g14365 nand P1_U2469 P1_U3265 P1_INSTQUEUE_REG_1__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U4403
g14366 nand P1_U2469 P1_U3266 P1_INSTQUEUE_REG_2__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U4404
g14367 nand P1_U4378 P1_U3270 P1_INSTQUEUE_REG_4__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U4405
g14368 nand P1_U3520 P1_U3521 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U4406
g14369 nand P1_U3522 P1_U3523 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U4407
g14370 nand P1_U3524 P1_U4380 ; P1_U4408
g14371 nand P1_U3525 P1_U3526 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U4409
g14372 nand P1_U3264 P1_INSTQUEUE_REG_11__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U4410
g14373 nand P1_U4378 P1_U3527 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U4411
g14374 nand P1_U3265 P1_INSTQUEUE_REG_13__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U4412
g14375 nand P1_U3266 P1_INSTQUEUE_REG_14__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U4413
g14376 nand P1_INSTQUEUE_REG_15__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U4414
g14377 not P1_U4173 ; P1_U4415
g14378 nand P1_U4382 P1_INSTQUEUE_REG_7__2__SCAN_IN ; P1_U4416
g14379 nand P1_U2472 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U4417
g14380 nand P1_U2471 P1_INSTQUEUE_REG_1__2__SCAN_IN ; P1_U4418
g14381 nand P1_U2470 P1_INSTQUEUE_REG_2__2__SCAN_IN ; P1_U4419
g14382 nand P1_U2468 P1_INSTQUEUE_REG_3__2__SCAN_IN ; P1_U4420
g14383 nand P1_U2467 P1_INSTQUEUE_REG_4__2__SCAN_IN ; P1_U4421
g14384 nand P1_U2466 P1_INSTQUEUE_REG_5__2__SCAN_IN ; P1_U4422
g14385 nand P1_U2465 P1_INSTQUEUE_REG_6__2__SCAN_IN ; P1_U4423
g14386 nand P1_U2464 P1_INSTQUEUE_REG_8__2__SCAN_IN ; P1_U4424
g14387 nand P1_U2463 P1_INSTQUEUE_REG_9__2__SCAN_IN ; P1_U4425
g14388 nand P1_U2461 P1_INSTQUEUE_REG_10__2__SCAN_IN ; P1_U4426
g14389 nand P1_U2459 P1_INSTQUEUE_REG_11__2__SCAN_IN ; P1_U4427
g14390 nand P1_U2458 P1_INSTQUEUE_REG_12__2__SCAN_IN ; P1_U4428
g14391 nand P1_U2457 P1_INSTQUEUE_REG_13__2__SCAN_IN ; P1_U4429
g14392 nand P1_U2455 P1_INSTQUEUE_REG_14__2__SCAN_IN ; P1_U4430
g14393 nand P1_U2453 P1_INSTQUEUE_REG_15__2__SCAN_IN ; P1_U4431
g14394 not P1_U4171 ; P1_U4432
g14395 nand P1_U4382 P1_INSTQUEUE_REG_7__7__SCAN_IN ; P1_U4433
g14396 nand P1_U2472 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U4434
g14397 nand P1_U2471 P1_INSTQUEUE_REG_1__7__SCAN_IN ; P1_U4435
g14398 nand P1_U2470 P1_INSTQUEUE_REG_2__7__SCAN_IN ; P1_U4436
g14399 nand P1_U2468 P1_INSTQUEUE_REG_3__7__SCAN_IN ; P1_U4437
g14400 nand P1_U2467 P1_INSTQUEUE_REG_4__7__SCAN_IN ; P1_U4438
g14401 nand P1_U2466 P1_INSTQUEUE_REG_5__7__SCAN_IN ; P1_U4439
g14402 nand P1_U2465 P1_INSTQUEUE_REG_6__7__SCAN_IN ; P1_U4440
g14403 nand P1_U2464 P1_INSTQUEUE_REG_8__7__SCAN_IN ; P1_U4441
g14404 nand P1_U2463 P1_INSTQUEUE_REG_9__7__SCAN_IN ; P1_U4442
g14405 nand P1_U2461 P1_INSTQUEUE_REG_10__7__SCAN_IN ; P1_U4443
g14406 nand P1_U2459 P1_INSTQUEUE_REG_11__7__SCAN_IN ; P1_U4444
g14407 nand P1_U2458 P1_INSTQUEUE_REG_12__7__SCAN_IN ; P1_U4445
g14408 nand P1_U2457 P1_INSTQUEUE_REG_13__7__SCAN_IN ; P1_U4446
g14409 nand P1_U2455 P1_INSTQUEUE_REG_14__7__SCAN_IN ; P1_U4447
g14410 nand P1_U2453 P1_INSTQUEUE_REG_15__7__SCAN_IN ; P1_U4448
g14411 not P1_U3391 ; P1_U4449
g14412 nand P1_U3498 P1_U4381 P1_INSTQUEUE_REG_7__6__SCAN_IN ; P1_U4450
g14413 nand P1_U2469 P1_U2456 P1_INSTQUEUE_REG_1__6__SCAN_IN ; P1_U4451
g14414 nand P1_U2469 P1_U2454 P1_INSTQUEUE_REG_2__6__SCAN_IN ; P1_U4452
g14415 nand P1_U4378 P1_U4381 P1_INSTQUEUE_REG_4__6__SCAN_IN ; P1_U4453
g14416 nand P1_U2456 P1_U4381 P1_INSTQUEUE_REG_5__6__SCAN_IN ; P1_U4454
g14417 nand P1_U2454 P1_U4381 P1_INSTQUEUE_REG_6__6__SCAN_IN ; P1_U4455
g14418 nand P1_U4378 P1_U3507 P1_INSTQUEUE_REG_12__6__SCAN_IN ; P1_U4456
g14419 nand P1_U3507 P1_U2456 P1_INSTQUEUE_REG_13__6__SCAN_IN ; P1_U4457
g14420 nand P1_U3507 P1_U2454 P1_INSTQUEUE_REG_14__6__SCAN_IN ; P1_U4458
g14421 nand P1_U3507 P1_U3498 P1_INSTQUEUE_REG_15__6__SCAN_IN ; P1_U4459
g14422 not P1_U3277 ; P1_U4460
g14423 nand P1_U4382 P1_INSTQUEUE_REG_7__1__SCAN_IN ; P1_U4461
g14424 nand P1_U2472 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U4462
g14425 nand P1_U2471 P1_INSTQUEUE_REG_1__1__SCAN_IN ; P1_U4463
g14426 nand P1_U2470 P1_INSTQUEUE_REG_2__1__SCAN_IN ; P1_U4464
g14427 nand P1_U2468 P1_INSTQUEUE_REG_3__1__SCAN_IN ; P1_U4465
g14428 nand P1_U2467 P1_INSTQUEUE_REG_4__1__SCAN_IN ; P1_U4466
g14429 nand P1_U2466 P1_INSTQUEUE_REG_5__1__SCAN_IN ; P1_U4467
g14430 nand P1_U2465 P1_INSTQUEUE_REG_6__1__SCAN_IN ; P1_U4468
g14431 nand P1_U2464 P1_INSTQUEUE_REG_8__1__SCAN_IN ; P1_U4469
g14432 nand P1_U2463 P1_INSTQUEUE_REG_9__1__SCAN_IN ; P1_U4470
g14433 nand P1_U2461 P1_INSTQUEUE_REG_10__1__SCAN_IN ; P1_U4471
g14434 nand P1_U2459 P1_INSTQUEUE_REG_11__1__SCAN_IN ; P1_U4472
g14435 nand P1_U2458 P1_INSTQUEUE_REG_12__1__SCAN_IN ; P1_U4473
g14436 nand P1_U2457 P1_INSTQUEUE_REG_13__1__SCAN_IN ; P1_U4474
g14437 nand P1_U2455 P1_INSTQUEUE_REG_14__1__SCAN_IN ; P1_U4475
g14438 nand P1_U2453 P1_INSTQUEUE_REG_15__1__SCAN_IN ; P1_U4476
g14439 not P1_U3271 ; P1_U4477
g14440 nand P1_U4382 P1_INSTQUEUE_REG_7__0__SCAN_IN ; P1_U4478
g14441 nand P1_U2472 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U4479
g14442 nand P1_U2471 P1_INSTQUEUE_REG_1__0__SCAN_IN ; P1_U4480
g14443 nand P1_U2470 P1_INSTQUEUE_REG_2__0__SCAN_IN ; P1_U4481
g14444 nand P1_U2468 P1_INSTQUEUE_REG_3__0__SCAN_IN ; P1_U4482
g14445 nand P1_U2467 P1_INSTQUEUE_REG_4__0__SCAN_IN ; P1_U4483
g14446 nand P1_U2466 P1_INSTQUEUE_REG_5__0__SCAN_IN ; P1_U4484
g14447 nand P1_U2465 P1_INSTQUEUE_REG_6__0__SCAN_IN ; P1_U4485
g14448 nand P1_U2464 P1_INSTQUEUE_REG_8__0__SCAN_IN ; P1_U4486
g14449 nand P1_U2463 P1_INSTQUEUE_REG_9__0__SCAN_IN ; P1_U4487
g14450 nand P1_U2461 P1_INSTQUEUE_REG_10__0__SCAN_IN ; P1_U4488
g14451 nand P1_U2459 P1_INSTQUEUE_REG_11__0__SCAN_IN ; P1_U4489
g14452 nand P1_U2458 P1_INSTQUEUE_REG_12__0__SCAN_IN ; P1_U4490
g14453 nand P1_U2457 P1_INSTQUEUE_REG_13__0__SCAN_IN ; P1_U4491
g14454 nand P1_U2455 P1_INSTQUEUE_REG_14__0__SCAN_IN ; P1_U4492
g14455 nand P1_U2453 P1_INSTQUEUE_REG_15__0__SCAN_IN ; P1_U4493
g14456 not P1_U3284 ; P1_U4494
g14457 nand P1_U3248 P1_STATE_REG_2__SCAN_IN ; P1_U4495
g14458 nand P1_U3254 P1_U4495 ; P1_U4496
g14459 not P1_U3272 ; P1_U4497
g14460 nand P1_U4477 P1_U3388 ; P1_U4498
g14461 not P1_U3437 ; P1_U4499
g14462 nand P1_U3272 P1_U3390 P1_U3287 ; P1_U4500
g14463 nand P1_U4500 P1_U3257 ; P1_U4501
g14464 not P1_U3285 ; P1_U4502
g14465 nand P1_U4460 P1_U4173 ; P1_U4503
g14466 nand P1_U4196 P1_U3286 ; P1_U4504
g14467 nand P1_U4504 P1_U3579 ; P1_U4505
g14468 nand P1_U3580 P1_U4505 ; P1_U4506
g14469 nand P1_U4215 P1_U3388 ; P1_U4507
g14470 nand P1_U7682 P1_U7681 P1_U4507 ; P1_U4508
g14471 nand P1_U2448 P1_U4262 ; P1_U4509
g14472 or P1_FLUSH_REG_SCAN_IN P1_MORE_REG_SCAN_IN ; P1_U4510
g14473 not P1_U3293 ; P1_U4511
g14474 nand P1_U4511 P1_U3262 ; P1_U4512
g14475 nand U210 P1_STATE2_REG_1__SCAN_IN ; P1_U4513
g14476 not P1_U3295 ; P1_U4514
g14477 nand P1_U7688 P1_U7687 P1_STATE2_REG_1__SCAN_IN ; P1_U4515
g14478 nand P1_U3295 P1_STATE2_REG_2__SCAN_IN ; P1_U4516
g14479 nand P1_U7604 P1_U4246 ; P1_U4517
g14480 nand P1_U3583 P1_U4514 ; P1_U4518
g14481 nand P1_U4517 P1_STATE2_REG_1__SCAN_IN ; P1_U4519
g14482 nand P1_U2368 P1_U7604 ; P1_U4520
g14483 nand P1_U4252 P1_U4261 ; P1_U4521
g14484 nand P1_U7604 P1_U4245 ; P1_U4522
g14485 nand P1_U2368 P1_U3293 ; P1_U4523
g14486 not P1_U3325 ; P1_U4524
g14487 not P1_U3331 ; P1_U4525
g14488 not P1_U3332 ; P1_U4526
g14489 not P1_U3314 ; P1_U4527
g14490 not P1_U3313 ; P1_U4528
g14491 not P1_U3342 ; P1_U4529
g14492 nand P1_R2144_U8 P1_U3313 ; P1_U4530
g14493 not P1_U3358 ; P1_U4531
g14494 not P1_U3315 ; P1_U4532
g14495 not P1_U3305 ; P1_U4533
g14496 not P1_U3306 ; P1_U4534
g14497 nand P1_U2438 P1_U2442 ; P1_U4535
g14498 not P1_U3321 ; P1_U4536
g14499 not P1_U3356 ; P1_U4537
g14500 not P1_U3340 ; P1_U4538
g14501 nand P1_U3305 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_U4539
g14502 not P1_U3360 ; P1_U4540
g14503 not P1_U3329 ; P1_U4541
g14504 not P1_U3323 ; P1_U4542
g14505 not P1_U3235 ; P1_U4543
g14506 nand P1_U2432 P1_U2436 ; P1_U4544
g14507 not P1_U3322 ; P1_U4545
g14508 nand P1_U3263 P1_STATE2_REG_1__SCAN_IN ; P1_U4546
g14509 nand P1_U4546 P1_U3297 P1_U3299 ; P1_U4547
g14510 nand P1_U4528 P1_U2476 ; P1_U4548
g14511 nand P1_U2480 P1_U2358 ; P1_U4549
g14512 nand P1_U3320 P1_U4549 ; P1_U4550
g14513 nand P1_U4536 P1_U4550 ; P1_U4551
g14514 nand P1_U3306 P1_STATE2_REG_3__SCAN_IN ; P1_U4552
g14515 nand P1_U4545 P1_STATE2_REG_2__SCAN_IN ; P1_U4553
g14516 nand P1_U4551 P1_U3587 ; P1_U4554
g14517 nand P1_U2480 P1_U2388 ; P1_U4555
g14518 nand P1_U3320 P1_U4555 ; P1_U4556
g14519 nand P1_U4556 P1_U3321 ; P1_U4557
g14520 nand P1_U3322 P1_STATE2_REG_2__SCAN_IN ; P1_U4558
g14521 nand P1_U4558 P1_U4557 ; P1_U4559
g14522 nand P1_U2415 P1_U4534 ; P1_U4560
g14523 nand P1_U2413 P1_U2477 ; P1_U4561
g14524 nand P1_U2412 P1_U4532 ; P1_U4562
g14525 nand P1_U2397 P1_U4559 ; P1_U4563
g14526 nand P1_U4554 P1_INSTQUEUE_REG_15__7__SCAN_IN ; P1_U4564
g14527 nand P1_U2416 P1_U4534 ; P1_U4565
g14528 nand P1_U2411 P1_U2477 ; P1_U4566
g14529 nand P1_U2410 P1_U4532 ; P1_U4567
g14530 nand P1_U2396 P1_U4559 ; P1_U4568
g14531 nand P1_U4554 P1_INSTQUEUE_REG_15__6__SCAN_IN ; P1_U4569
g14532 nand P1_U2420 P1_U4534 ; P1_U4570
g14533 nand P1_U2409 P1_U2477 ; P1_U4571
g14534 nand P1_U2408 P1_U4532 ; P1_U4572
g14535 nand P1_U2395 P1_U4559 ; P1_U4573
g14536 nand P1_U4554 P1_INSTQUEUE_REG_15__5__SCAN_IN ; P1_U4574
g14537 nand P1_U2419 P1_U4534 ; P1_U4575
g14538 nand P1_U2407 P1_U2477 ; P1_U4576
g14539 nand P1_U2406 P1_U4532 ; P1_U4577
g14540 nand P1_U2394 P1_U4559 ; P1_U4578
g14541 nand P1_U4554 P1_INSTQUEUE_REG_15__4__SCAN_IN ; P1_U4579
g14542 nand P1_U2418 P1_U4534 ; P1_U4580
g14543 nand P1_U2405 P1_U2477 ; P1_U4581
g14544 nand P1_U2404 P1_U4532 ; P1_U4582
g14545 nand P1_U2393 P1_U4559 ; P1_U4583
g14546 nand P1_U4554 P1_INSTQUEUE_REG_15__3__SCAN_IN ; P1_U4584
g14547 nand P1_U2421 P1_U4534 ; P1_U4585
g14548 nand P1_U2403 P1_U2477 ; P1_U4586
g14549 nand P1_U2402 P1_U4532 ; P1_U4587
g14550 nand P1_U2392 P1_U4559 ; P1_U4588
g14551 nand P1_U4554 P1_INSTQUEUE_REG_15__2__SCAN_IN ; P1_U4589
g14552 nand P1_U2414 P1_U4534 ; P1_U4590
g14553 nand P1_U2401 P1_U2477 ; P1_U4591
g14554 nand P1_U2400 P1_U4532 ; P1_U4592
g14555 nand P1_U2391 P1_U4559 ; P1_U4593
g14556 nand P1_U4554 P1_INSTQUEUE_REG_15__1__SCAN_IN ; P1_U4594
g14557 nand P1_U2417 P1_U4534 ; P1_U4595
g14558 nand P1_U2399 P1_U2477 ; P1_U4596
g14559 nand P1_U2398 P1_U4532 ; P1_U4597
g14560 nand P1_U2390 P1_U4559 ; P1_U4598
g14561 nand P1_U4554 P1_INSTQUEUE_REG_15__0__SCAN_IN ; P1_U4599
g14562 not P1_U3326 ; P1_U4600
g14563 not P1_U3327 ; P1_U4601
g14564 not P1_U3324 ; P1_U4602
g14565 nand P1_U2443 P1_U2438 ; P1_U4603
g14566 not P1_U3328 ; P1_U4604
g14567 not P1_U3236 ; P1_U4605
g14568 nand P1_U4524 P1_U2476 ; P1_U4606
g14569 nand P1_U2482 P1_U2358 ; P1_U4607
g14570 nand P1_U3320 P1_U4607 ; P1_U4608
g14571 nand P1_U4604 P1_U4608 ; P1_U4609
g14572 nand P1_U3324 P1_STATE2_REG_3__SCAN_IN ; P1_U4610
g14573 nand P1_U3236 P1_STATE2_REG_2__SCAN_IN ; P1_U4611
g14574 nand P1_U4609 P1_U3596 ; P1_U4612
g14575 nand P1_U2482 P1_U2388 ; P1_U4613
g14576 nand P1_U3320 P1_U4613 ; P1_U4614
g14577 nand P1_U4614 P1_U3328 ; P1_U4615
g14578 nand P1_U4605 P1_STATE2_REG_2__SCAN_IN ; P1_U4616
g14579 nand P1_U4616 P1_U4615 ; P1_U4617
g14580 nand P1_U4602 P1_U2415 ; P1_U4618
g14581 nand P1_U2481 P1_U2413 ; P1_U4619
g14582 nand P1_U4601 P1_U2412 ; P1_U4620
g14583 nand P1_U2397 P1_U4617 ; P1_U4621
g14584 nand P1_U4612 P1_INSTQUEUE_REG_14__7__SCAN_IN ; P1_U4622
g14585 nand P1_U4602 P1_U2416 ; P1_U4623
g14586 nand P1_U2481 P1_U2411 ; P1_U4624
g14587 nand P1_U4601 P1_U2410 ; P1_U4625
g14588 nand P1_U2396 P1_U4617 ; P1_U4626
g14589 nand P1_U4612 P1_INSTQUEUE_REG_14__6__SCAN_IN ; P1_U4627
g14590 nand P1_U4602 P1_U2420 ; P1_U4628
g14591 nand P1_U2481 P1_U2409 ; P1_U4629
g14592 nand P1_U4601 P1_U2408 ; P1_U4630
g14593 nand P1_U2395 P1_U4617 ; P1_U4631
g14594 nand P1_U4612 P1_INSTQUEUE_REG_14__5__SCAN_IN ; P1_U4632
g14595 nand P1_U4602 P1_U2419 ; P1_U4633
g14596 nand P1_U2481 P1_U2407 ; P1_U4634
g14597 nand P1_U4601 P1_U2406 ; P1_U4635
g14598 nand P1_U2394 P1_U4617 ; P1_U4636
g14599 nand P1_U4612 P1_INSTQUEUE_REG_14__4__SCAN_IN ; P1_U4637
g14600 nand P1_U4602 P1_U2418 ; P1_U4638
g14601 nand P1_U2481 P1_U2405 ; P1_U4639
g14602 nand P1_U4601 P1_U2404 ; P1_U4640
g14603 nand P1_U2393 P1_U4617 ; P1_U4641
g14604 nand P1_U4612 P1_INSTQUEUE_REG_14__3__SCAN_IN ; P1_U4642
g14605 nand P1_U4602 P1_U2421 ; P1_U4643
g14606 nand P1_U2481 P1_U2403 ; P1_U4644
g14607 nand P1_U4601 P1_U2402 ; P1_U4645
g14608 nand P1_U2392 P1_U4617 ; P1_U4646
g14609 nand P1_U4612 P1_INSTQUEUE_REG_14__2__SCAN_IN ; P1_U4647
g14610 nand P1_U4602 P1_U2414 ; P1_U4648
g14611 nand P1_U2481 P1_U2401 ; P1_U4649
g14612 nand P1_U4601 P1_U2400 ; P1_U4650
g14613 nand P1_U2391 P1_U4617 ; P1_U4651
g14614 nand P1_U4612 P1_INSTQUEUE_REG_14__1__SCAN_IN ; P1_U4652
g14615 nand P1_U4602 P1_U2417 ; P1_U4653
g14616 nand P1_U2481 P1_U2399 ; P1_U4654
g14617 nand P1_U4601 P1_U2398 ; P1_U4655
g14618 nand P1_U2390 P1_U4617 ; P1_U4656
g14619 nand P1_U4612 P1_INSTQUEUE_REG_14__0__SCAN_IN ; P1_U4657
g14620 not P1_U3333 ; P1_U4658
g14621 not P1_U3334 ; P1_U4659
g14622 not P1_U3330 ; P1_U4660
g14623 nand P1_U2444 P1_U2438 ; P1_U4661
g14624 not P1_U3335 ; P1_U4662
g14625 nand P1_U2437 P1_U2432 ; P1_U4663
g14626 not P1_U3336 ; P1_U4664
g14627 nand P1_U4525 P1_U2476 ; P1_U4665
g14628 nand P1_U2484 P1_U2358 ; P1_U4666
g14629 nand P1_U3320 P1_U4666 ; P1_U4667
g14630 nand P1_U4662 P1_U4667 ; P1_U4668
g14631 nand P1_U3330 P1_STATE2_REG_3__SCAN_IN ; P1_U4669
g14632 nand P1_U4664 P1_STATE2_REG_2__SCAN_IN ; P1_U4670
g14633 nand P1_U4668 P1_U3605 ; P1_U4671
g14634 nand P1_U2484 P1_U2388 ; P1_U4672
g14635 nand P1_U3320 P1_U4672 ; P1_U4673
g14636 nand P1_U4673 P1_U3335 ; P1_U4674
g14637 nand P1_U3336 P1_STATE2_REG_2__SCAN_IN ; P1_U4675
g14638 nand P1_U4675 P1_U4674 ; P1_U4676
g14639 nand P1_U4660 P1_U2415 ; P1_U4677
g14640 nand P1_U2483 P1_U2413 ; P1_U4678
g14641 nand P1_U4659 P1_U2412 ; P1_U4679
g14642 nand P1_U2397 P1_U4676 ; P1_U4680
g14643 nand P1_U4671 P1_INSTQUEUE_REG_13__7__SCAN_IN ; P1_U4681
g14644 nand P1_U4660 P1_U2416 ; P1_U4682
g14645 nand P1_U2483 P1_U2411 ; P1_U4683
g14646 nand P1_U4659 P1_U2410 ; P1_U4684
g14647 nand P1_U2396 P1_U4676 ; P1_U4685
g14648 nand P1_U4671 P1_INSTQUEUE_REG_13__6__SCAN_IN ; P1_U4686
g14649 nand P1_U4660 P1_U2420 ; P1_U4687
g14650 nand P1_U2483 P1_U2409 ; P1_U4688
g14651 nand P1_U4659 P1_U2408 ; P1_U4689
g14652 nand P1_U2395 P1_U4676 ; P1_U4690
g14653 nand P1_U4671 P1_INSTQUEUE_REG_13__5__SCAN_IN ; P1_U4691
g14654 nand P1_U4660 P1_U2419 ; P1_U4692
g14655 nand P1_U2483 P1_U2407 ; P1_U4693
g14656 nand P1_U4659 P1_U2406 ; P1_U4694
g14657 nand P1_U2394 P1_U4676 ; P1_U4695
g14658 nand P1_U4671 P1_INSTQUEUE_REG_13__4__SCAN_IN ; P1_U4696
g14659 nand P1_U4660 P1_U2418 ; P1_U4697
g14660 nand P1_U2483 P1_U2405 ; P1_U4698
g14661 nand P1_U4659 P1_U2404 ; P1_U4699
g14662 nand P1_U2393 P1_U4676 ; P1_U4700
g14663 nand P1_U4671 P1_INSTQUEUE_REG_13__3__SCAN_IN ; P1_U4701
g14664 nand P1_U4660 P1_U2421 ; P1_U4702
g14665 nand P1_U2483 P1_U2403 ; P1_U4703
g14666 nand P1_U4659 P1_U2402 ; P1_U4704
g14667 nand P1_U2392 P1_U4676 ; P1_U4705
g14668 nand P1_U4671 P1_INSTQUEUE_REG_13__2__SCAN_IN ; P1_U4706
g14669 nand P1_U4660 P1_U2414 ; P1_U4707
g14670 nand P1_U2483 P1_U2401 ; P1_U4708
g14671 nand P1_U4659 P1_U2400 ; P1_U4709
g14672 nand P1_U2391 P1_U4676 ; P1_U4710
g14673 nand P1_U4671 P1_INSTQUEUE_REG_13__1__SCAN_IN ; P1_U4711
g14674 nand P1_U4660 P1_U2417 ; P1_U4712
g14675 nand P1_U2483 P1_U2399 ; P1_U4713
g14676 nand P1_U4659 P1_U2398 ; P1_U4714
g14677 nand P1_U2390 P1_U4676 ; P1_U4715
g14678 nand P1_U4671 P1_INSTQUEUE_REG_13__0__SCAN_IN ; P1_U4716
g14679 not P1_U3338 ; P1_U4717
g14680 not P1_U3337 ; P1_U4718
g14681 nand P1_U2445 P1_U2438 ; P1_U4719
g14682 not P1_U3339 ; P1_U4720
g14683 not P1_U3237 ; P1_U4721
g14684 nand P1_U2486 P1_U2476 ; P1_U4722
g14685 nand P1_U2489 P1_U2358 ; P1_U4723
g14686 nand P1_U3320 P1_U4723 ; P1_U4724
g14687 nand P1_U4720 P1_U4724 ; P1_U4725
g14688 nand P1_U3337 P1_STATE2_REG_3__SCAN_IN ; P1_U4726
g14689 nand P1_U3237 P1_STATE2_REG_2__SCAN_IN ; P1_U4727
g14690 nand P1_U4725 P1_U3614 ; P1_U4728
g14691 nand P1_U2489 P1_U2388 ; P1_U4729
g14692 nand P1_U3320 P1_U4729 ; P1_U4730
g14693 nand P1_U4730 P1_U3339 ; P1_U4731
g14694 nand P1_U4721 P1_STATE2_REG_2__SCAN_IN ; P1_U4732
g14695 nand P1_U4732 P1_U4731 ; P1_U4733
g14696 nand P1_U4718 P1_U2415 ; P1_U4734
g14697 nand P1_U2487 P1_U2413 ; P1_U4735
g14698 nand P1_U4717 P1_U2412 ; P1_U4736
g14699 nand P1_U2397 P1_U4733 ; P1_U4737
g14700 nand P1_U4728 P1_INSTQUEUE_REG_12__7__SCAN_IN ; P1_U4738
g14701 nand P1_U4718 P1_U2416 ; P1_U4739
g14702 nand P1_U2487 P1_U2411 ; P1_U4740
g14703 nand P1_U4717 P1_U2410 ; P1_U4741
g14704 nand P1_U2396 P1_U4733 ; P1_U4742
g14705 nand P1_U4728 P1_INSTQUEUE_REG_12__6__SCAN_IN ; P1_U4743
g14706 nand P1_U4718 P1_U2420 ; P1_U4744
g14707 nand P1_U2487 P1_U2409 ; P1_U4745
g14708 nand P1_U4717 P1_U2408 ; P1_U4746
g14709 nand P1_U2395 P1_U4733 ; P1_U4747
g14710 nand P1_U4728 P1_INSTQUEUE_REG_12__5__SCAN_IN ; P1_U4748
g14711 nand P1_U4718 P1_U2419 ; P1_U4749
g14712 nand P1_U2487 P1_U2407 ; P1_U4750
g14713 nand P1_U4717 P1_U2406 ; P1_U4751
g14714 nand P1_U2394 P1_U4733 ; P1_U4752
g14715 nand P1_U4728 P1_INSTQUEUE_REG_12__4__SCAN_IN ; P1_U4753
g14716 nand P1_U4718 P1_U2418 ; P1_U4754
g14717 nand P1_U2487 P1_U2405 ; P1_U4755
g14718 nand P1_U4717 P1_U2404 ; P1_U4756
g14719 nand P1_U2393 P1_U4733 ; P1_U4757
g14720 nand P1_U4728 P1_INSTQUEUE_REG_12__3__SCAN_IN ; P1_U4758
g14721 nand P1_U4718 P1_U2421 ; P1_U4759
g14722 nand P1_U2487 P1_U2403 ; P1_U4760
g14723 nand P1_U4717 P1_U2402 ; P1_U4761
g14724 nand P1_U2392 P1_U4733 ; P1_U4762
g14725 nand P1_U4728 P1_INSTQUEUE_REG_12__2__SCAN_IN ; P1_U4763
g14726 nand P1_U4718 P1_U2414 ; P1_U4764
g14727 nand P1_U2487 P1_U2401 ; P1_U4765
g14728 nand P1_U4717 P1_U2400 ; P1_U4766
g14729 nand P1_U2391 P1_U4733 ; P1_U4767
g14730 nand P1_U4728 P1_INSTQUEUE_REG_12__1__SCAN_IN ; P1_U4768
g14731 nand P1_U4718 P1_U2417 ; P1_U4769
g14732 nand P1_U2487 P1_U2399 ; P1_U4770
g14733 nand P1_U4717 P1_U2398 ; P1_U4771
g14734 nand P1_U2390 P1_U4733 ; P1_U4772
g14735 nand P1_U4728 P1_INSTQUEUE_REG_12__0__SCAN_IN ; P1_U4773
g14736 not P1_U3343 ; P1_U4774
g14737 not P1_U3341 ; P1_U4775
g14738 nand P1_U2440 P1_U2442 ; P1_U4776
g14739 not P1_U3344 ; P1_U4777
g14740 nand P1_U2434 P1_U2436 ; P1_U4778
g14741 not P1_U3345 ; P1_U4779
g14742 nand P1_U4529 P1_U4528 ; P1_U4780
g14743 nand P1_U2492 P1_U2358 ; P1_U4781
g14744 nand P1_U3320 P1_U4781 ; P1_U4782
g14745 nand P1_U4777 P1_U4782 ; P1_U4783
g14746 nand P1_U3341 P1_STATE2_REG_3__SCAN_IN ; P1_U4784
g14747 nand P1_U4779 P1_STATE2_REG_2__SCAN_IN ; P1_U4785
g14748 nand P1_U4783 P1_U3623 ; P1_U4786
g14749 nand P1_U2492 P1_U2388 ; P1_U4787
g14750 nand P1_U3320 P1_U4787 ; P1_U4788
g14751 nand P1_U4788 P1_U3344 ; P1_U4789
g14752 nand P1_U3345 P1_STATE2_REG_2__SCAN_IN ; P1_U4790
g14753 nand P1_U4790 P1_U4789 ; P1_U4791
g14754 nand P1_U4775 P1_U2415 ; P1_U4792
g14755 nand P1_U2491 P1_U2413 ; P1_U4793
g14756 nand P1_U4774 P1_U2412 ; P1_U4794
g14757 nand P1_U2397 P1_U4791 ; P1_U4795
g14758 nand P1_U4786 P1_INSTQUEUE_REG_11__7__SCAN_IN ; P1_U4796
g14759 nand P1_U4775 P1_U2416 ; P1_U4797
g14760 nand P1_U2491 P1_U2411 ; P1_U4798
g14761 nand P1_U4774 P1_U2410 ; P1_U4799
g14762 nand P1_U2396 P1_U4791 ; P1_U4800
g14763 nand P1_U4786 P1_INSTQUEUE_REG_11__6__SCAN_IN ; P1_U4801
g14764 nand P1_U4775 P1_U2420 ; P1_U4802
g14765 nand P1_U2491 P1_U2409 ; P1_U4803
g14766 nand P1_U4774 P1_U2408 ; P1_U4804
g14767 nand P1_U2395 P1_U4791 ; P1_U4805
g14768 nand P1_U4786 P1_INSTQUEUE_REG_11__5__SCAN_IN ; P1_U4806
g14769 nand P1_U4775 P1_U2419 ; P1_U4807
g14770 nand P1_U2491 P1_U2407 ; P1_U4808
g14771 nand P1_U4774 P1_U2406 ; P1_U4809
g14772 nand P1_U2394 P1_U4791 ; P1_U4810
g14773 nand P1_U4786 P1_INSTQUEUE_REG_11__4__SCAN_IN ; P1_U4811
g14774 nand P1_U4775 P1_U2418 ; P1_U4812
g14775 nand P1_U2491 P1_U2405 ; P1_U4813
g14776 nand P1_U4774 P1_U2404 ; P1_U4814
g14777 nand P1_U2393 P1_U4791 ; P1_U4815
g14778 nand P1_U4786 P1_INSTQUEUE_REG_11__3__SCAN_IN ; P1_U4816
g14779 nand P1_U4775 P1_U2421 ; P1_U4817
g14780 nand P1_U2491 P1_U2403 ; P1_U4818
g14781 nand P1_U4774 P1_U2402 ; P1_U4819
g14782 nand P1_U2392 P1_U4791 ; P1_U4820
g14783 nand P1_U4786 P1_INSTQUEUE_REG_11__2__SCAN_IN ; P1_U4821
g14784 nand P1_U4775 P1_U2414 ; P1_U4822
g14785 nand P1_U2491 P1_U2401 ; P1_U4823
g14786 nand P1_U4774 P1_U2400 ; P1_U4824
g14787 nand P1_U2391 P1_U4791 ; P1_U4825
g14788 nand P1_U4786 P1_INSTQUEUE_REG_11__1__SCAN_IN ; P1_U4826
g14789 nand P1_U4775 P1_U2417 ; P1_U4827
g14790 nand P1_U2491 P1_U2399 ; P1_U4828
g14791 nand P1_U4774 P1_U2398 ; P1_U4829
g14792 nand P1_U2390 P1_U4791 ; P1_U4830
g14793 nand P1_U4786 P1_INSTQUEUE_REG_11__0__SCAN_IN ; P1_U4831
g14794 not P1_U3347 ; P1_U4832
g14795 not P1_U3346 ; P1_U4833
g14796 nand P1_U2440 P1_U2443 ; P1_U4834
g14797 not P1_U3348 ; P1_U4835
g14798 not P1_U3238 ; P1_U4836
g14799 nand P1_U4529 P1_U4524 ; P1_U4837
g14800 nand P1_U2494 P1_U2358 ; P1_U4838
g14801 nand P1_U3320 P1_U4838 ; P1_U4839
g14802 nand P1_U4835 P1_U4839 ; P1_U4840
g14803 nand P1_U3346 P1_STATE2_REG_3__SCAN_IN ; P1_U4841
g14804 nand P1_U3238 P1_STATE2_REG_2__SCAN_IN ; P1_U4842
g14805 nand P1_U4840 P1_U3632 ; P1_U4843
g14806 nand P1_U2494 P1_U2388 ; P1_U4844
g14807 nand P1_U3320 P1_U4844 ; P1_U4845
g14808 nand P1_U4845 P1_U3348 ; P1_U4846
g14809 nand P1_U4836 P1_STATE2_REG_2__SCAN_IN ; P1_U4847
g14810 nand P1_U4847 P1_U4846 ; P1_U4848
g14811 nand P1_U4833 P1_U2415 ; P1_U4849
g14812 nand P1_U2493 P1_U2413 ; P1_U4850
g14813 nand P1_U4832 P1_U2412 ; P1_U4851
g14814 nand P1_U2397 P1_U4848 ; P1_U4852
g14815 nand P1_U4843 P1_INSTQUEUE_REG_10__7__SCAN_IN ; P1_U4853
g14816 nand P1_U4833 P1_U2416 ; P1_U4854
g14817 nand P1_U2493 P1_U2411 ; P1_U4855
g14818 nand P1_U4832 P1_U2410 ; P1_U4856
g14819 nand P1_U2396 P1_U4848 ; P1_U4857
g14820 nand P1_U4843 P1_INSTQUEUE_REG_10__6__SCAN_IN ; P1_U4858
g14821 nand P1_U4833 P1_U2420 ; P1_U4859
g14822 nand P1_U2493 P1_U2409 ; P1_U4860
g14823 nand P1_U4832 P1_U2408 ; P1_U4861
g14824 nand P1_U2395 P1_U4848 ; P1_U4862
g14825 nand P1_U4843 P1_INSTQUEUE_REG_10__5__SCAN_IN ; P1_U4863
g14826 nand P1_U4833 P1_U2419 ; P1_U4864
g14827 nand P1_U2493 P1_U2407 ; P1_U4865
g14828 nand P1_U4832 P1_U2406 ; P1_U4866
g14829 nand P1_U2394 P1_U4848 ; P1_U4867
g14830 nand P1_U4843 P1_INSTQUEUE_REG_10__4__SCAN_IN ; P1_U4868
g14831 nand P1_U4833 P1_U2418 ; P1_U4869
g14832 nand P1_U2493 P1_U2405 ; P1_U4870
g14833 nand P1_U4832 P1_U2404 ; P1_U4871
g14834 nand P1_U2393 P1_U4848 ; P1_U4872
g14835 nand P1_U4843 P1_INSTQUEUE_REG_10__3__SCAN_IN ; P1_U4873
g14836 nand P1_U4833 P1_U2421 ; P1_U4874
g14837 nand P1_U2493 P1_U2403 ; P1_U4875
g14838 nand P1_U4832 P1_U2402 ; P1_U4876
g14839 nand P1_U2392 P1_U4848 ; P1_U4877
g14840 nand P1_U4843 P1_INSTQUEUE_REG_10__2__SCAN_IN ; P1_U4878
g14841 nand P1_U4833 P1_U2414 ; P1_U4879
g14842 nand P1_U2493 P1_U2401 ; P1_U4880
g14843 nand P1_U4832 P1_U2400 ; P1_U4881
g14844 nand P1_U2391 P1_U4848 ; P1_U4882
g14845 nand P1_U4843 P1_INSTQUEUE_REG_10__1__SCAN_IN ; P1_U4883
g14846 nand P1_U4833 P1_U2417 ; P1_U4884
g14847 nand P1_U2493 P1_U2399 ; P1_U4885
g14848 nand P1_U4832 P1_U2398 ; P1_U4886
g14849 nand P1_U2390 P1_U4848 ; P1_U4887
g14850 nand P1_U4843 P1_INSTQUEUE_REG_10__0__SCAN_IN ; P1_U4888
g14851 not P1_U3350 ; P1_U4889
g14852 not P1_U3349 ; P1_U4890
g14853 nand P1_U2440 P1_U2444 ; P1_U4891
g14854 not P1_U3351 ; P1_U4892
g14855 nand P1_U2434 P1_U2437 ; P1_U4893
g14856 not P1_U3352 ; P1_U4894
g14857 nand P1_U4529 P1_U4525 ; P1_U4895
g14858 nand P1_U2496 P1_U2358 ; P1_U4896
g14859 nand P1_U3320 P1_U4896 ; P1_U4897
g14860 nand P1_U4892 P1_U4897 ; P1_U4898
g14861 nand P1_U3349 P1_STATE2_REG_3__SCAN_IN ; P1_U4899
g14862 nand P1_U4894 P1_STATE2_REG_2__SCAN_IN ; P1_U4900
g14863 nand P1_U4898 P1_U3641 ; P1_U4901
g14864 nand P1_U2496 P1_U2388 ; P1_U4902
g14865 nand P1_U3320 P1_U4902 ; P1_U4903
g14866 nand P1_U4903 P1_U3351 ; P1_U4904
g14867 nand P1_U3352 P1_STATE2_REG_2__SCAN_IN ; P1_U4905
g14868 nand P1_U4905 P1_U4904 ; P1_U4906
g14869 nand P1_U4890 P1_U2415 ; P1_U4907
g14870 nand P1_U2495 P1_U2413 ; P1_U4908
g14871 nand P1_U4889 P1_U2412 ; P1_U4909
g14872 nand P1_U2397 P1_U4906 ; P1_U4910
g14873 nand P1_U4901 P1_INSTQUEUE_REG_9__7__SCAN_IN ; P1_U4911
g14874 nand P1_U4890 P1_U2416 ; P1_U4912
g14875 nand P1_U2495 P1_U2411 ; P1_U4913
g14876 nand P1_U4889 P1_U2410 ; P1_U4914
g14877 nand P1_U2396 P1_U4906 ; P1_U4915
g14878 nand P1_U4901 P1_INSTQUEUE_REG_9__6__SCAN_IN ; P1_U4916
g14879 nand P1_U4890 P1_U2420 ; P1_U4917
g14880 nand P1_U2495 P1_U2409 ; P1_U4918
g14881 nand P1_U4889 P1_U2408 ; P1_U4919
g14882 nand P1_U2395 P1_U4906 ; P1_U4920
g14883 nand P1_U4901 P1_INSTQUEUE_REG_9__5__SCAN_IN ; P1_U4921
g14884 nand P1_U4890 P1_U2419 ; P1_U4922
g14885 nand P1_U2495 P1_U2407 ; P1_U4923
g14886 nand P1_U4889 P1_U2406 ; P1_U4924
g14887 nand P1_U2394 P1_U4906 ; P1_U4925
g14888 nand P1_U4901 P1_INSTQUEUE_REG_9__4__SCAN_IN ; P1_U4926
g14889 nand P1_U4890 P1_U2418 ; P1_U4927
g14890 nand P1_U2495 P1_U2405 ; P1_U4928
g14891 nand P1_U4889 P1_U2404 ; P1_U4929
g14892 nand P1_U2393 P1_U4906 ; P1_U4930
g14893 nand P1_U4901 P1_INSTQUEUE_REG_9__3__SCAN_IN ; P1_U4931
g14894 nand P1_U4890 P1_U2421 ; P1_U4932
g14895 nand P1_U2495 P1_U2403 ; P1_U4933
g14896 nand P1_U4889 P1_U2402 ; P1_U4934
g14897 nand P1_U2392 P1_U4906 ; P1_U4935
g14898 nand P1_U4901 P1_INSTQUEUE_REG_9__2__SCAN_IN ; P1_U4936
g14899 nand P1_U4890 P1_U2414 ; P1_U4937
g14900 nand P1_U2495 P1_U2401 ; P1_U4938
g14901 nand P1_U4889 P1_U2400 ; P1_U4939
g14902 nand P1_U2391 P1_U4906 ; P1_U4940
g14903 nand P1_U4901 P1_INSTQUEUE_REG_9__1__SCAN_IN ; P1_U4941
g14904 nand P1_U4890 P1_U2417 ; P1_U4942
g14905 nand P1_U2495 P1_U2399 ; P1_U4943
g14906 nand P1_U4889 P1_U2398 ; P1_U4944
g14907 nand P1_U2390 P1_U4906 ; P1_U4945
g14908 nand P1_U4901 P1_INSTQUEUE_REG_9__0__SCAN_IN ; P1_U4946
g14909 not P1_U3354 ; P1_U4947
g14910 not P1_U3353 ; P1_U4948
g14911 nand P1_U2440 P1_U2445 ; P1_U4949
g14912 not P1_U3355 ; P1_U4950
g14913 not P1_U3239 ; P1_U4951
g14914 nand P1_U4529 P1_U2486 ; P1_U4952
g14915 nand P1_U2498 P1_U2358 ; P1_U4953
g14916 nand P1_U3320 P1_U4953 ; P1_U4954
g14917 nand P1_U4950 P1_U4954 ; P1_U4955
g14918 nand P1_U3353 P1_STATE2_REG_3__SCAN_IN ; P1_U4956
g14919 nand P1_U3239 P1_STATE2_REG_2__SCAN_IN ; P1_U4957
g14920 nand P1_U4955 P1_U3650 ; P1_U4958
g14921 nand P1_U2498 P1_U2388 ; P1_U4959
g14922 nand P1_U3320 P1_U4959 ; P1_U4960
g14923 nand P1_U4960 P1_U3355 ; P1_U4961
g14924 nand P1_U4951 P1_STATE2_REG_2__SCAN_IN ; P1_U4962
g14925 nand P1_U4962 P1_U4961 ; P1_U4963
g14926 nand P1_U4948 P1_U2415 ; P1_U4964
g14927 nand P1_U2497 P1_U2413 ; P1_U4965
g14928 nand P1_U4947 P1_U2412 ; P1_U4966
g14929 nand P1_U2397 P1_U4963 ; P1_U4967
g14930 nand P1_U4958 P1_INSTQUEUE_REG_8__7__SCAN_IN ; P1_U4968
g14931 nand P1_U4948 P1_U2416 ; P1_U4969
g14932 nand P1_U2497 P1_U2411 ; P1_U4970
g14933 nand P1_U4947 P1_U2410 ; P1_U4971
g14934 nand P1_U2396 P1_U4963 ; P1_U4972
g14935 nand P1_U4958 P1_INSTQUEUE_REG_8__6__SCAN_IN ; P1_U4973
g14936 nand P1_U4948 P1_U2420 ; P1_U4974
g14937 nand P1_U2497 P1_U2409 ; P1_U4975
g14938 nand P1_U4947 P1_U2408 ; P1_U4976
g14939 nand P1_U2395 P1_U4963 ; P1_U4977
g14940 nand P1_U4958 P1_INSTQUEUE_REG_8__5__SCAN_IN ; P1_U4978
g14941 nand P1_U4948 P1_U2419 ; P1_U4979
g14942 nand P1_U2497 P1_U2407 ; P1_U4980
g14943 nand P1_U4947 P1_U2406 ; P1_U4981
g14944 nand P1_U2394 P1_U4963 ; P1_U4982
g14945 nand P1_U4958 P1_INSTQUEUE_REG_8__4__SCAN_IN ; P1_U4983
g14946 nand P1_U4948 P1_U2418 ; P1_U4984
g14947 nand P1_U2497 P1_U2405 ; P1_U4985
g14948 nand P1_U4947 P1_U2404 ; P1_U4986
g14949 nand P1_U2393 P1_U4963 ; P1_U4987
g14950 nand P1_U4958 P1_INSTQUEUE_REG_8__3__SCAN_IN ; P1_U4988
g14951 nand P1_U4948 P1_U2421 ; P1_U4989
g14952 nand P1_U2497 P1_U2403 ; P1_U4990
g14953 nand P1_U4947 P1_U2402 ; P1_U4991
g14954 nand P1_U2392 P1_U4963 ; P1_U4992
g14955 nand P1_U4958 P1_INSTQUEUE_REG_8__2__SCAN_IN ; P1_U4993
g14956 nand P1_U4948 P1_U2414 ; P1_U4994
g14957 nand P1_U2497 P1_U2401 ; P1_U4995
g14958 nand P1_U4947 P1_U2400 ; P1_U4996
g14959 nand P1_U2391 P1_U4963 ; P1_U4997
g14960 nand P1_U4958 P1_INSTQUEUE_REG_8__1__SCAN_IN ; P1_U4998
g14961 nand P1_U4948 P1_U2417 ; P1_U4999
g14962 nand P1_U2497 P1_U2399 ; P1_U5000
g14963 nand P1_U4947 P1_U2398 ; P1_U5001
g14964 nand P1_U2390 P1_U4963 ; P1_U5002
g14965 nand P1_U4958 P1_INSTQUEUE_REG_8__0__SCAN_IN ; P1_U5003
g14966 not P1_U3359 ; P1_U5004
g14967 nand P1_U2439 P1_U2442 ; P1_U5005
g14968 not P1_U3361 ; P1_U5006
g14969 nand P1_U2433 P1_U2436 ; P1_U5007
g14970 not P1_U3362 ; P1_U5008
g14971 nand P1_U2500 P1_U2358 ; P1_U5009
g14972 nand P1_U3320 P1_U5009 ; P1_U5010
g14973 nand P1_U5006 P1_U5010 ; P1_U5011
g14974 nand P1_U3356 P1_STATE2_REG_3__SCAN_IN ; P1_U5012
g14975 nand P1_U5008 P1_STATE2_REG_2__SCAN_IN ; P1_U5013
g14976 nand P1_U5011 P1_U3659 ; P1_U5014
g14977 nand P1_U2500 P1_U2388 ; P1_U5015
g14978 nand P1_U3320 P1_U5015 ; P1_U5016
g14979 nand P1_U5016 P1_U3361 ; P1_U5017
g14980 nand P1_U3362 P1_STATE2_REG_2__SCAN_IN ; P1_U5018
g14981 nand P1_U5018 P1_U5017 ; P1_U5019
g14982 nand P1_U4537 P1_U2415 ; P1_U5020
g14983 nand P1_U4238 P1_U2413 ; P1_U5021
g14984 nand P1_U5004 P1_U2412 ; P1_U5022
g14985 nand P1_U2397 P1_U5019 ; P1_U5023
g14986 nand P1_U5014 P1_INSTQUEUE_REG_7__7__SCAN_IN ; P1_U5024
g14987 nand P1_U4537 P1_U2416 ; P1_U5025
g14988 nand P1_U4238 P1_U2411 ; P1_U5026
g14989 nand P1_U5004 P1_U2410 ; P1_U5027
g14990 nand P1_U2396 P1_U5019 ; P1_U5028
g14991 nand P1_U5014 P1_INSTQUEUE_REG_7__6__SCAN_IN ; P1_U5029
g14992 nand P1_U4537 P1_U2420 ; P1_U5030
g14993 nand P1_U4238 P1_U2409 ; P1_U5031
g14994 nand P1_U5004 P1_U2408 ; P1_U5032
g14995 nand P1_U2395 P1_U5019 ; P1_U5033
g14996 nand P1_U5014 P1_INSTQUEUE_REG_7__5__SCAN_IN ; P1_U5034
g14997 nand P1_U4537 P1_U2419 ; P1_U5035
g14998 nand P1_U4238 P1_U2407 ; P1_U5036
g14999 nand P1_U5004 P1_U2406 ; P1_U5037
g15000 nand P1_U2394 P1_U5019 ; P1_U5038
g15001 nand P1_U5014 P1_INSTQUEUE_REG_7__4__SCAN_IN ; P1_U5039
g15002 nand P1_U4537 P1_U2418 ; P1_U5040
g15003 nand P1_U4238 P1_U2405 ; P1_U5041
g15004 nand P1_U5004 P1_U2404 ; P1_U5042
g15005 nand P1_U2393 P1_U5019 ; P1_U5043
g15006 nand P1_U5014 P1_INSTQUEUE_REG_7__3__SCAN_IN ; P1_U5044
g15007 nand P1_U4537 P1_U2421 ; P1_U5045
g15008 nand P1_U4238 P1_U2403 ; P1_U5046
g15009 nand P1_U5004 P1_U2402 ; P1_U5047
g15010 nand P1_U2392 P1_U5019 ; P1_U5048
g15011 nand P1_U5014 P1_INSTQUEUE_REG_7__2__SCAN_IN ; P1_U5049
g15012 nand P1_U4537 P1_U2414 ; P1_U5050
g15013 nand P1_U4238 P1_U2401 ; P1_U5051
g15014 nand P1_U5004 P1_U2400 ; P1_U5052
g15015 nand P1_U2391 P1_U5019 ; P1_U5053
g15016 nand P1_U5014 P1_INSTQUEUE_REG_7__1__SCAN_IN ; P1_U5054
g15017 nand P1_U4537 P1_U2417 ; P1_U5055
g15018 nand P1_U4238 P1_U2399 ; P1_U5056
g15019 nand P1_U5004 P1_U2398 ; P1_U5057
g15020 nand P1_U2390 P1_U5019 ; P1_U5058
g15021 nand P1_U5014 P1_INSTQUEUE_REG_7__0__SCAN_IN ; P1_U5059
g15022 not P1_U3364 ; P1_U5060
g15023 not P1_U3363 ; P1_U5061
g15024 nand P1_U2439 P1_U2443 ; P1_U5062
g15025 not P1_U3365 ; P1_U5063
g15026 not P1_U3240 ; P1_U5064
g15027 nand P1_U4524 P1_U2474 ; P1_U5065
g15028 nand P1_U2502 P1_U2358 ; P1_U5066
g15029 nand P1_U3320 P1_U5066 ; P1_U5067
g15030 nand P1_U5063 P1_U5067 ; P1_U5068
g15031 nand P1_U3363 P1_STATE2_REG_3__SCAN_IN ; P1_U5069
g15032 nand P1_U3240 P1_STATE2_REG_2__SCAN_IN ; P1_U5070
g15033 nand P1_U5068 P1_U3668 ; P1_U5071
g15034 nand P1_U2502 P1_U2388 ; P1_U5072
g15035 nand P1_U3320 P1_U5072 ; P1_U5073
g15036 nand P1_U5073 P1_U3365 ; P1_U5074
g15037 nand P1_U5064 P1_STATE2_REG_2__SCAN_IN ; P1_U5075
g15038 nand P1_U5075 P1_U5074 ; P1_U5076
g15039 nand P1_U5061 P1_U2415 ; P1_U5077
g15040 nand P1_U2501 P1_U2413 ; P1_U5078
g15041 nand P1_U5060 P1_U2412 ; P1_U5079
g15042 nand P1_U2397 P1_U5076 ; P1_U5080
g15043 nand P1_U5071 P1_INSTQUEUE_REG_6__7__SCAN_IN ; P1_U5081
g15044 nand P1_U5061 P1_U2416 ; P1_U5082
g15045 nand P1_U2501 P1_U2411 ; P1_U5083
g15046 nand P1_U5060 P1_U2410 ; P1_U5084
g15047 nand P1_U2396 P1_U5076 ; P1_U5085
g15048 nand P1_U5071 P1_INSTQUEUE_REG_6__6__SCAN_IN ; P1_U5086
g15049 nand P1_U5061 P1_U2420 ; P1_U5087
g15050 nand P1_U2501 P1_U2409 ; P1_U5088
g15051 nand P1_U5060 P1_U2408 ; P1_U5089
g15052 nand P1_U2395 P1_U5076 ; P1_U5090
g15053 nand P1_U5071 P1_INSTQUEUE_REG_6__5__SCAN_IN ; P1_U5091
g15054 nand P1_U5061 P1_U2419 ; P1_U5092
g15055 nand P1_U2501 P1_U2407 ; P1_U5093
g15056 nand P1_U5060 P1_U2406 ; P1_U5094
g15057 nand P1_U2394 P1_U5076 ; P1_U5095
g15058 nand P1_U5071 P1_INSTQUEUE_REG_6__4__SCAN_IN ; P1_U5096
g15059 nand P1_U5061 P1_U2418 ; P1_U5097
g15060 nand P1_U2501 P1_U2405 ; P1_U5098
g15061 nand P1_U5060 P1_U2404 ; P1_U5099
g15062 nand P1_U2393 P1_U5076 ; P1_U5100
g15063 nand P1_U5071 P1_INSTQUEUE_REG_6__3__SCAN_IN ; P1_U5101
g15064 nand P1_U5061 P1_U2421 ; P1_U5102
g15065 nand P1_U2501 P1_U2403 ; P1_U5103
g15066 nand P1_U5060 P1_U2402 ; P1_U5104
g15067 nand P1_U2392 P1_U5076 ; P1_U5105
g15068 nand P1_U5071 P1_INSTQUEUE_REG_6__2__SCAN_IN ; P1_U5106
g15069 nand P1_U5061 P1_U2414 ; P1_U5107
g15070 nand P1_U2501 P1_U2401 ; P1_U5108
g15071 nand P1_U5060 P1_U2400 ; P1_U5109
g15072 nand P1_U2391 P1_U5076 ; P1_U5110
g15073 nand P1_U5071 P1_INSTQUEUE_REG_6__1__SCAN_IN ; P1_U5111
g15074 nand P1_U5061 P1_U2417 ; P1_U5112
g15075 nand P1_U2501 P1_U2399 ; P1_U5113
g15076 nand P1_U5060 P1_U2398 ; P1_U5114
g15077 nand P1_U2390 P1_U5076 ; P1_U5115
g15078 nand P1_U5071 P1_INSTQUEUE_REG_6__0__SCAN_IN ; P1_U5116
g15079 not P1_U3367 ; P1_U5117
g15080 not P1_U3366 ; P1_U5118
g15081 nand P1_U2439 P1_U2444 ; P1_U5119
g15082 not P1_U3368 ; P1_U5120
g15083 nand P1_U2433 P1_U2437 ; P1_U5121
g15084 not P1_U3369 ; P1_U5122
g15085 nand P1_U4525 P1_U2474 ; P1_U5123
g15086 nand P1_U2504 P1_U2358 ; P1_U5124
g15087 nand P1_U3320 P1_U5124 ; P1_U5125
g15088 nand P1_U5120 P1_U5125 ; P1_U5126
g15089 nand P1_U3366 P1_STATE2_REG_3__SCAN_IN ; P1_U5127
g15090 nand P1_U5122 P1_STATE2_REG_2__SCAN_IN ; P1_U5128
g15091 nand P1_U5126 P1_U3677 ; P1_U5129
g15092 nand P1_U2504 P1_U2388 ; P1_U5130
g15093 nand P1_U3320 P1_U5130 ; P1_U5131
g15094 nand P1_U5131 P1_U3368 ; P1_U5132
g15095 nand P1_U3369 P1_STATE2_REG_2__SCAN_IN ; P1_U5133
g15096 nand P1_U5133 P1_U5132 ; P1_U5134
g15097 nand P1_U5118 P1_U2415 ; P1_U5135
g15098 nand P1_U2503 P1_U2413 ; P1_U5136
g15099 nand P1_U5117 P1_U2412 ; P1_U5137
g15100 nand P1_U2397 P1_U5134 ; P1_U5138
g15101 nand P1_U5129 P1_INSTQUEUE_REG_5__7__SCAN_IN ; P1_U5139
g15102 nand P1_U5118 P1_U2416 ; P1_U5140
g15103 nand P1_U2503 P1_U2411 ; P1_U5141
g15104 nand P1_U5117 P1_U2410 ; P1_U5142
g15105 nand P1_U2396 P1_U5134 ; P1_U5143
g15106 nand P1_U5129 P1_INSTQUEUE_REG_5__6__SCAN_IN ; P1_U5144
g15107 nand P1_U5118 P1_U2420 ; P1_U5145
g15108 nand P1_U2503 P1_U2409 ; P1_U5146
g15109 nand P1_U5117 P1_U2408 ; P1_U5147
g15110 nand P1_U2395 P1_U5134 ; P1_U5148
g15111 nand P1_U5129 P1_INSTQUEUE_REG_5__5__SCAN_IN ; P1_U5149
g15112 nand P1_U5118 P1_U2419 ; P1_U5150
g15113 nand P1_U2503 P1_U2407 ; P1_U5151
g15114 nand P1_U5117 P1_U2406 ; P1_U5152
g15115 nand P1_U2394 P1_U5134 ; P1_U5153
g15116 nand P1_U5129 P1_INSTQUEUE_REG_5__4__SCAN_IN ; P1_U5154
g15117 nand P1_U5118 P1_U2418 ; P1_U5155
g15118 nand P1_U2503 P1_U2405 ; P1_U5156
g15119 nand P1_U5117 P1_U2404 ; P1_U5157
g15120 nand P1_U2393 P1_U5134 ; P1_U5158
g15121 nand P1_U5129 P1_INSTQUEUE_REG_5__3__SCAN_IN ; P1_U5159
g15122 nand P1_U5118 P1_U2421 ; P1_U5160
g15123 nand P1_U2503 P1_U2403 ; P1_U5161
g15124 nand P1_U5117 P1_U2402 ; P1_U5162
g15125 nand P1_U2392 P1_U5134 ; P1_U5163
g15126 nand P1_U5129 P1_INSTQUEUE_REG_5__2__SCAN_IN ; P1_U5164
g15127 nand P1_U5118 P1_U2414 ; P1_U5165
g15128 nand P1_U2503 P1_U2401 ; P1_U5166
g15129 nand P1_U5117 P1_U2400 ; P1_U5167
g15130 nand P1_U2391 P1_U5134 ; P1_U5168
g15131 nand P1_U5129 P1_INSTQUEUE_REG_5__1__SCAN_IN ; P1_U5169
g15132 nand P1_U5118 P1_U2417 ; P1_U5170
g15133 nand P1_U2503 P1_U2399 ; P1_U5171
g15134 nand P1_U5117 P1_U2398 ; P1_U5172
g15135 nand P1_U2390 P1_U5134 ; P1_U5173
g15136 nand P1_U5129 P1_INSTQUEUE_REG_5__0__SCAN_IN ; P1_U5174
g15137 not P1_U3371 ; P1_U5175
g15138 not P1_U3370 ; P1_U5176
g15139 nand P1_U2439 P1_U2445 ; P1_U5177
g15140 not P1_U3372 ; P1_U5178
g15141 not P1_U3241 ; P1_U5179
g15142 nand P1_U2486 P1_U2474 ; P1_U5180
g15143 nand P1_U2506 P1_U2358 ; P1_U5181
g15144 nand P1_U3320 P1_U5181 ; P1_U5182
g15145 nand P1_U5178 P1_U5182 ; P1_U5183
g15146 nand P1_U3370 P1_STATE2_REG_3__SCAN_IN ; P1_U5184
g15147 nand P1_U3241 P1_STATE2_REG_2__SCAN_IN ; P1_U5185
g15148 nand P1_U5183 P1_U3686 ; P1_U5186
g15149 nand P1_U2506 P1_U2388 ; P1_U5187
g15150 nand P1_U3320 P1_U5187 ; P1_U5188
g15151 nand P1_U5188 P1_U3372 ; P1_U5189
g15152 nand P1_U5179 P1_STATE2_REG_2__SCAN_IN ; P1_U5190
g15153 nand P1_U5190 P1_U5189 ; P1_U5191
g15154 nand P1_U5176 P1_U2415 ; P1_U5192
g15155 nand P1_U2505 P1_U2413 ; P1_U5193
g15156 nand P1_U5175 P1_U2412 ; P1_U5194
g15157 nand P1_U2397 P1_U5191 ; P1_U5195
g15158 nand P1_U5186 P1_INSTQUEUE_REG_4__7__SCAN_IN ; P1_U5196
g15159 nand P1_U5176 P1_U2416 ; P1_U5197
g15160 nand P1_U2505 P1_U2411 ; P1_U5198
g15161 nand P1_U5175 P1_U2410 ; P1_U5199
g15162 nand P1_U2396 P1_U5191 ; P1_U5200
g15163 nand P1_U5186 P1_INSTQUEUE_REG_4__6__SCAN_IN ; P1_U5201
g15164 nand P1_U5176 P1_U2420 ; P1_U5202
g15165 nand P1_U2505 P1_U2409 ; P1_U5203
g15166 nand P1_U5175 P1_U2408 ; P1_U5204
g15167 nand P1_U2395 P1_U5191 ; P1_U5205
g15168 nand P1_U5186 P1_INSTQUEUE_REG_4__5__SCAN_IN ; P1_U5206
g15169 nand P1_U5176 P1_U2419 ; P1_U5207
g15170 nand P1_U2505 P1_U2407 ; P1_U5208
g15171 nand P1_U5175 P1_U2406 ; P1_U5209
g15172 nand P1_U2394 P1_U5191 ; P1_U5210
g15173 nand P1_U5186 P1_INSTQUEUE_REG_4__4__SCAN_IN ; P1_U5211
g15174 nand P1_U5176 P1_U2418 ; P1_U5212
g15175 nand P1_U2505 P1_U2405 ; P1_U5213
g15176 nand P1_U5175 P1_U2404 ; P1_U5214
g15177 nand P1_U2393 P1_U5191 ; P1_U5215
g15178 nand P1_U5186 P1_INSTQUEUE_REG_4__3__SCAN_IN ; P1_U5216
g15179 nand P1_U5176 P1_U2421 ; P1_U5217
g15180 nand P1_U2505 P1_U2403 ; P1_U5218
g15181 nand P1_U5175 P1_U2402 ; P1_U5219
g15182 nand P1_U2392 P1_U5191 ; P1_U5220
g15183 nand P1_U5186 P1_INSTQUEUE_REG_4__2__SCAN_IN ; P1_U5221
g15184 nand P1_U5176 P1_U2414 ; P1_U5222
g15185 nand P1_U2505 P1_U2401 ; P1_U5223
g15186 nand P1_U5175 P1_U2400 ; P1_U5224
g15187 nand P1_U2391 P1_U5191 ; P1_U5225
g15188 nand P1_U5186 P1_INSTQUEUE_REG_4__1__SCAN_IN ; P1_U5226
g15189 nand P1_U5176 P1_U2417 ; P1_U5227
g15190 nand P1_U2505 P1_U2399 ; P1_U5228
g15191 nand P1_U5175 P1_U2398 ; P1_U5229
g15192 nand P1_U2390 P1_U5191 ; P1_U5230
g15193 nand P1_U5186 P1_INSTQUEUE_REG_4__0__SCAN_IN ; P1_U5231
g15194 not P1_U3374 ; P1_U5232
g15195 not P1_U3373 ; P1_U5233
g15196 nand P1_U2441 P1_U2442 ; P1_U5234
g15197 not P1_U3375 ; P1_U5235
g15198 nand P1_U2435 P1_U2436 ; P1_U5236
g15199 not P1_U3376 ; P1_U5237
g15200 nand P1_U2508 P1_U4528 ; P1_U5238
g15201 nand P1_U2511 P1_U2358 ; P1_U5239
g15202 nand P1_U3320 P1_U5239 ; P1_U5240
g15203 nand P1_U5235 P1_U5240 ; P1_U5241
g15204 nand P1_U3373 P1_STATE2_REG_3__SCAN_IN ; P1_U5242
g15205 nand P1_U5237 P1_STATE2_REG_2__SCAN_IN ; P1_U5243
g15206 nand P1_U5241 P1_U3695 ; P1_U5244
g15207 nand P1_U2511 P1_U2388 ; P1_U5245
g15208 nand P1_U3320 P1_U5245 ; P1_U5246
g15209 nand P1_U5246 P1_U3375 ; P1_U5247
g15210 nand P1_U3376 P1_STATE2_REG_2__SCAN_IN ; P1_U5248
g15211 nand P1_U5248 P1_U5247 ; P1_U5249
g15212 nand P1_U5233 P1_U2415 ; P1_U5250
g15213 nand P1_U2509 P1_U2413 ; P1_U5251
g15214 nand P1_U5232 P1_U2412 ; P1_U5252
g15215 nand P1_U2397 P1_U5249 ; P1_U5253
g15216 nand P1_U5244 P1_INSTQUEUE_REG_3__7__SCAN_IN ; P1_U5254
g15217 nand P1_U5233 P1_U2416 ; P1_U5255
g15218 nand P1_U2509 P1_U2411 ; P1_U5256
g15219 nand P1_U5232 P1_U2410 ; P1_U5257
g15220 nand P1_U2396 P1_U5249 ; P1_U5258
g15221 nand P1_U5244 P1_INSTQUEUE_REG_3__6__SCAN_IN ; P1_U5259
g15222 nand P1_U5233 P1_U2420 ; P1_U5260
g15223 nand P1_U2509 P1_U2409 ; P1_U5261
g15224 nand P1_U5232 P1_U2408 ; P1_U5262
g15225 nand P1_U2395 P1_U5249 ; P1_U5263
g15226 nand P1_U5244 P1_INSTQUEUE_REG_3__5__SCAN_IN ; P1_U5264
g15227 nand P1_U5233 P1_U2419 ; P1_U5265
g15228 nand P1_U2509 P1_U2407 ; P1_U5266
g15229 nand P1_U5232 P1_U2406 ; P1_U5267
g15230 nand P1_U2394 P1_U5249 ; P1_U5268
g15231 nand P1_U5244 P1_INSTQUEUE_REG_3__4__SCAN_IN ; P1_U5269
g15232 nand P1_U5233 P1_U2418 ; P1_U5270
g15233 nand P1_U2509 P1_U2405 ; P1_U5271
g15234 nand P1_U5232 P1_U2404 ; P1_U5272
g15235 nand P1_U2393 P1_U5249 ; P1_U5273
g15236 nand P1_U5244 P1_INSTQUEUE_REG_3__3__SCAN_IN ; P1_U5274
g15237 nand P1_U5233 P1_U2421 ; P1_U5275
g15238 nand P1_U2509 P1_U2403 ; P1_U5276
g15239 nand P1_U5232 P1_U2402 ; P1_U5277
g15240 nand P1_U2392 P1_U5249 ; P1_U5278
g15241 nand P1_U5244 P1_INSTQUEUE_REG_3__2__SCAN_IN ; P1_U5279
g15242 nand P1_U5233 P1_U2414 ; P1_U5280
g15243 nand P1_U2509 P1_U2401 ; P1_U5281
g15244 nand P1_U5232 P1_U2400 ; P1_U5282
g15245 nand P1_U2391 P1_U5249 ; P1_U5283
g15246 nand P1_U5244 P1_INSTQUEUE_REG_3__1__SCAN_IN ; P1_U5284
g15247 nand P1_U5233 P1_U2417 ; P1_U5285
g15248 nand P1_U2509 P1_U2399 ; P1_U5286
g15249 nand P1_U5232 P1_U2398 ; P1_U5287
g15250 nand P1_U2390 P1_U5249 ; P1_U5288
g15251 nand P1_U5244 P1_INSTQUEUE_REG_3__0__SCAN_IN ; P1_U5289
g15252 not P1_U3378 ; P1_U5290
g15253 not P1_U3377 ; P1_U5291
g15254 nand P1_U2441 P1_U2443 ; P1_U5292
g15255 not P1_U3379 ; P1_U5293
g15256 not P1_U3242 ; P1_U5294
g15257 nand P1_U2508 P1_U4524 ; P1_U5295
g15258 nand P1_U2513 P1_U2358 ; P1_U5296
g15259 nand P1_U3320 P1_U5296 ; P1_U5297
g15260 nand P1_U5293 P1_U5297 ; P1_U5298
g15261 nand P1_U3377 P1_STATE2_REG_3__SCAN_IN ; P1_U5299
g15262 nand P1_U3242 P1_STATE2_REG_2__SCAN_IN ; P1_U5300
g15263 nand P1_U5298 P1_U3704 ; P1_U5301
g15264 nand P1_U2513 P1_U2388 ; P1_U5302
g15265 nand P1_U3320 P1_U5302 ; P1_U5303
g15266 nand P1_U5303 P1_U3379 ; P1_U5304
g15267 nand P1_U5294 P1_STATE2_REG_2__SCAN_IN ; P1_U5305
g15268 nand P1_U5305 P1_U5304 ; P1_U5306
g15269 nand P1_U5291 P1_U2415 ; P1_U5307
g15270 nand P1_U2512 P1_U2413 ; P1_U5308
g15271 nand P1_U5290 P1_U2412 ; P1_U5309
g15272 nand P1_U2397 P1_U5306 ; P1_U5310
g15273 nand P1_U5301 P1_INSTQUEUE_REG_2__7__SCAN_IN ; P1_U5311
g15274 nand P1_U5291 P1_U2416 ; P1_U5312
g15275 nand P1_U2512 P1_U2411 ; P1_U5313
g15276 nand P1_U5290 P1_U2410 ; P1_U5314
g15277 nand P1_U2396 P1_U5306 ; P1_U5315
g15278 nand P1_U5301 P1_INSTQUEUE_REG_2__6__SCAN_IN ; P1_U5316
g15279 nand P1_U5291 P1_U2420 ; P1_U5317
g15280 nand P1_U2512 P1_U2409 ; P1_U5318
g15281 nand P1_U5290 P1_U2408 ; P1_U5319
g15282 nand P1_U2395 P1_U5306 ; P1_U5320
g15283 nand P1_U5301 P1_INSTQUEUE_REG_2__5__SCAN_IN ; P1_U5321
g15284 nand P1_U5291 P1_U2419 ; P1_U5322
g15285 nand P1_U2512 P1_U2407 ; P1_U5323
g15286 nand P1_U5290 P1_U2406 ; P1_U5324
g15287 nand P1_U2394 P1_U5306 ; P1_U5325
g15288 nand P1_U5301 P1_INSTQUEUE_REG_2__4__SCAN_IN ; P1_U5326
g15289 nand P1_U5291 P1_U2418 ; P1_U5327
g15290 nand P1_U2512 P1_U2405 ; P1_U5328
g15291 nand P1_U5290 P1_U2404 ; P1_U5329
g15292 nand P1_U2393 P1_U5306 ; P1_U5330
g15293 nand P1_U5301 P1_INSTQUEUE_REG_2__3__SCAN_IN ; P1_U5331
g15294 nand P1_U5291 P1_U2421 ; P1_U5332
g15295 nand P1_U2512 P1_U2403 ; P1_U5333
g15296 nand P1_U5290 P1_U2402 ; P1_U5334
g15297 nand P1_U2392 P1_U5306 ; P1_U5335
g15298 nand P1_U5301 P1_INSTQUEUE_REG_2__2__SCAN_IN ; P1_U5336
g15299 nand P1_U5291 P1_U2414 ; P1_U5337
g15300 nand P1_U2512 P1_U2401 ; P1_U5338
g15301 nand P1_U5290 P1_U2400 ; P1_U5339
g15302 nand P1_U2391 P1_U5306 ; P1_U5340
g15303 nand P1_U5301 P1_INSTQUEUE_REG_2__1__SCAN_IN ; P1_U5341
g15304 nand P1_U5291 P1_U2417 ; P1_U5342
g15305 nand P1_U2512 P1_U2399 ; P1_U5343
g15306 nand P1_U5290 P1_U2398 ; P1_U5344
g15307 nand P1_U2390 P1_U5306 ; P1_U5345
g15308 nand P1_U5301 P1_INSTQUEUE_REG_2__0__SCAN_IN ; P1_U5346
g15309 not P1_U3381 ; P1_U5347
g15310 not P1_U3380 ; P1_U5348
g15311 nand P1_U2441 P1_U2444 ; P1_U5349
g15312 not P1_U3382 ; P1_U5350
g15313 nand P1_U2435 P1_U2437 ; P1_U5351
g15314 not P1_U3383 ; P1_U5352
g15315 nand P1_U2508 P1_U4525 ; P1_U5353
g15316 nand P1_U2515 P1_U2358 ; P1_U5354
g15317 nand P1_U3320 P1_U5354 ; P1_U5355
g15318 nand P1_U5350 P1_U5355 ; P1_U5356
g15319 nand P1_U3380 P1_STATE2_REG_3__SCAN_IN ; P1_U5357
g15320 nand P1_U5352 P1_STATE2_REG_2__SCAN_IN ; P1_U5358
g15321 nand P1_U5356 P1_U3713 ; P1_U5359
g15322 nand P1_U2515 P1_U2388 ; P1_U5360
g15323 nand P1_U3320 P1_U5360 ; P1_U5361
g15324 nand P1_U5361 P1_U3382 ; P1_U5362
g15325 nand P1_U3383 P1_STATE2_REG_2__SCAN_IN ; P1_U5363
g15326 nand P1_U5363 P1_U5362 ; P1_U5364
g15327 nand P1_U5348 P1_U2415 ; P1_U5365
g15328 nand P1_U2514 P1_U2413 ; P1_U5366
g15329 nand P1_U5347 P1_U2412 ; P1_U5367
g15330 nand P1_U2397 P1_U5364 ; P1_U5368
g15331 nand P1_U5359 P1_INSTQUEUE_REG_1__7__SCAN_IN ; P1_U5369
g15332 nand P1_U5348 P1_U2416 ; P1_U5370
g15333 nand P1_U2514 P1_U2411 ; P1_U5371
g15334 nand P1_U5347 P1_U2410 ; P1_U5372
g15335 nand P1_U2396 P1_U5364 ; P1_U5373
g15336 nand P1_U5359 P1_INSTQUEUE_REG_1__6__SCAN_IN ; P1_U5374
g15337 nand P1_U5348 P1_U2420 ; P1_U5375
g15338 nand P1_U2514 P1_U2409 ; P1_U5376
g15339 nand P1_U5347 P1_U2408 ; P1_U5377
g15340 nand P1_U2395 P1_U5364 ; P1_U5378
g15341 nand P1_U5359 P1_INSTQUEUE_REG_1__5__SCAN_IN ; P1_U5379
g15342 nand P1_U5348 P1_U2419 ; P1_U5380
g15343 nand P1_U2514 P1_U2407 ; P1_U5381
g15344 nand P1_U5347 P1_U2406 ; P1_U5382
g15345 nand P1_U2394 P1_U5364 ; P1_U5383
g15346 nand P1_U5359 P1_INSTQUEUE_REG_1__4__SCAN_IN ; P1_U5384
g15347 nand P1_U5348 P1_U2418 ; P1_U5385
g15348 nand P1_U2514 P1_U2405 ; P1_U5386
g15349 nand P1_U5347 P1_U2404 ; P1_U5387
g15350 nand P1_U2393 P1_U5364 ; P1_U5388
g15351 nand P1_U5359 P1_INSTQUEUE_REG_1__3__SCAN_IN ; P1_U5389
g15352 nand P1_U5348 P1_U2421 ; P1_U5390
g15353 nand P1_U2514 P1_U2403 ; P1_U5391
g15354 nand P1_U5347 P1_U2402 ; P1_U5392
g15355 nand P1_U2392 P1_U5364 ; P1_U5393
g15356 nand P1_U5359 P1_INSTQUEUE_REG_1__2__SCAN_IN ; P1_U5394
g15357 nand P1_U5348 P1_U2414 ; P1_U5395
g15358 nand P1_U2514 P1_U2401 ; P1_U5396
g15359 nand P1_U5347 P1_U2400 ; P1_U5397
g15360 nand P1_U2391 P1_U5364 ; P1_U5398
g15361 nand P1_U5359 P1_INSTQUEUE_REG_1__1__SCAN_IN ; P1_U5399
g15362 nand P1_U5348 P1_U2417 ; P1_U5400
g15363 nand P1_U2514 P1_U2399 ; P1_U5401
g15364 nand P1_U5347 P1_U2398 ; P1_U5402
g15365 nand P1_U2390 P1_U5364 ; P1_U5403
g15366 nand P1_U5359 P1_INSTQUEUE_REG_1__0__SCAN_IN ; P1_U5404
g15367 not P1_U3385 ; P1_U5405
g15368 not P1_U3384 ; P1_U5406
g15369 nand P1_U2441 P1_U2445 ; P1_U5407
g15370 not P1_U3386 ; P1_U5408
g15371 not P1_U3243 ; P1_U5409
g15372 nand P1_U2508 P1_U2486 ; P1_U5410
g15373 nand P1_U2517 P1_U2358 ; P1_U5411
g15374 nand P1_U3320 P1_U5411 ; P1_U5412
g15375 nand P1_U5408 P1_U5412 ; P1_U5413
g15376 nand P1_U3384 P1_STATE2_REG_3__SCAN_IN ; P1_U5414
g15377 nand P1_U3243 P1_STATE2_REG_2__SCAN_IN ; P1_U5415
g15378 nand P1_U5413 P1_U3722 ; P1_U5416
g15379 nand P1_U2517 P1_U2388 ; P1_U5417
g15380 nand P1_U3320 P1_U5417 ; P1_U5418
g15381 nand P1_U5418 P1_U3386 ; P1_U5419
g15382 nand P1_U5409 P1_STATE2_REG_2__SCAN_IN ; P1_U5420
g15383 nand P1_U5420 P1_U5419 ; P1_U5421
g15384 nand P1_U5406 P1_U2415 ; P1_U5422
g15385 nand P1_U2516 P1_U2413 ; P1_U5423
g15386 nand P1_U5405 P1_U2412 ; P1_U5424
g15387 nand P1_U2397 P1_U5421 ; P1_U5425
g15388 nand P1_U5416 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U5426
g15389 nand P1_U5406 P1_U2416 ; P1_U5427
g15390 nand P1_U2516 P1_U2411 ; P1_U5428
g15391 nand P1_U5405 P1_U2410 ; P1_U5429
g15392 nand P1_U2396 P1_U5421 ; P1_U5430
g15393 nand P1_U5416 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U5431
g15394 nand P1_U5406 P1_U2420 ; P1_U5432
g15395 nand P1_U2516 P1_U2409 ; P1_U5433
g15396 nand P1_U5405 P1_U2408 ; P1_U5434
g15397 nand P1_U2395 P1_U5421 ; P1_U5435
g15398 nand P1_U5416 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U5436
g15399 nand P1_U5406 P1_U2419 ; P1_U5437
g15400 nand P1_U2516 P1_U2407 ; P1_U5438
g15401 nand P1_U5405 P1_U2406 ; P1_U5439
g15402 nand P1_U2394 P1_U5421 ; P1_U5440
g15403 nand P1_U5406 P1_U2418 ; P1_U5441
g15404 nand P1_U2516 P1_U2405 ; P1_U5442
g15405 nand P1_U5405 P1_U2404 ; P1_U5443
g15406 nand P1_U2393 P1_U5421 ; P1_U5444
g15407 nand P1_U5416 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U5445
g15408 nand P1_U5406 P1_U2421 ; P1_U5446
g15409 nand P1_U2516 P1_U2403 ; P1_U5447
g15410 nand P1_U5405 P1_U2402 ; P1_U5448
g15411 nand P1_U2392 P1_U5421 ; P1_U5449
g15412 nand P1_U5416 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U5450
g15413 nand P1_U5406 P1_U2414 ; P1_U5451
g15414 nand P1_U2516 P1_U2401 ; P1_U5452
g15415 nand P1_U5405 P1_U2400 ; P1_U5453
g15416 nand P1_U2391 P1_U5421 ; P1_U5454
g15417 nand P1_U5416 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U5455
g15418 nand P1_U5406 P1_U2417 ; P1_U5456
g15419 nand P1_U2516 P1_U2399 ; P1_U5457
g15420 nand P1_U5405 P1_U2398 ; P1_U5458
g15421 nand P1_U2390 P1_U5421 ; P1_U5459
g15422 nand P1_U5416 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U5460
g15423 not P1_U3423 ; P1_U5461
g15424 nand P1_U3391 P1_U3394 P1_U4503 ; P1_U5462
g15425 nand P1_U4400 P1_U4173 P1_U4460 ; P1_U5463
g15426 not P1_U3244 ; P1_U5464
g15427 nand P1_U4494 P1_U3289 ; P1_U5465
g15428 nand P1_U5465 P1_U3283 P1_U5464 ; P1_U5466
g15429 nand P1_U3732 P1_U2452 ; P1_U5467
g15430 nand P1_U4208 P1_U5462 ; P1_U5468
g15431 nand P1_U3733 P1_U7609 ; P1_U5469
g15432 nand P1_U4215 P1_U3257 P1_GTE_485_U6 ; P1_U5470
g15433 nand P1_U2449 P1_U7494 ; P1_U5471
g15434 nand P1_U4257 P1_U4503 ; P1_U5472
g15435 not P1_U4182 ; P1_U5473
g15436 nand P1_U2368 P1_U4182 ; P1_U5474
g15437 nand P1_U3294 P1_STATE2_REG_3__SCAN_IN ; P1_U5475
g15438 not P1_U4172 ; P1_U5476
g15439 nand P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U5477
g15440 nand P1_U5477 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U5478
g15441 nand P1_U4381 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U5479
g15442 not P1_U3442 ; P1_U5480
g15443 nand P1_U3498 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U5481
g15444 nand P1_U5481 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U5482
g15445 not P1_U3438 ; P1_U5483
g15446 nand P1_U3275 P1_U3264 ; P1_U5484
g15447 nand P1_U5484 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U5485
g15448 nand P1_U2469 P1_U3275 ; P1_U5486
g15449 nand P1_U4494 P1_U3290 ; P1_U5487
g15450 nand P1_U4400 P1_U2605 ; P1_U5488
g15451 nand P1_U7704 P1_U7703 P1_U7494 ; P1_U5489
g15452 nand P1_U4449 P1_U5488 ; P1_U5490
g15453 nand P1_U4400 P1_U3394 P1_U3409 ; P1_U5491
g15454 nand P1_U5491 P1_U4171 ; P1_U5492
g15455 nand P1_U7629 P1_U5492 ; P1_U5493
g15456 nand P1_U4460 P1_U4171 ; P1_U5494
g15457 nand P1_U3395 P1_U5494 ; P1_U5495
g15458 nand P1_U4208 P1_U5462 ; P1_U5496
g15459 nand P1_U4257 P1_U4503 ; P1_U5497
g15460 nand P1_U5495 P1_U3271 ; P1_U5498
g15461 nand P1_U4494 P1_U7707 ; P1_U5499
g15462 nand P1_U4190 P1_U3244 ; P1_U5500
g15463 nand P1_U3292 P1_U4217 ; P1_U5501
g15464 nand P1_U3740 P1_U5501 ; P1_U5502
g15465 nand P1_R2182_U25 P1_U7509 ; P1_U5503
g15466 nand P1_U4218 P1_U3438 ; P1_U5504
g15467 nand P1_U4214 P1_U3442 ; P1_U5505
g15468 nand P1_U5503 P1_U3747 ; P1_U5506
g15469 nand P1_U4252 P1_U3438 ; P1_U5507
g15470 nand P1_U2427 P1_U5506 ; P1_U5508
g15471 nand P1_U5508 P1_U5507 ; P1_U5509
g15472 nand P1_U3275 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U5510
g15473 not P1_U3401 ; P1_U5511
g15474 nand P1_R2182_U42 P1_U7509 ; P1_U5512
g15475 nand P1_U4214 P1_U3456 ; P1_U5513
g15476 nand P1_U3749 P1_U5512 ; P1_U5514
g15477 nand P1_U2446 P1_U3470 ; P1_U5515
g15478 nand P1_U4252 P1_U3401 ; P1_U5516
g15479 nand P1_U2427 P1_U5514 ; P1_U5517
g15480 nand P1_U5517 P1_U5515 P1_U5516 ; P1_U5518
g15481 not P1_U3402 ; P1_U5519
g15482 nand P1_U2431 P1_U4249 ; P1_U5520
g15483 nand P1_U3292 P1_U5520 ; P1_U5521
g15484 nand P1_U5519 P1_U5521 ; P1_U5522
g15485 nand P1_R2182_U33 P1_U7509 ; P1_U5523
g15486 nand P1_U4214 P1_U3265 ; P1_U5524
g15487 nand P1_U3750 P1_U5523 ; P1_U5525
g15488 nand P1_U7712 P1_U2446 ; P1_U5526
g15489 nand P1_U5519 P1_U4252 ; P1_U5527
g15490 nand P1_U2427 P1_U5525 ; P1_U5528
g15491 nand P1_U5528 P1_U5526 P1_U5527 ; P1_U5529
g15492 nand P1_R2182_U34 P1_U7509 ; P1_U5530
g15493 nand P1_U4175 P1_U5530 ; P1_U5531
g15494 nand P1_U4252 P1_U3266 ; P1_U5532
g15495 nand P1_U2427 P1_U5531 ; P1_U5533
g15496 nand P1_U7715 P1_STATE2_REG_1__SCAN_IN ; P1_U5534
g15497 nand P1_U5533 P1_U5534 P1_U5532 ; P1_U5535
g15498 nand P1_U2428 P1_LT_589_U6 P1_STATE2_REG_0__SCAN_IN ; P1_U5536
g15499 not P1_U3404 ; P1_U5537
g15500 nand P1_U3296 P1_STATE2_REG_1__SCAN_IN ; P1_U5538
g15501 nand P1_U4527 P1_U3454 ; P1_U5539
g15502 nand P1_U3358 P1_U5539 ; P1_U5540
g15503 nand P1_U3359 P1_U5540 ; P1_U5541
g15504 nand P1_U2388 P1_U5541 ; P1_U5542
g15505 nand P1_R2182_U25 P1_U5538 ; P1_U5543
g15506 nand P1_U4226 P1_R2144_U8 ; P1_U5544
g15507 nand P1_U3751 P1_U5542 ; P1_U5545
g15508 nand P1_U2388 P1_U7733 ; P1_U5546
g15509 nand P1_R2182_U42 P1_U5538 ; P1_U5547
g15510 nand P1_U4226 P1_R2144_U49 ; P1_U5548
g15511 nand P1_U3752 P1_U5546 ; P1_U5549
g15512 nand P1_U3326 P1_U3333 ; P1_U5550
g15513 nand P1_U2388 P1_U5550 ; P1_U5551
g15514 nand P1_R2182_U33 P1_U5538 ; P1_U5552
g15515 nand P1_U4226 P1_R2144_U50 ; P1_U5553
g15516 nand P1_U3753 P1_U5551 ; P1_U5554
g15517 nand P1_R2182_U34 P1_U5538 ; P1_U5555
g15518 nand P1_R2144_U43 P1_U4209 ; P1_U5556
g15519 nand P1_U5555 P1_U5556 P1_U4245 ; P1_U5557
g15520 nand P1_U4477 P1_U3272 ; P1_U5558
g15521 nand P1_U4260 P1_U2431 ; P1_U5559
g15522 nand P1_U2518 P1_U5559 P1_U7743 P1_U7742 ; P1_U5560
g15523 nand P1_U4235 P1_U4503 P1_U4192 ; P1_U5561
g15524 nand P1_U2368 P1_U5560 ; P1_U5562
g15525 nand P1_U4203 P1_U3263 ; P1_U5563
g15526 not P1_U3414 ; P1_U5564
g15527 nand P1_U4262 P1_U4208 ; P1_U5565
g15528 nand P1_U4256 P1_U2389 ; P1_U5566
g15529 nand P1_U4266 P1_U4250 ; P1_U5567
g15530 nand P1_U4264 P1_U4494 ; P1_U5568
g15531 nand P1_U3758 P1_U2519 ; P1_U5569
g15532 nand P1_R2099_U86 P1_U2380 ; P1_U5570
g15533 nand P1_R2027_U5 P1_U2378 ; P1_U5571
g15534 nand P1_R2278_U99 P1_U2377 ; P1_U5572
g15535 nand P1_ADD_405_U4 P1_U2375 ; P1_U5573
g15536 nand P1_U2374 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_U5574
g15537 nand P1_U2370 P1_REIP_REG_0__SCAN_IN ; P1_U5575
g15538 nand P1_U5564 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_U5576
g15539 nand P1_R2099_U87 P1_U2380 ; P1_U5577
g15540 nand P1_R2027_U71 P1_U2378 ; P1_U5578
g15541 nand P1_R2278_U19 P1_U2377 ; P1_U5579
g15542 nand P1_ADD_405_U85 P1_U2375 ; P1_U5580
g15543 nand P1_ADD_515_U4 P1_U2374 ; P1_U5581
g15544 nand P1_U2370 P1_REIP_REG_1__SCAN_IN ; P1_U5582
g15545 nand P1_U5564 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_U5583
g15546 nand P1_R2099_U138 P1_U2380 ; P1_U5584
g15547 nand P1_R2027_U60 P1_U2378 ; P1_U5585
g15548 nand P1_R2278_U107 P1_U2377 ; P1_U5586
g15549 nand P1_ADD_405_U5 P1_U2375 ; P1_U5587
g15550 nand P1_ADD_515_U67 P1_U2374 ; P1_U5588
g15551 nand P1_U2370 P1_REIP_REG_2__SCAN_IN ; P1_U5589
g15552 nand P1_U5564 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_U5590
g15553 nand P1_R2099_U42 P1_U2380 ; P1_U5591
g15554 nand P1_R2027_U57 P1_U2378 ; P1_U5592
g15555 nand P1_R2278_U105 P1_U2377 ; P1_U5593
g15556 nand P1_ADD_405_U95 P1_U2375 ; P1_U5594
g15557 nand P1_ADD_515_U85 P1_U2374 ; P1_U5595
g15558 nand P1_U2370 P1_REIP_REG_3__SCAN_IN ; P1_U5596
g15559 nand P1_U5564 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_U5597
g15560 nand P1_R2099_U41 P1_U2380 ; P1_U5598
g15561 nand P1_R2027_U56 P1_U2378 ; P1_U5599
g15562 nand P1_R2278_U104 P1_U2377 ; P1_U5600
g15563 nand P1_ADD_405_U76 P1_U2375 ; P1_U5601
g15564 nand P1_ADD_515_U76 P1_U2374 ; P1_U5602
g15565 nand P1_U2370 P1_REIP_REG_4__SCAN_IN ; P1_U5603
g15566 nand P1_U5564 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_U5604
g15567 nand P1_R2099_U40 P1_U2380 ; P1_U5605
g15568 nand P1_R2027_U55 P1_U2378 ; P1_U5606
g15569 nand P1_R2278_U17 P1_U2377 ; P1_U5607
g15570 nand P1_ADD_405_U79 P1_U2375 ; P1_U5608
g15571 nand P1_ADD_515_U79 P1_U2374 ; P1_U5609
g15572 nand P1_U2370 P1_REIP_REG_5__SCAN_IN ; P1_U5610
g15573 nand P1_U5564 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_U5611
g15574 nand P1_R2099_U39 P1_U2380 ; P1_U5612
g15575 nand P1_R2027_U54 P1_U2378 ; P1_U5613
g15576 nand P1_R2278_U103 P1_U2377 ; P1_U5614
g15577 nand P1_ADD_405_U63 P1_U2375 ; P1_U5615
g15578 nand P1_ADD_515_U62 P1_U2374 ; P1_U5616
g15579 nand P1_U2370 P1_REIP_REG_6__SCAN_IN ; P1_U5617
g15580 nand P1_U5564 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_U5618
g15581 nand P1_R2099_U38 P1_U2380 ; P1_U5619
g15582 nand P1_R2027_U53 P1_U2378 ; P1_U5620
g15583 nand P1_R2278_U18 P1_U2377 ; P1_U5621
g15584 nand P1_ADD_405_U89 P1_U2375 ; P1_U5622
g15585 nand P1_ADD_515_U89 P1_U2374 ; P1_U5623
g15586 nand P1_U2370 P1_REIP_REG_7__SCAN_IN ; P1_U5624
g15587 nand P1_U5564 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_U5625
g15588 nand P1_R2099_U37 P1_U2380 ; P1_U5626
g15589 nand P1_R2027_U52 P1_U2378 ; P1_U5627
g15590 nand P1_R2278_U102 P1_U2377 ; P1_U5628
g15591 nand P1_ADD_405_U80 P1_U2375 ; P1_U5629
g15592 nand P1_ADD_515_U80 P1_U2374 ; P1_U5630
g15593 nand P1_U2370 P1_REIP_REG_8__SCAN_IN ; P1_U5631
g15594 nand P1_U5564 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_U5632
g15595 nand P1_R2099_U36 P1_U2380 ; P1_U5633
g15596 nand P1_R2027_U51 P1_U2378 ; P1_U5634
g15597 nand P1_R2278_U101 P1_U2377 ; P1_U5635
g15598 nand P1_ADD_405_U70 P1_U2375 ; P1_U5636
g15599 nand P1_ADD_515_U70 P1_U2374 ; P1_U5637
g15600 nand P1_U2370 P1_REIP_REG_9__SCAN_IN ; P1_U5638
g15601 nand P1_U5564 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_U5639
g15602 nand P1_R2099_U85 P1_U2380 ; P1_U5640
g15603 nand P1_R2027_U81 P1_U2378 ; P1_U5641
g15604 nand P1_R2278_U126 P1_U2377 ; P1_U5642
g15605 nand P1_ADD_405_U83 P1_U2375 ; P1_U5643
g15606 nand P1_ADD_515_U83 P1_U2374 ; P1_U5644
g15607 nand P1_U2370 P1_REIP_REG_10__SCAN_IN ; P1_U5645
g15608 nand P1_U5564 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_U5646
g15609 nand P1_R2099_U84 P1_U2380 ; P1_U5647
g15610 nand P1_R2027_U80 P1_U2378 ; P1_U5648
g15611 nand P1_R2278_U15 P1_U2377 ; P1_U5649
g15612 nand P1_ADD_405_U73 P1_U2375 ; P1_U5650
g15613 nand P1_ADD_515_U73 P1_U2374 ; P1_U5651
g15614 nand P1_U2370 P1_REIP_REG_11__SCAN_IN ; P1_U5652
g15615 nand P1_U5564 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_U5653
g15616 nand P1_R2099_U83 P1_U2380 ; P1_U5654
g15617 nand P1_R2027_U79 P1_U2378 ; P1_U5655
g15618 nand P1_R2278_U125 P1_U2377 ; P1_U5656
g15619 nand P1_ADD_405_U88 P1_U2375 ; P1_U5657
g15620 nand P1_ADD_515_U88 P1_U2374 ; P1_U5658
g15621 nand P1_U2370 P1_REIP_REG_12__SCAN_IN ; P1_U5659
g15622 nand P1_U5564 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_U5660
g15623 nand P1_R2099_U82 P1_U2380 ; P1_U5661
g15624 nand P1_R2027_U78 P1_U2378 ; P1_U5662
g15625 nand P1_R2278_U123 P1_U2377 ; P1_U5663
g15626 nand P1_ADD_405_U69 P1_U2375 ; P1_U5664
g15627 nand P1_ADD_515_U69 P1_U2374 ; P1_U5665
g15628 nand P1_U2370 P1_REIP_REG_13__SCAN_IN ; P1_U5666
g15629 nand P1_U5564 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_U5667
g15630 nand P1_R2099_U81 P1_U2380 ; P1_U5668
g15631 nand P1_R2027_U77 P1_U2378 ; P1_U5669
g15632 nand P1_R2278_U122 P1_U2377 ; P1_U5670
g15633 nand P1_ADD_405_U78 P1_U2375 ; P1_U5671
g15634 nand P1_ADD_515_U78 P1_U2374 ; P1_U5672
g15635 nand P1_U2370 P1_REIP_REG_14__SCAN_IN ; P1_U5673
g15636 nand P1_U5564 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_U5674
g15637 nand P1_R2099_U80 P1_U2380 ; P1_U5675
g15638 nand P1_R2027_U76 P1_U2378 ; P1_U5676
g15639 nand P1_R2278_U20 P1_U2377 ; P1_U5677
g15640 nand P1_ADD_405_U75 P1_U2375 ; P1_U5678
g15641 nand P1_ADD_515_U75 P1_U2374 ; P1_U5679
g15642 nand P1_U2370 P1_REIP_REG_15__SCAN_IN ; P1_U5680
g15643 nand P1_U5564 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_U5681
g15644 nand P1_R2099_U79 P1_U2380 ; P1_U5682
g15645 nand P1_R2027_U75 P1_U2378 ; P1_U5683
g15646 nand P1_R2278_U121 P1_U2377 ; P1_U5684
g15647 nand P1_ADD_405_U91 P1_U2375 ; P1_U5685
g15648 nand P1_ADD_515_U91 P1_U2374 ; P1_U5686
g15649 nand P1_U2370 P1_REIP_REG_16__SCAN_IN ; P1_U5687
g15650 nand P1_U5564 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_U5688
g15651 nand P1_R2099_U78 P1_U2380 ; P1_U5689
g15652 nand P1_R2027_U74 P1_U2378 ; P1_U5690
g15653 nand P1_R2278_U120 P1_U2377 ; P1_U5691
g15654 nand P1_ADD_405_U67 P1_U2375 ; P1_U5692
g15655 nand P1_ADD_515_U66 P1_U2374 ; P1_U5693
g15656 nand P1_U2370 P1_REIP_REG_17__SCAN_IN ; P1_U5694
g15657 nand P1_U5564 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_U5695
g15658 nand P1_R2099_U77 P1_U2380 ; P1_U5696
g15659 nand P1_R2027_U73 P1_U2378 ; P1_U5697
g15660 nand P1_R2278_U119 P1_U2377 ; P1_U5698
g15661 nand P1_ADD_405_U72 P1_U2375 ; P1_U5699
g15662 nand P1_ADD_515_U72 P1_U2374 ; P1_U5700
g15663 nand P1_U2370 P1_REIP_REG_18__SCAN_IN ; P1_U5701
g15664 nand P1_U5564 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_U5702
g15665 nand P1_R2099_U76 P1_U2380 ; P1_U5703
g15666 nand P1_R2027_U72 P1_U2378 ; P1_U5704
g15667 nand P1_R2278_U118 P1_U2377 ; P1_U5705
g15668 nand P1_ADD_405_U82 P1_U2375 ; P1_U5706
g15669 nand P1_ADD_515_U82 P1_U2374 ; P1_U5707
g15670 nand P1_U2370 P1_REIP_REG_19__SCAN_IN ; P1_U5708
g15671 nand P1_U5564 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_U5709
g15672 nand P1_R2099_U75 P1_U2380 ; P1_U5710
g15673 nand P1_R2027_U70 P1_U2378 ; P1_U5711
g15674 nand P1_R2278_U117 P1_U2377 ; P1_U5712
g15675 nand P1_ADD_405_U68 P1_U2375 ; P1_U5713
g15676 nand P1_ADD_515_U68 P1_U2374 ; P1_U5714
g15677 nand P1_U2370 P1_REIP_REG_20__SCAN_IN ; P1_U5715
g15678 nand P1_U5564 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_U5716
g15679 nand P1_R2099_U74 P1_U2380 ; P1_U5717
g15680 nand P1_R2027_U69 P1_U2378 ; P1_U5718
g15681 nand P1_R2278_U116 P1_U2377 ; P1_U5719
g15682 nand P1_ADD_405_U87 P1_U2375 ; P1_U5720
g15683 nand P1_ADD_515_U87 P1_U2374 ; P1_U5721
g15684 nand P1_U2370 P1_REIP_REG_21__SCAN_IN ; P1_U5722
g15685 nand P1_U5564 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_U5723
g15686 nand P1_R2099_U73 P1_U2380 ; P1_U5724
g15687 nand P1_R2027_U68 P1_U2378 ; P1_U5725
g15688 nand P1_R2278_U115 P1_U2377 ; P1_U5726
g15689 nand P1_ADD_405_U71 P1_U2375 ; P1_U5727
g15690 nand P1_ADD_515_U71 P1_U2374 ; P1_U5728
g15691 nand P1_U2370 P1_REIP_REG_22__SCAN_IN ; P1_U5729
g15692 nand P1_U5564 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_U5730
g15693 nand P1_R2099_U72 P1_U2380 ; P1_U5731
g15694 nand P1_R2027_U67 P1_U2378 ; P1_U5732
g15695 nand P1_R2278_U114 P1_U2377 ; P1_U5733
g15696 nand P1_ADD_405_U81 P1_U2375 ; P1_U5734
g15697 nand P1_ADD_515_U81 P1_U2374 ; P1_U5735
g15698 nand P1_U2370 P1_REIP_REG_23__SCAN_IN ; P1_U5736
g15699 nand P1_U5564 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_U5737
g15700 nand P1_R2099_U71 P1_U2380 ; P1_U5738
g15701 nand P1_R2027_U66 P1_U2378 ; P1_U5739
g15702 nand P1_R2278_U113 P1_U2377 ; P1_U5740
g15703 nand P1_ADD_405_U66 P1_U2375 ; P1_U5741
g15704 nand P1_ADD_515_U65 P1_U2374 ; P1_U5742
g15705 nand P1_U2370 P1_REIP_REG_24__SCAN_IN ; P1_U5743
g15706 nand P1_U5564 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_U5744
g15707 nand P1_R2099_U70 P1_U2380 ; P1_U5745
g15708 nand P1_R2027_U65 P1_U2378 ; P1_U5746
g15709 nand P1_R2278_U112 P1_U2377 ; P1_U5747
g15710 nand P1_ADD_405_U90 P1_U2375 ; P1_U5748
g15711 nand P1_ADD_515_U90 P1_U2374 ; P1_U5749
g15712 nand P1_U2370 P1_REIP_REG_25__SCAN_IN ; P1_U5750
g15713 nand P1_U5564 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_U5751
g15714 nand P1_R2099_U69 P1_U2380 ; P1_U5752
g15715 nand P1_R2027_U64 P1_U2378 ; P1_U5753
g15716 nand P1_R2278_U111 P1_U2377 ; P1_U5754
g15717 nand P1_ADD_405_U74 P1_U2375 ; P1_U5755
g15718 nand P1_ADD_515_U74 P1_U2374 ; P1_U5756
g15719 nand P1_U2370 P1_REIP_REG_26__SCAN_IN ; P1_U5757
g15720 nand P1_U5564 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_U5758
g15721 nand P1_R2099_U68 P1_U2380 ; P1_U5759
g15722 nand P1_R2027_U63 P1_U2378 ; P1_U5760
g15723 nand P1_R2278_U110 P1_U2377 ; P1_U5761
g15724 nand P1_ADD_405_U77 P1_U2375 ; P1_U5762
g15725 nand P1_ADD_515_U77 P1_U2374 ; P1_U5763
g15726 nand P1_U2370 P1_REIP_REG_27__SCAN_IN ; P1_U5764
g15727 nand P1_U5564 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_U5765
g15728 nand P1_R2099_U67 P1_U2380 ; P1_U5766
g15729 nand P1_R2027_U62 P1_U2378 ; P1_U5767
g15730 nand P1_R2278_U109 P1_U2377 ; P1_U5768
g15731 nand P1_ADD_405_U86 P1_U2375 ; P1_U5769
g15732 nand P1_ADD_515_U86 P1_U2374 ; P1_U5770
g15733 nand P1_U2370 P1_REIP_REG_28__SCAN_IN ; P1_U5771
g15734 nand P1_U5564 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_U5772
g15735 nand P1_R2099_U66 P1_U2380 ; P1_U5773
g15736 nand P1_R2027_U61 P1_U2378 ; P1_U5774
g15737 nand P1_R2278_U108 P1_U2377 ; P1_U5775
g15738 nand P1_ADD_405_U65 P1_U2375 ; P1_U5776
g15739 nand P1_ADD_515_U64 P1_U2374 ; P1_U5777
g15740 nand P1_U2370 P1_REIP_REG_29__SCAN_IN ; P1_U5778
g15741 nand P1_U5564 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_U5779
g15742 nand P1_R2099_U65 P1_U2380 ; P1_U5780
g15743 nand P1_R2027_U59 P1_U2378 ; P1_U5781
g15744 nand P1_R2278_U106 P1_U2377 ; P1_U5782
g15745 nand P1_ADD_405_U64 P1_U2375 ; P1_U5783
g15746 nand P1_ADD_515_U63 P1_U2374 ; P1_U5784
g15747 nand P1_U2370 P1_REIP_REG_30__SCAN_IN ; P1_U5785
g15748 nand P1_U5564 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_U5786
g15749 nand P1_R2099_U64 P1_U2380 ; P1_U5787
g15750 nand P1_R2027_U58 P1_U2378 ; P1_U5788
g15751 nand P1_R2278_U16 P1_U2377 ; P1_U5789
g15752 nand P1_ADD_405_U84 P1_U2375 ; P1_U5790
g15753 nand P1_ADD_515_U84 P1_U2374 ; P1_U5791
g15754 nand P1_U2370 P1_REIP_REG_31__SCAN_IN ; P1_U5792
g15755 nand P1_U5564 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_U5793
g15756 nand P1_U4209 P1_U3294 ; P1_U5794
g15757 not P1_U3416 ; P1_U5795
g15758 nand P1_U3294 P1_STATE2_REG_2__SCAN_IN ; P1_U5796
g15759 nand P1_U3308 P1_STATE2_REG_1__SCAN_IN ; P1_U5797
g15760 nand P1_U5797 P1_U5796 ; P1_U5798
g15761 nand P1_U2376 P1_PHYADDRPOINTER_REG_0__SCAN_IN ; P1_U5799
g15762 nand P1_U2372 P1_R2278_U99 ; P1_U5800
g15763 nand P1_U2365 P1_REIP_REG_0__SCAN_IN ; P1_U5801
g15764 nand P1_R2358_U76 P1_U2364 ; P1_U5802
g15765 nand P1_U5795 P1_PHYADDRPOINTER_REG_0__SCAN_IN ; P1_U5803
g15766 nand P1_R2337_U4 P1_U2376 ; P1_U5804
g15767 nand P1_U2372 P1_R2278_U19 ; P1_U5805
g15768 nand P1_U2365 P1_REIP_REG_1__SCAN_IN ; P1_U5806
g15769 nand P1_R2358_U107 P1_U2364 ; P1_U5807
g15770 nand P1_U5795 P1_PHYADDRPOINTER_REG_1__SCAN_IN ; P1_U5808
g15771 nand P1_R2337_U71 P1_U2376 ; P1_U5809
g15772 nand P1_U2372 P1_R2278_U107 ; P1_U5810
g15773 nand P1_U2365 P1_REIP_REG_2__SCAN_IN ; P1_U5811
g15774 nand P1_R2358_U18 P1_U2364 ; P1_U5812
g15775 nand P1_U5795 P1_PHYADDRPOINTER_REG_2__SCAN_IN ; P1_U5813
g15776 nand P1_R2337_U68 P1_U2376 ; P1_U5814
g15777 nand P1_U2372 P1_R2278_U105 ; P1_U5815
g15778 nand P1_U2365 P1_REIP_REG_3__SCAN_IN ; P1_U5816
g15779 nand P1_R2358_U19 P1_U2364 ; P1_U5817
g15780 nand P1_U5795 P1_PHYADDRPOINTER_REG_3__SCAN_IN ; P1_U5818
g15781 nand P1_R2337_U67 P1_U2376 ; P1_U5819
g15782 nand P1_U2372 P1_R2278_U104 ; P1_U5820
g15783 nand P1_U2365 P1_REIP_REG_4__SCAN_IN ; P1_U5821
g15784 nand P1_R2358_U84 P1_U2364 ; P1_U5822
g15785 nand P1_U5795 P1_PHYADDRPOINTER_REG_4__SCAN_IN ; P1_U5823
g15786 nand P1_R2337_U66 P1_U2376 ; P1_U5824
g15787 nand P1_U2372 P1_R2278_U17 ; P1_U5825
g15788 nand P1_U2365 P1_REIP_REG_5__SCAN_IN ; P1_U5826
g15789 nand P1_R2358_U82 P1_U2364 ; P1_U5827
g15790 nand P1_U5795 P1_PHYADDRPOINTER_REG_5__SCAN_IN ; P1_U5828
g15791 nand P1_R2337_U65 P1_U2376 ; P1_U5829
g15792 nand P1_U2372 P1_R2278_U103 ; P1_U5830
g15793 nand P1_U2365 P1_REIP_REG_6__SCAN_IN ; P1_U5831
g15794 nand P1_R2358_U20 P1_U2364 ; P1_U5832
g15795 nand P1_U5795 P1_PHYADDRPOINTER_REG_6__SCAN_IN ; P1_U5833
g15796 nand P1_R2337_U64 P1_U2376 ; P1_U5834
g15797 nand P1_U2372 P1_R2278_U18 ; P1_U5835
g15798 nand P1_U2365 P1_REIP_REG_7__SCAN_IN ; P1_U5836
g15799 nand P1_R2358_U21 P1_U2364 ; P1_U5837
g15800 nand P1_U5795 P1_PHYADDRPOINTER_REG_7__SCAN_IN ; P1_U5838
g15801 nand P1_R2337_U63 P1_U2376 ; P1_U5839
g15802 nand P1_U2372 P1_R2278_U102 ; P1_U5840
g15803 nand P1_U2365 P1_REIP_REG_8__SCAN_IN ; P1_U5841
g15804 nand P1_R2358_U80 P1_U2364 ; P1_U5842
g15805 nand P1_U5795 P1_PHYADDRPOINTER_REG_8__SCAN_IN ; P1_U5843
g15806 nand P1_R2337_U62 P1_U2376 ; P1_U5844
g15807 nand P1_U2372 P1_R2278_U101 ; P1_U5845
g15808 nand P1_U2365 P1_REIP_REG_9__SCAN_IN ; P1_U5846
g15809 nand P1_R2358_U78 P1_U2364 ; P1_U5847
g15810 nand P1_U5795 P1_PHYADDRPOINTER_REG_9__SCAN_IN ; P1_U5848
g15811 nand P1_R2337_U91 P1_U2376 ; P1_U5849
g15812 nand P1_U2372 P1_R2278_U126 ; P1_U5850
g15813 nand P1_U2365 P1_REIP_REG_10__SCAN_IN ; P1_U5851
g15814 nand P1_R2358_U14 P1_U2364 ; P1_U5852
g15815 nand P1_U5795 P1_PHYADDRPOINTER_REG_10__SCAN_IN ; P1_U5853
g15816 nand P1_R2337_U90 P1_U2376 ; P1_U5854
g15817 nand P1_U2372 P1_R2278_U15 ; P1_U5855
g15818 nand P1_U2365 P1_REIP_REG_11__SCAN_IN ; P1_U5856
g15819 nand P1_R2358_U15 P1_U2364 ; P1_U5857
g15820 nand P1_U5795 P1_PHYADDRPOINTER_REG_11__SCAN_IN ; P1_U5858
g15821 nand P1_R2337_U89 P1_U2376 ; P1_U5859
g15822 nand P1_U2372 P1_R2278_U125 ; P1_U5860
g15823 nand P1_U2365 P1_REIP_REG_12__SCAN_IN ; P1_U5861
g15824 nand P1_R2358_U119 P1_U2364 ; P1_U5862
g15825 nand P1_U5795 P1_PHYADDRPOINTER_REG_12__SCAN_IN ; P1_U5863
g15826 nand P1_R2337_U88 P1_U2376 ; P1_U5864
g15827 nand P1_U2372 P1_R2278_U123 ; P1_U5865
g15828 nand P1_U2365 P1_REIP_REG_13__SCAN_IN ; P1_U5866
g15829 nand P1_R2358_U117 P1_U2364 ; P1_U5867
g15830 nand P1_U5795 P1_PHYADDRPOINTER_REG_13__SCAN_IN ; P1_U5868
g15831 nand P1_R2337_U87 P1_U2376 ; P1_U5869
g15832 nand P1_U2372 P1_R2278_U122 ; P1_U5870
g15833 nand P1_U2365 P1_REIP_REG_14__SCAN_IN ; P1_U5871
g15834 nand P1_R2358_U16 P1_U2364 ; P1_U5872
g15835 nand P1_U5795 P1_PHYADDRPOINTER_REG_14__SCAN_IN ; P1_U5873
g15836 nand P1_R2337_U86 P1_U2376 ; P1_U5874
g15837 nand P1_U2372 P1_R2278_U20 ; P1_U5875
g15838 nand P1_U2365 P1_REIP_REG_15__SCAN_IN ; P1_U5876
g15839 nand P1_R2358_U17 P1_U2364 ; P1_U5877
g15840 nand P1_U5795 P1_PHYADDRPOINTER_REG_15__SCAN_IN ; P1_U5878
g15841 nand P1_R2337_U85 P1_U2376 ; P1_U5879
g15842 nand P1_U2372 P1_R2278_U121 ; P1_U5880
g15843 nand P1_U2365 P1_REIP_REG_16__SCAN_IN ; P1_U5881
g15844 nand P1_R2358_U115 P1_U2364 ; P1_U5882
g15845 nand P1_U5795 P1_PHYADDRPOINTER_REG_16__SCAN_IN ; P1_U5883
g15846 nand P1_R2337_U84 P1_U2376 ; P1_U5884
g15847 nand P1_U2372 P1_R2278_U120 ; P1_U5885
g15848 nand P1_U2365 P1_REIP_REG_17__SCAN_IN ; P1_U5886
g15849 nand P1_R2358_U113 P1_U2364 ; P1_U5887
g15850 nand P1_U5795 P1_PHYADDRPOINTER_REG_17__SCAN_IN ; P1_U5888
g15851 nand P1_R2337_U83 P1_U2376 ; P1_U5889
g15852 nand P1_U2372 P1_R2278_U119 ; P1_U5890
g15853 nand P1_U2365 P1_REIP_REG_18__SCAN_IN ; P1_U5891
g15854 nand P1_R2358_U111 P1_U2364 ; P1_U5892
g15855 nand P1_U5795 P1_PHYADDRPOINTER_REG_18__SCAN_IN ; P1_U5893
g15856 nand P1_R2337_U82 P1_U2376 ; P1_U5894
g15857 nand P1_U2372 P1_R2278_U118 ; P1_U5895
g15858 nand P1_U2365 P1_REIP_REG_19__SCAN_IN ; P1_U5896
g15859 nand P1_R2358_U109 P1_U2364 ; P1_U5897
g15860 nand P1_U5795 P1_PHYADDRPOINTER_REG_19__SCAN_IN ; P1_U5898
g15861 nand P1_R2337_U81 P1_U2376 ; P1_U5899
g15862 nand P1_U2372 P1_R2278_U117 ; P1_U5900
g15863 nand P1_U2365 P1_REIP_REG_20__SCAN_IN ; P1_U5901
g15864 nand P1_R2358_U105 P1_U2364 ; P1_U5902
g15865 nand P1_U5795 P1_PHYADDRPOINTER_REG_20__SCAN_IN ; P1_U5903
g15866 nand P1_R2337_U80 P1_U2376 ; P1_U5904
g15867 nand P1_U2372 P1_R2278_U116 ; P1_U5905
g15868 nand P1_U2365 P1_REIP_REG_21__SCAN_IN ; P1_U5906
g15869 nand P1_R2358_U103 P1_U2364 ; P1_U5907
g15870 nand P1_U5795 P1_PHYADDRPOINTER_REG_21__SCAN_IN ; P1_U5908
g15871 nand P1_R2337_U79 P1_U2376 ; P1_U5909
g15872 nand P1_U2372 P1_R2278_U115 ; P1_U5910
g15873 nand P1_U2365 P1_REIP_REG_22__SCAN_IN ; P1_U5911
g15874 nand P1_R2358_U101 P1_U2364 ; P1_U5912
g15875 nand P1_U5795 P1_PHYADDRPOINTER_REG_22__SCAN_IN ; P1_U5913
g15876 nand P1_R2337_U78 P1_U2376 ; P1_U5914
g15877 nand P1_U2372 P1_R2278_U114 ; P1_U5915
g15878 nand P1_U2365 P1_REIP_REG_23__SCAN_IN ; P1_U5916
g15879 nand P1_R2358_U99 P1_U2364 ; P1_U5917
g15880 nand P1_U5795 P1_PHYADDRPOINTER_REG_23__SCAN_IN ; P1_U5918
g15881 nand P1_R2337_U77 P1_U2376 ; P1_U5919
g15882 nand P1_U2372 P1_R2278_U113 ; P1_U5920
g15883 nand P1_U2365 P1_REIP_REG_24__SCAN_IN ; P1_U5921
g15884 nand P1_R2358_U97 P1_U2364 ; P1_U5922
g15885 nand P1_U5795 P1_PHYADDRPOINTER_REG_24__SCAN_IN ; P1_U5923
g15886 nand P1_R2337_U76 P1_U2376 ; P1_U5924
g15887 nand P1_U2372 P1_R2278_U112 ; P1_U5925
g15888 nand P1_U2365 P1_REIP_REG_25__SCAN_IN ; P1_U5926
g15889 nand P1_R2358_U95 P1_U2364 ; P1_U5927
g15890 nand P1_U5795 P1_PHYADDRPOINTER_REG_25__SCAN_IN ; P1_U5928
g15891 nand P1_R2337_U75 P1_U2376 ; P1_U5929
g15892 nand P1_U2372 P1_R2278_U111 ; P1_U5930
g15893 nand P1_U2365 P1_REIP_REG_26__SCAN_IN ; P1_U5931
g15894 nand P1_R2358_U93 P1_U2364 ; P1_U5932
g15895 nand P1_U5795 P1_PHYADDRPOINTER_REG_26__SCAN_IN ; P1_U5933
g15896 nand P1_R2337_U74 P1_U2376 ; P1_U5934
g15897 nand P1_U2372 P1_R2278_U110 ; P1_U5935
g15898 nand P1_U2365 P1_REIP_REG_27__SCAN_IN ; P1_U5936
g15899 nand P1_R2358_U91 P1_U2364 ; P1_U5937
g15900 nand P1_U5795 P1_PHYADDRPOINTER_REG_27__SCAN_IN ; P1_U5938
g15901 nand P1_R2337_U73 P1_U2376 ; P1_U5939
g15902 nand P1_U2372 P1_R2278_U109 ; P1_U5940
g15903 nand P1_U2365 P1_REIP_REG_28__SCAN_IN ; P1_U5941
g15904 nand P1_R2358_U89 P1_U2364 ; P1_U5942
g15905 nand P1_U5795 P1_PHYADDRPOINTER_REG_28__SCAN_IN ; P1_U5943
g15906 nand P1_R2337_U72 P1_U2376 ; P1_U5944
g15907 nand P1_U2372 P1_R2278_U108 ; P1_U5945
g15908 nand P1_U2365 P1_REIP_REG_29__SCAN_IN ; P1_U5946
g15909 nand P1_R2358_U87 P1_U2364 ; P1_U5947
g15910 nand P1_U5795 P1_PHYADDRPOINTER_REG_29__SCAN_IN ; P1_U5948
g15911 nand P1_R2337_U70 P1_U2376 ; P1_U5949
g15912 nand P1_U2372 P1_R2278_U106 ; P1_U5950
g15913 nand P1_U2365 P1_REIP_REG_30__SCAN_IN ; P1_U5951
g15914 nand P1_R2358_U85 P1_U2364 ; P1_U5952
g15915 nand P1_U5795 P1_PHYADDRPOINTER_REG_30__SCAN_IN ; P1_U5953
g15916 nand P1_R2337_U69 P1_U2376 ; P1_U5954
g15917 nand P1_U2372 P1_R2278_U16 ; P1_U5955
g15918 nand P1_U2365 P1_REIP_REG_31__SCAN_IN ; P1_U5956
g15919 nand P1_R2358_U22 P1_U2364 ; P1_U5957
g15920 nand P1_U5795 P1_PHYADDRPOINTER_REG_31__SCAN_IN ; P1_U5958
g15921 nand U210 P1_U3282 ; P1_U5959
g15922 nand P1_U2382 P1_EAX_REG_15__SCAN_IN ; P1_U5960
g15923 nand U340 P1_U2381 ; P1_U5961
g15924 nand P1_U5961 P1_U5960 ; P1_U5962
g15925 nand P1_U2382 P1_EAX_REG_14__SCAN_IN ; P1_U5963
g15926 nand U341 P1_U2381 ; P1_U5964
g15927 nand P1_U5964 P1_U5963 ; P1_U5965
g15928 nand P1_U2382 P1_EAX_REG_13__SCAN_IN ; P1_U5966
g15929 nand U342 P1_U2381 ; P1_U5967
g15930 nand P1_U5967 P1_U5966 ; P1_U5968
g15931 nand P1_U2382 P1_EAX_REG_12__SCAN_IN ; P1_U5969
g15932 nand U343 P1_U2381 ; P1_U5970
g15933 nand P1_U5970 P1_U5969 ; P1_U5971
g15934 nand P1_U2382 P1_EAX_REG_11__SCAN_IN ; P1_U5972
g15935 nand U344 P1_U2381 ; P1_U5973
g15936 nand P1_U5973 P1_U5972 ; P1_U5974
g15937 nand P1_U2382 P1_EAX_REG_10__SCAN_IN ; P1_U5975
g15938 nand U345 P1_U2381 ; P1_U5976
g15939 nand P1_U5976 P1_U5975 ; P1_U5977
g15940 nand P1_U2382 P1_EAX_REG_9__SCAN_IN ; P1_U5978
g15941 nand U315 P1_U2381 ; P1_U5979
g15942 nand P1_U5979 P1_U5978 ; P1_U5980
g15943 nand P1_U2382 P1_EAX_REG_8__SCAN_IN ; P1_U5981
g15944 nand U316 P1_U2381 ; P1_U5982
g15945 nand P1_U5982 P1_U5981 ; P1_U5983
g15946 nand P1_U2382 P1_EAX_REG_7__SCAN_IN ; P1_U5984
g15947 nand P1_U2381 U317 ; P1_U5985
g15948 nand P1_U5985 P1_U5984 ; P1_U5986
g15949 nand P1_U2382 P1_EAX_REG_6__SCAN_IN ; P1_U5987
g15950 nand P1_U2381 U318 ; P1_U5988
g15951 nand P1_U5988 P1_U5987 ; P1_U5989
g15952 nand P1_U2382 P1_EAX_REG_5__SCAN_IN ; P1_U5990
g15953 nand P1_U2381 U319 ; P1_U5991
g15954 nand P1_U5991 P1_U5990 ; P1_U5992
g15955 nand P1_U2382 P1_EAX_REG_4__SCAN_IN ; P1_U5993
g15956 nand P1_U2381 U320 ; P1_U5994
g15957 nand P1_U5994 P1_U5993 ; P1_U5995
g15958 nand P1_U2382 P1_EAX_REG_3__SCAN_IN ; P1_U5996
g15959 nand P1_U2381 U321 ; P1_U5997
g15960 nand P1_U5997 P1_U5996 ; P1_U5998
g15961 nand P1_U2382 P1_EAX_REG_2__SCAN_IN ; P1_U5999
g15962 nand P1_U2381 U324 ; P1_U6000
g15963 nand P1_U6000 P1_U5999 ; P1_U6001
g15964 nand P1_U2382 P1_EAX_REG_1__SCAN_IN ; P1_U6002
g15965 nand P1_U2381 U335 ; P1_U6003
g15966 nand P1_U6003 P1_U6002 ; P1_U6004
g15967 nand P1_U2382 P1_EAX_REG_0__SCAN_IN ; P1_U6005
g15968 nand P1_U2381 U346 ; P1_U6006
g15969 nand P1_U6006 P1_U6005 ; P1_U6007
g15970 nand P1_U2382 P1_EAX_REG_30__SCAN_IN ; P1_U6008
g15971 nand U341 P1_U2381 ; P1_U6009
g15972 nand P1_U6009 P1_U6008 ; P1_U6010
g15973 nand P1_U2382 P1_EAX_REG_29__SCAN_IN ; P1_U6011
g15974 nand U342 P1_U2381 ; P1_U6012
g15975 nand P1_U6012 P1_U6011 ; P1_U6013
g15976 nand P1_U2382 P1_EAX_REG_28__SCAN_IN ; P1_U6014
g15977 nand U343 P1_U2381 ; P1_U6015
g15978 nand P1_U6015 P1_U6014 ; P1_U6016
g15979 nand P1_U2382 P1_EAX_REG_27__SCAN_IN ; P1_U6017
g15980 nand U344 P1_U2381 ; P1_U6018
g15981 nand P1_U6018 P1_U6017 ; P1_U6019
g15982 nand P1_U2382 P1_EAX_REG_26__SCAN_IN ; P1_U6020
g15983 nand U345 P1_U2381 ; P1_U6021
g15984 nand P1_U6021 P1_U6020 ; P1_U6022
g15985 nand P1_U2382 P1_EAX_REG_25__SCAN_IN ; P1_U6023
g15986 nand U315 P1_U2381 ; P1_U6024
g15987 nand P1_U6024 P1_U6023 ; P1_U6025
g15988 nand P1_U2382 P1_EAX_REG_24__SCAN_IN ; P1_U6026
g15989 nand U316 P1_U2381 ; P1_U6027
g15990 nand P1_U6027 P1_U6026 ; P1_U6028
g15991 nand P1_U2382 P1_EAX_REG_23__SCAN_IN ; P1_U6029
g15992 nand P1_U2381 U317 ; P1_U6030
g15993 nand P1_U6030 P1_U6029 ; P1_U6031
g15994 nand P1_U2382 P1_EAX_REG_22__SCAN_IN ; P1_U6032
g15995 nand P1_U2381 U318 ; P1_U6033
g15996 nand P1_U6033 P1_U6032 ; P1_U6034
g15997 nand P1_U2382 P1_EAX_REG_21__SCAN_IN ; P1_U6035
g15998 nand P1_U2381 U319 ; P1_U6036
g15999 nand P1_U6036 P1_U6035 ; P1_U6037
g16000 nand P1_U2382 P1_EAX_REG_20__SCAN_IN ; P1_U6038
g16001 nand P1_U2381 U320 ; P1_U6039
g16002 nand P1_U6039 P1_U6038 ; P1_U6040
g16003 nand P1_U2382 P1_EAX_REG_19__SCAN_IN ; P1_U6041
g16004 nand P1_U2381 U321 ; P1_U6042
g16005 nand P1_U6042 P1_U6041 ; P1_U6043
g16006 nand P1_U2382 P1_EAX_REG_18__SCAN_IN ; P1_U6044
g16007 nand P1_U2381 U324 ; P1_U6045
g16008 nand P1_U6045 P1_U6044 ; P1_U6046
g16009 nand P1_U2382 P1_EAX_REG_17__SCAN_IN ; P1_U6047
g16010 nand P1_U2381 U335 ; P1_U6048
g16011 nand P1_U6048 P1_U6047 ; P1_U6049
g16012 nand P1_U2382 P1_EAX_REG_16__SCAN_IN ; P1_U6050
g16013 nand P1_U2381 U346 ; P1_U6051
g16014 nand P1_U6051 P1_U6050 ; P1_U6052
g16015 nand P1_U4235 P1_U7606 P1_U4259 ; P1_U6053
g16016 nand P1_U2428 P1_U3294 ; P1_U6054
g16017 not P1_U3417 ; P1_U6055
g16018 nand P1_U2385 P1_LWORD_REG_0__SCAN_IN ; P1_U6056
g16019 nand P1_U2384 P1_EAX_REG_0__SCAN_IN ; P1_U6057
g16020 nand P1_U6055 P1_DATAO_REG_0__SCAN_IN ; P1_U6058
g16021 nand P1_U2385 P1_LWORD_REG_1__SCAN_IN ; P1_U6059
g16022 nand P1_U2384 P1_EAX_REG_1__SCAN_IN ; P1_U6060
g16023 nand P1_U6055 P1_DATAO_REG_1__SCAN_IN ; P1_U6061
g16024 nand P1_U2385 P1_LWORD_REG_2__SCAN_IN ; P1_U6062
g16025 nand P1_U2384 P1_EAX_REG_2__SCAN_IN ; P1_U6063
g16026 nand P1_U6055 P1_DATAO_REG_2__SCAN_IN ; P1_U6064
g16027 nand P1_U2385 P1_LWORD_REG_3__SCAN_IN ; P1_U6065
g16028 nand P1_U2384 P1_EAX_REG_3__SCAN_IN ; P1_U6066
g16029 nand P1_U6055 P1_DATAO_REG_3__SCAN_IN ; P1_U6067
g16030 nand P1_U2385 P1_LWORD_REG_4__SCAN_IN ; P1_U6068
g16031 nand P1_U2384 P1_EAX_REG_4__SCAN_IN ; P1_U6069
g16032 nand P1_U6055 P1_DATAO_REG_4__SCAN_IN ; P1_U6070
g16033 nand P1_U2385 P1_LWORD_REG_5__SCAN_IN ; P1_U6071
g16034 nand P1_U2384 P1_EAX_REG_5__SCAN_IN ; P1_U6072
g16035 nand P1_U6055 P1_DATAO_REG_5__SCAN_IN ; P1_U6073
g16036 nand P1_U2385 P1_LWORD_REG_6__SCAN_IN ; P1_U6074
g16037 nand P1_U2384 P1_EAX_REG_6__SCAN_IN ; P1_U6075
g16038 nand P1_U6055 P1_DATAO_REG_6__SCAN_IN ; P1_U6076
g16039 nand P1_U2385 P1_LWORD_REG_7__SCAN_IN ; P1_U6077
g16040 nand P1_U2384 P1_EAX_REG_7__SCAN_IN ; P1_U6078
g16041 nand P1_U6055 P1_DATAO_REG_7__SCAN_IN ; P1_U6079
g16042 nand P1_U2385 P1_LWORD_REG_8__SCAN_IN ; P1_U6080
g16043 nand P1_U2384 P1_EAX_REG_8__SCAN_IN ; P1_U6081
g16044 nand P1_U6055 P1_DATAO_REG_8__SCAN_IN ; P1_U6082
g16045 nand P1_U2385 P1_LWORD_REG_9__SCAN_IN ; P1_U6083
g16046 nand P1_U2384 P1_EAX_REG_9__SCAN_IN ; P1_U6084
g16047 nand P1_U6055 P1_DATAO_REG_9__SCAN_IN ; P1_U6085
g16048 nand P1_U2385 P1_LWORD_REG_10__SCAN_IN ; P1_U6086
g16049 nand P1_U2384 P1_EAX_REG_10__SCAN_IN ; P1_U6087
g16050 nand P1_U6055 P1_DATAO_REG_10__SCAN_IN ; P1_U6088
g16051 nand P1_U2385 P1_LWORD_REG_11__SCAN_IN ; P1_U6089
g16052 nand P1_U2384 P1_EAX_REG_11__SCAN_IN ; P1_U6090
g16053 nand P1_U6055 P1_DATAO_REG_11__SCAN_IN ; P1_U6091
g16054 nand P1_U2385 P1_LWORD_REG_12__SCAN_IN ; P1_U6092
g16055 nand P1_U2384 P1_EAX_REG_12__SCAN_IN ; P1_U6093
g16056 nand P1_U6055 P1_DATAO_REG_12__SCAN_IN ; P1_U6094
g16057 nand P1_U2385 P1_LWORD_REG_13__SCAN_IN ; P1_U6095
g16058 nand P1_U2384 P1_EAX_REG_13__SCAN_IN ; P1_U6096
g16059 nand P1_U6055 P1_DATAO_REG_13__SCAN_IN ; P1_U6097
g16060 nand P1_U2385 P1_LWORD_REG_14__SCAN_IN ; P1_U6098
g16061 nand P1_U2384 P1_EAX_REG_14__SCAN_IN ; P1_U6099
g16062 nand P1_U6055 P1_DATAO_REG_14__SCAN_IN ; P1_U6100
g16063 nand P1_U2385 P1_LWORD_REG_15__SCAN_IN ; P1_U6101
g16064 nand P1_U2384 P1_EAX_REG_15__SCAN_IN ; P1_U6102
g16065 nand P1_U6055 P1_DATAO_REG_15__SCAN_IN ; P1_U6103
g16066 nand P1_U2424 P1_EAX_REG_16__SCAN_IN ; P1_U6104
g16067 nand P1_U2385 P1_UWORD_REG_0__SCAN_IN ; P1_U6105
g16068 nand P1_U6055 P1_DATAO_REG_16__SCAN_IN ; P1_U6106
g16069 nand P1_U2424 P1_EAX_REG_17__SCAN_IN ; P1_U6107
g16070 nand P1_U2385 P1_UWORD_REG_1__SCAN_IN ; P1_U6108
g16071 nand P1_U6055 P1_DATAO_REG_17__SCAN_IN ; P1_U6109
g16072 nand P1_U2424 P1_EAX_REG_18__SCAN_IN ; P1_U6110
g16073 nand P1_U2385 P1_UWORD_REG_2__SCAN_IN ; P1_U6111
g16074 nand P1_U6055 P1_DATAO_REG_18__SCAN_IN ; P1_U6112
g16075 nand P1_U2424 P1_EAX_REG_19__SCAN_IN ; P1_U6113
g16076 nand P1_U2385 P1_UWORD_REG_3__SCAN_IN ; P1_U6114
g16077 nand P1_U6055 P1_DATAO_REG_19__SCAN_IN ; P1_U6115
g16078 nand P1_U2424 P1_EAX_REG_20__SCAN_IN ; P1_U6116
g16079 nand P1_U2385 P1_UWORD_REG_4__SCAN_IN ; P1_U6117
g16080 nand P1_U6055 P1_DATAO_REG_20__SCAN_IN ; P1_U6118
g16081 nand P1_U2424 P1_EAX_REG_21__SCAN_IN ; P1_U6119
g16082 nand P1_U2385 P1_UWORD_REG_5__SCAN_IN ; P1_U6120
g16083 nand P1_U6055 P1_DATAO_REG_21__SCAN_IN ; P1_U6121
g16084 nand P1_U2424 P1_EAX_REG_22__SCAN_IN ; P1_U6122
g16085 nand P1_U2385 P1_UWORD_REG_6__SCAN_IN ; P1_U6123
g16086 nand P1_U6055 P1_DATAO_REG_22__SCAN_IN ; P1_U6124
g16087 nand P1_U2424 P1_EAX_REG_23__SCAN_IN ; P1_U6125
g16088 nand P1_U2385 P1_UWORD_REG_7__SCAN_IN ; P1_U6126
g16089 nand P1_U6055 P1_DATAO_REG_23__SCAN_IN ; P1_U6127
g16090 nand P1_U2424 P1_EAX_REG_24__SCAN_IN ; P1_U6128
g16091 nand P1_U2385 P1_UWORD_REG_8__SCAN_IN ; P1_U6129
g16092 nand P1_U6055 P1_DATAO_REG_24__SCAN_IN ; P1_U6130
g16093 nand P1_U2424 P1_EAX_REG_25__SCAN_IN ; P1_U6131
g16094 nand P1_U2385 P1_UWORD_REG_9__SCAN_IN ; P1_U6132
g16095 nand P1_U6055 P1_DATAO_REG_25__SCAN_IN ; P1_U6133
g16096 nand P1_U2424 P1_EAX_REG_26__SCAN_IN ; P1_U6134
g16097 nand P1_U2385 P1_UWORD_REG_10__SCAN_IN ; P1_U6135
g16098 nand P1_U6055 P1_DATAO_REG_26__SCAN_IN ; P1_U6136
g16099 nand P1_U2424 P1_EAX_REG_27__SCAN_IN ; P1_U6137
g16100 nand P1_U2385 P1_UWORD_REG_11__SCAN_IN ; P1_U6138
g16101 nand P1_U6055 P1_DATAO_REG_27__SCAN_IN ; P1_U6139
g16102 nand P1_U2424 P1_EAX_REG_28__SCAN_IN ; P1_U6140
g16103 nand P1_U2385 P1_UWORD_REG_12__SCAN_IN ; P1_U6141
g16104 nand P1_U6055 P1_DATAO_REG_28__SCAN_IN ; P1_U6142
g16105 nand P1_U2424 P1_EAX_REG_29__SCAN_IN ; P1_U6143
g16106 nand P1_U2385 P1_UWORD_REG_13__SCAN_IN ; P1_U6144
g16107 nand P1_U6055 P1_DATAO_REG_29__SCAN_IN ; P1_U6145
g16108 nand P1_U2424 P1_EAX_REG_30__SCAN_IN ; P1_U6146
g16109 nand P1_U2385 P1_UWORD_REG_14__SCAN_IN ; P1_U6147
g16110 nand P1_U6055 P1_DATAO_REG_30__SCAN_IN ; P1_U6148
g16111 nand P1_U4194 P1_U2447 P1_GTE_485_U6 ; P1_U6149
g16112 nand P1_U4254 P1_U4197 P1_U4194 ; P1_U6150
g16113 nand P1_U4200 P1_U3283 P1_R2167_U17 ; P1_U6151
g16114 nand P1_U7503 P1_U3257 ; P1_U6152
g16115 nand P1_U3883 P1_U6152 ; P1_U6153
g16116 nand P1_U2422 U346 ; P1_U6154
g16117 nand P1_U2386 P1_R2358_U76 ; P1_U6155
g16118 nand P1_U3424 P1_EAX_REG_0__SCAN_IN ; P1_U6156
g16119 nand P1_U2422 U335 ; P1_U6157
g16120 nand P1_U2386 P1_R2358_U107 ; P1_U6158
g16121 nand P1_U3424 P1_EAX_REG_1__SCAN_IN ; P1_U6159
g16122 nand P1_U2422 U324 ; P1_U6160
g16123 nand P1_U2386 P1_R2358_U18 ; P1_U6161
g16124 nand P1_U3424 P1_EAX_REG_2__SCAN_IN ; P1_U6162
g16125 nand P1_U2422 U321 ; P1_U6163
g16126 nand P1_U2386 P1_R2358_U19 ; P1_U6164
g16127 nand P1_U3424 P1_EAX_REG_3__SCAN_IN ; P1_U6165
g16128 nand P1_U2422 U320 ; P1_U6166
g16129 nand P1_U2386 P1_R2358_U84 ; P1_U6167
g16130 nand P1_U3424 P1_EAX_REG_4__SCAN_IN ; P1_U6168
g16131 nand P1_U2422 U319 ; P1_U6169
g16132 nand P1_U2386 P1_R2358_U82 ; P1_U6170
g16133 nand P1_U3424 P1_EAX_REG_5__SCAN_IN ; P1_U6171
g16134 nand P1_U2422 U318 ; P1_U6172
g16135 nand P1_U2386 P1_R2358_U20 ; P1_U6173
g16136 nand P1_U3424 P1_EAX_REG_6__SCAN_IN ; P1_U6174
g16137 nand P1_U2422 U317 ; P1_U6175
g16138 nand P1_U2386 P1_R2358_U21 ; P1_U6176
g16139 nand P1_U3424 P1_EAX_REG_7__SCAN_IN ; P1_U6177
g16140 nand P1_U2422 U316 ; P1_U6178
g16141 nand P1_U2386 P1_R2358_U80 ; P1_U6179
g16142 nand P1_U3424 P1_EAX_REG_8__SCAN_IN ; P1_U6180
g16143 nand P1_U2422 U315 ; P1_U6181
g16144 nand P1_U2386 P1_R2358_U78 ; P1_U6182
g16145 nand P1_U3424 P1_EAX_REG_9__SCAN_IN ; P1_U6183
g16146 nand P1_U2422 U345 ; P1_U6184
g16147 nand P1_U2386 P1_R2358_U14 ; P1_U6185
g16148 nand P1_U3424 P1_EAX_REG_10__SCAN_IN ; P1_U6186
g16149 nand P1_U2422 U344 ; P1_U6187
g16150 nand P1_U2386 P1_R2358_U15 ; P1_U6188
g16151 nand P1_U3424 P1_EAX_REG_11__SCAN_IN ; P1_U6189
g16152 nand P1_U2422 U343 ; P1_U6190
g16153 nand P1_U2386 P1_R2358_U119 ; P1_U6191
g16154 nand P1_U3424 P1_EAX_REG_12__SCAN_IN ; P1_U6192
g16155 nand P1_U2422 U342 ; P1_U6193
g16156 nand P1_U2386 P1_R2358_U117 ; P1_U6194
g16157 nand P1_U3424 P1_EAX_REG_13__SCAN_IN ; P1_U6195
g16158 nand P1_U2422 U341 ; P1_U6196
g16159 nand P1_U2386 P1_R2358_U16 ; P1_U6197
g16160 nand P1_U3424 P1_EAX_REG_14__SCAN_IN ; P1_U6198
g16161 nand P1_U2422 U340 ; P1_U6199
g16162 nand P1_U2386 P1_R2358_U17 ; P1_U6200
g16163 nand P1_U3424 P1_EAX_REG_15__SCAN_IN ; P1_U6201
g16164 nand P1_U2423 U339 ; P1_U6202
g16165 nand P1_U2387 U346 ; P1_U6203
g16166 nand P1_U2386 P1_R2358_U115 ; P1_U6204
g16167 nand P1_U3424 P1_EAX_REG_16__SCAN_IN ; P1_U6205
g16168 nand P1_U2423 U338 ; P1_U6206
g16169 nand P1_U2387 U335 ; P1_U6207
g16170 nand P1_U2386 P1_R2358_U113 ; P1_U6208
g16171 nand P1_U3424 P1_EAX_REG_17__SCAN_IN ; P1_U6209
g16172 nand P1_U2423 U337 ; P1_U6210
g16173 nand P1_U2387 U324 ; P1_U6211
g16174 nand P1_U2386 P1_R2358_U111 ; P1_U6212
g16175 nand P1_U3424 P1_EAX_REG_18__SCAN_IN ; P1_U6213
g16176 nand P1_U2423 U336 ; P1_U6214
g16177 nand P1_U2387 U321 ; P1_U6215
g16178 nand P1_U2386 P1_R2358_U109 ; P1_U6216
g16179 nand P1_U3424 P1_EAX_REG_19__SCAN_IN ; P1_U6217
g16180 nand P1_U2423 U334 ; P1_U6218
g16181 nand P1_U2387 U320 ; P1_U6219
g16182 nand P1_U2386 P1_R2358_U105 ; P1_U6220
g16183 nand P1_U3424 P1_EAX_REG_20__SCAN_IN ; P1_U6221
g16184 nand P1_U2423 U333 ; P1_U6222
g16185 nand P1_U2387 U319 ; P1_U6223
g16186 nand P1_U2386 P1_R2358_U103 ; P1_U6224
g16187 nand P1_U3424 P1_EAX_REG_21__SCAN_IN ; P1_U6225
g16188 nand P1_U2423 U332 ; P1_U6226
g16189 nand P1_U2387 U318 ; P1_U6227
g16190 nand P1_U2386 P1_R2358_U101 ; P1_U6228
g16191 nand P1_U3424 P1_EAX_REG_22__SCAN_IN ; P1_U6229
g16192 nand P1_U2423 U331 ; P1_U6230
g16193 nand P1_U2387 U317 ; P1_U6231
g16194 nand P1_U2386 P1_R2358_U99 ; P1_U6232
g16195 nand P1_U3424 P1_EAX_REG_23__SCAN_IN ; P1_U6233
g16196 nand P1_U2423 U330 ; P1_U6234
g16197 nand P1_U2387 U316 ; P1_U6235
g16198 nand P1_U2386 P1_R2358_U97 ; P1_U6236
g16199 nand P1_U3424 P1_EAX_REG_24__SCAN_IN ; P1_U6237
g16200 nand P1_U2423 U329 ; P1_U6238
g16201 nand P1_U2387 U315 ; P1_U6239
g16202 nand P1_U2386 P1_R2358_U95 ; P1_U6240
g16203 nand P1_U3424 P1_EAX_REG_25__SCAN_IN ; P1_U6241
g16204 nand P1_U2423 U328 ; P1_U6242
g16205 nand P1_U2387 U345 ; P1_U6243
g16206 nand P1_U2386 P1_R2358_U93 ; P1_U6244
g16207 nand P1_U3424 P1_EAX_REG_26__SCAN_IN ; P1_U6245
g16208 nand P1_U2423 U327 ; P1_U6246
g16209 nand P1_U2387 U344 ; P1_U6247
g16210 nand P1_U2386 P1_R2358_U91 ; P1_U6248
g16211 nand P1_U3424 P1_EAX_REG_27__SCAN_IN ; P1_U6249
g16212 nand P1_U2423 U326 ; P1_U6250
g16213 nand P1_U2387 U343 ; P1_U6251
g16214 nand P1_U2386 P1_R2358_U89 ; P1_U6252
g16215 nand P1_U3424 P1_EAX_REG_28__SCAN_IN ; P1_U6253
g16216 nand P1_U2423 U325 ; P1_U6254
g16217 nand P1_U2387 U342 ; P1_U6255
g16218 nand P1_U2386 P1_R2358_U87 ; P1_U6256
g16219 nand P1_U3424 P1_EAX_REG_29__SCAN_IN ; P1_U6257
g16220 nand P1_U2423 U323 ; P1_U6258
g16221 nand P1_U2387 U341 ; P1_U6259
g16222 nand P1_U2386 P1_R2358_U85 ; P1_U6260
g16223 nand P1_U3424 P1_EAX_REG_30__SCAN_IN ; P1_U6261
g16224 nand P1_U2423 U322 ; P1_U6262
g16225 nand P1_U4198 P1_U3273 ; P1_U6263
g16226 nand P1_U4205 P1_U6263 ; P1_U6264
g16227 nand P1_U2383 P1_R2358_U76 ; P1_U6265
g16228 nand P1_U2371 P1_R2099_U86 ; P1_U6266
g16229 nand P1_U3426 P1_EBX_REG_0__SCAN_IN ; P1_U6267
g16230 nand P1_U2383 P1_R2358_U107 ; P1_U6268
g16231 nand P1_U2371 P1_R2099_U87 ; P1_U6269
g16232 nand P1_U3426 P1_EBX_REG_1__SCAN_IN ; P1_U6270
g16233 nand P1_U2383 P1_R2358_U18 ; P1_U6271
g16234 nand P1_U2371 P1_R2099_U138 ; P1_U6272
g16235 nand P1_U3426 P1_EBX_REG_2__SCAN_IN ; P1_U6273
g16236 nand P1_U2383 P1_R2358_U19 ; P1_U6274
g16237 nand P1_U2371 P1_R2099_U42 ; P1_U6275
g16238 nand P1_U3426 P1_EBX_REG_3__SCAN_IN ; P1_U6276
g16239 nand P1_U2383 P1_R2358_U84 ; P1_U6277
g16240 nand P1_U2371 P1_R2099_U41 ; P1_U6278
g16241 nand P1_U3426 P1_EBX_REG_4__SCAN_IN ; P1_U6279
g16242 nand P1_U2383 P1_R2358_U82 ; P1_U6280
g16243 nand P1_U2371 P1_R2099_U40 ; P1_U6281
g16244 nand P1_U3426 P1_EBX_REG_5__SCAN_IN ; P1_U6282
g16245 nand P1_U2383 P1_R2358_U20 ; P1_U6283
g16246 nand P1_U2371 P1_R2099_U39 ; P1_U6284
g16247 nand P1_U3426 P1_EBX_REG_6__SCAN_IN ; P1_U6285
g16248 nand P1_U2383 P1_R2358_U21 ; P1_U6286
g16249 nand P1_U2371 P1_R2099_U38 ; P1_U6287
g16250 nand P1_U3426 P1_EBX_REG_7__SCAN_IN ; P1_U6288
g16251 nand P1_U2383 P1_R2358_U80 ; P1_U6289
g16252 nand P1_U2371 P1_R2099_U37 ; P1_U6290
g16253 nand P1_U3426 P1_EBX_REG_8__SCAN_IN ; P1_U6291
g16254 nand P1_U2383 P1_R2358_U78 ; P1_U6292
g16255 nand P1_U2371 P1_R2099_U36 ; P1_U6293
g16256 nand P1_U3426 P1_EBX_REG_9__SCAN_IN ; P1_U6294
g16257 nand P1_U2383 P1_R2358_U14 ; P1_U6295
g16258 nand P1_U2371 P1_R2099_U85 ; P1_U6296
g16259 nand P1_U3426 P1_EBX_REG_10__SCAN_IN ; P1_U6297
g16260 nand P1_U2383 P1_R2358_U15 ; P1_U6298
g16261 nand P1_U2371 P1_R2099_U84 ; P1_U6299
g16262 nand P1_U3426 P1_EBX_REG_11__SCAN_IN ; P1_U6300
g16263 nand P1_U2383 P1_R2358_U119 ; P1_U6301
g16264 nand P1_U2371 P1_R2099_U83 ; P1_U6302
g16265 nand P1_U3426 P1_EBX_REG_12__SCAN_IN ; P1_U6303
g16266 nand P1_U2383 P1_R2358_U117 ; P1_U6304
g16267 nand P1_U2371 P1_R2099_U82 ; P1_U6305
g16268 nand P1_U3426 P1_EBX_REG_13__SCAN_IN ; P1_U6306
g16269 nand P1_U2383 P1_R2358_U16 ; P1_U6307
g16270 nand P1_U2371 P1_R2099_U81 ; P1_U6308
g16271 nand P1_U3426 P1_EBX_REG_14__SCAN_IN ; P1_U6309
g16272 nand P1_U2383 P1_R2358_U17 ; P1_U6310
g16273 nand P1_U2371 P1_R2099_U80 ; P1_U6311
g16274 nand P1_U3426 P1_EBX_REG_15__SCAN_IN ; P1_U6312
g16275 nand P1_U2383 P1_R2358_U115 ; P1_U6313
g16276 nand P1_U2371 P1_R2099_U79 ; P1_U6314
g16277 nand P1_U3426 P1_EBX_REG_16__SCAN_IN ; P1_U6315
g16278 nand P1_U2383 P1_R2358_U113 ; P1_U6316
g16279 nand P1_U2371 P1_R2099_U78 ; P1_U6317
g16280 nand P1_U3426 P1_EBX_REG_17__SCAN_IN ; P1_U6318
g16281 nand P1_U2383 P1_R2358_U111 ; P1_U6319
g16282 nand P1_U2371 P1_R2099_U77 ; P1_U6320
g16283 nand P1_U3426 P1_EBX_REG_18__SCAN_IN ; P1_U6321
g16284 nand P1_U2383 P1_R2358_U109 ; P1_U6322
g16285 nand P1_U2371 P1_R2099_U76 ; P1_U6323
g16286 nand P1_U3426 P1_EBX_REG_19__SCAN_IN ; P1_U6324
g16287 nand P1_U2383 P1_R2358_U105 ; P1_U6325
g16288 nand P1_U2371 P1_R2099_U75 ; P1_U6326
g16289 nand P1_U3426 P1_EBX_REG_20__SCAN_IN ; P1_U6327
g16290 nand P1_U2383 P1_R2358_U103 ; P1_U6328
g16291 nand P1_U2371 P1_R2099_U74 ; P1_U6329
g16292 nand P1_U3426 P1_EBX_REG_21__SCAN_IN ; P1_U6330
g16293 nand P1_U2383 P1_R2358_U101 ; P1_U6331
g16294 nand P1_U2371 P1_R2099_U73 ; P1_U6332
g16295 nand P1_U3426 P1_EBX_REG_22__SCAN_IN ; P1_U6333
g16296 nand P1_U2383 P1_R2358_U99 ; P1_U6334
g16297 nand P1_U2371 P1_R2099_U72 ; P1_U6335
g16298 nand P1_U3426 P1_EBX_REG_23__SCAN_IN ; P1_U6336
g16299 nand P1_U2383 P1_R2358_U97 ; P1_U6337
g16300 nand P1_U2371 P1_R2099_U71 ; P1_U6338
g16301 nand P1_U3426 P1_EBX_REG_24__SCAN_IN ; P1_U6339
g16302 nand P1_U2383 P1_R2358_U95 ; P1_U6340
g16303 nand P1_U2371 P1_R2099_U70 ; P1_U6341
g16304 nand P1_U3426 P1_EBX_REG_25__SCAN_IN ; P1_U6342
g16305 nand P1_U2383 P1_R2358_U93 ; P1_U6343
g16306 nand P1_U2371 P1_R2099_U69 ; P1_U6344
g16307 nand P1_U3426 P1_EBX_REG_26__SCAN_IN ; P1_U6345
g16308 nand P1_U2383 P1_R2358_U91 ; P1_U6346
g16309 nand P1_U2371 P1_R2099_U68 ; P1_U6347
g16310 nand P1_U3426 P1_EBX_REG_27__SCAN_IN ; P1_U6348
g16311 nand P1_U2383 P1_R2358_U89 ; P1_U6349
g16312 nand P1_U2371 P1_R2099_U67 ; P1_U6350
g16313 nand P1_U3426 P1_EBX_REG_28__SCAN_IN ; P1_U6351
g16314 nand P1_U2383 P1_R2358_U87 ; P1_U6352
g16315 nand P1_U2371 P1_R2099_U66 ; P1_U6353
g16316 nand P1_U3426 P1_EBX_REG_29__SCAN_IN ; P1_U6354
g16317 nand P1_U2383 P1_R2358_U85 ; P1_U6355
g16318 nand P1_U2371 P1_R2099_U65 ; P1_U6356
g16319 nand P1_U3426 P1_EBX_REG_30__SCAN_IN ; P1_U6357
g16320 nand P1_U2371 P1_R2099_U64 ; P1_U6358
g16321 nand P1_U3426 P1_EBX_REG_31__SCAN_IN ; P1_U6359
g16322 nand P1_U4204 P1_GTE_485_U6 ; P1_U6360
g16323 nand P1_U4202 P1_R2167_U17 ; P1_U6361
g16324 nand P1_U4203 P1_U3263 ; P1_U6362
g16325 not P1_U3431 ; P1_U6363
g16326 nand P1_U4249 P1_STATE2_REG_2__SCAN_IN ; P1_U6364
g16327 nand P1_R2337_U69 P1_STATE2_REG_1__SCAN_IN ; P1_U6365
g16328 nand P1_U6365 P1_U6364 ; P1_U6366
g16329 or U210 P1_STATEBS16_REG_SCAN_IN ; P1_U6367
g16330 nand P1_U2604 P1_R2099_U86 ; P1_U6368
g16331 nand P1_U7485 P1_REIP_REG_0__SCAN_IN ; P1_U6369
g16332 nand P1_U7484 P1_EBX_REG_0__SCAN_IN ; P1_U6370
g16333 nand P1_U2429 P1_R2358_U76 ; P1_U6371
g16334 nand P1_U2426 P1_R2182_U34 ; P1_U6372
g16335 nand P1_U2373 P1_PHYADDRPOINTER_REG_0__SCAN_IN ; P1_U6373
g16336 nand P1_U2366 P1_PHYADDRPOINTER_REG_0__SCAN_IN ; P1_U6374
g16337 nand P1_U6363 P1_REIP_REG_0__SCAN_IN ; P1_U6375
g16338 nand P1_U2604 P1_R2099_U87 ; P1_U6376
g16339 nand P1_R2096_U4 P1_U7485 ; P1_U6377
g16340 nand P1_U7484 P1_EBX_REG_1__SCAN_IN ; P1_U6378
g16341 nand P1_U2429 P1_R2358_U107 ; P1_U6379
g16342 nand P1_U2426 P1_R2182_U33 ; P1_U6380
g16343 nand P1_U2373 P1_PHYADDRPOINTER_REG_1__SCAN_IN ; P1_U6381
g16344 nand P1_U2366 P1_R2337_U4 ; P1_U6382
g16345 nand P1_U6363 P1_REIP_REG_1__SCAN_IN ; P1_U6383
g16346 nand P1_U2604 P1_R2099_U138 ; P1_U6384
g16347 nand P1_R2096_U71 P1_U7485 ; P1_U6385
g16348 nand P1_U7484 P1_EBX_REG_2__SCAN_IN ; P1_U6386
g16349 nand P1_U2429 P1_R2358_U18 ; P1_U6387
g16350 nand P1_U2426 P1_R2182_U42 ; P1_U6388
g16351 nand P1_U2373 P1_PHYADDRPOINTER_REG_2__SCAN_IN ; P1_U6389
g16352 nand P1_U2366 P1_R2337_U71 ; P1_U6390
g16353 nand P1_U6363 P1_REIP_REG_2__SCAN_IN ; P1_U6391
g16354 nand P1_U2604 P1_R2099_U42 ; P1_U6392
g16355 nand P1_R2096_U68 P1_U7485 ; P1_U6393
g16356 nand P1_U7484 P1_EBX_REG_3__SCAN_IN ; P1_U6394
g16357 nand P1_U2429 P1_R2358_U19 ; P1_U6395
g16358 nand P1_U2426 P1_R2182_U25 ; P1_U6396
g16359 nand P1_U2373 P1_PHYADDRPOINTER_REG_3__SCAN_IN ; P1_U6397
g16360 nand P1_U2366 P1_R2337_U68 ; P1_U6398
g16361 nand P1_U6363 P1_REIP_REG_3__SCAN_IN ; P1_U6399
g16362 nand P1_U2604 P1_R2099_U41 ; P1_U6400
g16363 nand P1_R2096_U67 P1_U7485 ; P1_U6401
g16364 nand P1_U7484 P1_EBX_REG_4__SCAN_IN ; P1_U6402
g16365 nand P1_U2429 P1_R2358_U84 ; P1_U6403
g16366 nand P1_U2426 P1_R2182_U24 ; P1_U6404
g16367 nand P1_U2373 P1_PHYADDRPOINTER_REG_4__SCAN_IN ; P1_U6405
g16368 nand P1_U2366 P1_R2337_U67 ; P1_U6406
g16369 nand P1_U6363 P1_REIP_REG_4__SCAN_IN ; P1_U6407
g16370 nand P1_U2604 P1_R2099_U40 ; P1_U6408
g16371 nand P1_R2096_U66 P1_U7485 ; P1_U6409
g16372 nand P1_U7484 P1_EBX_REG_5__SCAN_IN ; P1_U6410
g16373 nand P1_U2429 P1_R2358_U82 ; P1_U6411
g16374 nand P1_R2182_U5 P1_U2426 ; P1_U6412
g16375 nand P1_U2373 P1_PHYADDRPOINTER_REG_5__SCAN_IN ; P1_U6413
g16376 nand P1_U2366 P1_R2337_U66 ; P1_U6414
g16377 nand P1_U6363 P1_REIP_REG_5__SCAN_IN ; P1_U6415
g16378 nand P1_U2604 P1_R2099_U39 ; P1_U6416
g16379 nand P1_R2096_U65 P1_U7485 ; P1_U6417
g16380 nand P1_U7484 P1_EBX_REG_6__SCAN_IN ; P1_U6418
g16381 nand P1_U2373 P1_PHYADDRPOINTER_REG_6__SCAN_IN ; P1_U6419
g16382 nand P1_U2367 P1_R2358_U20 ; P1_U6420
g16383 nand P1_U2366 P1_R2337_U65 ; P1_U6421
g16384 nand P1_U6363 P1_REIP_REG_6__SCAN_IN ; P1_U6422
g16385 nand P1_U2604 P1_R2099_U38 ; P1_U6423
g16386 nand P1_R2096_U64 P1_U7485 ; P1_U6424
g16387 nand P1_U7484 P1_EBX_REG_7__SCAN_IN ; P1_U6425
g16388 nand P1_U2373 P1_PHYADDRPOINTER_REG_7__SCAN_IN ; P1_U6426
g16389 nand P1_U2367 P1_R2358_U21 ; P1_U6427
g16390 nand P1_U2366 P1_R2337_U64 ; P1_U6428
g16391 nand P1_U6363 P1_REIP_REG_7__SCAN_IN ; P1_U6429
g16392 nand P1_U2604 P1_R2099_U37 ; P1_U6430
g16393 nand P1_R2096_U63 P1_U7485 ; P1_U6431
g16394 nand P1_U7484 P1_EBX_REG_8__SCAN_IN ; P1_U6432
g16395 nand P1_U2373 P1_PHYADDRPOINTER_REG_8__SCAN_IN ; P1_U6433
g16396 nand P1_U2367 P1_R2358_U80 ; P1_U6434
g16397 nand P1_U2366 P1_R2337_U63 ; P1_U6435
g16398 nand P1_U6363 P1_REIP_REG_8__SCAN_IN ; P1_U6436
g16399 nand P1_U2604 P1_R2099_U36 ; P1_U6437
g16400 nand P1_R2096_U62 P1_U7485 ; P1_U6438
g16401 nand P1_U7484 P1_EBX_REG_9__SCAN_IN ; P1_U6439
g16402 nand P1_U2373 P1_PHYADDRPOINTER_REG_9__SCAN_IN ; P1_U6440
g16403 nand P1_U2367 P1_R2358_U78 ; P1_U6441
g16404 nand P1_U2366 P1_R2337_U62 ; P1_U6442
g16405 nand P1_U6363 P1_REIP_REG_9__SCAN_IN ; P1_U6443
g16406 nand P1_U2604 P1_R2099_U85 ; P1_U6444
g16407 nand P1_R2096_U91 P1_U7485 ; P1_U6445
g16408 nand P1_U7484 P1_EBX_REG_10__SCAN_IN ; P1_U6446
g16409 nand P1_U2373 P1_PHYADDRPOINTER_REG_10__SCAN_IN ; P1_U6447
g16410 nand P1_U2367 P1_R2358_U14 ; P1_U6448
g16411 nand P1_U2366 P1_R2337_U91 ; P1_U6449
g16412 nand P1_U6363 P1_REIP_REG_10__SCAN_IN ; P1_U6450
g16413 nand P1_U2604 P1_R2099_U84 ; P1_U6451
g16414 nand P1_R2096_U90 P1_U7485 ; P1_U6452
g16415 nand P1_U7484 P1_EBX_REG_11__SCAN_IN ; P1_U6453
g16416 nand P1_U2373 P1_PHYADDRPOINTER_REG_11__SCAN_IN ; P1_U6454
g16417 nand P1_U2367 P1_R2358_U15 ; P1_U6455
g16418 nand P1_U2366 P1_R2337_U90 ; P1_U6456
g16419 nand P1_U6363 P1_REIP_REG_11__SCAN_IN ; P1_U6457
g16420 nand P1_U2604 P1_R2099_U83 ; P1_U6458
g16421 nand P1_R2096_U89 P1_U7485 ; P1_U6459
g16422 nand P1_U7484 P1_EBX_REG_12__SCAN_IN ; P1_U6460
g16423 nand P1_U2373 P1_PHYADDRPOINTER_REG_12__SCAN_IN ; P1_U6461
g16424 nand P1_U2367 P1_R2358_U119 ; P1_U6462
g16425 nand P1_U2366 P1_R2337_U89 ; P1_U6463
g16426 nand P1_U6363 P1_REIP_REG_12__SCAN_IN ; P1_U6464
g16427 nand P1_U2604 P1_R2099_U82 ; P1_U6465
g16428 nand P1_R2096_U88 P1_U7485 ; P1_U6466
g16429 nand P1_U7484 P1_EBX_REG_13__SCAN_IN ; P1_U6467
g16430 nand P1_U2373 P1_PHYADDRPOINTER_REG_13__SCAN_IN ; P1_U6468
g16431 nand P1_U2367 P1_R2358_U117 ; P1_U6469
g16432 nand P1_U2366 P1_R2337_U88 ; P1_U6470
g16433 nand P1_U6363 P1_REIP_REG_13__SCAN_IN ; P1_U6471
g16434 nand P1_U2604 P1_R2099_U81 ; P1_U6472
g16435 nand P1_R2096_U87 P1_U7485 ; P1_U6473
g16436 nand P1_U7484 P1_EBX_REG_14__SCAN_IN ; P1_U6474
g16437 nand P1_U2373 P1_PHYADDRPOINTER_REG_14__SCAN_IN ; P1_U6475
g16438 nand P1_U2367 P1_R2358_U16 ; P1_U6476
g16439 nand P1_U2366 P1_R2337_U87 ; P1_U6477
g16440 nand P1_U6363 P1_REIP_REG_14__SCAN_IN ; P1_U6478
g16441 nand P1_U2604 P1_R2099_U80 ; P1_U6479
g16442 nand P1_R2096_U86 P1_U7485 ; P1_U6480
g16443 nand P1_U7484 P1_EBX_REG_15__SCAN_IN ; P1_U6481
g16444 nand P1_U2373 P1_PHYADDRPOINTER_REG_15__SCAN_IN ; P1_U6482
g16445 nand P1_U2367 P1_R2358_U17 ; P1_U6483
g16446 nand P1_U2366 P1_R2337_U86 ; P1_U6484
g16447 nand P1_U6363 P1_REIP_REG_15__SCAN_IN ; P1_U6485
g16448 nand P1_U2604 P1_R2099_U79 ; P1_U6486
g16449 nand P1_R2096_U85 P1_U7485 ; P1_U6487
g16450 nand P1_U7484 P1_EBX_REG_16__SCAN_IN ; P1_U6488
g16451 nand P1_U2373 P1_PHYADDRPOINTER_REG_16__SCAN_IN ; P1_U6489
g16452 nand P1_U2367 P1_R2358_U115 ; P1_U6490
g16453 nand P1_U2366 P1_R2337_U85 ; P1_U6491
g16454 nand P1_U6363 P1_REIP_REG_16__SCAN_IN ; P1_U6492
g16455 nand P1_U2604 P1_R2099_U78 ; P1_U6493
g16456 nand P1_R2096_U84 P1_U7485 ; P1_U6494
g16457 nand P1_U7484 P1_EBX_REG_17__SCAN_IN ; P1_U6495
g16458 nand P1_U2373 P1_PHYADDRPOINTER_REG_17__SCAN_IN ; P1_U6496
g16459 nand P1_U2367 P1_R2358_U113 ; P1_U6497
g16460 nand P1_U2366 P1_R2337_U84 ; P1_U6498
g16461 nand P1_U6363 P1_REIP_REG_17__SCAN_IN ; P1_U6499
g16462 nand P1_U2604 P1_R2099_U77 ; P1_U6500
g16463 nand P1_R2096_U83 P1_U7485 ; P1_U6501
g16464 nand P1_U7484 P1_EBX_REG_18__SCAN_IN ; P1_U6502
g16465 nand P1_U2373 P1_PHYADDRPOINTER_REG_18__SCAN_IN ; P1_U6503
g16466 nand P1_U2367 P1_R2358_U111 ; P1_U6504
g16467 nand P1_U2366 P1_R2337_U83 ; P1_U6505
g16468 nand P1_U6363 P1_REIP_REG_18__SCAN_IN ; P1_U6506
g16469 nand P1_U2604 P1_R2099_U76 ; P1_U6507
g16470 nand P1_R2096_U82 P1_U7485 ; P1_U6508
g16471 nand P1_U7484 P1_EBX_REG_19__SCAN_IN ; P1_U6509
g16472 nand P1_U2373 P1_PHYADDRPOINTER_REG_19__SCAN_IN ; P1_U6510
g16473 nand P1_U2367 P1_R2358_U109 ; P1_U6511
g16474 nand P1_U2366 P1_R2337_U82 ; P1_U6512
g16475 nand P1_U6363 P1_REIP_REG_19__SCAN_IN ; P1_U6513
g16476 nand P1_U2604 P1_R2099_U75 ; P1_U6514
g16477 nand P1_R2096_U81 P1_U7485 ; P1_U6515
g16478 nand P1_U7484 P1_EBX_REG_20__SCAN_IN ; P1_U6516
g16479 nand P1_U2373 P1_PHYADDRPOINTER_REG_20__SCAN_IN ; P1_U6517
g16480 nand P1_U2367 P1_R2358_U105 ; P1_U6518
g16481 nand P1_U2366 P1_R2337_U81 ; P1_U6519
g16482 nand P1_U6363 P1_REIP_REG_20__SCAN_IN ; P1_U6520
g16483 nand P1_U2604 P1_R2099_U74 ; P1_U6521
g16484 nand P1_R2096_U80 P1_U7485 ; P1_U6522
g16485 nand P1_U7484 P1_EBX_REG_21__SCAN_IN ; P1_U6523
g16486 nand P1_U2373 P1_PHYADDRPOINTER_REG_21__SCAN_IN ; P1_U6524
g16487 nand P1_U2367 P1_R2358_U103 ; P1_U6525
g16488 nand P1_U2366 P1_R2337_U80 ; P1_U6526
g16489 nand P1_U6363 P1_REIP_REG_21__SCAN_IN ; P1_U6527
g16490 nand P1_U2604 P1_R2099_U73 ; P1_U6528
g16491 nand P1_R2096_U79 P1_U7485 ; P1_U6529
g16492 nand P1_U7484 P1_EBX_REG_22__SCAN_IN ; P1_U6530
g16493 nand P1_U2373 P1_PHYADDRPOINTER_REG_22__SCAN_IN ; P1_U6531
g16494 nand P1_U2367 P1_R2358_U101 ; P1_U6532
g16495 nand P1_U2366 P1_R2337_U79 ; P1_U6533
g16496 nand P1_U6363 P1_REIP_REG_22__SCAN_IN ; P1_U6534
g16497 nand P1_U2604 P1_R2099_U72 ; P1_U6535
g16498 nand P1_R2096_U78 P1_U7485 ; P1_U6536
g16499 nand P1_U7484 P1_EBX_REG_23__SCAN_IN ; P1_U6537
g16500 nand P1_U2373 P1_PHYADDRPOINTER_REG_23__SCAN_IN ; P1_U6538
g16501 nand P1_U2367 P1_R2358_U99 ; P1_U6539
g16502 nand P1_U2366 P1_R2337_U78 ; P1_U6540
g16503 nand P1_U6363 P1_REIP_REG_23__SCAN_IN ; P1_U6541
g16504 nand P1_U2604 P1_R2099_U71 ; P1_U6542
g16505 nand P1_R2096_U77 P1_U7485 ; P1_U6543
g16506 nand P1_U7484 P1_EBX_REG_24__SCAN_IN ; P1_U6544
g16507 nand P1_U2373 P1_PHYADDRPOINTER_REG_24__SCAN_IN ; P1_U6545
g16508 nand P1_U2367 P1_R2358_U97 ; P1_U6546
g16509 nand P1_U2366 P1_R2337_U77 ; P1_U6547
g16510 nand P1_U6363 P1_REIP_REG_24__SCAN_IN ; P1_U6548
g16511 nand P1_U2604 P1_R2099_U70 ; P1_U6549
g16512 nand P1_R2096_U76 P1_U7485 ; P1_U6550
g16513 nand P1_U7484 P1_EBX_REG_25__SCAN_IN ; P1_U6551
g16514 nand P1_U2373 P1_PHYADDRPOINTER_REG_25__SCAN_IN ; P1_U6552
g16515 nand P1_U2367 P1_R2358_U95 ; P1_U6553
g16516 nand P1_U2366 P1_R2337_U76 ; P1_U6554
g16517 nand P1_U6363 P1_REIP_REG_25__SCAN_IN ; P1_U6555
g16518 nand P1_U2604 P1_R2099_U69 ; P1_U6556
g16519 nand P1_R2096_U75 P1_U7485 ; P1_U6557
g16520 nand P1_U7484 P1_EBX_REG_26__SCAN_IN ; P1_U6558
g16521 nand P1_U2373 P1_PHYADDRPOINTER_REG_26__SCAN_IN ; P1_U6559
g16522 nand P1_U2367 P1_R2358_U93 ; P1_U6560
g16523 nand P1_U2366 P1_R2337_U75 ; P1_U6561
g16524 nand P1_U6363 P1_REIP_REG_26__SCAN_IN ; P1_U6562
g16525 nand P1_U2604 P1_R2099_U68 ; P1_U6563
g16526 nand P1_R2096_U74 P1_U7485 ; P1_U6564
g16527 nand P1_U7484 P1_EBX_REG_27__SCAN_IN ; P1_U6565
g16528 nand P1_U2373 P1_PHYADDRPOINTER_REG_27__SCAN_IN ; P1_U6566
g16529 nand P1_U2367 P1_R2358_U91 ; P1_U6567
g16530 nand P1_U2366 P1_R2337_U74 ; P1_U6568
g16531 nand P1_U6363 P1_REIP_REG_27__SCAN_IN ; P1_U6569
g16532 nand P1_U2604 P1_R2099_U67 ; P1_U6570
g16533 nand P1_R2096_U73 P1_U7485 ; P1_U6571
g16534 nand P1_U7484 P1_EBX_REG_28__SCAN_IN ; P1_U6572
g16535 nand P1_U2373 P1_PHYADDRPOINTER_REG_28__SCAN_IN ; P1_U6573
g16536 nand P1_U2367 P1_R2358_U89 ; P1_U6574
g16537 nand P1_U2366 P1_R2337_U73 ; P1_U6575
g16538 nand P1_U6363 P1_REIP_REG_28__SCAN_IN ; P1_U6576
g16539 nand P1_U2604 P1_R2099_U66 ; P1_U6577
g16540 nand P1_R2096_U72 P1_U7485 ; P1_U6578
g16541 nand P1_U7484 P1_EBX_REG_29__SCAN_IN ; P1_U6579
g16542 nand P1_U2373 P1_PHYADDRPOINTER_REG_29__SCAN_IN ; P1_U6580
g16543 nand P1_U2367 P1_R2358_U87 ; P1_U6581
g16544 nand P1_U2366 P1_R2337_U72 ; P1_U6582
g16545 nand P1_U6363 P1_REIP_REG_29__SCAN_IN ; P1_U6583
g16546 nand P1_U2604 P1_R2099_U65 ; P1_U6584
g16547 nand P1_R2096_U70 P1_U7485 ; P1_U6585
g16548 nand P1_U7484 P1_EBX_REG_30__SCAN_IN ; P1_U6586
g16549 nand P1_U2373 P1_PHYADDRPOINTER_REG_30__SCAN_IN ; P1_U6587
g16550 nand P1_U2367 P1_R2358_U85 ; P1_U6588
g16551 nand P1_U2366 P1_R2337_U70 ; P1_U6589
g16552 nand P1_U6363 P1_REIP_REG_30__SCAN_IN ; P1_U6590
g16553 nand P1_U2604 P1_R2099_U64 ; P1_U6591
g16554 nand P1_R2096_U69 P1_U7485 ; P1_U6592
g16555 nand P1_U7484 P1_EBX_REG_31__SCAN_IN ; P1_U6593
g16556 nand P1_U2373 P1_PHYADDRPOINTER_REG_31__SCAN_IN ; P1_U6594
g16557 nand P1_U2367 P1_R2358_U22 ; P1_U6595
g16558 nand P1_U2366 P1_R2337_U69 ; P1_U6596
g16559 nand P1_U6363 P1_REIP_REG_31__SCAN_IN ; P1_U6597
g16560 nand P1_DATAWIDTH_REG_0__SCAN_IN P1_DATAWIDTH_REG_1__SCAN_IN ; P1_U6598
g16561 or P1_REIP_REG_0__SCAN_IN P1_REIP_REG_1__SCAN_IN ; P1_U6599
g16562 not P1_U4177 ; P1_U6600
g16563 nand P1_U4177 P1_FLUSH_REG_SCAN_IN ; P1_U6601
g16564 nand P1_U3966 P1_U2428 ; P1_U6602
g16565 not P1_U4180 ; P1_U6603
g16566 nand P1_U4497 P1_STATEBS16_REG_SCAN_IN ; P1_U6604
g16567 nand P1_U4208 P1_U6604 ; P1_U6605
g16568 nand P1_U3964 P1_U6605 ; P1_U6606
g16569 nand P1_U6606 P1_STATE2_REG_0__SCAN_IN ; P1_U6607
g16570 nand P1_U4193 P1_U3272 ; P1_U6608
g16571 nand P1_U3965 P1_U6607 ; P1_U6609
g16572 nand P1_U2368 P1_U2473 ; P1_U6610
g16573 nand P1_U6610 P1_CODEFETCH_REG_SCAN_IN ; P1_U6611
g16574 nand P1_U4255 P1_STATE2_REG_0__SCAN_IN ; P1_U6612
g16575 nand P1_STATE_REG_0__SCAN_IN P1_ADS_N_REG_SCAN_IN ; P1_U6613
g16576 not P1_U4181 ; P1_U6614
g16577 nand P1_U3968 P1_U3291 ; P1_U6615
g16578 nand P1_U4499 P1_U3969 P1_U3406 ; P1_U6616
g16579 nand P1_U6616 P1_MEMORYFETCH_REG_SCAN_IN ; P1_U6617
g16580 nand P1_U2544 P1_INSTQUEUE_REG_15__7__SCAN_IN ; P1_U6618
g16581 nand P1_U2543 P1_INSTQUEUE_REG_14__7__SCAN_IN ; P1_U6619
g16582 nand P1_U2542 P1_INSTQUEUE_REG_13__7__SCAN_IN ; P1_U6620
g16583 nand P1_U2541 P1_INSTQUEUE_REG_12__7__SCAN_IN ; P1_U6621
g16584 nand P1_U2539 P1_INSTQUEUE_REG_11__7__SCAN_IN ; P1_U6622
g16585 nand P1_U2538 P1_INSTQUEUE_REG_10__7__SCAN_IN ; P1_U6623
g16586 nand P1_U2537 P1_INSTQUEUE_REG_9__7__SCAN_IN ; P1_U6624
g16587 nand P1_U2536 P1_INSTQUEUE_REG_8__7__SCAN_IN ; P1_U6625
g16588 nand P1_U2534 P1_INSTQUEUE_REG_7__7__SCAN_IN ; P1_U6626
g16589 nand P1_U2533 P1_INSTQUEUE_REG_6__7__SCAN_IN ; P1_U6627
g16590 nand P1_U2532 P1_INSTQUEUE_REG_5__7__SCAN_IN ; P1_U6628
g16591 nand P1_U2531 P1_INSTQUEUE_REG_4__7__SCAN_IN ; P1_U6629
g16592 nand P1_U2529 P1_INSTQUEUE_REG_3__7__SCAN_IN ; P1_U6630
g16593 nand P1_U2527 P1_INSTQUEUE_REG_2__7__SCAN_IN ; P1_U6631
g16594 nand P1_U2525 P1_INSTQUEUE_REG_1__7__SCAN_IN ; P1_U6632
g16595 nand P1_U2523 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U6633
g16596 nand P1_U2544 P1_INSTQUEUE_REG_15__6__SCAN_IN ; P1_U6634
g16597 nand P1_U2543 P1_INSTQUEUE_REG_14__6__SCAN_IN ; P1_U6635
g16598 nand P1_U2542 P1_INSTQUEUE_REG_13__6__SCAN_IN ; P1_U6636
g16599 nand P1_U2541 P1_INSTQUEUE_REG_12__6__SCAN_IN ; P1_U6637
g16600 nand P1_U2539 P1_INSTQUEUE_REG_11__6__SCAN_IN ; P1_U6638
g16601 nand P1_U2538 P1_INSTQUEUE_REG_10__6__SCAN_IN ; P1_U6639
g16602 nand P1_U2537 P1_INSTQUEUE_REG_9__6__SCAN_IN ; P1_U6640
g16603 nand P1_U2536 P1_INSTQUEUE_REG_8__6__SCAN_IN ; P1_U6641
g16604 nand P1_U2534 P1_INSTQUEUE_REG_7__6__SCAN_IN ; P1_U6642
g16605 nand P1_U2533 P1_INSTQUEUE_REG_6__6__SCAN_IN ; P1_U6643
g16606 nand P1_U2532 P1_INSTQUEUE_REG_5__6__SCAN_IN ; P1_U6644
g16607 nand P1_U2531 P1_INSTQUEUE_REG_4__6__SCAN_IN ; P1_U6645
g16608 nand P1_U2529 P1_INSTQUEUE_REG_3__6__SCAN_IN ; P1_U6646
g16609 nand P1_U2527 P1_INSTQUEUE_REG_2__6__SCAN_IN ; P1_U6647
g16610 nand P1_U2525 P1_INSTQUEUE_REG_1__6__SCAN_IN ; P1_U6648
g16611 nand P1_U2523 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U6649
g16612 nand P1_U2544 P1_INSTQUEUE_REG_15__5__SCAN_IN ; P1_U6650
g16613 nand P1_U2543 P1_INSTQUEUE_REG_14__5__SCAN_IN ; P1_U6651
g16614 nand P1_U2542 P1_INSTQUEUE_REG_13__5__SCAN_IN ; P1_U6652
g16615 nand P1_U2541 P1_INSTQUEUE_REG_12__5__SCAN_IN ; P1_U6653
g16616 nand P1_U2539 P1_INSTQUEUE_REG_11__5__SCAN_IN ; P1_U6654
g16617 nand P1_U2538 P1_INSTQUEUE_REG_10__5__SCAN_IN ; P1_U6655
g16618 nand P1_U2537 P1_INSTQUEUE_REG_9__5__SCAN_IN ; P1_U6656
g16619 nand P1_U2536 P1_INSTQUEUE_REG_8__5__SCAN_IN ; P1_U6657
g16620 nand P1_U2534 P1_INSTQUEUE_REG_7__5__SCAN_IN ; P1_U6658
g16621 nand P1_U2533 P1_INSTQUEUE_REG_6__5__SCAN_IN ; P1_U6659
g16622 nand P1_U2532 P1_INSTQUEUE_REG_5__5__SCAN_IN ; P1_U6660
g16623 nand P1_U2531 P1_INSTQUEUE_REG_4__5__SCAN_IN ; P1_U6661
g16624 nand P1_U2529 P1_INSTQUEUE_REG_3__5__SCAN_IN ; P1_U6662
g16625 nand P1_U2527 P1_INSTQUEUE_REG_2__5__SCAN_IN ; P1_U6663
g16626 nand P1_U2525 P1_INSTQUEUE_REG_1__5__SCAN_IN ; P1_U6664
g16627 nand P1_U2523 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U6665
g16628 nand P1_U2544 P1_INSTQUEUE_REG_15__4__SCAN_IN ; P1_U6666
g16629 nand P1_U2543 P1_INSTQUEUE_REG_14__4__SCAN_IN ; P1_U6667
g16630 nand P1_U2542 P1_INSTQUEUE_REG_13__4__SCAN_IN ; P1_U6668
g16631 nand P1_U2541 P1_INSTQUEUE_REG_12__4__SCAN_IN ; P1_U6669
g16632 nand P1_U2539 P1_INSTQUEUE_REG_11__4__SCAN_IN ; P1_U6670
g16633 nand P1_U2538 P1_INSTQUEUE_REG_10__4__SCAN_IN ; P1_U6671
g16634 nand P1_U2537 P1_INSTQUEUE_REG_9__4__SCAN_IN ; P1_U6672
g16635 nand P1_U2536 P1_INSTQUEUE_REG_8__4__SCAN_IN ; P1_U6673
g16636 nand P1_U2534 P1_INSTQUEUE_REG_7__4__SCAN_IN ; P1_U6674
g16637 nand P1_U2533 P1_INSTQUEUE_REG_6__4__SCAN_IN ; P1_U6675
g16638 nand P1_U2532 P1_INSTQUEUE_REG_5__4__SCAN_IN ; P1_U6676
g16639 nand P1_U2531 P1_INSTQUEUE_REG_4__4__SCAN_IN ; P1_U6677
g16640 nand P1_U2529 P1_INSTQUEUE_REG_3__4__SCAN_IN ; P1_U6678
g16641 nand P1_U2527 P1_INSTQUEUE_REG_2__4__SCAN_IN ; P1_U6679
g16642 nand P1_U2525 P1_INSTQUEUE_REG_1__4__SCAN_IN ; P1_U6680
g16643 nand P1_U2544 P1_INSTQUEUE_REG_15__3__SCAN_IN ; P1_U6681
g16644 nand P1_U2543 P1_INSTQUEUE_REG_14__3__SCAN_IN ; P1_U6682
g16645 nand P1_U2542 P1_INSTQUEUE_REG_13__3__SCAN_IN ; P1_U6683
g16646 nand P1_U2541 P1_INSTQUEUE_REG_12__3__SCAN_IN ; P1_U6684
g16647 nand P1_U2539 P1_INSTQUEUE_REG_11__3__SCAN_IN ; P1_U6685
g16648 nand P1_U2538 P1_INSTQUEUE_REG_10__3__SCAN_IN ; P1_U6686
g16649 nand P1_U2537 P1_INSTQUEUE_REG_9__3__SCAN_IN ; P1_U6687
g16650 nand P1_U2536 P1_INSTQUEUE_REG_8__3__SCAN_IN ; P1_U6688
g16651 nand P1_U2534 P1_INSTQUEUE_REG_7__3__SCAN_IN ; P1_U6689
g16652 nand P1_U2533 P1_INSTQUEUE_REG_6__3__SCAN_IN ; P1_U6690
g16653 nand P1_U2532 P1_INSTQUEUE_REG_5__3__SCAN_IN ; P1_U6691
g16654 nand P1_U2531 P1_INSTQUEUE_REG_4__3__SCAN_IN ; P1_U6692
g16655 nand P1_U2529 P1_INSTQUEUE_REG_3__3__SCAN_IN ; P1_U6693
g16656 nand P1_U2527 P1_INSTQUEUE_REG_2__3__SCAN_IN ; P1_U6694
g16657 nand P1_U2525 P1_INSTQUEUE_REG_1__3__SCAN_IN ; P1_U6695
g16658 nand P1_U2523 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U6696
g16659 nand P1_U2544 P1_INSTQUEUE_REG_15__2__SCAN_IN ; P1_U6697
g16660 nand P1_U2543 P1_INSTQUEUE_REG_14__2__SCAN_IN ; P1_U6698
g16661 nand P1_U2542 P1_INSTQUEUE_REG_13__2__SCAN_IN ; P1_U6699
g16662 nand P1_U2541 P1_INSTQUEUE_REG_12__2__SCAN_IN ; P1_U6700
g16663 nand P1_U2539 P1_INSTQUEUE_REG_11__2__SCAN_IN ; P1_U6701
g16664 nand P1_U2538 P1_INSTQUEUE_REG_10__2__SCAN_IN ; P1_U6702
g16665 nand P1_U2537 P1_INSTQUEUE_REG_9__2__SCAN_IN ; P1_U6703
g16666 nand P1_U2536 P1_INSTQUEUE_REG_8__2__SCAN_IN ; P1_U6704
g16667 nand P1_U2534 P1_INSTQUEUE_REG_7__2__SCAN_IN ; P1_U6705
g16668 nand P1_U2533 P1_INSTQUEUE_REG_6__2__SCAN_IN ; P1_U6706
g16669 nand P1_U2532 P1_INSTQUEUE_REG_5__2__SCAN_IN ; P1_U6707
g16670 nand P1_U2531 P1_INSTQUEUE_REG_4__2__SCAN_IN ; P1_U6708
g16671 nand P1_U2529 P1_INSTQUEUE_REG_3__2__SCAN_IN ; P1_U6709
g16672 nand P1_U2527 P1_INSTQUEUE_REG_2__2__SCAN_IN ; P1_U6710
g16673 nand P1_U2525 P1_INSTQUEUE_REG_1__2__SCAN_IN ; P1_U6711
g16674 nand P1_U2523 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U6712
g16675 nand P1_U2544 P1_INSTQUEUE_REG_15__1__SCAN_IN ; P1_U6713
g16676 nand P1_U2543 P1_INSTQUEUE_REG_14__1__SCAN_IN ; P1_U6714
g16677 nand P1_U2542 P1_INSTQUEUE_REG_13__1__SCAN_IN ; P1_U6715
g16678 nand P1_U2541 P1_INSTQUEUE_REG_12__1__SCAN_IN ; P1_U6716
g16679 nand P1_U2539 P1_INSTQUEUE_REG_11__1__SCAN_IN ; P1_U6717
g16680 nand P1_U2538 P1_INSTQUEUE_REG_10__1__SCAN_IN ; P1_U6718
g16681 nand P1_U2537 P1_INSTQUEUE_REG_9__1__SCAN_IN ; P1_U6719
g16682 nand P1_U2536 P1_INSTQUEUE_REG_8__1__SCAN_IN ; P1_U6720
g16683 nand P1_U2534 P1_INSTQUEUE_REG_7__1__SCAN_IN ; P1_U6721
g16684 nand P1_U2533 P1_INSTQUEUE_REG_6__1__SCAN_IN ; P1_U6722
g16685 nand P1_U2532 P1_INSTQUEUE_REG_5__1__SCAN_IN ; P1_U6723
g16686 nand P1_U2531 P1_INSTQUEUE_REG_4__1__SCAN_IN ; P1_U6724
g16687 nand P1_U2529 P1_INSTQUEUE_REG_3__1__SCAN_IN ; P1_U6725
g16688 nand P1_U2527 P1_INSTQUEUE_REG_2__1__SCAN_IN ; P1_U6726
g16689 nand P1_U2525 P1_INSTQUEUE_REG_1__1__SCAN_IN ; P1_U6727
g16690 nand P1_U2523 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U6728
g16691 nand P1_U2544 P1_INSTQUEUE_REG_15__0__SCAN_IN ; P1_U6729
g16692 nand P1_U2543 P1_INSTQUEUE_REG_14__0__SCAN_IN ; P1_U6730
g16693 nand P1_U2542 P1_INSTQUEUE_REG_13__0__SCAN_IN ; P1_U6731
g16694 nand P1_U2541 P1_INSTQUEUE_REG_12__0__SCAN_IN ; P1_U6732
g16695 nand P1_U2539 P1_INSTQUEUE_REG_11__0__SCAN_IN ; P1_U6733
g16696 nand P1_U2538 P1_INSTQUEUE_REG_10__0__SCAN_IN ; P1_U6734
g16697 nand P1_U2537 P1_INSTQUEUE_REG_9__0__SCAN_IN ; P1_U6735
g16698 nand P1_U2536 P1_INSTQUEUE_REG_8__0__SCAN_IN ; P1_U6736
g16699 nand P1_U2534 P1_INSTQUEUE_REG_7__0__SCAN_IN ; P1_U6737
g16700 nand P1_U2533 P1_INSTQUEUE_REG_6__0__SCAN_IN ; P1_U6738
g16701 nand P1_U2532 P1_INSTQUEUE_REG_5__0__SCAN_IN ; P1_U6739
g16702 nand P1_U2531 P1_INSTQUEUE_REG_4__0__SCAN_IN ; P1_U6740
g16703 nand P1_U2529 P1_INSTQUEUE_REG_3__0__SCAN_IN ; P1_U6741
g16704 nand P1_U2527 P1_INSTQUEUE_REG_2__0__SCAN_IN ; P1_U6742
g16705 nand P1_U2525 P1_INSTQUEUE_REG_1__0__SCAN_IN ; P1_U6743
g16706 nand P1_U2523 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U6744
g16707 nand P1_U4460 P1_STATE2_REG_2__SCAN_IN ; P1_U6745
g16708 nand P1_U3412 P1_U6745 ; P1_U6746
g16709 nand P1_U4188 P1_EAX_REG_9__SCAN_IN ; P1_U6747
g16710 nand P1_U4187 P1_PHYADDRPOINTER_REG_9__SCAN_IN ; P1_U6748
g16711 nand P1_R2337_U62 P1_U2352 ; P1_U6749
g16712 nand P1_U4188 P1_EAX_REG_8__SCAN_IN ; P1_U6750
g16713 nand P1_U4187 P1_PHYADDRPOINTER_REG_8__SCAN_IN ; P1_U6751
g16714 nand P1_R2337_U63 P1_U2352 ; P1_U6752
g16715 nand P1_U4188 P1_EAX_REG_7__SCAN_IN ; P1_U6753
g16716 nand P1_U4187 P1_PHYADDRPOINTER_REG_7__SCAN_IN ; P1_U6754
g16717 nand P1_R2337_U64 P1_U2352 ; P1_U6755
g16718 nand P1_U4188 P1_EAX_REG_6__SCAN_IN ; P1_U6756
g16719 nand P1_U4187 P1_PHYADDRPOINTER_REG_6__SCAN_IN ; P1_U6757
g16720 nand P1_R2337_U65 P1_U2352 ; P1_U6758
g16721 nand P1_R2182_U5 P1_U6746 ; P1_U6759
g16722 nand P1_U4188 P1_EAX_REG_5__SCAN_IN ; P1_U6760
g16723 nand P1_U4187 P1_PHYADDRPOINTER_REG_5__SCAN_IN ; P1_U6761
g16724 nand P1_R2337_U66 P1_U2352 ; P1_U6762
g16725 nand P1_R2182_U24 P1_U6746 ; P1_U6763
g16726 nand P1_U4188 P1_EAX_REG_4__SCAN_IN ; P1_U6764
g16727 nand P1_U4187 P1_PHYADDRPOINTER_REG_4__SCAN_IN ; P1_U6765
g16728 nand P1_R2337_U67 P1_U2352 ; P1_U6766
g16729 nand P1_U2353 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_U6767
g16730 nand P1_U4188 P1_EAX_REG_31__SCAN_IN ; P1_U6768
g16731 nand P1_U4187 P1_PHYADDRPOINTER_REG_31__SCAN_IN ; P1_U6769
g16732 nand P1_R2337_U69 P1_U2352 ; P1_U6770
g16733 nand P1_R2182_U26 P1_U6746 ; P1_U6771
g16734 nand P1_U4188 P1_EAX_REG_30__SCAN_IN ; P1_U6772
g16735 nand P1_U4187 P1_PHYADDRPOINTER_REG_30__SCAN_IN ; P1_U6773
g16736 nand P1_R2337_U70 P1_U2352 ; P1_U6774
g16737 nand P1_R2182_U25 P1_U6746 ; P1_U6775
g16738 nand P1_U4188 P1_EAX_REG_3__SCAN_IN ; P1_U6776
g16739 nand P1_U4187 P1_PHYADDRPOINTER_REG_3__SCAN_IN ; P1_U6777
g16740 nand P1_R2337_U68 P1_U2352 ; P1_U6778
g16741 nand P1_U2353 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U6779
g16742 nand P1_R2182_U27 P1_U6746 ; P1_U6780
g16743 nand P1_U4188 P1_EAX_REG_29__SCAN_IN ; P1_U6781
g16744 nand P1_U4187 P1_PHYADDRPOINTER_REG_29__SCAN_IN ; P1_U6782
g16745 nand P1_R2337_U72 P1_U2352 ; P1_U6783
g16746 nand P1_R2182_U28 P1_U6746 ; P1_U6784
g16747 nand P1_U4188 P1_EAX_REG_28__SCAN_IN ; P1_U6785
g16748 nand P1_U4187 P1_PHYADDRPOINTER_REG_28__SCAN_IN ; P1_U6786
g16749 nand P1_R2337_U73 P1_U2352 ; P1_U6787
g16750 nand P1_R2182_U29 P1_U6746 ; P1_U6788
g16751 nand P1_U4188 P1_EAX_REG_27__SCAN_IN ; P1_U6789
g16752 nand P1_U4187 P1_PHYADDRPOINTER_REG_27__SCAN_IN ; P1_U6790
g16753 nand P1_R2337_U74 P1_U2352 ; P1_U6791
g16754 nand P1_R2182_U30 P1_U6746 ; P1_U6792
g16755 nand P1_U4188 P1_EAX_REG_26__SCAN_IN ; P1_U6793
g16756 nand P1_U4187 P1_PHYADDRPOINTER_REG_26__SCAN_IN ; P1_U6794
g16757 nand P1_R2337_U75 P1_U2352 ; P1_U6795
g16758 nand P1_R2182_U31 P1_U6746 ; P1_U6796
g16759 nand P1_U4188 P1_EAX_REG_25__SCAN_IN ; P1_U6797
g16760 nand P1_U4187 P1_PHYADDRPOINTER_REG_25__SCAN_IN ; P1_U6798
g16761 nand P1_R2337_U76 P1_U2352 ; P1_U6799
g16762 nand P1_R2182_U32 P1_U6746 ; P1_U6800
g16763 nand P1_U4188 P1_EAX_REG_24__SCAN_IN ; P1_U6801
g16764 nand P1_U4187 P1_PHYADDRPOINTER_REG_24__SCAN_IN ; P1_U6802
g16765 nand P1_R2337_U77 P1_U2352 ; P1_U6803
g16766 nand P1_R2182_U6 P1_U6746 ; P1_U6804
g16767 nand P1_U4188 P1_EAX_REG_23__SCAN_IN ; P1_U6805
g16768 nand P1_U4187 P1_PHYADDRPOINTER_REG_23__SCAN_IN ; P1_U6806
g16769 nand P1_R2337_U78 P1_U2352 ; P1_U6807
g16770 nand P1_U2724 P1_U6746 ; P1_U6808
g16771 nand P1_U4188 P1_EAX_REG_22__SCAN_IN ; P1_U6809
g16772 nand P1_U4187 P1_PHYADDRPOINTER_REG_22__SCAN_IN ; P1_U6810
g16773 nand P1_R2337_U79 P1_U2352 ; P1_U6811
g16774 nand P1_U2725 P1_U6746 ; P1_U6812
g16775 nand P1_U4188 P1_EAX_REG_21__SCAN_IN ; P1_U6813
g16776 nand P1_U4187 P1_PHYADDRPOINTER_REG_21__SCAN_IN ; P1_U6814
g16777 nand P1_R2337_U80 P1_U2352 ; P1_U6815
g16778 nand P1_U2726 P1_U6746 ; P1_U6816
g16779 nand P1_U4188 P1_EAX_REG_20__SCAN_IN ; P1_U6817
g16780 nand P1_U4187 P1_PHYADDRPOINTER_REG_20__SCAN_IN ; P1_U6818
g16781 nand P1_R2337_U81 P1_U2352 ; P1_U6819
g16782 nand P1_R2182_U42 P1_U6746 ; P1_U6820
g16783 nand P1_U4188 P1_EAX_REG_2__SCAN_IN ; P1_U6821
g16784 nand P1_U4187 P1_PHYADDRPOINTER_REG_2__SCAN_IN ; P1_U6822
g16785 nand P1_R2337_U71 P1_U2352 ; P1_U6823
g16786 nand P1_U2353 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U6824
g16787 nand P1_U2727 P1_U6746 ; P1_U6825
g16788 nand P1_U4188 P1_EAX_REG_19__SCAN_IN ; P1_U6826
g16789 nand P1_U4187 P1_PHYADDRPOINTER_REG_19__SCAN_IN ; P1_U6827
g16790 nand P1_R2337_U82 P1_U2352 ; P1_U6828
g16791 nand P1_U2728 P1_U6746 ; P1_U6829
g16792 nand P1_U4188 P1_EAX_REG_18__SCAN_IN ; P1_U6830
g16793 nand P1_U4187 P1_PHYADDRPOINTER_REG_18__SCAN_IN ; P1_U6831
g16794 nand P1_R2337_U83 P1_U2352 ; P1_U6832
g16795 nand P1_U2729 P1_U6746 ; P1_U6833
g16796 nand P1_U4188 P1_EAX_REG_17__SCAN_IN ; P1_U6834
g16797 nand P1_U4187 P1_PHYADDRPOINTER_REG_17__SCAN_IN ; P1_U6835
g16798 nand P1_R2337_U84 P1_U2352 ; P1_U6836
g16799 nand P1_U2730 P1_U6746 ; P1_U6837
g16800 nand P1_U4188 P1_EAX_REG_16__SCAN_IN ; P1_U6838
g16801 nand P1_U4187 P1_PHYADDRPOINTER_REG_16__SCAN_IN ; P1_U6839
g16802 nand P1_R2337_U85 P1_U2352 ; P1_U6840
g16803 nand P1_U4188 P1_EAX_REG_15__SCAN_IN ; P1_U6841
g16804 nand P1_U4187 P1_PHYADDRPOINTER_REG_15__SCAN_IN ; P1_U6842
g16805 nand P1_R2337_U86 P1_U2352 ; P1_U6843
g16806 nand P1_U4188 P1_EAX_REG_14__SCAN_IN ; P1_U6844
g16807 nand P1_U4187 P1_PHYADDRPOINTER_REG_14__SCAN_IN ; P1_U6845
g16808 nand P1_R2337_U87 P1_U2352 ; P1_U6846
g16809 nand P1_U4188 P1_EAX_REG_13__SCAN_IN ; P1_U6847
g16810 nand P1_U4187 P1_PHYADDRPOINTER_REG_13__SCAN_IN ; P1_U6848
g16811 nand P1_R2337_U88 P1_U2352 ; P1_U6849
g16812 nand P1_U4188 P1_EAX_REG_12__SCAN_IN ; P1_U6850
g16813 nand P1_U4187 P1_PHYADDRPOINTER_REG_12__SCAN_IN ; P1_U6851
g16814 nand P1_R2337_U89 P1_U2352 ; P1_U6852
g16815 nand P1_U4188 P1_EAX_REG_11__SCAN_IN ; P1_U6853
g16816 nand P1_U4187 P1_PHYADDRPOINTER_REG_11__SCAN_IN ; P1_U6854
g16817 nand P1_R2337_U90 P1_U2352 ; P1_U6855
g16818 nand P1_U4188 P1_EAX_REG_10__SCAN_IN ; P1_U6856
g16819 nand P1_U4187 P1_PHYADDRPOINTER_REG_10__SCAN_IN ; P1_U6857
g16820 nand P1_R2337_U91 P1_U2352 ; P1_U6858
g16821 nand P1_R2182_U33 P1_U6746 ; P1_U6859
g16822 nand P1_U4188 P1_EAX_REG_1__SCAN_IN ; P1_U6860
g16823 nand P1_U4187 P1_PHYADDRPOINTER_REG_1__SCAN_IN ; P1_U6861
g16824 nand P1_R2337_U4 P1_U2352 ; P1_U6862
g16825 nand P1_U2353 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U6863
g16826 nand P1_R2182_U34 P1_U6746 ; P1_U6864
g16827 nand P1_U4188 P1_EAX_REG_0__SCAN_IN ; P1_U6865
g16828 nand P1_U4187 P1_PHYADDRPOINTER_REG_0__SCAN_IN ; P1_U6866
g16829 nand P1_U2352 P1_PHYADDRPOINTER_REG_0__SCAN_IN ; P1_U6867
g16830 nand P1_U2353 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U6868
g16831 nand P1_R2144_U49 P1_U6746 ; P1_U6869
g16832 nand P1_U3439 P1_U4460 P1_U3309 ; P1_U6870
g16833 nand P1_U4159 P1_R2144_U80 ; P1_U6871
g16834 nand P1_ADD_371_U6 P1_U4208 ; P1_U6872
g16835 nand P1_U4159 P1_R2144_U10 ; P1_U6873
g16836 nand P1_ADD_371_U21 P1_U4208 ; P1_U6874
g16837 nand P1_U4159 P1_R2144_U9 ; P1_U6875
g16838 nand P1_ADD_371_U17 P1_U4208 ; P1_U6876
g16839 nand P1_U4159 P1_R2144_U45 ; P1_U6877
g16840 nand P1_ADD_371_U19 P1_U4208 ; P1_U6878
g16841 nand P1_U4159 P1_R2144_U47 ; P1_U6879
g16842 nand P1_ADD_371_U18 P1_U4208 ; P1_U6880
g16843 nand P1_U4159 P1_R2144_U8 ; P1_U6881
g16844 nand P1_ADD_371_U24 P1_U4208 ; P1_U6882
g16845 nand P1_U4159 P1_R2144_U49 ; P1_U6883
g16846 nand P1_ADD_371_U5 P1_U4208 ; P1_U6884
g16847 nand P1_U4494 P1_U3283 ; P1_U6885
g16848 nand P1_U4159 P1_R2144_U50 ; P1_U6886
g16849 nand P1_ADD_371_U20 P1_U4208 ; P1_U6887
g16850 nand P1_U2605 P1_U3284 ; P1_U6888
g16851 nand P1_U4159 P1_R2144_U43 ; P1_U6889
g16852 nand P1_ADD_371_U4 P1_U4208 ; P1_U6890
g16853 nand P1_U4494 P1_U3283 ; P1_U6891
g16854 nand P1_U2564 P1_INSTQUEUE_REG_15__1__SCAN_IN ; P1_U6892
g16855 nand P1_U2563 P1_INSTQUEUE_REG_14__1__SCAN_IN ; P1_U6893
g16856 nand P1_U2562 P1_INSTQUEUE_REG_13__1__SCAN_IN ; P1_U6894
g16857 nand P1_U2561 P1_INSTQUEUE_REG_12__1__SCAN_IN ; P1_U6895
g16858 nand P1_U2559 P1_INSTQUEUE_REG_11__1__SCAN_IN ; P1_U6896
g16859 nand P1_U2558 P1_INSTQUEUE_REG_10__1__SCAN_IN ; P1_U6897
g16860 nand P1_U2557 P1_INSTQUEUE_REG_9__1__SCAN_IN ; P1_U6898
g16861 nand P1_U2556 P1_INSTQUEUE_REG_8__1__SCAN_IN ; P1_U6899
g16862 nand P1_U2554 P1_INSTQUEUE_REG_7__1__SCAN_IN ; P1_U6900
g16863 nand P1_U2553 P1_INSTQUEUE_REG_6__1__SCAN_IN ; P1_U6901
g16864 nand P1_U2552 P1_INSTQUEUE_REG_5__1__SCAN_IN ; P1_U6902
g16865 nand P1_U2551 P1_INSTQUEUE_REG_4__1__SCAN_IN ; P1_U6903
g16866 nand P1_U2549 P1_INSTQUEUE_REG_3__1__SCAN_IN ; P1_U6904
g16867 nand P1_U2548 P1_INSTQUEUE_REG_2__1__SCAN_IN ; P1_U6905
g16868 nand P1_U2547 P1_INSTQUEUE_REG_1__1__SCAN_IN ; P1_U6906
g16869 nand P1_U2546 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U6907
g16870 nand P1_U4032 P1_U4031 P1_U4030 P1_U4029 ; P1_U6908
g16871 nand P1_U3405 P1_U3418 ; P1_U6909
g16872 nand P1_U2564 P1_INSTQUEUE_REG_15__0__SCAN_IN ; P1_U6910
g16873 nand P1_U2563 P1_INSTQUEUE_REG_14__0__SCAN_IN ; P1_U6911
g16874 nand P1_U2562 P1_INSTQUEUE_REG_13__0__SCAN_IN ; P1_U6912
g16875 nand P1_U2561 P1_INSTQUEUE_REG_12__0__SCAN_IN ; P1_U6913
g16876 nand P1_U2559 P1_INSTQUEUE_REG_11__0__SCAN_IN ; P1_U6914
g16877 nand P1_U2558 P1_INSTQUEUE_REG_10__0__SCAN_IN ; P1_U6915
g16878 nand P1_U2557 P1_INSTQUEUE_REG_9__0__SCAN_IN ; P1_U6916
g16879 nand P1_U2556 P1_INSTQUEUE_REG_8__0__SCAN_IN ; P1_U6917
g16880 nand P1_U2554 P1_INSTQUEUE_REG_7__0__SCAN_IN ; P1_U6918
g16881 nand P1_U2553 P1_INSTQUEUE_REG_6__0__SCAN_IN ; P1_U6919
g16882 nand P1_U2552 P1_INSTQUEUE_REG_5__0__SCAN_IN ; P1_U6920
g16883 nand P1_U2551 P1_INSTQUEUE_REG_4__0__SCAN_IN ; P1_U6921
g16884 nand P1_U2549 P1_INSTQUEUE_REG_3__0__SCAN_IN ; P1_U6922
g16885 nand P1_U2548 P1_INSTQUEUE_REG_2__0__SCAN_IN ; P1_U6923
g16886 nand P1_U2547 P1_INSTQUEUE_REG_1__0__SCAN_IN ; P1_U6924
g16887 nand P1_U2546 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U6925
g16888 nand P1_U4036 P1_U4035 P1_U4034 P1_U4033 ; P1_U6926
g16889 nand P1_U4207 P1_U3234 ; P1_U6927
g16890 nand P1_U2355 P1_SUB_357_U8 ; P1_U6928
g16891 nand P1_U4207 P1_U3233 ; P1_U6929
g16892 nand P1_SUB_357_U6 P1_U2355 ; P1_U6930
g16893 nand P1_U4207 P1_U3232 ; P1_U6931
g16894 nand P1_SUB_357_U9 P1_U2355 ; P1_U6932
g16895 nand P1_U4207 P1_U3231 ; P1_U6933
g16896 nand P1_SUB_357_U13 P1_U2355 ; P1_U6934
g16897 nand P1_U4207 P1_U3230 ; P1_U6935
g16898 nand P1_SUB_357_U11 P1_U2355 ; P1_U6936
g16899 nand P1_R2182_U25 P1_U3294 ; P1_U6937
g16900 nand P1_U4207 P1_U3229 ; P1_U6938
g16901 nand P1_SUB_357_U12 P1_U2355 ; P1_U6939
g16902 nand P1_R2182_U42 P1_U3294 ; P1_U6940
g16903 nand P1_U2564 P1_INSTQUEUE_REG_15__7__SCAN_IN ; P1_U6941
g16904 nand P1_U2563 P1_INSTQUEUE_REG_14__7__SCAN_IN ; P1_U6942
g16905 nand P1_U2562 P1_INSTQUEUE_REG_13__7__SCAN_IN ; P1_U6943
g16906 nand P1_U2561 P1_INSTQUEUE_REG_12__7__SCAN_IN ; P1_U6944
g16907 nand P1_U2559 P1_INSTQUEUE_REG_11__7__SCAN_IN ; P1_U6945
g16908 nand P1_U2558 P1_INSTQUEUE_REG_10__7__SCAN_IN ; P1_U6946
g16909 nand P1_U2557 P1_INSTQUEUE_REG_9__7__SCAN_IN ; P1_U6947
g16910 nand P1_U2556 P1_INSTQUEUE_REG_8__7__SCAN_IN ; P1_U6948
g16911 nand P1_U2554 P1_INSTQUEUE_REG_7__7__SCAN_IN ; P1_U6949
g16912 nand P1_U2553 P1_INSTQUEUE_REG_6__7__SCAN_IN ; P1_U6950
g16913 nand P1_U2552 P1_INSTQUEUE_REG_5__7__SCAN_IN ; P1_U6951
g16914 nand P1_U2551 P1_INSTQUEUE_REG_4__7__SCAN_IN ; P1_U6952
g16915 nand P1_U2549 P1_INSTQUEUE_REG_3__7__SCAN_IN ; P1_U6953
g16916 nand P1_U2548 P1_INSTQUEUE_REG_2__7__SCAN_IN ; P1_U6954
g16917 nand P1_U2547 P1_INSTQUEUE_REG_1__7__SCAN_IN ; P1_U6955
g16918 nand P1_U2546 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U6956
g16919 nand P1_U4040 P1_U4039 P1_U4038 P1_U4037 ; P1_U6957
g16920 nand P1_U2564 P1_INSTQUEUE_REG_15__6__SCAN_IN ; P1_U6958
g16921 nand P1_U2563 P1_INSTQUEUE_REG_14__6__SCAN_IN ; P1_U6959
g16922 nand P1_U2562 P1_INSTQUEUE_REG_13__6__SCAN_IN ; P1_U6960
g16923 nand P1_U2561 P1_INSTQUEUE_REG_12__6__SCAN_IN ; P1_U6961
g16924 nand P1_U2559 P1_INSTQUEUE_REG_11__6__SCAN_IN ; P1_U6962
g16925 nand P1_U2558 P1_INSTQUEUE_REG_10__6__SCAN_IN ; P1_U6963
g16926 nand P1_U2557 P1_INSTQUEUE_REG_9__6__SCAN_IN ; P1_U6964
g16927 nand P1_U2556 P1_INSTQUEUE_REG_8__6__SCAN_IN ; P1_U6965
g16928 nand P1_U2554 P1_INSTQUEUE_REG_7__6__SCAN_IN ; P1_U6966
g16929 nand P1_U2553 P1_INSTQUEUE_REG_6__6__SCAN_IN ; P1_U6967
g16930 nand P1_U2552 P1_INSTQUEUE_REG_5__6__SCAN_IN ; P1_U6968
g16931 nand P1_U2551 P1_INSTQUEUE_REG_4__6__SCAN_IN ; P1_U6969
g16932 nand P1_U2549 P1_INSTQUEUE_REG_3__6__SCAN_IN ; P1_U6970
g16933 nand P1_U2548 P1_INSTQUEUE_REG_2__6__SCAN_IN ; P1_U6971
g16934 nand P1_U2547 P1_INSTQUEUE_REG_1__6__SCAN_IN ; P1_U6972
g16935 nand P1_U2546 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U6973
g16936 nand P1_U4044 P1_U4043 P1_U4042 P1_U4041 ; P1_U6974
g16937 nand P1_U2564 P1_INSTQUEUE_REG_15__5__SCAN_IN ; P1_U6975
g16938 nand P1_U2563 P1_INSTQUEUE_REG_14__5__SCAN_IN ; P1_U6976
g16939 nand P1_U2562 P1_INSTQUEUE_REG_13__5__SCAN_IN ; P1_U6977
g16940 nand P1_U2561 P1_INSTQUEUE_REG_12__5__SCAN_IN ; P1_U6978
g16941 nand P1_U2559 P1_INSTQUEUE_REG_11__5__SCAN_IN ; P1_U6979
g16942 nand P1_U2558 P1_INSTQUEUE_REG_10__5__SCAN_IN ; P1_U6980
g16943 nand P1_U2557 P1_INSTQUEUE_REG_9__5__SCAN_IN ; P1_U6981
g16944 nand P1_U2556 P1_INSTQUEUE_REG_8__5__SCAN_IN ; P1_U6982
g16945 nand P1_U2554 P1_INSTQUEUE_REG_7__5__SCAN_IN ; P1_U6983
g16946 nand P1_U2553 P1_INSTQUEUE_REG_6__5__SCAN_IN ; P1_U6984
g16947 nand P1_U2552 P1_INSTQUEUE_REG_5__5__SCAN_IN ; P1_U6985
g16948 nand P1_U2551 P1_INSTQUEUE_REG_4__5__SCAN_IN ; P1_U6986
g16949 nand P1_U2549 P1_INSTQUEUE_REG_3__5__SCAN_IN ; P1_U6987
g16950 nand P1_U2548 P1_INSTQUEUE_REG_2__5__SCAN_IN ; P1_U6988
g16951 nand P1_U2547 P1_INSTQUEUE_REG_1__5__SCAN_IN ; P1_U6989
g16952 nand P1_U2546 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U6990
g16953 nand P1_U4048 P1_U4047 P1_U4046 P1_U4045 ; P1_U6991
g16954 nand P1_U2564 P1_INSTQUEUE_REG_15__4__SCAN_IN ; P1_U6992
g16955 nand P1_U2563 P1_INSTQUEUE_REG_14__4__SCAN_IN ; P1_U6993
g16956 nand P1_U2562 P1_INSTQUEUE_REG_13__4__SCAN_IN ; P1_U6994
g16957 nand P1_U2561 P1_INSTQUEUE_REG_12__4__SCAN_IN ; P1_U6995
g16958 nand P1_U2559 P1_INSTQUEUE_REG_11__4__SCAN_IN ; P1_U6996
g16959 nand P1_U2558 P1_INSTQUEUE_REG_10__4__SCAN_IN ; P1_U6997
g16960 nand P1_U2557 P1_INSTQUEUE_REG_9__4__SCAN_IN ; P1_U6998
g16961 nand P1_U2556 P1_INSTQUEUE_REG_8__4__SCAN_IN ; P1_U6999
g16962 nand P1_U2554 P1_INSTQUEUE_REG_7__4__SCAN_IN ; P1_U7000
g16963 nand P1_U2553 P1_INSTQUEUE_REG_6__4__SCAN_IN ; P1_U7001
g16964 nand P1_U2552 P1_INSTQUEUE_REG_5__4__SCAN_IN ; P1_U7002
g16965 nand P1_U2551 P1_INSTQUEUE_REG_4__4__SCAN_IN ; P1_U7003
g16966 nand P1_U2549 P1_INSTQUEUE_REG_3__4__SCAN_IN ; P1_U7004
g16967 nand P1_U2548 P1_INSTQUEUE_REG_2__4__SCAN_IN ; P1_U7005
g16968 nand P1_U2547 P1_INSTQUEUE_REG_1__4__SCAN_IN ; P1_U7006
g16969 nand P1_U2564 P1_INSTQUEUE_REG_15__3__SCAN_IN ; P1_U7007
g16970 nand P1_U2563 P1_INSTQUEUE_REG_14__3__SCAN_IN ; P1_U7008
g16971 nand P1_U2562 P1_INSTQUEUE_REG_13__3__SCAN_IN ; P1_U7009
g16972 nand P1_U2561 P1_INSTQUEUE_REG_12__3__SCAN_IN ; P1_U7010
g16973 nand P1_U2559 P1_INSTQUEUE_REG_11__3__SCAN_IN ; P1_U7011
g16974 nand P1_U2558 P1_INSTQUEUE_REG_10__3__SCAN_IN ; P1_U7012
g16975 nand P1_U2557 P1_INSTQUEUE_REG_9__3__SCAN_IN ; P1_U7013
g16976 nand P1_U2556 P1_INSTQUEUE_REG_8__3__SCAN_IN ; P1_U7014
g16977 nand P1_U2554 P1_INSTQUEUE_REG_7__3__SCAN_IN ; P1_U7015
g16978 nand P1_U2553 P1_INSTQUEUE_REG_6__3__SCAN_IN ; P1_U7016
g16979 nand P1_U2552 P1_INSTQUEUE_REG_5__3__SCAN_IN ; P1_U7017
g16980 nand P1_U2551 P1_INSTQUEUE_REG_4__3__SCAN_IN ; P1_U7018
g16981 nand P1_U2549 P1_INSTQUEUE_REG_3__3__SCAN_IN ; P1_U7019
g16982 nand P1_U2548 P1_INSTQUEUE_REG_2__3__SCAN_IN ; P1_U7020
g16983 nand P1_U2547 P1_INSTQUEUE_REG_1__3__SCAN_IN ; P1_U7021
g16984 nand P1_U2546 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U7022
g16985 nand P1_U4056 P1_U4055 P1_U4054 P1_U4053 ; P1_U7023
g16986 nand P1_U2564 P1_INSTQUEUE_REG_15__2__SCAN_IN ; P1_U7024
g16987 nand P1_U2563 P1_INSTQUEUE_REG_14__2__SCAN_IN ; P1_U7025
g16988 nand P1_U2562 P1_INSTQUEUE_REG_13__2__SCAN_IN ; P1_U7026
g16989 nand P1_U2561 P1_INSTQUEUE_REG_12__2__SCAN_IN ; P1_U7027
g16990 nand P1_U2559 P1_INSTQUEUE_REG_11__2__SCAN_IN ; P1_U7028
g16991 nand P1_U2558 P1_INSTQUEUE_REG_10__2__SCAN_IN ; P1_U7029
g16992 nand P1_U2557 P1_INSTQUEUE_REG_9__2__SCAN_IN ; P1_U7030
g16993 nand P1_U2556 P1_INSTQUEUE_REG_8__2__SCAN_IN ; P1_U7031
g16994 nand P1_U2554 P1_INSTQUEUE_REG_7__2__SCAN_IN ; P1_U7032
g16995 nand P1_U2553 P1_INSTQUEUE_REG_6__2__SCAN_IN ; P1_U7033
g16996 nand P1_U2552 P1_INSTQUEUE_REG_5__2__SCAN_IN ; P1_U7034
g16997 nand P1_U2551 P1_INSTQUEUE_REG_4__2__SCAN_IN ; P1_U7035
g16998 nand P1_U2549 P1_INSTQUEUE_REG_3__2__SCAN_IN ; P1_U7036
g16999 nand P1_U2548 P1_INSTQUEUE_REG_2__2__SCAN_IN ; P1_U7037
g17000 nand P1_U2547 P1_INSTQUEUE_REG_1__2__SCAN_IN ; P1_U7038
g17001 nand P1_U2546 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U7039
g17002 nand P1_U4060 P1_U4059 P1_U4058 P1_U4057 ; P1_U7040
g17003 nand P1_U4207 P1_U3228 ; P1_U7041
g17004 nand P1_SUB_357_U7 P1_U2355 ; P1_U7042
g17005 nand P1_R2182_U33 P1_U3294 ; P1_U7043
g17006 nand P1_U4207 P1_U3227 ; P1_U7044
g17007 nand P1_SUB_357_U10 P1_U2355 ; P1_U7045
g17008 nand P1_R2182_U34 P1_U3294 ; P1_U7046
g17009 nand P1_U4206 P1_U3234 ; P1_U7047
g17010 nand P1_U4192 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U7048
g17011 nand P1_U4206 P1_U3233 ; P1_U7049
g17012 nand P1_U4192 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U7050
g17013 nand P1_U4206 P1_U3232 ; P1_U7051
g17014 nand P1_U4192 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U7052
g17015 nand P1_U4206 P1_U3231 ; P1_U7053
g17016 nand P1_U4206 P1_U3230 ; P1_U7054
g17017 nand P1_U4192 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U7055
g17018 nand P1_U4206 P1_U3229 ; P1_U7056
g17019 nand P1_U4192 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U7057
g17020 nand P1_U4206 P1_U3228 ; P1_U7058
g17021 nand P1_U4192 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U7059
g17022 nand P1_U4206 P1_U3227 ; P1_U7060
g17023 nand P1_U3234 P1_U4400 ; P1_U7061
g17024 nand P1_U4192 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U7062
g17025 nand P1_U3428 P1_U3427 ; P1_U7063
g17026 nand P1_U3264 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7064
g17027 not P1_U3445 ; P1_U7065
g17028 nand P1_U2582 P1_INSTQUEUE_REG_8__7__SCAN_IN ; P1_U7066
g17029 nand P1_U2581 P1_INSTQUEUE_REG_9__7__SCAN_IN ; P1_U7067
g17030 nand P1_U2580 P1_INSTQUEUE_REG_10__7__SCAN_IN ; P1_U7068
g17031 nand P1_U2579 P1_INSTQUEUE_REG_11__7__SCAN_IN ; P1_U7069
g17032 nand P1_U2577 P1_INSTQUEUE_REG_12__7__SCAN_IN ; P1_U7070
g17033 nand P1_U2576 P1_INSTQUEUE_REG_13__7__SCAN_IN ; P1_U7071
g17034 nand P1_U2575 P1_INSTQUEUE_REG_14__7__SCAN_IN ; P1_U7072
g17035 nand P1_U2574 P1_INSTQUEUE_REG_15__7__SCAN_IN ; P1_U7073
g17036 nand P1_U2573 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U7074
g17037 nand P1_U2572 P1_INSTQUEUE_REG_1__7__SCAN_IN ; P1_U7075
g17038 nand P1_U2571 P1_INSTQUEUE_REG_2__7__SCAN_IN ; P1_U7076
g17039 nand P1_U2570 P1_INSTQUEUE_REG_3__7__SCAN_IN ; P1_U7077
g17040 nand P1_U2568 P1_INSTQUEUE_REG_4__7__SCAN_IN ; P1_U7078
g17041 nand P1_U2567 P1_INSTQUEUE_REG_5__7__SCAN_IN ; P1_U7079
g17042 nand P1_U2566 P1_INSTQUEUE_REG_6__7__SCAN_IN ; P1_U7080
g17043 nand P1_U2565 P1_INSTQUEUE_REG_7__7__SCAN_IN ; P1_U7081
g17044 nand P1_U4066 P1_U4065 P1_U4064 P1_U4063 ; P1_U7082
g17045 nand P1_U3425 P1_U3421 ; P1_U7083
g17046 nand P1_U4073 P1_U4191 ; P1_U7084
g17047 nand P1_U7084 P1_U3422 ; P1_U7085
g17048 nand P1_U4503 P1_U3278 ; P1_U7086
g17049 not P1_U3245 ; P1_U7087
g17050 nand P1_U4400 P1_U4503 P1_U4154 P1_U3394 ; P1_U7088
g17051 nand P1_U4189 P1_STATE2_REG_0__SCAN_IN ; P1_U7089
g17052 nand P1_U4067 P1_U3245 ; P1_U7090
g17053 not P1_U3451 ; P1_U7091
g17054 nand P1_U3451 P1_U5492 P1_U7629 ; P1_U7092
g17055 nand P1_U4194 P1_U7092 ; P1_U7093
g17056 not P1_U3450 ; P1_U7094
g17057 nand P1_U3297 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_U7095
g17058 nand P1_U3450 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7096
g17059 nand P1_U4203 P1_U3360 ; P1_U7097
g17060 nand P1_U2582 P1_INSTQUEUE_REG_8__6__SCAN_IN ; P1_U7098
g17061 nand P1_U2581 P1_INSTQUEUE_REG_9__6__SCAN_IN ; P1_U7099
g17062 nand P1_U2580 P1_INSTQUEUE_REG_10__6__SCAN_IN ; P1_U7100
g17063 nand P1_U2579 P1_INSTQUEUE_REG_11__6__SCAN_IN ; P1_U7101
g17064 nand P1_U2577 P1_INSTQUEUE_REG_12__6__SCAN_IN ; P1_U7102
g17065 nand P1_U2576 P1_INSTQUEUE_REG_13__6__SCAN_IN ; P1_U7103
g17066 nand P1_U2575 P1_INSTQUEUE_REG_14__6__SCAN_IN ; P1_U7104
g17067 nand P1_U2574 P1_INSTQUEUE_REG_15__6__SCAN_IN ; P1_U7105
g17068 nand P1_U2573 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U7106
g17069 nand P1_U2572 P1_INSTQUEUE_REG_1__6__SCAN_IN ; P1_U7107
g17070 nand P1_U2571 P1_INSTQUEUE_REG_2__6__SCAN_IN ; P1_U7108
g17071 nand P1_U2570 P1_INSTQUEUE_REG_3__6__SCAN_IN ; P1_U7109
g17072 nand P1_U2568 P1_INSTQUEUE_REG_4__6__SCAN_IN ; P1_U7110
g17073 nand P1_U2567 P1_INSTQUEUE_REG_5__6__SCAN_IN ; P1_U7111
g17074 nand P1_U2566 P1_INSTQUEUE_REG_6__6__SCAN_IN ; P1_U7112
g17075 nand P1_U2565 P1_INSTQUEUE_REG_7__6__SCAN_IN ; P1_U7113
g17076 nand P1_U4082 P1_U4081 P1_U4080 P1_U4079 ; P1_U7114
g17077 nand P1_U2582 P1_INSTQUEUE_REG_8__5__SCAN_IN ; P1_U7115
g17078 nand P1_U2581 P1_INSTQUEUE_REG_9__5__SCAN_IN ; P1_U7116
g17079 nand P1_U2580 P1_INSTQUEUE_REG_10__5__SCAN_IN ; P1_U7117
g17080 nand P1_U2579 P1_INSTQUEUE_REG_11__5__SCAN_IN ; P1_U7118
g17081 nand P1_U2577 P1_INSTQUEUE_REG_12__5__SCAN_IN ; P1_U7119
g17082 nand P1_U2576 P1_INSTQUEUE_REG_13__5__SCAN_IN ; P1_U7120
g17083 nand P1_U2575 P1_INSTQUEUE_REG_14__5__SCAN_IN ; P1_U7121
g17084 nand P1_U2574 P1_INSTQUEUE_REG_15__5__SCAN_IN ; P1_U7122
g17085 nand P1_U2573 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U7123
g17086 nand P1_U2572 P1_INSTQUEUE_REG_1__5__SCAN_IN ; P1_U7124
g17087 nand P1_U2571 P1_INSTQUEUE_REG_2__5__SCAN_IN ; P1_U7125
g17088 nand P1_U2570 P1_INSTQUEUE_REG_3__5__SCAN_IN ; P1_U7126
g17089 nand P1_U2568 P1_INSTQUEUE_REG_4__5__SCAN_IN ; P1_U7127
g17090 nand P1_U2567 P1_INSTQUEUE_REG_5__5__SCAN_IN ; P1_U7128
g17091 nand P1_U2566 P1_INSTQUEUE_REG_6__5__SCAN_IN ; P1_U7129
g17092 nand P1_U2565 P1_INSTQUEUE_REG_7__5__SCAN_IN ; P1_U7130
g17093 nand P1_U4086 P1_U4085 P1_U4084 P1_U4083 ; P1_U7131
g17094 nand P1_U2582 P1_INSTQUEUE_REG_8__4__SCAN_IN ; P1_U7132
g17095 nand P1_U2581 P1_INSTQUEUE_REG_9__4__SCAN_IN ; P1_U7133
g17096 nand P1_U2580 P1_INSTQUEUE_REG_10__4__SCAN_IN ; P1_U7134
g17097 nand P1_U2579 P1_INSTQUEUE_REG_11__4__SCAN_IN ; P1_U7135
g17098 nand P1_U2577 P1_INSTQUEUE_REG_12__4__SCAN_IN ; P1_U7136
g17099 nand P1_U2576 P1_INSTQUEUE_REG_13__4__SCAN_IN ; P1_U7137
g17100 nand P1_U2575 P1_INSTQUEUE_REG_14__4__SCAN_IN ; P1_U7138
g17101 nand P1_U2574 P1_INSTQUEUE_REG_15__4__SCAN_IN ; P1_U7139
g17102 nand P1_U2572 P1_INSTQUEUE_REG_1__4__SCAN_IN ; P1_U7140
g17103 nand P1_U2571 P1_INSTQUEUE_REG_2__4__SCAN_IN ; P1_U7141
g17104 nand P1_U2570 P1_INSTQUEUE_REG_3__4__SCAN_IN ; P1_U7142
g17105 nand P1_U2568 P1_INSTQUEUE_REG_4__4__SCAN_IN ; P1_U7143
g17106 nand P1_U2567 P1_INSTQUEUE_REG_5__4__SCAN_IN ; P1_U7144
g17107 nand P1_U2566 P1_INSTQUEUE_REG_6__4__SCAN_IN ; P1_U7145
g17108 nand P1_U2565 P1_INSTQUEUE_REG_7__4__SCAN_IN ; P1_U7146
g17109 nand P1_U2582 P1_INSTQUEUE_REG_8__3__SCAN_IN ; P1_U7147
g17110 nand P1_U2581 P1_INSTQUEUE_REG_9__3__SCAN_IN ; P1_U7148
g17111 nand P1_U2580 P1_INSTQUEUE_REG_10__3__SCAN_IN ; P1_U7149
g17112 nand P1_U2579 P1_INSTQUEUE_REG_11__3__SCAN_IN ; P1_U7150
g17113 nand P1_U2577 P1_INSTQUEUE_REG_12__3__SCAN_IN ; P1_U7151
g17114 nand P1_U2576 P1_INSTQUEUE_REG_13__3__SCAN_IN ; P1_U7152
g17115 nand P1_U2575 P1_INSTQUEUE_REG_14__3__SCAN_IN ; P1_U7153
g17116 nand P1_U2574 P1_INSTQUEUE_REG_15__3__SCAN_IN ; P1_U7154
g17117 nand P1_U2573 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U7155
g17118 nand P1_U2572 P1_INSTQUEUE_REG_1__3__SCAN_IN ; P1_U7156
g17119 nand P1_U2571 P1_INSTQUEUE_REG_2__3__SCAN_IN ; P1_U7157
g17120 nand P1_U2570 P1_INSTQUEUE_REG_3__3__SCAN_IN ; P1_U7158
g17121 nand P1_U2568 P1_INSTQUEUE_REG_4__3__SCAN_IN ; P1_U7159
g17122 nand P1_U2567 P1_INSTQUEUE_REG_5__3__SCAN_IN ; P1_U7160
g17123 nand P1_U2566 P1_INSTQUEUE_REG_6__3__SCAN_IN ; P1_U7161
g17124 nand P1_U2565 P1_INSTQUEUE_REG_7__3__SCAN_IN ; P1_U7162
g17125 nand P1_U4095 P1_U4094 P1_U4093 P1_U4092 ; P1_U7163
g17126 nand P1_U2582 P1_INSTQUEUE_REG_8__2__SCAN_IN ; P1_U7164
g17127 nand P1_U2581 P1_INSTQUEUE_REG_9__2__SCAN_IN ; P1_U7165
g17128 nand P1_U2580 P1_INSTQUEUE_REG_10__2__SCAN_IN ; P1_U7166
g17129 nand P1_U2579 P1_INSTQUEUE_REG_11__2__SCAN_IN ; P1_U7167
g17130 nand P1_U2577 P1_INSTQUEUE_REG_12__2__SCAN_IN ; P1_U7168
g17131 nand P1_U2576 P1_INSTQUEUE_REG_13__2__SCAN_IN ; P1_U7169
g17132 nand P1_U2575 P1_INSTQUEUE_REG_14__2__SCAN_IN ; P1_U7170
g17133 nand P1_U2574 P1_INSTQUEUE_REG_15__2__SCAN_IN ; P1_U7171
g17134 nand P1_U2573 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U7172
g17135 nand P1_U2572 P1_INSTQUEUE_REG_1__2__SCAN_IN ; P1_U7173
g17136 nand P1_U2571 P1_INSTQUEUE_REG_2__2__SCAN_IN ; P1_U7174
g17137 nand P1_U2570 P1_INSTQUEUE_REG_3__2__SCAN_IN ; P1_U7175
g17138 nand P1_U2568 P1_INSTQUEUE_REG_4__2__SCAN_IN ; P1_U7176
g17139 nand P1_U2567 P1_INSTQUEUE_REG_5__2__SCAN_IN ; P1_U7177
g17140 nand P1_U2566 P1_INSTQUEUE_REG_6__2__SCAN_IN ; P1_U7178
g17141 nand P1_U2565 P1_INSTQUEUE_REG_7__2__SCAN_IN ; P1_U7179
g17142 nand P1_U4099 P1_U4098 P1_U4097 P1_U4096 ; P1_U7180
g17143 nand P1_U2582 P1_INSTQUEUE_REG_8__1__SCAN_IN ; P1_U7181
g17144 nand P1_U2581 P1_INSTQUEUE_REG_9__1__SCAN_IN ; P1_U7182
g17145 nand P1_U2580 P1_INSTQUEUE_REG_10__1__SCAN_IN ; P1_U7183
g17146 nand P1_U2579 P1_INSTQUEUE_REG_11__1__SCAN_IN ; P1_U7184
g17147 nand P1_U2577 P1_INSTQUEUE_REG_12__1__SCAN_IN ; P1_U7185
g17148 nand P1_U2576 P1_INSTQUEUE_REG_13__1__SCAN_IN ; P1_U7186
g17149 nand P1_U2575 P1_INSTQUEUE_REG_14__1__SCAN_IN ; P1_U7187
g17150 nand P1_U2574 P1_INSTQUEUE_REG_15__1__SCAN_IN ; P1_U7188
g17151 nand P1_U2573 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U7189
g17152 nand P1_U2572 P1_INSTQUEUE_REG_1__1__SCAN_IN ; P1_U7190
g17153 nand P1_U2571 P1_INSTQUEUE_REG_2__1__SCAN_IN ; P1_U7191
g17154 nand P1_U2570 P1_INSTQUEUE_REG_3__1__SCAN_IN ; P1_U7192
g17155 nand P1_U2568 P1_INSTQUEUE_REG_4__1__SCAN_IN ; P1_U7193
g17156 nand P1_U2567 P1_INSTQUEUE_REG_5__1__SCAN_IN ; P1_U7194
g17157 nand P1_U2566 P1_INSTQUEUE_REG_6__1__SCAN_IN ; P1_U7195
g17158 nand P1_U2565 P1_INSTQUEUE_REG_7__1__SCAN_IN ; P1_U7196
g17159 nand P1_U4103 P1_U4102 P1_U4101 P1_U4100 ; P1_U7197
g17160 nand P1_U2582 P1_INSTQUEUE_REG_8__0__SCAN_IN ; P1_U7198
g17161 nand P1_U2581 P1_INSTQUEUE_REG_9__0__SCAN_IN ; P1_U7199
g17162 nand P1_U2580 P1_INSTQUEUE_REG_10__0__SCAN_IN ; P1_U7200
g17163 nand P1_U2579 P1_INSTQUEUE_REG_11__0__SCAN_IN ; P1_U7201
g17164 nand P1_U2577 P1_INSTQUEUE_REG_12__0__SCAN_IN ; P1_U7202
g17165 nand P1_U2576 P1_INSTQUEUE_REG_13__0__SCAN_IN ; P1_U7203
g17166 nand P1_U2575 P1_INSTQUEUE_REG_14__0__SCAN_IN ; P1_U7204
g17167 nand P1_U2574 P1_INSTQUEUE_REG_15__0__SCAN_IN ; P1_U7205
g17168 nand P1_U2573 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U7206
g17169 nand P1_U2572 P1_INSTQUEUE_REG_1__0__SCAN_IN ; P1_U7207
g17170 nand P1_U2571 P1_INSTQUEUE_REG_2__0__SCAN_IN ; P1_U7208
g17171 nand P1_U2570 P1_INSTQUEUE_REG_3__0__SCAN_IN ; P1_U7209
g17172 nand P1_U2568 P1_INSTQUEUE_REG_4__0__SCAN_IN ; P1_U7210
g17173 nand P1_U2567 P1_INSTQUEUE_REG_5__0__SCAN_IN ; P1_U7211
g17174 nand P1_U2566 P1_INSTQUEUE_REG_6__0__SCAN_IN ; P1_U7212
g17175 nand P1_U2565 P1_INSTQUEUE_REG_7__0__SCAN_IN ; P1_U7213
g17176 nand P1_U4107 P1_U4106 P1_U4105 P1_U4104 ; P1_U7214
g17177 nand P1_U3297 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U7215
g17178 nand P1_U4203 P1_U3455 ; P1_U7216
g17179 nand P1_U3297 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_U7217
g17180 nand P1_U4203 P1_U3235 ; P1_U7218
g17181 not P1_U4183 ; P1_U7219
g17182 nand P1_U2602 P1_INSTQUEUE_REG_8__7__SCAN_IN ; P1_U7220
g17183 nand P1_U2601 P1_INSTQUEUE_REG_9__7__SCAN_IN ; P1_U7221
g17184 nand P1_U2600 P1_INSTQUEUE_REG_10__7__SCAN_IN ; P1_U7222
g17185 nand P1_U2599 P1_INSTQUEUE_REG_11__7__SCAN_IN ; P1_U7223
g17186 nand P1_U2597 P1_INSTQUEUE_REG_12__7__SCAN_IN ; P1_U7224
g17187 nand P1_U2596 P1_INSTQUEUE_REG_13__7__SCAN_IN ; P1_U7225
g17188 nand P1_U2595 P1_INSTQUEUE_REG_14__7__SCAN_IN ; P1_U7226
g17189 nand P1_U2594 P1_INSTQUEUE_REG_15__7__SCAN_IN ; P1_U7227
g17190 nand P1_U2592 P1_INSTQUEUE_REG_0__7__SCAN_IN ; P1_U7228
g17191 nand P1_U2591 P1_INSTQUEUE_REG_1__7__SCAN_IN ; P1_U7229
g17192 nand P1_U2590 P1_INSTQUEUE_REG_2__7__SCAN_IN ; P1_U7230
g17193 nand P1_U2589 P1_INSTQUEUE_REG_3__7__SCAN_IN ; P1_U7231
g17194 nand P1_U2587 P1_INSTQUEUE_REG_4__7__SCAN_IN ; P1_U7232
g17195 nand P1_U2586 P1_INSTQUEUE_REG_5__7__SCAN_IN ; P1_U7233
g17196 nand P1_U2585 P1_INSTQUEUE_REG_6__7__SCAN_IN ; P1_U7234
g17197 nand P1_U2584 P1_INSTQUEUE_REG_7__7__SCAN_IN ; P1_U7235
g17198 nand P1_U4124 P1_U4123 P1_U4122 P1_U4121 ; P1_U7236
g17199 nand P1_U2602 P1_INSTQUEUE_REG_8__6__SCAN_IN ; P1_U7237
g17200 nand P1_U2601 P1_INSTQUEUE_REG_9__6__SCAN_IN ; P1_U7238
g17201 nand P1_U2600 P1_INSTQUEUE_REG_10__6__SCAN_IN ; P1_U7239
g17202 nand P1_U2599 P1_INSTQUEUE_REG_11__6__SCAN_IN ; P1_U7240
g17203 nand P1_U2597 P1_INSTQUEUE_REG_12__6__SCAN_IN ; P1_U7241
g17204 nand P1_U2596 P1_INSTQUEUE_REG_13__6__SCAN_IN ; P1_U7242
g17205 nand P1_U2595 P1_INSTQUEUE_REG_14__6__SCAN_IN ; P1_U7243
g17206 nand P1_U2594 P1_INSTQUEUE_REG_15__6__SCAN_IN ; P1_U7244
g17207 nand P1_U2592 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U7245
g17208 nand P1_U2591 P1_INSTQUEUE_REG_1__6__SCAN_IN ; P1_U7246
g17209 nand P1_U2590 P1_INSTQUEUE_REG_2__6__SCAN_IN ; P1_U7247
g17210 nand P1_U2589 P1_INSTQUEUE_REG_3__6__SCAN_IN ; P1_U7248
g17211 nand P1_U2587 P1_INSTQUEUE_REG_4__6__SCAN_IN ; P1_U7249
g17212 nand P1_U2586 P1_INSTQUEUE_REG_5__6__SCAN_IN ; P1_U7250
g17213 nand P1_U2585 P1_INSTQUEUE_REG_6__6__SCAN_IN ; P1_U7251
g17214 nand P1_U2584 P1_INSTQUEUE_REG_7__6__SCAN_IN ; P1_U7252
g17215 nand P1_U4128 P1_U4127 P1_U4126 P1_U4125 ; P1_U7253
g17216 nand P1_U2602 P1_INSTQUEUE_REG_8__5__SCAN_IN ; P1_U7254
g17217 nand P1_U2601 P1_INSTQUEUE_REG_9__5__SCAN_IN ; P1_U7255
g17218 nand P1_U2600 P1_INSTQUEUE_REG_10__5__SCAN_IN ; P1_U7256
g17219 nand P1_U2599 P1_INSTQUEUE_REG_11__5__SCAN_IN ; P1_U7257
g17220 nand P1_U2597 P1_INSTQUEUE_REG_12__5__SCAN_IN ; P1_U7258
g17221 nand P1_U2596 P1_INSTQUEUE_REG_13__5__SCAN_IN ; P1_U7259
g17222 nand P1_U2595 P1_INSTQUEUE_REG_14__5__SCAN_IN ; P1_U7260
g17223 nand P1_U2594 P1_INSTQUEUE_REG_15__5__SCAN_IN ; P1_U7261
g17224 nand P1_U2592 P1_INSTQUEUE_REG_0__5__SCAN_IN ; P1_U7262
g17225 nand P1_U2591 P1_INSTQUEUE_REG_1__5__SCAN_IN ; P1_U7263
g17226 nand P1_U2590 P1_INSTQUEUE_REG_2__5__SCAN_IN ; P1_U7264
g17227 nand P1_U2589 P1_INSTQUEUE_REG_3__5__SCAN_IN ; P1_U7265
g17228 nand P1_U2587 P1_INSTQUEUE_REG_4__5__SCAN_IN ; P1_U7266
g17229 nand P1_U2586 P1_INSTQUEUE_REG_5__5__SCAN_IN ; P1_U7267
g17230 nand P1_U2585 P1_INSTQUEUE_REG_6__5__SCAN_IN ; P1_U7268
g17231 nand P1_U2584 P1_INSTQUEUE_REG_7__5__SCAN_IN ; P1_U7269
g17232 nand P1_U4132 P1_U4131 P1_U4130 P1_U4129 ; P1_U7270
g17233 nand P1_U2602 P1_INSTQUEUE_REG_8__4__SCAN_IN ; P1_U7271
g17234 nand P1_U2601 P1_INSTQUEUE_REG_9__4__SCAN_IN ; P1_U7272
g17235 nand P1_U2600 P1_INSTQUEUE_REG_10__4__SCAN_IN ; P1_U7273
g17236 nand P1_U2599 P1_INSTQUEUE_REG_11__4__SCAN_IN ; P1_U7274
g17237 nand P1_U2597 P1_INSTQUEUE_REG_12__4__SCAN_IN ; P1_U7275
g17238 nand P1_U2596 P1_INSTQUEUE_REG_13__4__SCAN_IN ; P1_U7276
g17239 nand P1_U2595 P1_INSTQUEUE_REG_14__4__SCAN_IN ; P1_U7277
g17240 nand P1_U2594 P1_INSTQUEUE_REG_15__4__SCAN_IN ; P1_U7278
g17241 nand P1_U2591 P1_INSTQUEUE_REG_1__4__SCAN_IN ; P1_U7279
g17242 nand P1_U2590 P1_INSTQUEUE_REG_2__4__SCAN_IN ; P1_U7280
g17243 nand P1_U2589 P1_INSTQUEUE_REG_3__4__SCAN_IN ; P1_U7281
g17244 nand P1_U2587 P1_INSTQUEUE_REG_4__4__SCAN_IN ; P1_U7282
g17245 nand P1_U2586 P1_INSTQUEUE_REG_5__4__SCAN_IN ; P1_U7283
g17246 nand P1_U2585 P1_INSTQUEUE_REG_6__4__SCAN_IN ; P1_U7284
g17247 nand P1_U2584 P1_INSTQUEUE_REG_7__4__SCAN_IN ; P1_U7285
g17248 nand P1_U2602 P1_INSTQUEUE_REG_8__3__SCAN_IN ; P1_U7286
g17249 nand P1_U2601 P1_INSTQUEUE_REG_9__3__SCAN_IN ; P1_U7287
g17250 nand P1_U2600 P1_INSTQUEUE_REG_10__3__SCAN_IN ; P1_U7288
g17251 nand P1_U2599 P1_INSTQUEUE_REG_11__3__SCAN_IN ; P1_U7289
g17252 nand P1_U2597 P1_INSTQUEUE_REG_12__3__SCAN_IN ; P1_U7290
g17253 nand P1_U2596 P1_INSTQUEUE_REG_13__3__SCAN_IN ; P1_U7291
g17254 nand P1_U2595 P1_INSTQUEUE_REG_14__3__SCAN_IN ; P1_U7292
g17255 nand P1_U2594 P1_INSTQUEUE_REG_15__3__SCAN_IN ; P1_U7293
g17256 nand P1_U2592 P1_INSTQUEUE_REG_0__3__SCAN_IN ; P1_U7294
g17257 nand P1_U2591 P1_INSTQUEUE_REG_1__3__SCAN_IN ; P1_U7295
g17258 nand P1_U2590 P1_INSTQUEUE_REG_2__3__SCAN_IN ; P1_U7296
g17259 nand P1_U2589 P1_INSTQUEUE_REG_3__3__SCAN_IN ; P1_U7297
g17260 nand P1_U2587 P1_INSTQUEUE_REG_4__3__SCAN_IN ; P1_U7298
g17261 nand P1_U2586 P1_INSTQUEUE_REG_5__3__SCAN_IN ; P1_U7299
g17262 nand P1_U2585 P1_INSTQUEUE_REG_6__3__SCAN_IN ; P1_U7300
g17263 nand P1_U2584 P1_INSTQUEUE_REG_7__3__SCAN_IN ; P1_U7301
g17264 nand P1_U4140 P1_U4139 P1_U4138 P1_U4137 ; P1_U7302
g17265 nand P1_U2602 P1_INSTQUEUE_REG_8__2__SCAN_IN ; P1_U7303
g17266 nand P1_U2601 P1_INSTQUEUE_REG_9__2__SCAN_IN ; P1_U7304
g17267 nand P1_U2600 P1_INSTQUEUE_REG_10__2__SCAN_IN ; P1_U7305
g17268 nand P1_U2599 P1_INSTQUEUE_REG_11__2__SCAN_IN ; P1_U7306
g17269 nand P1_U2597 P1_INSTQUEUE_REG_12__2__SCAN_IN ; P1_U7307
g17270 nand P1_U2596 P1_INSTQUEUE_REG_13__2__SCAN_IN ; P1_U7308
g17271 nand P1_U2595 P1_INSTQUEUE_REG_14__2__SCAN_IN ; P1_U7309
g17272 nand P1_U2594 P1_INSTQUEUE_REG_15__2__SCAN_IN ; P1_U7310
g17273 nand P1_U2592 P1_INSTQUEUE_REG_0__2__SCAN_IN ; P1_U7311
g17274 nand P1_U2591 P1_INSTQUEUE_REG_1__2__SCAN_IN ; P1_U7312
g17275 nand P1_U2590 P1_INSTQUEUE_REG_2__2__SCAN_IN ; P1_U7313
g17276 nand P1_U2589 P1_INSTQUEUE_REG_3__2__SCAN_IN ; P1_U7314
g17277 nand P1_U2587 P1_INSTQUEUE_REG_4__2__SCAN_IN ; P1_U7315
g17278 nand P1_U2586 P1_INSTQUEUE_REG_5__2__SCAN_IN ; P1_U7316
g17279 nand P1_U2585 P1_INSTQUEUE_REG_6__2__SCAN_IN ; P1_U7317
g17280 nand P1_U2584 P1_INSTQUEUE_REG_7__2__SCAN_IN ; P1_U7318
g17281 nand P1_U4144 P1_U4143 P1_U4142 P1_U4141 ; P1_U7319
g17282 nand P1_U2602 P1_INSTQUEUE_REG_8__1__SCAN_IN ; P1_U7320
g17283 nand P1_U2601 P1_INSTQUEUE_REG_9__1__SCAN_IN ; P1_U7321
g17284 nand P1_U2600 P1_INSTQUEUE_REG_10__1__SCAN_IN ; P1_U7322
g17285 nand P1_U2599 P1_INSTQUEUE_REG_11__1__SCAN_IN ; P1_U7323
g17286 nand P1_U2597 P1_INSTQUEUE_REG_12__1__SCAN_IN ; P1_U7324
g17287 nand P1_U2596 P1_INSTQUEUE_REG_13__1__SCAN_IN ; P1_U7325
g17288 nand P1_U2595 P1_INSTQUEUE_REG_14__1__SCAN_IN ; P1_U7326
g17289 nand P1_U2594 P1_INSTQUEUE_REG_15__1__SCAN_IN ; P1_U7327
g17290 nand P1_U2592 P1_INSTQUEUE_REG_0__1__SCAN_IN ; P1_U7328
g17291 nand P1_U2591 P1_INSTQUEUE_REG_1__1__SCAN_IN ; P1_U7329
g17292 nand P1_U2590 P1_INSTQUEUE_REG_2__1__SCAN_IN ; P1_U7330
g17293 nand P1_U2589 P1_INSTQUEUE_REG_3__1__SCAN_IN ; P1_U7331
g17294 nand P1_U2587 P1_INSTQUEUE_REG_4__1__SCAN_IN ; P1_U7332
g17295 nand P1_U2586 P1_INSTQUEUE_REG_5__1__SCAN_IN ; P1_U7333
g17296 nand P1_U2585 P1_INSTQUEUE_REG_6__1__SCAN_IN ; P1_U7334
g17297 nand P1_U2584 P1_INSTQUEUE_REG_7__1__SCAN_IN ; P1_U7335
g17298 nand P1_U4148 P1_U4147 P1_U4146 P1_U4145 ; P1_U7336
g17299 nand P1_U2602 P1_INSTQUEUE_REG_8__0__SCAN_IN ; P1_U7337
g17300 nand P1_U2601 P1_INSTQUEUE_REG_9__0__SCAN_IN ; P1_U7338
g17301 nand P1_U2600 P1_INSTQUEUE_REG_10__0__SCAN_IN ; P1_U7339
g17302 nand P1_U2599 P1_INSTQUEUE_REG_11__0__SCAN_IN ; P1_U7340
g17303 nand P1_U2597 P1_INSTQUEUE_REG_12__0__SCAN_IN ; P1_U7341
g17304 nand P1_U2596 P1_INSTQUEUE_REG_13__0__SCAN_IN ; P1_U7342
g17305 nand P1_U2595 P1_INSTQUEUE_REG_14__0__SCAN_IN ; P1_U7343
g17306 nand P1_U2594 P1_INSTQUEUE_REG_15__0__SCAN_IN ; P1_U7344
g17307 nand P1_U2592 P1_INSTQUEUE_REG_0__0__SCAN_IN ; P1_U7345
g17308 nand P1_U2591 P1_INSTQUEUE_REG_1__0__SCAN_IN ; P1_U7346
g17309 nand P1_U2590 P1_INSTQUEUE_REG_2__0__SCAN_IN ; P1_U7347
g17310 nand P1_U2589 P1_INSTQUEUE_REG_3__0__SCAN_IN ; P1_U7348
g17311 nand P1_U2587 P1_INSTQUEUE_REG_4__0__SCAN_IN ; P1_U7349
g17312 nand P1_U2586 P1_INSTQUEUE_REG_5__0__SCAN_IN ; P1_U7350
g17313 nand P1_U2585 P1_INSTQUEUE_REG_6__0__SCAN_IN ; P1_U7351
g17314 nand P1_U2584 P1_INSTQUEUE_REG_7__0__SCAN_IN ; P1_U7352
g17315 nand P1_U4152 P1_U4151 P1_U4150 P1_U4149 ; P1_U7353
g17316 nand P1_U4231 P1_U2354 P1_U4234 ; P1_U7354
g17317 nand P1_U4153 P1_U7087 ; P1_U7355
g17318 nand P1_U3396 P1_U3410 ; P1_U7356
g17319 nand P1_U4234 P1_U7356 ; P1_U7357
g17320 nand P1_U4190 P1_U2452 ; P1_U7358
g17321 nand P1_U7355 P1_U3271 ; P1_U7359
g17322 nand P1_U4208 P1_U7088 ; P1_U7360
g17323 nand P1_U4160 P1_U4208 ; P1_U7361
g17324 nand P1_U2451 P1_U4210 ; P1_U7362
g17325 nand P1_U3420 P1_U3434 P1_U4195 P1_U7362 P1_U7361 ; P1_U7363
g17326 nand P1_R2238_U6 P1_U7363 ; P1_U7364
g17327 nand P1_SUB_450_U6 P1_U2354 ; P1_U7365
g17328 nand P1_R2238_U19 P1_U7363 ; P1_U7366
g17329 nand P1_SUB_450_U19 P1_U2354 ; P1_U7367
g17330 nand P1_R2238_U20 P1_U7363 ; P1_U7368
g17331 nand P1_SUB_450_U20 P1_U2354 ; P1_U7369
g17332 nand P1_R2238_U21 P1_U7363 ; P1_U7370
g17333 nand P1_SUB_450_U21 P1_U2354 ; P1_U7371
g17334 nand P1_R2238_U22 P1_U7363 ; P1_U7372
g17335 nand P1_SUB_450_U22 P1_U2354 ; P1_U7373
g17336 nand P1_R2238_U7 P1_U7363 ; P1_U7374
g17337 nand P1_SUB_450_U7 P1_U2354 ; P1_U7375
g17338 nand P1_R2238_U19 P1_U4192 ; P1_U7376
g17339 nand P1_U3294 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_U7377
g17340 nand P1_R2238_U20 P1_U4192 ; P1_U7378
g17341 nand P1_U3294 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7379
g17342 nand P1_U4173 P1_STATE2_REG_0__SCAN_IN ; P1_U7380
g17343 nand P1_U3420 P1_U7380 ; P1_U7381
g17344 nand P1_R2238_U21 P1_U4192 ; P1_U7382
g17345 nand P1_U3294 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U7383
g17346 nand P1_U2450 P1_U3271 ; P1_U7384
g17347 nand P1_R2238_U22 P1_U4192 ; P1_U7385
g17348 nand P1_U3294 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7386
g17349 nand P1_U2451 P1_U3284 ; P1_U7387
g17350 nand P1_R2238_U7 P1_U4192 ; P1_U7388
g17351 nand P1_U3294 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7389
g17352 nand P1_U3393 P1_U3290 ; P1_U7390
g17353 nand P1_U3284 P1_U3449 ; P1_U7391
g17354 nand P1_U7391 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_U7392
g17355 nand P1_U7390 P1_EBX_REG_9__SCAN_IN ; P1_U7393
g17356 nand P1_U7391 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_U7394
g17357 nand P1_U7390 P1_EBX_REG_8__SCAN_IN ; P1_U7395
g17358 nand P1_U7391 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_U7396
g17359 nand P1_U7390 P1_EBX_REG_7__SCAN_IN ; P1_U7397
g17360 nand P1_U7391 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_U7398
g17361 nand P1_U7390 P1_EBX_REG_6__SCAN_IN ; P1_U7399
g17362 nand P1_U7391 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_U7400
g17363 nand P1_U7390 P1_EBX_REG_5__SCAN_IN ; P1_U7401
g17364 nand P1_U7391 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_U7402
g17365 nand P1_U7390 P1_EBX_REG_4__SCAN_IN ; P1_U7403
g17366 nand P1_U7391 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_U7404
g17367 nand P1_U7390 P1_EBX_REG_31__SCAN_IN ; P1_U7405
g17368 nand P1_U7391 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_U7406
g17369 nand P1_U7390 P1_EBX_REG_30__SCAN_IN ; P1_U7407
g17370 nand P1_U7391 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_U7408
g17371 nand P1_U7390 P1_EBX_REG_3__SCAN_IN ; P1_U7409
g17372 nand P1_U7391 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_U7410
g17373 nand P1_U7390 P1_EBX_REG_29__SCAN_IN ; P1_U7411
g17374 nand P1_U7391 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_U7412
g17375 nand P1_U7390 P1_EBX_REG_28__SCAN_IN ; P1_U7413
g17376 nand P1_U7391 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_U7414
g17377 nand P1_U7390 P1_EBX_REG_27__SCAN_IN ; P1_U7415
g17378 nand P1_U7391 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_U7416
g17379 nand P1_U7390 P1_EBX_REG_26__SCAN_IN ; P1_U7417
g17380 nand P1_U7391 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_U7418
g17381 nand P1_U7390 P1_EBX_REG_25__SCAN_IN ; P1_U7419
g17382 nand P1_U7391 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_U7420
g17383 nand P1_U7390 P1_EBX_REG_24__SCAN_IN ; P1_U7421
g17384 nand P1_U7391 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_U7422
g17385 nand P1_U7390 P1_EBX_REG_23__SCAN_IN ; P1_U7423
g17386 nand P1_U7391 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_U7424
g17387 nand P1_U7390 P1_EBX_REG_22__SCAN_IN ; P1_U7425
g17388 nand P1_U7391 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_U7426
g17389 nand P1_U7390 P1_EBX_REG_21__SCAN_IN ; P1_U7427
g17390 nand P1_U7391 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_U7428
g17391 nand P1_U7390 P1_EBX_REG_20__SCAN_IN ; P1_U7429
g17392 nand P1_U7391 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_U7430
g17393 nand P1_U7390 P1_EBX_REG_2__SCAN_IN ; P1_U7431
g17394 nand P1_U7391 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_U7432
g17395 nand P1_U7390 P1_EBX_REG_19__SCAN_IN ; P1_U7433
g17396 nand P1_U7391 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_U7434
g17397 nand P1_U7390 P1_EBX_REG_18__SCAN_IN ; P1_U7435
g17398 nand P1_U7391 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_U7436
g17399 nand P1_U7390 P1_EBX_REG_17__SCAN_IN ; P1_U7437
g17400 nand P1_U7391 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_U7438
g17401 nand P1_U7390 P1_EBX_REG_16__SCAN_IN ; P1_U7439
g17402 nand P1_U7391 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_U7440
g17403 nand P1_U7390 P1_EBX_REG_15__SCAN_IN ; P1_U7441
g17404 nand P1_U7391 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_U7442
g17405 nand P1_U7390 P1_EBX_REG_14__SCAN_IN ; P1_U7443
g17406 nand P1_U7391 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_U7444
g17407 nand P1_U7390 P1_EBX_REG_13__SCAN_IN ; P1_U7445
g17408 nand P1_U7391 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_U7446
g17409 nand P1_U7390 P1_EBX_REG_12__SCAN_IN ; P1_U7447
g17410 nand P1_U7391 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_U7448
g17411 nand P1_U7390 P1_EBX_REG_11__SCAN_IN ; P1_U7449
g17412 nand P1_U7391 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_U7450
g17413 nand P1_U7390 P1_EBX_REG_10__SCAN_IN ; P1_U7451
g17414 nand P1_U7391 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_U7452
g17415 nand P1_U7390 P1_EBX_REG_1__SCAN_IN ; P1_U7453
g17416 nand P1_U7391 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_U7454
g17417 nand P1_U7390 P1_EBX_REG_0__SCAN_IN ; P1_U7455
g17418 nand P1_U4477 P1_U4496 ; P1_U7456
g17419 nand P1_U2430 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_U7457
g17420 nand P1_U3489 P1_U3262 ; P1_U7458
g17421 nand P1_U2430 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7459
g17422 nand P1_U3490 P1_U3262 ; P1_U7460
g17423 nand P1_U2446 P1_U3470 P1_FLUSH_REG_SCAN_IN ; P1_U7461
g17424 nand P1_U2430 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U7462
g17425 nand P1_U3491 P1_U3262 ; P1_U7463
g17426 nand P1_U2446 P1_U7712 P1_FLUSH_REG_SCAN_IN ; P1_U7464
g17427 nand P1_U2430 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7465
g17428 nand P1_U3492 P1_U3262 ; P1_U7466
g17429 nand P1_U2430 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7467
g17430 nand P1_U4185 P1_STATE_REG_0__SCAN_IN ; P1_U7468
g17431 or U210 P1_STATE2_REG_2__SCAN_IN ; P1_U7469
g17432 nand P1_U4110 P1_U7218 ; P1_U7470
g17433 nand P1_U7084 P1_U3422 ; P1_U7471
g17434 nand P1_U4211 P1_STATE2_REG_0__SCAN_IN ; P1_U7472
g17435 nand P1_U4212 P1_STATE2_REG_0__SCAN_IN ; P1_U7473
g17436 nand P1_U4213 P1_STATE2_REG_0__SCAN_IN ; P1_U7474
g17437 nand P1_U4236 P1_STATE2_REG_0__SCAN_IN ; P1_U7475
g17438 nand P1_U4264 P1_STATE2_REG_0__SCAN_IN ; P1_U7476
g17439 nand P1_U7632 P1_STATE2_REG_0__SCAN_IN ; P1_U7477
g17440 nand P1_U2608 P1_U3266 ; P1_U7478
g17441 nand P1_U4117 P1_U7093 P1_U4118 P1_U4120 ; P1_U7479
g17442 nand P1_U7632 P1_STATE2_REG_0__SCAN_IN ; P1_U7480
g17443 nand P1_U2379 P1_U3429 ; P1_U7481
g17444 nand P1_U2369 P1_U6367 ; P1_U7482
g17445 nand P1_U3888 P1_U2369 ; P1_U7483
g17446 nand P1_U7481 P1_U4229 P1_U7482 ; P1_U7484
g17447 nand P1_U7483 P1_U4230 ; P1_U7485
g17448 nand P1_U5491 P1_U4171 P1_U4194 ; P1_U7486
g17449 nand P1_U7091 P1_U4194 ; P1_U7487
g17450 nand P1_U4194 P1_U3392 ; P1_U7488
g17451 nand P1_U4236 P1_STATE2_REG_0__SCAN_IN ; P1_U7489
g17452 nand P1_U7785 P1_U7784 P1_U4072 ; P1_U7490
g17453 nand P1_U4108 P1_U7216 ; P1_U7491
g17454 nand P1_U4109 P1_U7094 ; P1_U7492
g17455 not P1_U3279 ; P1_U7493
g17456 not P1_U3276 ; P1_U7494
g17457 nand P1_U4071 P1_U2607 P1_U4070 P1_U4069 P1_U4068 ; P1_U7495
g17458 nand P1_U3734 P1_U7493 ; P1_U7496
g17459 nand P1_U3735 P1_U5469 ; P1_U7497
g17460 nand P1_U2425 P1_U7493 ; P1_U7498
g17461 nand P1_U2425 P1_U7493 ; P1_U7499
g17462 nand P1_U6361 P1_U6360 P1_U7499 ; P1_U7500
g17463 nand P1_U7493 P1_R2167_U17 ; P1_U7501
g17464 nand P1_U7493 P1_U4201 P1_R2167_U17 ; P1_U7502
g17465 nand P1_U7502 P1_U6149 ; P1_U7503
g17466 nand P1_U7493 P1_U7085 ; P1_U7504
g17467 nand P1_U7493 P1_U7471 ; P1_U7505
g17468 nand P1_U4116 P1_U4115 P1_U4114 ; P1_U7506
g17469 nand P1_U3759 P1_U7493 ; P1_U7507
g17470 nand P1_U3761 P1_U5565 P1_U3760 ; P1_U7508
g17471 nand P1_U3746 P1_U2519 ; P1_U7509
g17472 nand P1_U7493 P1_U5962 ; P1_U7510
g17473 nand P1_U7493 P1_U5965 ; P1_U7511
g17474 nand P1_U7493 P1_U5968 ; P1_U7512
g17475 nand P1_U7493 P1_U5971 ; P1_U7513
g17476 nand P1_U7493 P1_U5974 ; P1_U7514
g17477 nand P1_U7493 P1_U5977 ; P1_U7515
g17478 nand P1_U7493 P1_U5980 ; P1_U7516
g17479 nand P1_U7493 P1_U5983 ; P1_U7517
g17480 nand P1_U7493 P1_U5986 ; P1_U7518
g17481 nand P1_U7493 P1_U5989 ; P1_U7519
g17482 nand P1_U7493 P1_U5992 ; P1_U7520
g17483 nand P1_U7493 P1_U5995 ; P1_U7521
g17484 nand P1_U7493 P1_U5998 ; P1_U7522
g17485 nand P1_U7493 P1_U6001 ; P1_U7523
g17486 nand P1_U7493 P1_U6004 ; P1_U7524
g17487 nand P1_U7493 P1_U6007 ; P1_U7525
g17488 nand P1_U7493 P1_U6010 ; P1_U7526
g17489 nand P1_U7493 P1_U6013 ; P1_U7527
g17490 nand P1_U7493 P1_U6016 ; P1_U7528
g17491 nand P1_U7493 P1_U6019 ; P1_U7529
g17492 nand P1_U7493 P1_U6022 ; P1_U7530
g17493 nand P1_U7493 P1_U6025 ; P1_U7531
g17494 nand P1_U7493 P1_U6028 ; P1_U7532
g17495 nand P1_U7493 P1_U6031 ; P1_U7533
g17496 nand P1_U7493 P1_U6034 ; P1_U7534
g17497 nand P1_U7493 P1_U6037 ; P1_U7535
g17498 nand P1_U7493 P1_U6040 ; P1_U7536
g17499 nand P1_U7493 P1_U6043 ; P1_U7537
g17500 nand P1_U7493 P1_U6046 ; P1_U7538
g17501 nand P1_U7493 P1_U6049 ; P1_U7539
g17502 nand P1_U7493 P1_U6052 ; P1_U7540
g17503 nand P1_U2357 P1_U7493 ; P1_U7541
g17504 nand P1_U7541 P1_UWORD_REG_0__SCAN_IN ; P1_U7542
g17505 nand P1_U2357 P1_U7493 ; P1_U7543
g17506 nand P1_U7543 P1_UWORD_REG_1__SCAN_IN ; P1_U7544
g17507 nand P1_U2357 P1_U7493 ; P1_U7545
g17508 nand P1_U7545 P1_UWORD_REG_2__SCAN_IN ; P1_U7546
g17509 nand P1_U2357 P1_U7493 ; P1_U7547
g17510 nand P1_U7547 P1_UWORD_REG_3__SCAN_IN ; P1_U7548
g17511 nand P1_U2357 P1_U7493 ; P1_U7549
g17512 nand P1_U7549 P1_UWORD_REG_4__SCAN_IN ; P1_U7550
g17513 nand P1_U2357 P1_U7493 ; P1_U7551
g17514 nand P1_U7551 P1_UWORD_REG_5__SCAN_IN ; P1_U7552
g17515 nand P1_U2357 P1_U7493 ; P1_U7553
g17516 nand P1_U7553 P1_UWORD_REG_6__SCAN_IN ; P1_U7554
g17517 nand P1_U2357 P1_U7493 ; P1_U7555
g17518 nand P1_U7555 P1_UWORD_REG_7__SCAN_IN ; P1_U7556
g17519 nand P1_U2357 P1_U7493 ; P1_U7557
g17520 nand P1_U7557 P1_UWORD_REG_8__SCAN_IN ; P1_U7558
g17521 nand P1_U2357 P1_U7493 ; P1_U7559
g17522 nand P1_U7559 P1_UWORD_REG_9__SCAN_IN ; P1_U7560
g17523 nand P1_U2357 P1_U7493 ; P1_U7561
g17524 nand P1_U7561 P1_UWORD_REG_10__SCAN_IN ; P1_U7562
g17525 nand P1_U2357 P1_U7493 ; P1_U7563
g17526 nand P1_U7563 P1_UWORD_REG_11__SCAN_IN ; P1_U7564
g17527 nand P1_U2357 P1_U7493 ; P1_U7565
g17528 nand P1_U7565 P1_UWORD_REG_12__SCAN_IN ; P1_U7566
g17529 nand P1_U2357 P1_U7493 ; P1_U7567
g17530 nand P1_U7567 P1_UWORD_REG_13__SCAN_IN ; P1_U7568
g17531 nand P1_U2357 P1_U7493 ; P1_U7569
g17532 nand P1_U7569 P1_UWORD_REG_14__SCAN_IN ; P1_U7570
g17533 nand P1_U2357 P1_U7493 ; P1_U7571
g17534 nand P1_U7571 P1_LWORD_REG_0__SCAN_IN ; P1_U7572
g17535 nand P1_U2357 P1_U7493 ; P1_U7573
g17536 nand P1_U7573 P1_LWORD_REG_1__SCAN_IN ; P1_U7574
g17537 nand P1_U2357 P1_U7493 ; P1_U7575
g17538 nand P1_U7575 P1_LWORD_REG_2__SCAN_IN ; P1_U7576
g17539 nand P1_U2357 P1_U7493 ; P1_U7577
g17540 nand P1_U7577 P1_LWORD_REG_3__SCAN_IN ; P1_U7578
g17541 nand P1_U2357 P1_U7493 ; P1_U7579
g17542 nand P1_U7579 P1_LWORD_REG_4__SCAN_IN ; P1_U7580
g17543 nand P1_U2357 P1_U7493 ; P1_U7581
g17544 nand P1_U7581 P1_LWORD_REG_5__SCAN_IN ; P1_U7582
g17545 nand P1_U2357 P1_U7493 ; P1_U7583
g17546 nand P1_U7583 P1_LWORD_REG_6__SCAN_IN ; P1_U7584
g17547 nand P1_U2357 P1_U7493 ; P1_U7585
g17548 nand P1_U7585 P1_LWORD_REG_7__SCAN_IN ; P1_U7586
g17549 nand P1_U2357 P1_U7493 ; P1_U7587
g17550 nand P1_U7587 P1_LWORD_REG_8__SCAN_IN ; P1_U7588
g17551 nand P1_U2357 P1_U7493 ; P1_U7589
g17552 nand P1_U7589 P1_LWORD_REG_9__SCAN_IN ; P1_U7590
g17553 nand P1_U2357 P1_U7493 ; P1_U7591
g17554 nand P1_U7591 P1_LWORD_REG_10__SCAN_IN ; P1_U7592
g17555 nand P1_U2357 P1_U7493 ; P1_U7593
g17556 nand P1_U7593 P1_LWORD_REG_11__SCAN_IN ; P1_U7594
g17557 nand P1_U2357 P1_U7493 ; P1_U7595
g17558 nand P1_U7595 P1_LWORD_REG_12__SCAN_IN ; P1_U7596
g17559 nand P1_U2357 P1_U7493 ; P1_U7597
g17560 nand P1_U7597 P1_LWORD_REG_13__SCAN_IN ; P1_U7598
g17561 nand P1_U2357 P1_U7493 ; P1_U7599
g17562 nand P1_U7599 P1_LWORD_REG_14__SCAN_IN ; P1_U7600
g17563 nand P1_U2357 P1_U7493 ; P1_U7601
g17564 nand P1_U7601 P1_LWORD_REG_15__SCAN_IN ; P1_U7602
g17565 nand P1_U7493 P1_U3568 P1_U4259 ; P1_U7603
g17566 nand P1_U7684 P1_U7683 P1_U3581 ; P1_U7604
g17567 nand P1_U3867 P1_U7493 ; P1_U7605
g17568 nand P1_U7605 P1_U3428 ; P1_U7606
g17569 nand P1_U4208 P1_U7493 ; P1_U7607
g17570 nand P1_U7607 P1_U3447 ; P1_U7608
g17571 nand P1_U3279 P1_U3400 ; P1_U7609
g17572 nand P1_U3754 P1_U7493 ; P1_U7610
g17573 nand P1_U3755 P1_U7610 ; P1_U7611
g17574 nand P1_U5416 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7612
g17575 nand P1_U2523 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7613
g17576 nand P1_U2546 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7614
g17577 nand P1_U4052 P1_U4051 P1_U4050 P1_U4049 ; P1_U7615
g17578 nand P1_U4192 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7616
g17579 nand P1_U2573 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7617
g17580 nand P1_U4091 P1_U4089 P1_U4088 P1_U4087 ; P1_U7618
g17581 nand P1_U2592 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7619
g17582 nand P1_U4136 P1_U4135 P1_U4134 P1_U4133 ; P1_U7620
g17583 not P1_U3259 ; P1_U7621
g17584 nand P1_U7621 P1_U3261 ; P1_U7622
g17585 nand P1_U4361 P1_U4358 P1_STATE_REG_1__SCAN_IN ; P1_U7623
g17586 nand P1_U7468 P1_STATE_REG_2__SCAN_IN ; P1_U7624
g17587 nand P1_U4358 P1_STATE_REG_1__SCAN_IN ; P1_U7625
g17588 nand P1_U4502 P1_U4510 ; P1_U7626
g17589 nand P1_U5487 P1_U4171 ; P1_U7627
g17590 nand P1_U3283 P1_U3289 ; P1_U7628
g17591 not P1_U3392 ; P1_U7629
g17592 nand P1_U4208 P1_U7490 ; P1_U7630
g17593 nand P1_U5487 P1_U4171 ; P1_U7631
g17594 nand P1_U7631 P1_U7630 ; P1_U7632
g17595 nand P1_U3249 P1_BE_N_REG_3__SCAN_IN ; P1_U7633
g17596 nand P1_U4221 P1_BYTEENABLE_REG_3__SCAN_IN ; P1_U7634
g17597 nand P1_U3249 P1_BE_N_REG_2__SCAN_IN ; P1_U7635
g17598 nand P1_U4221 P1_BYTEENABLE_REG_2__SCAN_IN ; P1_U7636
g17599 nand P1_U3249 P1_BE_N_REG_1__SCAN_IN ; P1_U7637
g17600 nand P1_U4221 P1_BYTEENABLE_REG_1__SCAN_IN ; P1_U7638
g17601 nand P1_U3249 P1_BE_N_REG_0__SCAN_IN ; P1_U7639
g17602 nand P1_U4221 P1_BYTEENABLE_REG_0__SCAN_IN ; P1_U7640
g17603 nand P1_U3251 P1_STATE_REG_0__SCAN_IN P1_REQUESTPENDING_REG_SCAN_IN ; P1_U7641
g17604 nand P1_U3259 P1_STATE_REG_2__SCAN_IN ; P1_U7642
g17605 nand P1_U7642 P1_U7641 ; P1_U7643
g17606 nand P1_U7624 P1_U4361 P1_STATE_REG_1__SCAN_IN ; P1_U7644
g17607 nand P1_U7643 P1_U3248 ; P1_U7645
g17608 nand P1_U3260 P1_STATE_REG_2__SCAN_IN P1_STATE_REG_0__SCAN_IN ; P1_U7646
g17609 nand P1_U4371 P1_U3251 ; P1_U7647
g17610 or P1_STATE_REG_1__SCAN_IN P1_STATE_REG_0__SCAN_IN ; P1_U7648
g17611 nand P1_U4258 P1_STATE_REG_0__SCAN_IN ; P1_U7649
g17612 not P1_U3462 ; P1_U7650
g17613 nand P1_U7650 P1_DATAWIDTH_REG_0__SCAN_IN ; P1_U7651
g17614 nand P1_U3463 P1_U3462 ; P1_U7652
g17615 nand P1_U3462 P1_U4376 ; P1_U7653
g17616 nand P1_U7650 P1_DATAWIDTH_REG_1__SCAN_IN ; P1_U7654
g17617 nand P1_U3541 P1_U3540 P1_U3265 ; P1_U7655
g17618 nand P1_U3270 P1_INSTQUEUE_REG_7__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7656
g17619 nand P1_U3270 P1_U3265 P1_INSTQUEUE_REG_5__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7657
g17620 nand P1_U3270 P1_U3264 P1_U3266 P1_INSTQUEUE_REG_2__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7658
g17621 nand P1_U3543 P1_U3542 P1_U3270 ; P1_U7659
g17622 nand P1_U3545 P1_U3544 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7660
g17623 nand P1_U3547 P1_U3546 P1_U3265 ; P1_U7661
g17624 nand P1_U3549 P1_U3548 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7662
g17625 nand P1_U3551 P1_U3550 P1_U3266 ; P1_U7663
g17626 nand P1_INSTQUEUE_REG_15__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7664
g17627 nand P1_U3264 P1_U3265 P1_U3266 P1_U3270 P1_INSTQUEUE_REG_0__4__SCAN_IN ; P1_U7665
g17628 nand P1_U3264 P1_U3265 P1_U3266 P1_INSTQUEUE_REG_8__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7666
g17629 nand P1_U3264 P1_U3266 P1_INSTQUEUE_REG_10__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7667
g17630 nand P1_U3553 P1_U3552 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7668
g17631 nand P1_U3264 P1_U3270 P1_INSTQUEUE_REG_3__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7669
g17632 nand P1_U3264 P1_INSTQUEUE_REG_11__4__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7670
g17633 nand P1_U3264 P1_U3270 P1_INSTQUEUE_REG_3__5__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7671
g17634 nand P1_U3529 P1_U3528 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7672
g17635 nand P1_U3264 P1_U3265 P1_INSTQUEUE_REG_9__6__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7673
g17636 nand P1_U3535 P1_U3534 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7674
g17637 nand P1_U3264 P1_U3266 P1_INSTQUEUE_REG_10__6__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7675
g17638 nand P1_U3264 P1_INSTQUEUE_REG_11__6__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7676
g17639 nand P1_U3264 P1_U3265 P1_U3266 P1_U3270 P1_INSTQUEUE_REG_0__6__SCAN_IN ; P1_U7677
g17640 nand P1_U3264 P1_U3265 P1_U3266 P1_INSTQUEUE_REG_8__6__SCAN_IN P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7678
g17641 nand P1_U4494 P1_U3437 ; P1_U7679
g17642 nand P1_U7501 P1_U3284 ; P1_U7680
g17643 nand P1_U4216 P1_R2167_U17 ; P1_U7681
g17644 nand P1_U4506 P1_U3273 ; P1_U7682
g17645 nand P1_U4512 P1_STATE2_REG_0__SCAN_IN ; P1_U7683
g17646 nand P1_U4513 P1_U3294 ; P1_U7684
g17647 nand P1_U3295 P1_STATE2_REG_3__SCAN_IN ; P1_U7685
g17648 nand P1_U2428 P1_U4514 ; P1_U7686
g17649 or P1_STATE2_REG_0__SCAN_IN P1_STATEBS16_REG_SCAN_IN ; P1_U7687
g17650 nand P1_U7469 P1_STATE2_REG_0__SCAN_IN ; P1_U7688
g17651 nand P1_U4522 P1_STATE2_REG_0__SCAN_IN ; P1_U7689
g17652 nand P1_U7604 P1_U4521 P1_U3294 ; P1_U7690
g17653 nand P1_R2144_U49 P1_U3313 ; P1_U7691
g17654 nand P1_U4528 P1_U3311 ; P1_U7692
g17655 not P1_U3454 ; P1_U7693
g17656 nand P1_U3305 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U7694
g17657 nand P1_U4533 P1_U3304 ; P1_U7695
g17658 not P1_U3455 ; P1_U7696
g17659 nand P1_U4216 P1_U3273 ; P1_U7697
g17660 nand P1_R2167_U17 P1_U7497 ; P1_U7698
g17661 nand P1_U4432 P1_U5466 ; P1_U7699
g17662 nand P1_U5467 P1_U4171 ; P1_U7700
g17663 nand P1_U3467 P1_U4172 ; P1_U7701
g17664 nand P1_U5476 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_U7702
g17665 nand P1_U4460 P1_U3278 ; P1_U7703
g17666 nand P1_U4415 P1_U3277 ; P1_U7704
g17667 nand P1_U3271 P1_U3415 ; P1_U7705
g17668 nand P1_U4477 P1_U5493 ; P1_U7706
g17669 nand P1_U7706 P1_U7705 ; P1_U7707
g17670 nand P1_U5476 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7708
g17671 nand P1_U5509 P1_U4172 ; P1_U7709
g17672 nand P1_U4174 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_U7710
g17673 nand P1_SUB_580_U6 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_U7711
g17674 not P1_U3470 ; P1_U7712
g17675 nand P1_U4174 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_U7713
g17676 nand P1_INSTADDRPOINTER_REG_0__SCAN_IN P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_U7714
g17677 not P1_U3471 ; P1_U7715
g17678 nand P1_U5511 P1_U5501 ; P1_U7716
g17679 nand P1_U4218 P1_U3401 ; P1_U7717
g17680 nand P1_U3264 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7718
g17681 nand P1_U3265 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U7719
g17682 not P1_U3456 ; P1_U7720
g17683 nand P1_U5476 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U7721
g17684 nand P1_U5518 P1_U4172 ; P1_U7722
g17685 nand P1_U5476 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7723
g17686 nand P1_U5529 P1_U4172 ; P1_U7724
g17687 nand P1_U4214 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7725
g17688 nand P1_U5521 P1_U3266 ; P1_U7726
g17689 nand P1_U5476 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7727
g17690 nand P1_U5535 P1_U4172 ; P1_U7728
g17691 nand P1_U5537 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_U7729
g17692 nand P1_U5545 P1_U3404 ; P1_U7730
g17693 nand P1_U7693 P1_U4527 ; P1_U7731
g17694 nand P1_U3454 P1_U3314 ; P1_U7732
g17695 nand P1_U7732 P1_U7731 ; P1_U7733
g17696 nand P1_U5537 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_U7734
g17697 nand P1_U5549 P1_U3404 ; P1_U7735
g17698 nand P1_U5537 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_U7736
g17699 nand P1_U5554 P1_U3404 ; P1_U7737
g17700 nand P1_U5537 P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_U7738
g17701 nand P1_U5557 P1_U3404 ; P1_U7739
g17702 nand P1_U4477 P1_U3388 ; P1_U7740
g17703 nand P1_U3271 P1_U3281 ; P1_U7741
g17704 nand P1_U7741 P1_U7740 P1_U3257 P1_U4171 ; P1_U7742
g17705 nand P1_R2167_U17 P1_U7611 P1_U4432 ; P1_U7743
g17706 nand P1_U3424 P1_EAX_REG_31__SCAN_IN ; P1_U7744
g17707 nand P1_U3479 P1_U4223 ; P1_U7745
g17708 nand P1_U3433 P1_BYTEENABLE_REG_3__SCAN_IN ; P1_U7746
g17709 nand P1_U3480 P1_U4220 ; P1_U7747
g17710 or P1_DATAWIDTH_REG_0__SCAN_IN P1_DATAWIDTH_REG_1__SCAN_IN ; P1_U7748
g17711 nand P1_U3413 P1_DATAWIDTH_REG_0__SCAN_IN ; P1_U7749
g17712 nand P1_U7749 P1_U7748 ; P1_U7750
g17713 nand P1_U7750 P1_U3253 ; P1_U7751
g17714 nand P1_REIP_REG_0__SCAN_IN P1_REIP_REG_1__SCAN_IN ; P1_U7752
g17715 nand P1_U7752 P1_U7751 ; P1_U7753
g17716 nand P1_U3433 P1_BYTEENABLE_REG_2__SCAN_IN ; P1_U7754
g17717 nand P1_U7753 P1_U4220 ; P1_U7755
g17718 nand P1_U3433 P1_BYTEENABLE_REG_1__SCAN_IN ; P1_U7756
g17719 nand P1_U4220 P1_REIP_REG_1__SCAN_IN ; P1_U7757
g17720 nand P1_U3433 P1_BYTEENABLE_REG_0__SCAN_IN ; P1_U7758
g17721 nand P1_U4220 P1_U6599 ; P1_U7759
g17722 nand P1_U4221 P1_U3436 ; P1_U7760
g17723 nand P1_U3249 P1_W_R_N_REG_SCAN_IN ; P1_U7761
g17724 nand P1_U4177 P1_MORE_REG_SCAN_IN ; P1_U7762
g17725 nand P1_U4237 P1_U6600 ; P1_U7763
g17726 nand P1_U7650 P1_STATEBS16_REG_SCAN_IN ; P1_U7764
g17727 nand BS16 P1_U3462 ; P1_U7765
g17728 nand P1_U6603 P1_REQUESTPENDING_REG_SCAN_IN ; P1_U7766
g17729 nand P1_U6609 P1_U4180 ; P1_U7767
g17730 nand P1_U4221 P1_U3435 ; P1_U7768
g17731 nand P1_U3249 P1_D_C_N_REG_SCAN_IN ; P1_U7769
g17732 nand P1_U3249 P1_M_IO_N_REG_SCAN_IN ; P1_U7770
g17733 nand P1_U4221 P1_MEMORYFETCH_REG_SCAN_IN ; P1_U7771
g17734 nand P1_U6614 P1_READREQUEST_REG_SCAN_IN ; P1_U7772
g17735 nand P1_U6615 P1_U4181 ; P1_U7773
g17736 nand P1_U3488 P1_U4182 ; P1_U7774
g17737 nand P1_U5473 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_U7775
g17738 nand P1_U5473 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7776
g17739 nand P1_U5506 P1_U4182 ; P1_U7777
g17740 nand P1_U5473 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_U7778
g17741 nand P1_U5514 P1_U4182 ; P1_U7779
g17742 nand P1_U5473 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_U7780
g17743 nand P1_U5525 P1_U4182 ; P1_U7781
g17744 nand P1_U5473 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_U7782
g17745 nand P1_U5531 P1_U4182 ; P1_U7783
g17746 nand P1_U2605 P1_U3277 ; P1_U7784
g17747 nand P1_U4460 P1_U7495 ; P1_U7785
g17748 nand P1_U4203 P1_U3301 ; P1_U7786
g17749 nand P1_U3297 P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_U7787
g17750 nand P1_U4183 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_U7788
g17751 nand P1_U7219 P1_U3270 ; P1_U7789
g17752 not P1_U3457 ; P1_U7790
g17753 nand P1_U3276 P1_U3284 ; P1_U7791
g17754 nand P1_U7707 P1_U4494 ; P1_U7792
g17755 nand P1_U3493 P1_U3262 ; P1_U7793
g17756 nand P1_U7715 P1_STATE2_REG_1__SCAN_IN P1_FLUSH_REG_SCAN_IN ; P1_U7794
g17757 nand LT_782_120_U7 P3_DATAO_REG_30__SCAN_IN ; LT_782_120_U6
g17758 not P3_DATAO_REG_31__SCAN_IN ; LT_782_120_U7
g17759 nand LT_782_U7 P1_DATAO_REG_30__SCAN_IN ; LT_782_U6
g17760 not P1_DATAO_REG_31__SCAN_IN ; LT_782_U7
g17761 not P2_ADDRESS_REG_29__SCAN_IN ; LT_748_U6
g17762 and R170_U15 P2_ADDRESS_REG_29__SCAN_IN ; R170_U6
g17763 or P2_ADDRESS_REG_22__SCAN_IN P2_ADDRESS_REG_17__SCAN_IN P2_ADDRESS_REG_9__SCAN_IN P2_ADDRESS_REG_7__SCAN_IN ; R170_U7
g17764 nor R170_U7 P2_ADDRESS_REG_25__SCAN_IN P2_ADDRESS_REG_24__SCAN_IN P2_ADDRESS_REG_19__SCAN_IN P2_ADDRESS_REG_10__SCAN_IN ; R170_U8
g17765 or P2_ADDRESS_REG_18__SCAN_IN P2_ADDRESS_REG_16__SCAN_IN P2_ADDRESS_REG_8__SCAN_IN P2_ADDRESS_REG_0__SCAN_IN ; R170_U9
g17766 nor R170_U9 P2_ADDRESS_REG_23__SCAN_IN P2_ADDRESS_REG_11__SCAN_IN P2_ADDRESS_REG_1__SCAN_IN ; R170_U10
g17767 or P2_ADDRESS_REG_28__SCAN_IN P2_ADDRESS_REG_26__SCAN_IN P2_ADDRESS_REG_21__SCAN_IN P2_ADDRESS_REG_6__SCAN_IN ; R170_U11
g17768 nor R170_U11 P2_ADDRESS_REG_14__SCAN_IN P2_ADDRESS_REG_12__SCAN_IN P2_ADDRESS_REG_4__SCAN_IN ; R170_U12
g17769 or P2_ADDRESS_REG_27__SCAN_IN P2_ADDRESS_REG_20__SCAN_IN P2_ADDRESS_REG_13__SCAN_IN P2_ADDRESS_REG_3__SCAN_IN ; R170_U13
g17770 nor R170_U13 P2_ADDRESS_REG_15__SCAN_IN P2_ADDRESS_REG_5__SCAN_IN P2_ADDRESS_REG_2__SCAN_IN ; R170_U14
g17771 nand R170_U14 R170_U12 R170_U10 R170_U8 ; R170_U15
g17772 and R165_U15 P1_ADDRESS_REG_29__SCAN_IN ; R165_U6
g17773 or P1_ADDRESS_REG_22__SCAN_IN P1_ADDRESS_REG_17__SCAN_IN P1_ADDRESS_REG_9__SCAN_IN P1_ADDRESS_REG_7__SCAN_IN ; R165_U7
g17774 nor R165_U7 P1_ADDRESS_REG_25__SCAN_IN P1_ADDRESS_REG_24__SCAN_IN P1_ADDRESS_REG_19__SCAN_IN P1_ADDRESS_REG_10__SCAN_IN ; R165_U8
g17775 or P1_ADDRESS_REG_18__SCAN_IN P1_ADDRESS_REG_16__SCAN_IN P1_ADDRESS_REG_8__SCAN_IN P1_ADDRESS_REG_0__SCAN_IN ; R165_U9
g17776 nor R165_U9 P1_ADDRESS_REG_23__SCAN_IN P1_ADDRESS_REG_11__SCAN_IN P1_ADDRESS_REG_1__SCAN_IN ; R165_U10
g17777 or P1_ADDRESS_REG_28__SCAN_IN P1_ADDRESS_REG_26__SCAN_IN P1_ADDRESS_REG_21__SCAN_IN P1_ADDRESS_REG_6__SCAN_IN ; R165_U11
g17778 nor R165_U11 P1_ADDRESS_REG_14__SCAN_IN P1_ADDRESS_REG_12__SCAN_IN P1_ADDRESS_REG_4__SCAN_IN ; R165_U12
g17779 or P1_ADDRESS_REG_27__SCAN_IN P1_ADDRESS_REG_20__SCAN_IN P1_ADDRESS_REG_13__SCAN_IN P1_ADDRESS_REG_3__SCAN_IN ; R165_U13
g17780 nor R165_U13 P1_ADDRESS_REG_15__SCAN_IN P1_ADDRESS_REG_5__SCAN_IN P1_ADDRESS_REG_2__SCAN_IN ; R165_U14
g17781 nand R165_U14 R165_U12 R165_U10 R165_U8 ; R165_U15
g17782 nand LT_782_119_U7 P2_DATAO_REG_30__SCAN_IN ; LT_782_119_U6
g17783 not P2_DATAO_REG_31__SCAN_IN ; LT_782_119_U7
g17784 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_526_U5
g17785 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_526_U6
g17786 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_526_U7
g17787 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_526_U8
g17788 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_526_U9
g17789 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_526_U10
g17790 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_526_U11
g17791 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_526_U12
g17792 nand P3_ADD_526_U82 P3_ADD_526_U111 ; P3_ADD_526_U13
g17793 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_526_U14
g17794 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_526_U15
g17795 nand P3_ADD_526_U83 P3_ADD_526_U112 ; P3_ADD_526_U16
g17796 nand P3_ADD_526_U84 P3_ADD_526_U118 ; P3_ADD_526_U17
g17797 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_526_U18
g17798 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_526_U19
g17799 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_526_U20
g17800 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_526_U21
g17801 nand P3_ADD_526_U85 P3_ADD_526_U120 ; P3_ADD_526_U22
g17802 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_526_U23
g17803 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_526_U24
g17804 nand P3_ADD_526_U86 P3_ADD_526_U113 ; P3_ADD_526_U25
g17805 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_526_U26
g17806 nand P3_ADD_526_U87 P3_ADD_526_U119 ; P3_ADD_526_U27
g17807 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_526_U28
g17808 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_526_U29
g17809 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_526_U30
g17810 nand P3_ADD_526_U88 P3_ADD_526_U124 ; P3_ADD_526_U31
g17811 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_526_U32
g17812 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_526_U33
g17813 nand P3_ADD_526_U89 P3_ADD_526_U117 ; P3_ADD_526_U34
g17814 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_526_U35
g17815 nand P3_ADD_526_U90 P3_ADD_526_U114 ; P3_ADD_526_U36
g17816 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_526_U37
g17817 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_526_U38
g17818 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_526_U39
g17819 nand P3_ADD_526_U91 P3_ADD_526_U121 ; P3_ADD_526_U40
g17820 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_526_U41
g17821 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_526_U42
g17822 nand P3_ADD_526_U92 P3_ADD_526_U115 ; P3_ADD_526_U43
g17823 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_526_U44
g17824 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_526_U45
g17825 nand P3_ADD_526_U93 P3_ADD_526_U116 ; P3_ADD_526_U46
g17826 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_526_U47
g17827 nand P3_ADD_526_U94 P3_ADD_526_U122 ; P3_ADD_526_U48
g17828 nand P3_ADD_526_U123 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_526_U49
g17829 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_526_U50
g17830 nand P3_ADD_526_U142 P3_ADD_526_U141 ; P3_ADD_526_U51
g17831 nand P3_ADD_526_U144 P3_ADD_526_U143 ; P3_ADD_526_U52
g17832 nand P3_ADD_526_U146 P3_ADD_526_U145 ; P3_ADD_526_U53
g17833 nand P3_ADD_526_U148 P3_ADD_526_U147 ; P3_ADD_526_U54
g17834 nand P3_ADD_526_U150 P3_ADD_526_U149 ; P3_ADD_526_U55
g17835 nand P3_ADD_526_U152 P3_ADD_526_U151 ; P3_ADD_526_U56
g17836 nand P3_ADD_526_U154 P3_ADD_526_U153 ; P3_ADD_526_U57
g17837 nand P3_ADD_526_U156 P3_ADD_526_U155 ; P3_ADD_526_U58
g17838 nand P3_ADD_526_U158 P3_ADD_526_U157 ; P3_ADD_526_U59
g17839 nand P3_ADD_526_U160 P3_ADD_526_U159 ; P3_ADD_526_U60
g17840 nand P3_ADD_526_U162 P3_ADD_526_U161 ; P3_ADD_526_U61
g17841 nand P3_ADD_526_U164 P3_ADD_526_U163 ; P3_ADD_526_U62
g17842 nand P3_ADD_526_U166 P3_ADD_526_U165 ; P3_ADD_526_U63
g17843 nand P3_ADD_526_U168 P3_ADD_526_U167 ; P3_ADD_526_U64
g17844 nand P3_ADD_526_U170 P3_ADD_526_U169 ; P3_ADD_526_U65
g17845 nand P3_ADD_526_U172 P3_ADD_526_U171 ; P3_ADD_526_U66
g17846 nand P3_ADD_526_U174 P3_ADD_526_U173 ; P3_ADD_526_U67
g17847 nand P3_ADD_526_U176 P3_ADD_526_U175 ; P3_ADD_526_U68
g17848 nand P3_ADD_526_U178 P3_ADD_526_U177 ; P3_ADD_526_U69
g17849 nand P3_ADD_526_U180 P3_ADD_526_U179 ; P3_ADD_526_U70
g17850 nand P3_ADD_526_U182 P3_ADD_526_U181 ; P3_ADD_526_U71
g17851 nand P3_ADD_526_U184 P3_ADD_526_U183 ; P3_ADD_526_U72
g17852 nand P3_ADD_526_U186 P3_ADD_526_U185 ; P3_ADD_526_U73
g17853 nand P3_ADD_526_U188 P3_ADD_526_U187 ; P3_ADD_526_U74
g17854 nand P3_ADD_526_U190 P3_ADD_526_U189 ; P3_ADD_526_U75
g17855 nand P3_ADD_526_U192 P3_ADD_526_U191 ; P3_ADD_526_U76
g17856 nand P3_ADD_526_U194 P3_ADD_526_U193 ; P3_ADD_526_U77
g17857 nand P3_ADD_526_U196 P3_ADD_526_U195 ; P3_ADD_526_U78
g17858 nand P3_ADD_526_U198 P3_ADD_526_U197 ; P3_ADD_526_U79
g17859 nand P3_ADD_526_U200 P3_ADD_526_U199 ; P3_ADD_526_U80
g17860 nand P3_ADD_526_U202 P3_ADD_526_U201 ; P3_ADD_526_U81
g17861 and P3_INSTADDRPOINTER_REG_3__SCAN_IN P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_526_U82
g17862 and P3_INSTADDRPOINTER_REG_5__SCAN_IN P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_526_U83
g17863 and P3_INSTADDRPOINTER_REG_7__SCAN_IN P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_526_U84
g17864 and P3_INSTADDRPOINTER_REG_9__SCAN_IN P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_526_U85
g17865 and P3_INSTADDRPOINTER_REG_11__SCAN_IN P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_526_U86
g17866 and P3_INSTADDRPOINTER_REG_13__SCAN_IN P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_526_U87
g17867 and P3_INSTADDRPOINTER_REG_15__SCAN_IN P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_526_U88
g17868 and P3_INSTADDRPOINTER_REG_17__SCAN_IN P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_526_U89
g17869 and P3_INSTADDRPOINTER_REG_19__SCAN_IN P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_526_U90
g17870 and P3_INSTADDRPOINTER_REG_21__SCAN_IN P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_526_U91
g17871 and P3_INSTADDRPOINTER_REG_23__SCAN_IN P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_526_U92
g17872 and P3_INSTADDRPOINTER_REG_25__SCAN_IN P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_526_U93
g17873 and P3_INSTADDRPOINTER_REG_27__SCAN_IN P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_526_U94
g17874 nand P3_ADD_526_U118 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_526_U95
g17875 nand P3_ADD_526_U112 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_526_U96
g17876 nand P3_ADD_526_U111 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_526_U97
g17877 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_526_U98
g17878 nand P3_ADD_526_U128 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_526_U99
g17879 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_526_U100
g17880 nand P3_ADD_526_U122 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_526_U101
g17881 nand P3_ADD_526_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_526_U102
g17882 nand P3_ADD_526_U115 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_526_U103
g17883 nand P3_ADD_526_U121 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_526_U104
g17884 nand P3_ADD_526_U114 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_526_U105
g17885 nand P3_ADD_526_U117 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_526_U106
g17886 nand P3_ADD_526_U124 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_526_U107
g17887 nand P3_ADD_526_U119 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_526_U108
g17888 nand P3_ADD_526_U113 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_526_U109
g17889 nand P3_ADD_526_U120 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_526_U110
g17890 not P3_ADD_526_U10 ; P3_ADD_526_U111
g17891 not P3_ADD_526_U13 ; P3_ADD_526_U112
g17892 not P3_ADD_526_U22 ; P3_ADD_526_U113
g17893 not P3_ADD_526_U34 ; P3_ADD_526_U114
g17894 not P3_ADD_526_U40 ; P3_ADD_526_U115
g17895 not P3_ADD_526_U43 ; P3_ADD_526_U116
g17896 not P3_ADD_526_U31 ; P3_ADD_526_U117
g17897 not P3_ADD_526_U16 ; P3_ADD_526_U118
g17898 not P3_ADD_526_U25 ; P3_ADD_526_U119
g17899 not P3_ADD_526_U17 ; P3_ADD_526_U120
g17900 not P3_ADD_526_U36 ; P3_ADD_526_U121
g17901 not P3_ADD_526_U46 ; P3_ADD_526_U122
g17902 not P3_ADD_526_U48 ; P3_ADD_526_U123
g17903 not P3_ADD_526_U27 ; P3_ADD_526_U124
g17904 not P3_ADD_526_U95 ; P3_ADD_526_U125
g17905 not P3_ADD_526_U96 ; P3_ADD_526_U126
g17906 not P3_ADD_526_U97 ; P3_ADD_526_U127
g17907 not P3_ADD_526_U49 ; P3_ADD_526_U128
g17908 not P3_ADD_526_U99 ; P3_ADD_526_U129
g17909 not P3_ADD_526_U100 ; P3_ADD_526_U130
g17910 not P3_ADD_526_U101 ; P3_ADD_526_U131
g17911 not P3_ADD_526_U102 ; P3_ADD_526_U132
g17912 not P3_ADD_526_U103 ; P3_ADD_526_U133
g17913 not P3_ADD_526_U104 ; P3_ADD_526_U134
g17914 not P3_ADD_526_U105 ; P3_ADD_526_U135
g17915 not P3_ADD_526_U106 ; P3_ADD_526_U136
g17916 not P3_ADD_526_U107 ; P3_ADD_526_U137
g17917 not P3_ADD_526_U108 ; P3_ADD_526_U138
g17918 not P3_ADD_526_U109 ; P3_ADD_526_U139
g17919 not P3_ADD_526_U110 ; P3_ADD_526_U140
g17920 nand P3_ADD_526_U120 P3_ADD_526_U18 ; P3_ADD_526_U141
g17921 nand P3_ADD_526_U17 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_526_U142
g17922 nand P3_ADD_526_U95 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_526_U143
g17923 nand P3_ADD_526_U125 P3_ADD_526_U14 ; P3_ADD_526_U144
g17924 nand P3_ADD_526_U118 P3_ADD_526_U15 ; P3_ADD_526_U145
g17925 nand P3_ADD_526_U16 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_526_U146
g17926 nand P3_ADD_526_U96 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_526_U147
g17927 nand P3_ADD_526_U126 P3_ADD_526_U11 ; P3_ADD_526_U148
g17928 nand P3_ADD_526_U112 P3_ADD_526_U12 ; P3_ADD_526_U149
g17929 nand P3_ADD_526_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_526_U150
g17930 nand P3_ADD_526_U97 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_526_U151
g17931 nand P3_ADD_526_U127 P3_ADD_526_U8 ; P3_ADD_526_U152
g17932 nand P3_ADD_526_U111 P3_ADD_526_U9 ; P3_ADD_526_U153
g17933 nand P3_ADD_526_U10 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_526_U154
g17934 nand P3_ADD_526_U99 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_526_U155
g17935 nand P3_ADD_526_U129 P3_ADD_526_U98 ; P3_ADD_526_U156
g17936 nand P3_ADD_526_U49 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_526_U157
g17937 nand P3_ADD_526_U128 P3_ADD_526_U50 ; P3_ADD_526_U158
g17938 nand P3_ADD_526_U100 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_526_U159
g17939 nand P3_ADD_526_U130 P3_ADD_526_U6 ; P3_ADD_526_U160
g17940 nand P3_ADD_526_U123 P3_ADD_526_U47 ; P3_ADD_526_U161
g17941 nand P3_ADD_526_U48 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_526_U162
g17942 nand P3_ADD_526_U101 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_526_U163
g17943 nand P3_ADD_526_U131 P3_ADD_526_U45 ; P3_ADD_526_U164
g17944 nand P3_ADD_526_U122 P3_ADD_526_U44 ; P3_ADD_526_U165
g17945 nand P3_ADD_526_U46 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_526_U166
g17946 nand P3_ADD_526_U102 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_526_U167
g17947 nand P3_ADD_526_U132 P3_ADD_526_U41 ; P3_ADD_526_U168
g17948 nand P3_ADD_526_U116 P3_ADD_526_U42 ; P3_ADD_526_U169
g17949 nand P3_ADD_526_U43 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_526_U170
g17950 nand P3_ADD_526_U103 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_526_U171
g17951 nand P3_ADD_526_U133 P3_ADD_526_U38 ; P3_ADD_526_U172
g17952 nand P3_ADD_526_U115 P3_ADD_526_U39 ; P3_ADD_526_U173
g17953 nand P3_ADD_526_U40 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_526_U174
g17954 nand P3_ADD_526_U104 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_526_U175
g17955 nand P3_ADD_526_U134 P3_ADD_526_U37 ; P3_ADD_526_U176
g17956 nand P3_ADD_526_U121 P3_ADD_526_U35 ; P3_ADD_526_U177
g17957 nand P3_ADD_526_U36 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_526_U178
g17958 nand P3_ADD_526_U105 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_526_U179
g17959 nand P3_ADD_526_U135 P3_ADD_526_U32 ; P3_ADD_526_U180
g17960 nand P3_ADD_526_U7 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_526_U181
g17961 nand P3_ADD_526_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_526_U182
g17962 nand P3_ADD_526_U114 P3_ADD_526_U33 ; P3_ADD_526_U183
g17963 nand P3_ADD_526_U34 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_526_U184
g17964 nand P3_ADD_526_U106 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_526_U185
g17965 nand P3_ADD_526_U136 P3_ADD_526_U29 ; P3_ADD_526_U186
g17966 nand P3_ADD_526_U117 P3_ADD_526_U30 ; P3_ADD_526_U187
g17967 nand P3_ADD_526_U31 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_526_U188
g17968 nand P3_ADD_526_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_526_U189
g17969 nand P3_ADD_526_U137 P3_ADD_526_U28 ; P3_ADD_526_U190
g17970 nand P3_ADD_526_U124 P3_ADD_526_U26 ; P3_ADD_526_U191
g17971 nand P3_ADD_526_U27 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_526_U192
g17972 nand P3_ADD_526_U108 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_526_U193
g17973 nand P3_ADD_526_U138 P3_ADD_526_U23 ; P3_ADD_526_U194
g17974 nand P3_ADD_526_U119 P3_ADD_526_U24 ; P3_ADD_526_U195
g17975 nand P3_ADD_526_U25 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_526_U196
g17976 nand P3_ADD_526_U109 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_526_U197
g17977 nand P3_ADD_526_U139 P3_ADD_526_U20 ; P3_ADD_526_U198
g17978 nand P3_ADD_526_U113 P3_ADD_526_U21 ; P3_ADD_526_U199
g17979 nand P3_ADD_526_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_526_U200
g17980 nand P3_ADD_526_U110 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_526_U201
g17981 nand P3_ADD_526_U140 P3_ADD_526_U19 ; P3_ADD_526_U202
g17982 not P3_EBX_REG_0__SCAN_IN ; P3_ADD_552_U5
g17983 not P3_EBX_REG_2__SCAN_IN ; P3_ADD_552_U6
g17984 not P3_EBX_REG_1__SCAN_IN ; P3_ADD_552_U7
g17985 not P3_EBX_REG_4__SCAN_IN ; P3_ADD_552_U8
g17986 not P3_EBX_REG_3__SCAN_IN ; P3_ADD_552_U9
g17987 nand P3_EBX_REG_0__SCAN_IN P3_EBX_REG_1__SCAN_IN P3_EBX_REG_2__SCAN_IN ; P3_ADD_552_U10
g17988 not P3_EBX_REG_6__SCAN_IN ; P3_ADD_552_U11
g17989 not P3_EBX_REG_5__SCAN_IN ; P3_ADD_552_U12
g17990 nand P3_ADD_552_U82 P3_ADD_552_U111 ; P3_ADD_552_U13
g17991 not P3_EBX_REG_8__SCAN_IN ; P3_ADD_552_U14
g17992 not P3_EBX_REG_7__SCAN_IN ; P3_ADD_552_U15
g17993 nand P3_ADD_552_U83 P3_ADD_552_U112 ; P3_ADD_552_U16
g17994 nand P3_ADD_552_U84 P3_ADD_552_U118 ; P3_ADD_552_U17
g17995 not P3_EBX_REG_9__SCAN_IN ; P3_ADD_552_U18
g17996 not P3_EBX_REG_10__SCAN_IN ; P3_ADD_552_U19
g17997 not P3_EBX_REG_12__SCAN_IN ; P3_ADD_552_U20
g17998 not P3_EBX_REG_11__SCAN_IN ; P3_ADD_552_U21
g17999 nand P3_ADD_552_U85 P3_ADD_552_U120 ; P3_ADD_552_U22
g18000 not P3_EBX_REG_14__SCAN_IN ; P3_ADD_552_U23
g18001 not P3_EBX_REG_13__SCAN_IN ; P3_ADD_552_U24
g18002 nand P3_ADD_552_U86 P3_ADD_552_U113 ; P3_ADD_552_U25
g18003 not P3_EBX_REG_15__SCAN_IN ; P3_ADD_552_U26
g18004 nand P3_ADD_552_U87 P3_ADD_552_U119 ; P3_ADD_552_U27
g18005 not P3_EBX_REG_16__SCAN_IN ; P3_ADD_552_U28
g18006 not P3_EBX_REG_18__SCAN_IN ; P3_ADD_552_U29
g18007 not P3_EBX_REG_17__SCAN_IN ; P3_ADD_552_U30
g18008 nand P3_ADD_552_U88 P3_ADD_552_U124 ; P3_ADD_552_U31
g18009 not P3_EBX_REG_20__SCAN_IN ; P3_ADD_552_U32
g18010 not P3_EBX_REG_19__SCAN_IN ; P3_ADD_552_U33
g18011 nand P3_ADD_552_U89 P3_ADD_552_U117 ; P3_ADD_552_U34
g18012 not P3_EBX_REG_21__SCAN_IN ; P3_ADD_552_U35
g18013 nand P3_ADD_552_U90 P3_ADD_552_U114 ; P3_ADD_552_U36
g18014 not P3_EBX_REG_22__SCAN_IN ; P3_ADD_552_U37
g18015 not P3_EBX_REG_24__SCAN_IN ; P3_ADD_552_U38
g18016 not P3_EBX_REG_23__SCAN_IN ; P3_ADD_552_U39
g18017 nand P3_ADD_552_U91 P3_ADD_552_U121 ; P3_ADD_552_U40
g18018 not P3_EBX_REG_26__SCAN_IN ; P3_ADD_552_U41
g18019 not P3_EBX_REG_25__SCAN_IN ; P3_ADD_552_U42
g18020 nand P3_ADD_552_U92 P3_ADD_552_U115 ; P3_ADD_552_U43
g18021 not P3_EBX_REG_27__SCAN_IN ; P3_ADD_552_U44
g18022 not P3_EBX_REG_28__SCAN_IN ; P3_ADD_552_U45
g18023 nand P3_ADD_552_U93 P3_ADD_552_U116 ; P3_ADD_552_U46
g18024 not P3_EBX_REG_29__SCAN_IN ; P3_ADD_552_U47
g18025 nand P3_ADD_552_U94 P3_ADD_552_U122 ; P3_ADD_552_U48
g18026 nand P3_ADD_552_U123 P3_EBX_REG_29__SCAN_IN ; P3_ADD_552_U49
g18027 not P3_EBX_REG_30__SCAN_IN ; P3_ADD_552_U50
g18028 nand P3_ADD_552_U142 P3_ADD_552_U141 ; P3_ADD_552_U51
g18029 nand P3_ADD_552_U144 P3_ADD_552_U143 ; P3_ADD_552_U52
g18030 nand P3_ADD_552_U146 P3_ADD_552_U145 ; P3_ADD_552_U53
g18031 nand P3_ADD_552_U148 P3_ADD_552_U147 ; P3_ADD_552_U54
g18032 nand P3_ADD_552_U150 P3_ADD_552_U149 ; P3_ADD_552_U55
g18033 nand P3_ADD_552_U152 P3_ADD_552_U151 ; P3_ADD_552_U56
g18034 nand P3_ADD_552_U154 P3_ADD_552_U153 ; P3_ADD_552_U57
g18035 nand P3_ADD_552_U156 P3_ADD_552_U155 ; P3_ADD_552_U58
g18036 nand P3_ADD_552_U158 P3_ADD_552_U157 ; P3_ADD_552_U59
g18037 nand P3_ADD_552_U160 P3_ADD_552_U159 ; P3_ADD_552_U60
g18038 nand P3_ADD_552_U162 P3_ADD_552_U161 ; P3_ADD_552_U61
g18039 nand P3_ADD_552_U164 P3_ADD_552_U163 ; P3_ADD_552_U62
g18040 nand P3_ADD_552_U166 P3_ADD_552_U165 ; P3_ADD_552_U63
g18041 nand P3_ADD_552_U168 P3_ADD_552_U167 ; P3_ADD_552_U64
g18042 nand P3_ADD_552_U170 P3_ADD_552_U169 ; P3_ADD_552_U65
g18043 nand P3_ADD_552_U172 P3_ADD_552_U171 ; P3_ADD_552_U66
g18044 nand P3_ADD_552_U174 P3_ADD_552_U173 ; P3_ADD_552_U67
g18045 nand P3_ADD_552_U176 P3_ADD_552_U175 ; P3_ADD_552_U68
g18046 nand P3_ADD_552_U178 P3_ADD_552_U177 ; P3_ADD_552_U69
g18047 nand P3_ADD_552_U180 P3_ADD_552_U179 ; P3_ADD_552_U70
g18048 nand P3_ADD_552_U182 P3_ADD_552_U181 ; P3_ADD_552_U71
g18049 nand P3_ADD_552_U184 P3_ADD_552_U183 ; P3_ADD_552_U72
g18050 nand P3_ADD_552_U186 P3_ADD_552_U185 ; P3_ADD_552_U73
g18051 nand P3_ADD_552_U188 P3_ADD_552_U187 ; P3_ADD_552_U74
g18052 nand P3_ADD_552_U190 P3_ADD_552_U189 ; P3_ADD_552_U75
g18053 nand P3_ADD_552_U192 P3_ADD_552_U191 ; P3_ADD_552_U76
g18054 nand P3_ADD_552_U194 P3_ADD_552_U193 ; P3_ADD_552_U77
g18055 nand P3_ADD_552_U196 P3_ADD_552_U195 ; P3_ADD_552_U78
g18056 nand P3_ADD_552_U198 P3_ADD_552_U197 ; P3_ADD_552_U79
g18057 nand P3_ADD_552_U200 P3_ADD_552_U199 ; P3_ADD_552_U80
g18058 nand P3_ADD_552_U202 P3_ADD_552_U201 ; P3_ADD_552_U81
g18059 and P3_EBX_REG_3__SCAN_IN P3_EBX_REG_4__SCAN_IN ; P3_ADD_552_U82
g18060 and P3_EBX_REG_5__SCAN_IN P3_EBX_REG_6__SCAN_IN ; P3_ADD_552_U83
g18061 and P3_EBX_REG_7__SCAN_IN P3_EBX_REG_8__SCAN_IN ; P3_ADD_552_U84
g18062 and P3_EBX_REG_9__SCAN_IN P3_EBX_REG_10__SCAN_IN ; P3_ADD_552_U85
g18063 and P3_EBX_REG_11__SCAN_IN P3_EBX_REG_12__SCAN_IN ; P3_ADD_552_U86
g18064 and P3_EBX_REG_13__SCAN_IN P3_EBX_REG_14__SCAN_IN ; P3_ADD_552_U87
g18065 and P3_EBX_REG_15__SCAN_IN P3_EBX_REG_16__SCAN_IN ; P3_ADD_552_U88
g18066 and P3_EBX_REG_17__SCAN_IN P3_EBX_REG_18__SCAN_IN ; P3_ADD_552_U89
g18067 and P3_EBX_REG_19__SCAN_IN P3_EBX_REG_20__SCAN_IN ; P3_ADD_552_U90
g18068 and P3_EBX_REG_21__SCAN_IN P3_EBX_REG_22__SCAN_IN ; P3_ADD_552_U91
g18069 and P3_EBX_REG_23__SCAN_IN P3_EBX_REG_24__SCAN_IN ; P3_ADD_552_U92
g18070 and P3_EBX_REG_25__SCAN_IN P3_EBX_REG_26__SCAN_IN ; P3_ADD_552_U93
g18071 and P3_EBX_REG_27__SCAN_IN P3_EBX_REG_28__SCAN_IN ; P3_ADD_552_U94
g18072 nand P3_ADD_552_U118 P3_EBX_REG_7__SCAN_IN ; P3_ADD_552_U95
g18073 nand P3_ADD_552_U112 P3_EBX_REG_5__SCAN_IN ; P3_ADD_552_U96
g18074 nand P3_ADD_552_U111 P3_EBX_REG_3__SCAN_IN ; P3_ADD_552_U97
g18075 not P3_EBX_REG_31__SCAN_IN ; P3_ADD_552_U98
g18076 nand P3_ADD_552_U128 P3_EBX_REG_30__SCAN_IN ; P3_ADD_552_U99
g18077 nand P3_EBX_REG_0__SCAN_IN P3_EBX_REG_1__SCAN_IN ; P3_ADD_552_U100
g18078 nand P3_ADD_552_U122 P3_EBX_REG_27__SCAN_IN ; P3_ADD_552_U101
g18079 nand P3_ADD_552_U116 P3_EBX_REG_25__SCAN_IN ; P3_ADD_552_U102
g18080 nand P3_ADD_552_U115 P3_EBX_REG_23__SCAN_IN ; P3_ADD_552_U103
g18081 nand P3_ADD_552_U121 P3_EBX_REG_21__SCAN_IN ; P3_ADD_552_U104
g18082 nand P3_ADD_552_U114 P3_EBX_REG_19__SCAN_IN ; P3_ADD_552_U105
g18083 nand P3_ADD_552_U117 P3_EBX_REG_17__SCAN_IN ; P3_ADD_552_U106
g18084 nand P3_ADD_552_U124 P3_EBX_REG_15__SCAN_IN ; P3_ADD_552_U107
g18085 nand P3_ADD_552_U119 P3_EBX_REG_13__SCAN_IN ; P3_ADD_552_U108
g18086 nand P3_ADD_552_U113 P3_EBX_REG_11__SCAN_IN ; P3_ADD_552_U109
g18087 nand P3_ADD_552_U120 P3_EBX_REG_9__SCAN_IN ; P3_ADD_552_U110
g18088 not P3_ADD_552_U10 ; P3_ADD_552_U111
g18089 not P3_ADD_552_U13 ; P3_ADD_552_U112
g18090 not P3_ADD_552_U22 ; P3_ADD_552_U113
g18091 not P3_ADD_552_U34 ; P3_ADD_552_U114
g18092 not P3_ADD_552_U40 ; P3_ADD_552_U115
g18093 not P3_ADD_552_U43 ; P3_ADD_552_U116
g18094 not P3_ADD_552_U31 ; P3_ADD_552_U117
g18095 not P3_ADD_552_U16 ; P3_ADD_552_U118
g18096 not P3_ADD_552_U25 ; P3_ADD_552_U119
g18097 not P3_ADD_552_U17 ; P3_ADD_552_U120
g18098 not P3_ADD_552_U36 ; P3_ADD_552_U121
g18099 not P3_ADD_552_U46 ; P3_ADD_552_U122
g18100 not P3_ADD_552_U48 ; P3_ADD_552_U123
g18101 not P3_ADD_552_U27 ; P3_ADD_552_U124
g18102 not P3_ADD_552_U95 ; P3_ADD_552_U125
g18103 not P3_ADD_552_U96 ; P3_ADD_552_U126
g18104 not P3_ADD_552_U97 ; P3_ADD_552_U127
g18105 not P3_ADD_552_U49 ; P3_ADD_552_U128
g18106 not P3_ADD_552_U99 ; P3_ADD_552_U129
g18107 not P3_ADD_552_U100 ; P3_ADD_552_U130
g18108 not P3_ADD_552_U101 ; P3_ADD_552_U131
g18109 not P3_ADD_552_U102 ; P3_ADD_552_U132
g18110 not P3_ADD_552_U103 ; P3_ADD_552_U133
g18111 not P3_ADD_552_U104 ; P3_ADD_552_U134
g18112 not P3_ADD_552_U105 ; P3_ADD_552_U135
g18113 not P3_ADD_552_U106 ; P3_ADD_552_U136
g18114 not P3_ADD_552_U107 ; P3_ADD_552_U137
g18115 not P3_ADD_552_U108 ; P3_ADD_552_U138
g18116 not P3_ADD_552_U109 ; P3_ADD_552_U139
g18117 not P3_ADD_552_U110 ; P3_ADD_552_U140
g18118 nand P3_ADD_552_U120 P3_ADD_552_U18 ; P3_ADD_552_U141
g18119 nand P3_ADD_552_U17 P3_EBX_REG_9__SCAN_IN ; P3_ADD_552_U142
g18120 nand P3_ADD_552_U95 P3_EBX_REG_8__SCAN_IN ; P3_ADD_552_U143
g18121 nand P3_ADD_552_U125 P3_ADD_552_U14 ; P3_ADD_552_U144
g18122 nand P3_ADD_552_U118 P3_ADD_552_U15 ; P3_ADD_552_U145
g18123 nand P3_ADD_552_U16 P3_EBX_REG_7__SCAN_IN ; P3_ADD_552_U146
g18124 nand P3_ADD_552_U96 P3_EBX_REG_6__SCAN_IN ; P3_ADD_552_U147
g18125 nand P3_ADD_552_U126 P3_ADD_552_U11 ; P3_ADD_552_U148
g18126 nand P3_ADD_552_U112 P3_ADD_552_U12 ; P3_ADD_552_U149
g18127 nand P3_ADD_552_U13 P3_EBX_REG_5__SCAN_IN ; P3_ADD_552_U150
g18128 nand P3_ADD_552_U97 P3_EBX_REG_4__SCAN_IN ; P3_ADD_552_U151
g18129 nand P3_ADD_552_U127 P3_ADD_552_U8 ; P3_ADD_552_U152
g18130 nand P3_ADD_552_U111 P3_ADD_552_U9 ; P3_ADD_552_U153
g18131 nand P3_ADD_552_U10 P3_EBX_REG_3__SCAN_IN ; P3_ADD_552_U154
g18132 nand P3_ADD_552_U99 P3_EBX_REG_31__SCAN_IN ; P3_ADD_552_U155
g18133 nand P3_ADD_552_U129 P3_ADD_552_U98 ; P3_ADD_552_U156
g18134 nand P3_ADD_552_U49 P3_EBX_REG_30__SCAN_IN ; P3_ADD_552_U157
g18135 nand P3_ADD_552_U128 P3_ADD_552_U50 ; P3_ADD_552_U158
g18136 nand P3_ADD_552_U100 P3_EBX_REG_2__SCAN_IN ; P3_ADD_552_U159
g18137 nand P3_ADD_552_U130 P3_ADD_552_U6 ; P3_ADD_552_U160
g18138 nand P3_ADD_552_U123 P3_ADD_552_U47 ; P3_ADD_552_U161
g18139 nand P3_ADD_552_U48 P3_EBX_REG_29__SCAN_IN ; P3_ADD_552_U162
g18140 nand P3_ADD_552_U101 P3_EBX_REG_28__SCAN_IN ; P3_ADD_552_U163
g18141 nand P3_ADD_552_U131 P3_ADD_552_U45 ; P3_ADD_552_U164
g18142 nand P3_ADD_552_U122 P3_ADD_552_U44 ; P3_ADD_552_U165
g18143 nand P3_ADD_552_U46 P3_EBX_REG_27__SCAN_IN ; P3_ADD_552_U166
g18144 nand P3_ADD_552_U102 P3_EBX_REG_26__SCAN_IN ; P3_ADD_552_U167
g18145 nand P3_ADD_552_U132 P3_ADD_552_U41 ; P3_ADD_552_U168
g18146 nand P3_ADD_552_U116 P3_ADD_552_U42 ; P3_ADD_552_U169
g18147 nand P3_ADD_552_U43 P3_EBX_REG_25__SCAN_IN ; P3_ADD_552_U170
g18148 nand P3_ADD_552_U103 P3_EBX_REG_24__SCAN_IN ; P3_ADD_552_U171
g18149 nand P3_ADD_552_U133 P3_ADD_552_U38 ; P3_ADD_552_U172
g18150 nand P3_ADD_552_U115 P3_ADD_552_U39 ; P3_ADD_552_U173
g18151 nand P3_ADD_552_U40 P3_EBX_REG_23__SCAN_IN ; P3_ADD_552_U174
g18152 nand P3_ADD_552_U104 P3_EBX_REG_22__SCAN_IN ; P3_ADD_552_U175
g18153 nand P3_ADD_552_U134 P3_ADD_552_U37 ; P3_ADD_552_U176
g18154 nand P3_ADD_552_U121 P3_ADD_552_U35 ; P3_ADD_552_U177
g18155 nand P3_ADD_552_U36 P3_EBX_REG_21__SCAN_IN ; P3_ADD_552_U178
g18156 nand P3_ADD_552_U105 P3_EBX_REG_20__SCAN_IN ; P3_ADD_552_U179
g18157 nand P3_ADD_552_U135 P3_ADD_552_U32 ; P3_ADD_552_U180
g18158 nand P3_ADD_552_U7 P3_EBX_REG_0__SCAN_IN ; P3_ADD_552_U181
g18159 nand P3_ADD_552_U5 P3_EBX_REG_1__SCAN_IN ; P3_ADD_552_U182
g18160 nand P3_ADD_552_U114 P3_ADD_552_U33 ; P3_ADD_552_U183
g18161 nand P3_ADD_552_U34 P3_EBX_REG_19__SCAN_IN ; P3_ADD_552_U184
g18162 nand P3_ADD_552_U106 P3_EBX_REG_18__SCAN_IN ; P3_ADD_552_U185
g18163 nand P3_ADD_552_U136 P3_ADD_552_U29 ; P3_ADD_552_U186
g18164 nand P3_ADD_552_U117 P3_ADD_552_U30 ; P3_ADD_552_U187
g18165 nand P3_ADD_552_U31 P3_EBX_REG_17__SCAN_IN ; P3_ADD_552_U188
g18166 nand P3_ADD_552_U107 P3_EBX_REG_16__SCAN_IN ; P3_ADD_552_U189
g18167 nand P3_ADD_552_U137 P3_ADD_552_U28 ; P3_ADD_552_U190
g18168 nand P3_ADD_552_U124 P3_ADD_552_U26 ; P3_ADD_552_U191
g18169 nand P3_ADD_552_U27 P3_EBX_REG_15__SCAN_IN ; P3_ADD_552_U192
g18170 nand P3_ADD_552_U108 P3_EBX_REG_14__SCAN_IN ; P3_ADD_552_U193
g18171 nand P3_ADD_552_U138 P3_ADD_552_U23 ; P3_ADD_552_U194
g18172 nand P3_ADD_552_U119 P3_ADD_552_U24 ; P3_ADD_552_U195
g18173 nand P3_ADD_552_U25 P3_EBX_REG_13__SCAN_IN ; P3_ADD_552_U196
g18174 nand P3_ADD_552_U109 P3_EBX_REG_12__SCAN_IN ; P3_ADD_552_U197
g18175 nand P3_ADD_552_U139 P3_ADD_552_U20 ; P3_ADD_552_U198
g18176 nand P3_ADD_552_U113 P3_ADD_552_U21 ; P3_ADD_552_U199
g18177 nand P3_ADD_552_U22 P3_EBX_REG_11__SCAN_IN ; P3_ADD_552_U200
g18178 nand P3_ADD_552_U110 P3_EBX_REG_10__SCAN_IN ; P3_ADD_552_U201
g18179 nand P3_ADD_552_U140 P3_ADD_552_U19 ; P3_ADD_552_U202
g18180 not P3_EAX_REG_0__SCAN_IN ; P3_ADD_546_U5
g18181 not P3_EAX_REG_2__SCAN_IN ; P3_ADD_546_U6
g18182 not P3_EAX_REG_1__SCAN_IN ; P3_ADD_546_U7
g18183 not P3_EAX_REG_4__SCAN_IN ; P3_ADD_546_U8
g18184 not P3_EAX_REG_3__SCAN_IN ; P3_ADD_546_U9
g18185 nand P3_EAX_REG_0__SCAN_IN P3_EAX_REG_1__SCAN_IN P3_EAX_REG_2__SCAN_IN ; P3_ADD_546_U10
g18186 not P3_EAX_REG_6__SCAN_IN ; P3_ADD_546_U11
g18187 not P3_EAX_REG_5__SCAN_IN ; P3_ADD_546_U12
g18188 nand P3_ADD_546_U82 P3_ADD_546_U111 ; P3_ADD_546_U13
g18189 not P3_EAX_REG_8__SCAN_IN ; P3_ADD_546_U14
g18190 not P3_EAX_REG_7__SCAN_IN ; P3_ADD_546_U15
g18191 nand P3_ADD_546_U83 P3_ADD_546_U112 ; P3_ADD_546_U16
g18192 nand P3_ADD_546_U84 P3_ADD_546_U118 ; P3_ADD_546_U17
g18193 not P3_EAX_REG_9__SCAN_IN ; P3_ADD_546_U18
g18194 not P3_EAX_REG_10__SCAN_IN ; P3_ADD_546_U19
g18195 not P3_EAX_REG_12__SCAN_IN ; P3_ADD_546_U20
g18196 not P3_EAX_REG_11__SCAN_IN ; P3_ADD_546_U21
g18197 nand P3_ADD_546_U85 P3_ADD_546_U120 ; P3_ADD_546_U22
g18198 not P3_EAX_REG_14__SCAN_IN ; P3_ADD_546_U23
g18199 not P3_EAX_REG_13__SCAN_IN ; P3_ADD_546_U24
g18200 nand P3_ADD_546_U86 P3_ADD_546_U113 ; P3_ADD_546_U25
g18201 not P3_EAX_REG_15__SCAN_IN ; P3_ADD_546_U26
g18202 nand P3_ADD_546_U87 P3_ADD_546_U119 ; P3_ADD_546_U27
g18203 not P3_EAX_REG_16__SCAN_IN ; P3_ADD_546_U28
g18204 not P3_EAX_REG_18__SCAN_IN ; P3_ADD_546_U29
g18205 not P3_EAX_REG_17__SCAN_IN ; P3_ADD_546_U30
g18206 nand P3_ADD_546_U88 P3_ADD_546_U124 ; P3_ADD_546_U31
g18207 not P3_EAX_REG_20__SCAN_IN ; P3_ADD_546_U32
g18208 not P3_EAX_REG_19__SCAN_IN ; P3_ADD_546_U33
g18209 nand P3_ADD_546_U89 P3_ADD_546_U117 ; P3_ADD_546_U34
g18210 not P3_EAX_REG_21__SCAN_IN ; P3_ADD_546_U35
g18211 nand P3_ADD_546_U90 P3_ADD_546_U114 ; P3_ADD_546_U36
g18212 not P3_EAX_REG_22__SCAN_IN ; P3_ADD_546_U37
g18213 not P3_EAX_REG_24__SCAN_IN ; P3_ADD_546_U38
g18214 not P3_EAX_REG_23__SCAN_IN ; P3_ADD_546_U39
g18215 nand P3_ADD_546_U91 P3_ADD_546_U121 ; P3_ADD_546_U40
g18216 not P3_EAX_REG_26__SCAN_IN ; P3_ADD_546_U41
g18217 not P3_EAX_REG_25__SCAN_IN ; P3_ADD_546_U42
g18218 nand P3_ADD_546_U92 P3_ADD_546_U115 ; P3_ADD_546_U43
g18219 not P3_EAX_REG_27__SCAN_IN ; P3_ADD_546_U44
g18220 not P3_EAX_REG_28__SCAN_IN ; P3_ADD_546_U45
g18221 nand P3_ADD_546_U93 P3_ADD_546_U116 ; P3_ADD_546_U46
g18222 not P3_EAX_REG_29__SCAN_IN ; P3_ADD_546_U47
g18223 nand P3_ADD_546_U94 P3_ADD_546_U122 ; P3_ADD_546_U48
g18224 nand P3_ADD_546_U123 P3_EAX_REG_29__SCAN_IN ; P3_ADD_546_U49
g18225 not P3_EAX_REG_30__SCAN_IN ; P3_ADD_546_U50
g18226 nand P3_ADD_546_U142 P3_ADD_546_U141 ; P3_ADD_546_U51
g18227 nand P3_ADD_546_U144 P3_ADD_546_U143 ; P3_ADD_546_U52
g18228 nand P3_ADD_546_U146 P3_ADD_546_U145 ; P3_ADD_546_U53
g18229 nand P3_ADD_546_U148 P3_ADD_546_U147 ; P3_ADD_546_U54
g18230 nand P3_ADD_546_U150 P3_ADD_546_U149 ; P3_ADD_546_U55
g18231 nand P3_ADD_546_U152 P3_ADD_546_U151 ; P3_ADD_546_U56
g18232 nand P3_ADD_546_U154 P3_ADD_546_U153 ; P3_ADD_546_U57
g18233 nand P3_ADD_546_U156 P3_ADD_546_U155 ; P3_ADD_546_U58
g18234 nand P3_ADD_546_U158 P3_ADD_546_U157 ; P3_ADD_546_U59
g18235 nand P3_ADD_546_U160 P3_ADD_546_U159 ; P3_ADD_546_U60
g18236 nand P3_ADD_546_U162 P3_ADD_546_U161 ; P3_ADD_546_U61
g18237 nand P3_ADD_546_U164 P3_ADD_546_U163 ; P3_ADD_546_U62
g18238 nand P3_ADD_546_U166 P3_ADD_546_U165 ; P3_ADD_546_U63
g18239 nand P3_ADD_546_U168 P3_ADD_546_U167 ; P3_ADD_546_U64
g18240 nand P3_ADD_546_U170 P3_ADD_546_U169 ; P3_ADD_546_U65
g18241 nand P3_ADD_546_U172 P3_ADD_546_U171 ; P3_ADD_546_U66
g18242 nand P3_ADD_546_U174 P3_ADD_546_U173 ; P3_ADD_546_U67
g18243 nand P3_ADD_546_U176 P3_ADD_546_U175 ; P3_ADD_546_U68
g18244 nand P3_ADD_546_U178 P3_ADD_546_U177 ; P3_ADD_546_U69
g18245 nand P3_ADD_546_U180 P3_ADD_546_U179 ; P3_ADD_546_U70
g18246 nand P3_ADD_546_U182 P3_ADD_546_U181 ; P3_ADD_546_U71
g18247 nand P3_ADD_546_U184 P3_ADD_546_U183 ; P3_ADD_546_U72
g18248 nand P3_ADD_546_U186 P3_ADD_546_U185 ; P3_ADD_546_U73
g18249 nand P3_ADD_546_U188 P3_ADD_546_U187 ; P3_ADD_546_U74
g18250 nand P3_ADD_546_U190 P3_ADD_546_U189 ; P3_ADD_546_U75
g18251 nand P3_ADD_546_U192 P3_ADD_546_U191 ; P3_ADD_546_U76
g18252 nand P3_ADD_546_U194 P3_ADD_546_U193 ; P3_ADD_546_U77
g18253 nand P3_ADD_546_U196 P3_ADD_546_U195 ; P3_ADD_546_U78
g18254 nand P3_ADD_546_U198 P3_ADD_546_U197 ; P3_ADD_546_U79
g18255 nand P3_ADD_546_U200 P3_ADD_546_U199 ; P3_ADD_546_U80
g18256 nand P3_ADD_546_U202 P3_ADD_546_U201 ; P3_ADD_546_U81
g18257 and P3_EAX_REG_3__SCAN_IN P3_EAX_REG_4__SCAN_IN ; P3_ADD_546_U82
g18258 and P3_EAX_REG_5__SCAN_IN P3_EAX_REG_6__SCAN_IN ; P3_ADD_546_U83
g18259 and P3_EAX_REG_7__SCAN_IN P3_EAX_REG_8__SCAN_IN ; P3_ADD_546_U84
g18260 and P3_EAX_REG_9__SCAN_IN P3_EAX_REG_10__SCAN_IN ; P3_ADD_546_U85
g18261 and P3_EAX_REG_11__SCAN_IN P3_EAX_REG_12__SCAN_IN ; P3_ADD_546_U86
g18262 and P3_EAX_REG_13__SCAN_IN P3_EAX_REG_14__SCAN_IN ; P3_ADD_546_U87
g18263 and P3_EAX_REG_15__SCAN_IN P3_EAX_REG_16__SCAN_IN ; P3_ADD_546_U88
g18264 and P3_EAX_REG_17__SCAN_IN P3_EAX_REG_18__SCAN_IN ; P3_ADD_546_U89
g18265 and P3_EAX_REG_19__SCAN_IN P3_EAX_REG_20__SCAN_IN ; P3_ADD_546_U90
g18266 and P3_EAX_REG_21__SCAN_IN P3_EAX_REG_22__SCAN_IN ; P3_ADD_546_U91
g18267 and P3_EAX_REG_23__SCAN_IN P3_EAX_REG_24__SCAN_IN ; P3_ADD_546_U92
g18268 and P3_EAX_REG_25__SCAN_IN P3_EAX_REG_26__SCAN_IN ; P3_ADD_546_U93
g18269 and P3_EAX_REG_27__SCAN_IN P3_EAX_REG_28__SCAN_IN ; P3_ADD_546_U94
g18270 nand P3_ADD_546_U118 P3_EAX_REG_7__SCAN_IN ; P3_ADD_546_U95
g18271 nand P3_ADD_546_U112 P3_EAX_REG_5__SCAN_IN ; P3_ADD_546_U96
g18272 nand P3_ADD_546_U111 P3_EAX_REG_3__SCAN_IN ; P3_ADD_546_U97
g18273 not P3_EAX_REG_31__SCAN_IN ; P3_ADD_546_U98
g18274 nand P3_ADD_546_U128 P3_EAX_REG_30__SCAN_IN ; P3_ADD_546_U99
g18275 nand P3_EAX_REG_0__SCAN_IN P3_EAX_REG_1__SCAN_IN ; P3_ADD_546_U100
g18276 nand P3_ADD_546_U122 P3_EAX_REG_27__SCAN_IN ; P3_ADD_546_U101
g18277 nand P3_ADD_546_U116 P3_EAX_REG_25__SCAN_IN ; P3_ADD_546_U102
g18278 nand P3_ADD_546_U115 P3_EAX_REG_23__SCAN_IN ; P3_ADD_546_U103
g18279 nand P3_ADD_546_U121 P3_EAX_REG_21__SCAN_IN ; P3_ADD_546_U104
g18280 nand P3_ADD_546_U114 P3_EAX_REG_19__SCAN_IN ; P3_ADD_546_U105
g18281 nand P3_ADD_546_U117 P3_EAX_REG_17__SCAN_IN ; P3_ADD_546_U106
g18282 nand P3_ADD_546_U124 P3_EAX_REG_15__SCAN_IN ; P3_ADD_546_U107
g18283 nand P3_ADD_546_U119 P3_EAX_REG_13__SCAN_IN ; P3_ADD_546_U108
g18284 nand P3_ADD_546_U113 P3_EAX_REG_11__SCAN_IN ; P3_ADD_546_U109
g18285 nand P3_ADD_546_U120 P3_EAX_REG_9__SCAN_IN ; P3_ADD_546_U110
g18286 not P3_ADD_546_U10 ; P3_ADD_546_U111
g18287 not P3_ADD_546_U13 ; P3_ADD_546_U112
g18288 not P3_ADD_546_U22 ; P3_ADD_546_U113
g18289 not P3_ADD_546_U34 ; P3_ADD_546_U114
g18290 not P3_ADD_546_U40 ; P3_ADD_546_U115
g18291 not P3_ADD_546_U43 ; P3_ADD_546_U116
g18292 not P3_ADD_546_U31 ; P3_ADD_546_U117
g18293 not P3_ADD_546_U16 ; P3_ADD_546_U118
g18294 not P3_ADD_546_U25 ; P3_ADD_546_U119
g18295 not P3_ADD_546_U17 ; P3_ADD_546_U120
g18296 not P3_ADD_546_U36 ; P3_ADD_546_U121
g18297 not P3_ADD_546_U46 ; P3_ADD_546_U122
g18298 not P3_ADD_546_U48 ; P3_ADD_546_U123
g18299 not P3_ADD_546_U27 ; P3_ADD_546_U124
g18300 not P3_ADD_546_U95 ; P3_ADD_546_U125
g18301 not P3_ADD_546_U96 ; P3_ADD_546_U126
g18302 not P3_ADD_546_U97 ; P3_ADD_546_U127
g18303 not P3_ADD_546_U49 ; P3_ADD_546_U128
g18304 not P3_ADD_546_U99 ; P3_ADD_546_U129
g18305 not P3_ADD_546_U100 ; P3_ADD_546_U130
g18306 not P3_ADD_546_U101 ; P3_ADD_546_U131
g18307 not P3_ADD_546_U102 ; P3_ADD_546_U132
g18308 not P3_ADD_546_U103 ; P3_ADD_546_U133
g18309 not P3_ADD_546_U104 ; P3_ADD_546_U134
g18310 not P3_ADD_546_U105 ; P3_ADD_546_U135
g18311 not P3_ADD_546_U106 ; P3_ADD_546_U136
g18312 not P3_ADD_546_U107 ; P3_ADD_546_U137
g18313 not P3_ADD_546_U108 ; P3_ADD_546_U138
g18314 not P3_ADD_546_U109 ; P3_ADD_546_U139
g18315 not P3_ADD_546_U110 ; P3_ADD_546_U140
g18316 nand P3_ADD_546_U120 P3_ADD_546_U18 ; P3_ADD_546_U141
g18317 nand P3_ADD_546_U17 P3_EAX_REG_9__SCAN_IN ; P3_ADD_546_U142
g18318 nand P3_ADD_546_U95 P3_EAX_REG_8__SCAN_IN ; P3_ADD_546_U143
g18319 nand P3_ADD_546_U125 P3_ADD_546_U14 ; P3_ADD_546_U144
g18320 nand P3_ADD_546_U118 P3_ADD_546_U15 ; P3_ADD_546_U145
g18321 nand P3_ADD_546_U16 P3_EAX_REG_7__SCAN_IN ; P3_ADD_546_U146
g18322 nand P3_ADD_546_U96 P3_EAX_REG_6__SCAN_IN ; P3_ADD_546_U147
g18323 nand P3_ADD_546_U126 P3_ADD_546_U11 ; P3_ADD_546_U148
g18324 nand P3_ADD_546_U112 P3_ADD_546_U12 ; P3_ADD_546_U149
g18325 nand P3_ADD_546_U13 P3_EAX_REG_5__SCAN_IN ; P3_ADD_546_U150
g18326 nand P3_ADD_546_U97 P3_EAX_REG_4__SCAN_IN ; P3_ADD_546_U151
g18327 nand P3_ADD_546_U127 P3_ADD_546_U8 ; P3_ADD_546_U152
g18328 nand P3_ADD_546_U111 P3_ADD_546_U9 ; P3_ADD_546_U153
g18329 nand P3_ADD_546_U10 P3_EAX_REG_3__SCAN_IN ; P3_ADD_546_U154
g18330 nand P3_ADD_546_U99 P3_EAX_REG_31__SCAN_IN ; P3_ADD_546_U155
g18331 nand P3_ADD_546_U129 P3_ADD_546_U98 ; P3_ADD_546_U156
g18332 nand P3_ADD_546_U49 P3_EAX_REG_30__SCAN_IN ; P3_ADD_546_U157
g18333 nand P3_ADD_546_U128 P3_ADD_546_U50 ; P3_ADD_546_U158
g18334 nand P3_ADD_546_U100 P3_EAX_REG_2__SCAN_IN ; P3_ADD_546_U159
g18335 nand P3_ADD_546_U130 P3_ADD_546_U6 ; P3_ADD_546_U160
g18336 nand P3_ADD_546_U123 P3_ADD_546_U47 ; P3_ADD_546_U161
g18337 nand P3_ADD_546_U48 P3_EAX_REG_29__SCAN_IN ; P3_ADD_546_U162
g18338 nand P3_ADD_546_U101 P3_EAX_REG_28__SCAN_IN ; P3_ADD_546_U163
g18339 nand P3_ADD_546_U131 P3_ADD_546_U45 ; P3_ADD_546_U164
g18340 nand P3_ADD_546_U122 P3_ADD_546_U44 ; P3_ADD_546_U165
g18341 nand P3_ADD_546_U46 P3_EAX_REG_27__SCAN_IN ; P3_ADD_546_U166
g18342 nand P3_ADD_546_U102 P3_EAX_REG_26__SCAN_IN ; P3_ADD_546_U167
g18343 nand P3_ADD_546_U132 P3_ADD_546_U41 ; P3_ADD_546_U168
g18344 nand P3_ADD_546_U116 P3_ADD_546_U42 ; P3_ADD_546_U169
g18345 nand P3_ADD_546_U43 P3_EAX_REG_25__SCAN_IN ; P3_ADD_546_U170
g18346 nand P3_ADD_546_U103 P3_EAX_REG_24__SCAN_IN ; P3_ADD_546_U171
g18347 nand P3_ADD_546_U133 P3_ADD_546_U38 ; P3_ADD_546_U172
g18348 nand P3_ADD_546_U115 P3_ADD_546_U39 ; P3_ADD_546_U173
g18349 nand P3_ADD_546_U40 P3_EAX_REG_23__SCAN_IN ; P3_ADD_546_U174
g18350 nand P3_ADD_546_U104 P3_EAX_REG_22__SCAN_IN ; P3_ADD_546_U175
g18351 nand P3_ADD_546_U134 P3_ADD_546_U37 ; P3_ADD_546_U176
g18352 nand P3_ADD_546_U121 P3_ADD_546_U35 ; P3_ADD_546_U177
g18353 nand P3_ADD_546_U36 P3_EAX_REG_21__SCAN_IN ; P3_ADD_546_U178
g18354 nand P3_ADD_546_U105 P3_EAX_REG_20__SCAN_IN ; P3_ADD_546_U179
g18355 nand P3_ADD_546_U135 P3_ADD_546_U32 ; P3_ADD_546_U180
g18356 nand P3_ADD_546_U7 P3_EAX_REG_0__SCAN_IN ; P3_ADD_546_U181
g18357 nand P3_ADD_546_U5 P3_EAX_REG_1__SCAN_IN ; P3_ADD_546_U182
g18358 nand P3_ADD_546_U114 P3_ADD_546_U33 ; P3_ADD_546_U183
g18359 nand P3_ADD_546_U34 P3_EAX_REG_19__SCAN_IN ; P3_ADD_546_U184
g18360 nand P3_ADD_546_U106 P3_EAX_REG_18__SCAN_IN ; P3_ADD_546_U185
g18361 nand P3_ADD_546_U136 P3_ADD_546_U29 ; P3_ADD_546_U186
g18362 nand P3_ADD_546_U117 P3_ADD_546_U30 ; P3_ADD_546_U187
g18363 nand P3_ADD_546_U31 P3_EAX_REG_17__SCAN_IN ; P3_ADD_546_U188
g18364 nand P3_ADD_546_U107 P3_EAX_REG_16__SCAN_IN ; P3_ADD_546_U189
g18365 nand P3_ADD_546_U137 P3_ADD_546_U28 ; P3_ADD_546_U190
g18366 nand P3_ADD_546_U124 P3_ADD_546_U26 ; P3_ADD_546_U191
g18367 nand P3_ADD_546_U27 P3_EAX_REG_15__SCAN_IN ; P3_ADD_546_U192
g18368 nand P3_ADD_546_U108 P3_EAX_REG_14__SCAN_IN ; P3_ADD_546_U193
g18369 nand P3_ADD_546_U138 P3_ADD_546_U23 ; P3_ADD_546_U194
g18370 nand P3_ADD_546_U119 P3_ADD_546_U24 ; P3_ADD_546_U195
g18371 nand P3_ADD_546_U25 P3_EAX_REG_13__SCAN_IN ; P3_ADD_546_U196
g18372 nand P3_ADD_546_U109 P3_EAX_REG_12__SCAN_IN ; P3_ADD_546_U197
g18373 nand P3_ADD_546_U139 P3_ADD_546_U20 ; P3_ADD_546_U198
g18374 nand P3_ADD_546_U113 P3_ADD_546_U21 ; P3_ADD_546_U199
g18375 nand P3_ADD_546_U22 P3_EAX_REG_11__SCAN_IN ; P3_ADD_546_U200
g18376 nand P3_ADD_546_U110 P3_EAX_REG_10__SCAN_IN ; P3_ADD_546_U201
g18377 nand P3_ADD_546_U140 P3_ADD_546_U19 ; P3_ADD_546_U202
g18378 nor P3_SUB_401_U6 P3_GTE_401_U8 ; P3_GTE_401_U6
g18379 and P3_SUB_401_U21 P3_GTE_401_U9 ; P3_GTE_401_U7
g18380 nor P3_SUB_401_U19 P3_SUB_401_U20 P3_GTE_401_U7 ; P3_GTE_401_U8
g18381 or P3_SUB_401_U7 P3_SUB_401_U22 ; P3_GTE_401_U9
g18382 not P3_U2613 ; P3_ADD_391_1180_U4
g18383 not P3_U3069 ; P3_ADD_391_1180_U5
g18384 nand P3_U3069 P3_U2613 ; P3_ADD_391_1180_U6
g18385 not P3_U2614 ; P3_ADD_391_1180_U7
g18386 nand P3_U2614 P3_ADD_391_1180_U28 ; P3_ADD_391_1180_U8
g18387 not P3_U2615 ; P3_ADD_391_1180_U9
g18388 nand P3_U2615 P3_ADD_391_1180_U29 ; P3_ADD_391_1180_U10
g18389 not P3_U2616 ; P3_ADD_391_1180_U11
g18390 nand P3_U2616 P3_ADD_391_1180_U30 ; P3_ADD_391_1180_U12
g18391 not P3_U2617 ; P3_ADD_391_1180_U13
g18392 nand P3_U2617 P3_ADD_391_1180_U31 ; P3_ADD_391_1180_U14
g18393 not P3_U2618 ; P3_ADD_391_1180_U15
g18394 nand P3_U2618 P3_ADD_391_1180_U32 ; P3_ADD_391_1180_U16
g18395 not P3_U2619 ; P3_ADD_391_1180_U17
g18396 nand P3_ADD_391_1180_U36 P3_ADD_391_1180_U35 ; P3_ADD_391_1180_U18
g18397 nand P3_ADD_391_1180_U38 P3_ADD_391_1180_U37 ; P3_ADD_391_1180_U19
g18398 nand P3_ADD_391_1180_U40 P3_ADD_391_1180_U39 ; P3_ADD_391_1180_U20
g18399 nand P3_ADD_391_1180_U42 P3_ADD_391_1180_U41 ; P3_ADD_391_1180_U21
g18400 nand P3_ADD_391_1180_U44 P3_ADD_391_1180_U43 ; P3_ADD_391_1180_U22
g18401 nand P3_ADD_391_1180_U46 P3_ADD_391_1180_U45 ; P3_ADD_391_1180_U23
g18402 nand P3_ADD_391_1180_U48 P3_ADD_391_1180_U47 ; P3_ADD_391_1180_U24
g18403 nand P3_ADD_391_1180_U50 P3_ADD_391_1180_U49 ; P3_ADD_391_1180_U25
g18404 not P3_U2620 ; P3_ADD_391_1180_U26
g18405 nand P3_U2619 P3_ADD_391_1180_U33 ; P3_ADD_391_1180_U27
g18406 not P3_ADD_391_1180_U6 ; P3_ADD_391_1180_U28
g18407 not P3_ADD_391_1180_U8 ; P3_ADD_391_1180_U29
g18408 not P3_ADD_391_1180_U10 ; P3_ADD_391_1180_U30
g18409 not P3_ADD_391_1180_U12 ; P3_ADD_391_1180_U31
g18410 not P3_ADD_391_1180_U14 ; P3_ADD_391_1180_U32
g18411 not P3_ADD_391_1180_U16 ; P3_ADD_391_1180_U33
g18412 not P3_ADD_391_1180_U27 ; P3_ADD_391_1180_U34
g18413 nand P3_U2620 P3_ADD_391_1180_U27 ; P3_ADD_391_1180_U35
g18414 nand P3_ADD_391_1180_U34 P3_ADD_391_1180_U26 ; P3_ADD_391_1180_U36
g18415 nand P3_U2619 P3_ADD_391_1180_U16 ; P3_ADD_391_1180_U37
g18416 nand P3_ADD_391_1180_U33 P3_ADD_391_1180_U17 ; P3_ADD_391_1180_U38
g18417 nand P3_U2618 P3_ADD_391_1180_U14 ; P3_ADD_391_1180_U39
g18418 nand P3_ADD_391_1180_U32 P3_ADD_391_1180_U15 ; P3_ADD_391_1180_U40
g18419 nand P3_U2617 P3_ADD_391_1180_U12 ; P3_ADD_391_1180_U41
g18420 nand P3_ADD_391_1180_U31 P3_ADD_391_1180_U13 ; P3_ADD_391_1180_U42
g18421 nand P3_U2616 P3_ADD_391_1180_U10 ; P3_ADD_391_1180_U43
g18422 nand P3_ADD_391_1180_U30 P3_ADD_391_1180_U11 ; P3_ADD_391_1180_U44
g18423 nand P3_U2615 P3_ADD_391_1180_U8 ; P3_ADD_391_1180_U45
g18424 nand P3_ADD_391_1180_U29 P3_ADD_391_1180_U9 ; P3_ADD_391_1180_U46
g18425 nand P3_U2614 P3_ADD_391_1180_U6 ; P3_ADD_391_1180_U47
g18426 nand P3_ADD_391_1180_U28 P3_ADD_391_1180_U7 ; P3_ADD_391_1180_U48
g18427 nand P3_U3069 P3_ADD_391_1180_U4 ; P3_ADD_391_1180_U49
g18428 nand P3_U2613 P3_ADD_391_1180_U5 ; P3_ADD_391_1180_U50
g18429 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_476_U4
g18430 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_476_U5
g18431 nand P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_476_U6
g18432 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_476_U7
g18433 nand P3_ADD_476_U94 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_476_U8
g18434 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_476_U9
g18435 nand P3_ADD_476_U95 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_476_U10
g18436 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_476_U11
g18437 nand P3_ADD_476_U96 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_476_U12
g18438 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_476_U13
g18439 nand P3_ADD_476_U97 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_476_U14
g18440 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_476_U15
g18441 nand P3_ADD_476_U98 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_476_U16
g18442 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_476_U17
g18443 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_476_U18
g18444 nand P3_ADD_476_U99 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_476_U19
g18445 nand P3_ADD_476_U100 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_476_U20
g18446 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_476_U21
g18447 nand P3_ADD_476_U101 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_476_U22
g18448 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_476_U23
g18449 nand P3_ADD_476_U102 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_476_U24
g18450 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_476_U25
g18451 nand P3_ADD_476_U103 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_476_U26
g18452 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_476_U27
g18453 nand P3_ADD_476_U104 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_476_U28
g18454 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_476_U29
g18455 nand P3_ADD_476_U105 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_476_U30
g18456 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_476_U31
g18457 nand P3_ADD_476_U106 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_476_U32
g18458 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_476_U33
g18459 nand P3_ADD_476_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_476_U34
g18460 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_476_U35
g18461 nand P3_ADD_476_U108 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_476_U36
g18462 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_476_U37
g18463 nand P3_ADD_476_U109 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_476_U38
g18464 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_476_U39
g18465 nand P3_ADD_476_U110 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_476_U40
g18466 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_476_U41
g18467 nand P3_ADD_476_U111 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_476_U42
g18468 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_476_U43
g18469 nand P3_ADD_476_U112 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_476_U44
g18470 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_476_U45
g18471 nand P3_ADD_476_U113 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_476_U46
g18472 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_476_U47
g18473 nand P3_ADD_476_U114 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_476_U48
g18474 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_476_U49
g18475 nand P3_ADD_476_U115 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_476_U50
g18476 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_476_U51
g18477 nand P3_ADD_476_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_476_U52
g18478 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_476_U53
g18479 nand P3_ADD_476_U117 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_476_U54
g18480 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_476_U55
g18481 nand P3_ADD_476_U118 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_476_U56
g18482 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_476_U57
g18483 nand P3_ADD_476_U119 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_476_U58
g18484 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_476_U59
g18485 nand P3_ADD_476_U120 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_476_U60
g18486 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_476_U61
g18487 nand P3_ADD_476_U124 P3_ADD_476_U123 ; P3_ADD_476_U62
g18488 nand P3_ADD_476_U126 P3_ADD_476_U125 ; P3_ADD_476_U63
g18489 nand P3_ADD_476_U128 P3_ADD_476_U127 ; P3_ADD_476_U64
g18490 nand P3_ADD_476_U130 P3_ADD_476_U129 ; P3_ADD_476_U65
g18491 nand P3_ADD_476_U132 P3_ADD_476_U131 ; P3_ADD_476_U66
g18492 nand P3_ADD_476_U134 P3_ADD_476_U133 ; P3_ADD_476_U67
g18493 nand P3_ADD_476_U136 P3_ADD_476_U135 ; P3_ADD_476_U68
g18494 nand P3_ADD_476_U138 P3_ADD_476_U137 ; P3_ADD_476_U69
g18495 nand P3_ADD_476_U140 P3_ADD_476_U139 ; P3_ADD_476_U70
g18496 nand P3_ADD_476_U142 P3_ADD_476_U141 ; P3_ADD_476_U71
g18497 nand P3_ADD_476_U144 P3_ADD_476_U143 ; P3_ADD_476_U72
g18498 nand P3_ADD_476_U146 P3_ADD_476_U145 ; P3_ADD_476_U73
g18499 nand P3_ADD_476_U148 P3_ADD_476_U147 ; P3_ADD_476_U74
g18500 nand P3_ADD_476_U150 P3_ADD_476_U149 ; P3_ADD_476_U75
g18501 nand P3_ADD_476_U152 P3_ADD_476_U151 ; P3_ADD_476_U76
g18502 nand P3_ADD_476_U154 P3_ADD_476_U153 ; P3_ADD_476_U77
g18503 nand P3_ADD_476_U156 P3_ADD_476_U155 ; P3_ADD_476_U78
g18504 nand P3_ADD_476_U158 P3_ADD_476_U157 ; P3_ADD_476_U79
g18505 nand P3_ADD_476_U160 P3_ADD_476_U159 ; P3_ADD_476_U80
g18506 nand P3_ADD_476_U162 P3_ADD_476_U161 ; P3_ADD_476_U81
g18507 nand P3_ADD_476_U164 P3_ADD_476_U163 ; P3_ADD_476_U82
g18508 nand P3_ADD_476_U166 P3_ADD_476_U165 ; P3_ADD_476_U83
g18509 nand P3_ADD_476_U168 P3_ADD_476_U167 ; P3_ADD_476_U84
g18510 nand P3_ADD_476_U170 P3_ADD_476_U169 ; P3_ADD_476_U85
g18511 nand P3_ADD_476_U172 P3_ADD_476_U171 ; P3_ADD_476_U86
g18512 nand P3_ADD_476_U174 P3_ADD_476_U173 ; P3_ADD_476_U87
g18513 nand P3_ADD_476_U176 P3_ADD_476_U175 ; P3_ADD_476_U88
g18514 nand P3_ADD_476_U178 P3_ADD_476_U177 ; P3_ADD_476_U89
g18515 nand P3_ADD_476_U180 P3_ADD_476_U179 ; P3_ADD_476_U90
g18516 nand P3_ADD_476_U182 P3_ADD_476_U181 ; P3_ADD_476_U91
g18517 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_476_U92
g18518 nand P3_ADD_476_U121 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_476_U93
g18519 not P3_ADD_476_U6 ; P3_ADD_476_U94
g18520 not P3_ADD_476_U8 ; P3_ADD_476_U95
g18521 not P3_ADD_476_U10 ; P3_ADD_476_U96
g18522 not P3_ADD_476_U12 ; P3_ADD_476_U97
g18523 not P3_ADD_476_U14 ; P3_ADD_476_U98
g18524 not P3_ADD_476_U16 ; P3_ADD_476_U99
g18525 not P3_ADD_476_U19 ; P3_ADD_476_U100
g18526 not P3_ADD_476_U20 ; P3_ADD_476_U101
g18527 not P3_ADD_476_U22 ; P3_ADD_476_U102
g18528 not P3_ADD_476_U24 ; P3_ADD_476_U103
g18529 not P3_ADD_476_U26 ; P3_ADD_476_U104
g18530 not P3_ADD_476_U28 ; P3_ADD_476_U105
g18531 not P3_ADD_476_U30 ; P3_ADD_476_U106
g18532 not P3_ADD_476_U32 ; P3_ADD_476_U107
g18533 not P3_ADD_476_U34 ; P3_ADD_476_U108
g18534 not P3_ADD_476_U36 ; P3_ADD_476_U109
g18535 not P3_ADD_476_U38 ; P3_ADD_476_U110
g18536 not P3_ADD_476_U40 ; P3_ADD_476_U111
g18537 not P3_ADD_476_U42 ; P3_ADD_476_U112
g18538 not P3_ADD_476_U44 ; P3_ADD_476_U113
g18539 not P3_ADD_476_U46 ; P3_ADD_476_U114
g18540 not P3_ADD_476_U48 ; P3_ADD_476_U115
g18541 not P3_ADD_476_U50 ; P3_ADD_476_U116
g18542 not P3_ADD_476_U52 ; P3_ADD_476_U117
g18543 not P3_ADD_476_U54 ; P3_ADD_476_U118
g18544 not P3_ADD_476_U56 ; P3_ADD_476_U119
g18545 not P3_ADD_476_U58 ; P3_ADD_476_U120
g18546 not P3_ADD_476_U60 ; P3_ADD_476_U121
g18547 not P3_ADD_476_U93 ; P3_ADD_476_U122
g18548 nand P3_ADD_476_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_476_U123
g18549 nand P3_ADD_476_U100 P3_ADD_476_U18 ; P3_ADD_476_U124
g18550 nand P3_ADD_476_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_476_U125
g18551 nand P3_ADD_476_U99 P3_ADD_476_U17 ; P3_ADD_476_U126
g18552 nand P3_ADD_476_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_476_U127
g18553 nand P3_ADD_476_U98 P3_ADD_476_U15 ; P3_ADD_476_U128
g18554 nand P3_ADD_476_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_476_U129
g18555 nand P3_ADD_476_U97 P3_ADD_476_U13 ; P3_ADD_476_U130
g18556 nand P3_ADD_476_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_476_U131
g18557 nand P3_ADD_476_U96 P3_ADD_476_U11 ; P3_ADD_476_U132
g18558 nand P3_ADD_476_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_476_U133
g18559 nand P3_ADD_476_U95 P3_ADD_476_U9 ; P3_ADD_476_U134
g18560 nand P3_ADD_476_U6 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_476_U135
g18561 nand P3_ADD_476_U94 P3_ADD_476_U7 ; P3_ADD_476_U136
g18562 nand P3_ADD_476_U93 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_476_U137
g18563 nand P3_ADD_476_U122 P3_ADD_476_U92 ; P3_ADD_476_U138
g18564 nand P3_ADD_476_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_476_U139
g18565 nand P3_ADD_476_U121 P3_ADD_476_U61 ; P3_ADD_476_U140
g18566 nand P3_ADD_476_U4 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_476_U141
g18567 nand P3_ADD_476_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_476_U142
g18568 nand P3_ADD_476_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_476_U143
g18569 nand P3_ADD_476_U120 P3_ADD_476_U59 ; P3_ADD_476_U144
g18570 nand P3_ADD_476_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_476_U145
g18571 nand P3_ADD_476_U119 P3_ADD_476_U57 ; P3_ADD_476_U146
g18572 nand P3_ADD_476_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_476_U147
g18573 nand P3_ADD_476_U118 P3_ADD_476_U55 ; P3_ADD_476_U148
g18574 nand P3_ADD_476_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_476_U149
g18575 nand P3_ADD_476_U117 P3_ADD_476_U53 ; P3_ADD_476_U150
g18576 nand P3_ADD_476_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_476_U151
g18577 nand P3_ADD_476_U116 P3_ADD_476_U51 ; P3_ADD_476_U152
g18578 nand P3_ADD_476_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_476_U153
g18579 nand P3_ADD_476_U115 P3_ADD_476_U49 ; P3_ADD_476_U154
g18580 nand P3_ADD_476_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_476_U155
g18581 nand P3_ADD_476_U114 P3_ADD_476_U47 ; P3_ADD_476_U156
g18582 nand P3_ADD_476_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_476_U157
g18583 nand P3_ADD_476_U113 P3_ADD_476_U45 ; P3_ADD_476_U158
g18584 nand P3_ADD_476_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_476_U159
g18585 nand P3_ADD_476_U112 P3_ADD_476_U43 ; P3_ADD_476_U160
g18586 nand P3_ADD_476_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_476_U161
g18587 nand P3_ADD_476_U111 P3_ADD_476_U41 ; P3_ADD_476_U162
g18588 nand P3_ADD_476_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_476_U163
g18589 nand P3_ADD_476_U110 P3_ADD_476_U39 ; P3_ADD_476_U164
g18590 nand P3_ADD_476_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_476_U165
g18591 nand P3_ADD_476_U109 P3_ADD_476_U37 ; P3_ADD_476_U166
g18592 nand P3_ADD_476_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_476_U167
g18593 nand P3_ADD_476_U108 P3_ADD_476_U35 ; P3_ADD_476_U168
g18594 nand P3_ADD_476_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_476_U169
g18595 nand P3_ADD_476_U107 P3_ADD_476_U33 ; P3_ADD_476_U170
g18596 nand P3_ADD_476_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_476_U171
g18597 nand P3_ADD_476_U106 P3_ADD_476_U31 ; P3_ADD_476_U172
g18598 nand P3_ADD_476_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_476_U173
g18599 nand P3_ADD_476_U105 P3_ADD_476_U29 ; P3_ADD_476_U174
g18600 nand P3_ADD_476_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_476_U175
g18601 nand P3_ADD_476_U104 P3_ADD_476_U27 ; P3_ADD_476_U176
g18602 nand P3_ADD_476_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_476_U177
g18603 nand P3_ADD_476_U103 P3_ADD_476_U25 ; P3_ADD_476_U178
g18604 nand P3_ADD_476_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_476_U179
g18605 nand P3_ADD_476_U102 P3_ADD_476_U23 ; P3_ADD_476_U180
g18606 nand P3_ADD_476_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_476_U181
g18607 nand P3_ADD_476_U101 P3_ADD_476_U21 ; P3_ADD_476_U182
g18608 nor P3_SUB_390_U6 P3_GTE_390_U8 ; P3_GTE_390_U6
g18609 and P3_SUB_390_U21 P3_GTE_390_U9 ; P3_GTE_390_U7
g18610 nor P3_SUB_390_U19 P3_SUB_390_U20 P3_GTE_390_U7 ; P3_GTE_390_U8
g18611 or P3_SUB_390_U7 P3_SUB_390_U22 ; P3_GTE_390_U9
g18612 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_531_U5
g18613 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_531_U6
g18614 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_531_U7
g18615 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_531_U8
g18616 nand P3_ADD_531_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_531_U9
g18617 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_531_U10
g18618 nand P3_ADD_531_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_531_U11
g18619 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_531_U12
g18620 nand P3_ADD_531_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_531_U13
g18621 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_531_U14
g18622 nand P3_ADD_531_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_531_U15
g18623 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_531_U16
g18624 nand P3_ADD_531_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_531_U17
g18625 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_531_U18
g18626 nand P3_ADD_531_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_531_U19
g18627 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_531_U20
g18628 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_531_U21
g18629 nand P3_ADD_531_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_531_U22
g18630 nand P3_ADD_531_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_531_U23
g18631 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_531_U24
g18632 nand P3_ADD_531_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_531_U25
g18633 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_531_U26
g18634 nand P3_ADD_531_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_531_U27
g18635 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_531_U28
g18636 nand P3_ADD_531_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_531_U29
g18637 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_531_U30
g18638 nand P3_ADD_531_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_531_U31
g18639 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_531_U32
g18640 nand P3_ADD_531_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_531_U33
g18641 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_531_U34
g18642 nand P3_ADD_531_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_531_U35
g18643 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_531_U36
g18644 nand P3_ADD_531_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_531_U37
g18645 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_531_U38
g18646 nand P3_ADD_531_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_531_U39
g18647 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_531_U40
g18648 nand P3_ADD_531_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_531_U41
g18649 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_531_U42
g18650 nand P3_ADD_531_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_531_U43
g18651 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_531_U44
g18652 nand P3_ADD_531_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_531_U45
g18653 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_531_U46
g18654 nand P3_ADD_531_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_531_U47
g18655 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_531_U48
g18656 nand P3_ADD_531_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_531_U49
g18657 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_531_U50
g18658 nand P3_ADD_531_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_531_U51
g18659 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_531_U52
g18660 nand P3_ADD_531_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_531_U53
g18661 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_531_U54
g18662 nand P3_ADD_531_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_531_U55
g18663 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_531_U56
g18664 nand P3_ADD_531_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_531_U57
g18665 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_531_U58
g18666 nand P3_ADD_531_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_531_U59
g18667 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_531_U60
g18668 nand P3_ADD_531_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_531_U61
g18669 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_531_U62
g18670 nand P3_ADD_531_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_531_U63
g18671 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_531_U64
g18672 nand P3_ADD_531_U129 P3_ADD_531_U128 ; P3_ADD_531_U65
g18673 nand P3_ADD_531_U131 P3_ADD_531_U130 ; P3_ADD_531_U66
g18674 nand P3_ADD_531_U133 P3_ADD_531_U132 ; P3_ADD_531_U67
g18675 nand P3_ADD_531_U135 P3_ADD_531_U134 ; P3_ADD_531_U68
g18676 nand P3_ADD_531_U137 P3_ADD_531_U136 ; P3_ADD_531_U69
g18677 nand P3_ADD_531_U139 P3_ADD_531_U138 ; P3_ADD_531_U70
g18678 nand P3_ADD_531_U141 P3_ADD_531_U140 ; P3_ADD_531_U71
g18679 nand P3_ADD_531_U143 P3_ADD_531_U142 ; P3_ADD_531_U72
g18680 nand P3_ADD_531_U145 P3_ADD_531_U144 ; P3_ADD_531_U73
g18681 nand P3_ADD_531_U147 P3_ADD_531_U146 ; P3_ADD_531_U74
g18682 nand P3_ADD_531_U149 P3_ADD_531_U148 ; P3_ADD_531_U75
g18683 nand P3_ADD_531_U151 P3_ADD_531_U150 ; P3_ADD_531_U76
g18684 nand P3_ADD_531_U153 P3_ADD_531_U152 ; P3_ADD_531_U77
g18685 nand P3_ADD_531_U155 P3_ADD_531_U154 ; P3_ADD_531_U78
g18686 nand P3_ADD_531_U157 P3_ADD_531_U156 ; P3_ADD_531_U79
g18687 nand P3_ADD_531_U159 P3_ADD_531_U158 ; P3_ADD_531_U80
g18688 nand P3_ADD_531_U161 P3_ADD_531_U160 ; P3_ADD_531_U81
g18689 nand P3_ADD_531_U163 P3_ADD_531_U162 ; P3_ADD_531_U82
g18690 nand P3_ADD_531_U165 P3_ADD_531_U164 ; P3_ADD_531_U83
g18691 nand P3_ADD_531_U167 P3_ADD_531_U166 ; P3_ADD_531_U84
g18692 nand P3_ADD_531_U169 P3_ADD_531_U168 ; P3_ADD_531_U85
g18693 nand P3_ADD_531_U171 P3_ADD_531_U170 ; P3_ADD_531_U86
g18694 nand P3_ADD_531_U173 P3_ADD_531_U172 ; P3_ADD_531_U87
g18695 nand P3_ADD_531_U175 P3_ADD_531_U174 ; P3_ADD_531_U88
g18696 nand P3_ADD_531_U177 P3_ADD_531_U176 ; P3_ADD_531_U89
g18697 nand P3_ADD_531_U179 P3_ADD_531_U178 ; P3_ADD_531_U90
g18698 nand P3_ADD_531_U181 P3_ADD_531_U180 ; P3_ADD_531_U91
g18699 nand P3_ADD_531_U183 P3_ADD_531_U182 ; P3_ADD_531_U92
g18700 nand P3_ADD_531_U185 P3_ADD_531_U184 ; P3_ADD_531_U93
g18701 nand P3_ADD_531_U187 P3_ADD_531_U186 ; P3_ADD_531_U94
g18702 nand P3_ADD_531_U189 P3_ADD_531_U188 ; P3_ADD_531_U95
g18703 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_531_U96
g18704 nand P3_ADD_531_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_531_U97
g18705 not P3_ADD_531_U7 ; P3_ADD_531_U98
g18706 not P3_ADD_531_U9 ; P3_ADD_531_U99
g18707 not P3_ADD_531_U11 ; P3_ADD_531_U100
g18708 not P3_ADD_531_U13 ; P3_ADD_531_U101
g18709 not P3_ADD_531_U15 ; P3_ADD_531_U102
g18710 not P3_ADD_531_U17 ; P3_ADD_531_U103
g18711 not P3_ADD_531_U19 ; P3_ADD_531_U104
g18712 not P3_ADD_531_U22 ; P3_ADD_531_U105
g18713 not P3_ADD_531_U23 ; P3_ADD_531_U106
g18714 not P3_ADD_531_U25 ; P3_ADD_531_U107
g18715 not P3_ADD_531_U27 ; P3_ADD_531_U108
g18716 not P3_ADD_531_U29 ; P3_ADD_531_U109
g18717 not P3_ADD_531_U31 ; P3_ADD_531_U110
g18718 not P3_ADD_531_U33 ; P3_ADD_531_U111
g18719 not P3_ADD_531_U35 ; P3_ADD_531_U112
g18720 not P3_ADD_531_U37 ; P3_ADD_531_U113
g18721 not P3_ADD_531_U39 ; P3_ADD_531_U114
g18722 not P3_ADD_531_U41 ; P3_ADD_531_U115
g18723 not P3_ADD_531_U43 ; P3_ADD_531_U116
g18724 not P3_ADD_531_U45 ; P3_ADD_531_U117
g18725 not P3_ADD_531_U47 ; P3_ADD_531_U118
g18726 not P3_ADD_531_U49 ; P3_ADD_531_U119
g18727 not P3_ADD_531_U51 ; P3_ADD_531_U120
g18728 not P3_ADD_531_U53 ; P3_ADD_531_U121
g18729 not P3_ADD_531_U55 ; P3_ADD_531_U122
g18730 not P3_ADD_531_U57 ; P3_ADD_531_U123
g18731 not P3_ADD_531_U59 ; P3_ADD_531_U124
g18732 not P3_ADD_531_U61 ; P3_ADD_531_U125
g18733 not P3_ADD_531_U63 ; P3_ADD_531_U126
g18734 not P3_ADD_531_U97 ; P3_ADD_531_U127
g18735 nand P3_ADD_531_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_531_U128
g18736 nand P3_ADD_531_U105 P3_ADD_531_U21 ; P3_ADD_531_U129
g18737 nand P3_ADD_531_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_531_U130
g18738 nand P3_ADD_531_U104 P3_ADD_531_U20 ; P3_ADD_531_U131
g18739 nand P3_ADD_531_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_531_U132
g18740 nand P3_ADD_531_U103 P3_ADD_531_U18 ; P3_ADD_531_U133
g18741 nand P3_ADD_531_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_531_U134
g18742 nand P3_ADD_531_U102 P3_ADD_531_U16 ; P3_ADD_531_U135
g18743 nand P3_ADD_531_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_531_U136
g18744 nand P3_ADD_531_U101 P3_ADD_531_U14 ; P3_ADD_531_U137
g18745 nand P3_ADD_531_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_531_U138
g18746 nand P3_ADD_531_U100 P3_ADD_531_U12 ; P3_ADD_531_U139
g18747 nand P3_ADD_531_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_531_U140
g18748 nand P3_ADD_531_U99 P3_ADD_531_U10 ; P3_ADD_531_U141
g18749 nand P3_ADD_531_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_531_U142
g18750 nand P3_ADD_531_U127 P3_ADD_531_U96 ; P3_ADD_531_U143
g18751 nand P3_ADD_531_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_531_U144
g18752 nand P3_ADD_531_U126 P3_ADD_531_U64 ; P3_ADD_531_U145
g18753 nand P3_ADD_531_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_531_U146
g18754 nand P3_ADD_531_U98 P3_ADD_531_U8 ; P3_ADD_531_U147
g18755 nand P3_ADD_531_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_531_U148
g18756 nand P3_ADD_531_U125 P3_ADD_531_U62 ; P3_ADD_531_U149
g18757 nand P3_ADD_531_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_531_U150
g18758 nand P3_ADD_531_U124 P3_ADD_531_U60 ; P3_ADD_531_U151
g18759 nand P3_ADD_531_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_531_U152
g18760 nand P3_ADD_531_U123 P3_ADD_531_U58 ; P3_ADD_531_U153
g18761 nand P3_ADD_531_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_531_U154
g18762 nand P3_ADD_531_U122 P3_ADD_531_U56 ; P3_ADD_531_U155
g18763 nand P3_ADD_531_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_531_U156
g18764 nand P3_ADD_531_U121 P3_ADD_531_U54 ; P3_ADD_531_U157
g18765 nand P3_ADD_531_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_531_U158
g18766 nand P3_ADD_531_U120 P3_ADD_531_U52 ; P3_ADD_531_U159
g18767 nand P3_ADD_531_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_531_U160
g18768 nand P3_ADD_531_U119 P3_ADD_531_U50 ; P3_ADD_531_U161
g18769 nand P3_ADD_531_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_531_U162
g18770 nand P3_ADD_531_U118 P3_ADD_531_U48 ; P3_ADD_531_U163
g18771 nand P3_ADD_531_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_531_U164
g18772 nand P3_ADD_531_U117 P3_ADD_531_U46 ; P3_ADD_531_U165
g18773 nand P3_ADD_531_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_531_U166
g18774 nand P3_ADD_531_U116 P3_ADD_531_U44 ; P3_ADD_531_U167
g18775 nand P3_ADD_531_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_531_U168
g18776 nand P3_ADD_531_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_531_U169
g18777 nand P3_ADD_531_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_531_U170
g18778 nand P3_ADD_531_U115 P3_ADD_531_U42 ; P3_ADD_531_U171
g18779 nand P3_ADD_531_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_531_U172
g18780 nand P3_ADD_531_U114 P3_ADD_531_U40 ; P3_ADD_531_U173
g18781 nand P3_ADD_531_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_531_U174
g18782 nand P3_ADD_531_U113 P3_ADD_531_U38 ; P3_ADD_531_U175
g18783 nand P3_ADD_531_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_531_U176
g18784 nand P3_ADD_531_U112 P3_ADD_531_U36 ; P3_ADD_531_U177
g18785 nand P3_ADD_531_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_531_U178
g18786 nand P3_ADD_531_U111 P3_ADD_531_U34 ; P3_ADD_531_U179
g18787 nand P3_ADD_531_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_531_U180
g18788 nand P3_ADD_531_U110 P3_ADD_531_U32 ; P3_ADD_531_U181
g18789 nand P3_ADD_531_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_531_U182
g18790 nand P3_ADD_531_U109 P3_ADD_531_U30 ; P3_ADD_531_U183
g18791 nand P3_ADD_531_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_531_U184
g18792 nand P3_ADD_531_U108 P3_ADD_531_U28 ; P3_ADD_531_U185
g18793 nand P3_ADD_531_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_531_U186
g18794 nand P3_ADD_531_U107 P3_ADD_531_U26 ; P3_ADD_531_U187
g18795 nand P3_ADD_531_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_531_U188
g18796 nand P3_ADD_531_U106 P3_ADD_531_U24 ; P3_ADD_531_U189
g18797 and P3_SUB_320_U126 P3_SUB_320_U28 ; P3_SUB_320_U6
g18798 and P3_SUB_320_U124 P3_SUB_320_U29 ; P3_SUB_320_U7
g18799 and P3_SUB_320_U122 P3_SUB_320_U30 ; P3_SUB_320_U8
g18800 and P3_SUB_320_U120 P3_SUB_320_U31 ; P3_SUB_320_U9
g18801 and P3_SUB_320_U118 P3_SUB_320_U32 ; P3_SUB_320_U10
g18802 and P3_SUB_320_U116 P3_SUB_320_U33 ; P3_SUB_320_U11
g18803 and P3_SUB_320_U114 P3_SUB_320_U34 ; P3_SUB_320_U12
g18804 and P3_SUB_320_U112 P3_SUB_320_U35 ; P3_SUB_320_U13
g18805 and P3_SUB_320_U110 P3_SUB_320_U36 ; P3_SUB_320_U14
g18806 and P3_SUB_320_U108 P3_SUB_320_U37 ; P3_SUB_320_U15
g18807 and P3_SUB_320_U106 P3_SUB_320_U38 ; P3_SUB_320_U16
g18808 and P3_SUB_320_U105 P3_SUB_320_U21 ; P3_SUB_320_U17
g18809 and P3_SUB_320_U92 P3_SUB_320_U22 ; P3_SUB_320_U18
g18810 and P3_SUB_320_U90 P3_SUB_320_U23 ; P3_SUB_320_U19
g18811 and P3_SUB_320_U88 P3_SUB_320_U24 ; P3_SUB_320_U20
g18812 or P3_ADD_318_U4 P3_ADD_318_U71 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_320_U21
g18813 nand P3_SUB_320_U27 P3_SUB_320_U58 P3_SUB_320_U83 ; P3_SUB_320_U22
g18814 nand P3_SUB_320_U26 P3_SUB_320_U56 P3_SUB_320_U84 ; P3_SUB_320_U23
g18815 nand P3_SUB_320_U25 P3_SUB_320_U54 P3_SUB_320_U85 ; P3_SUB_320_U24
g18816 not P3_ADD_318_U63 ; P3_SUB_320_U25
g18817 not P3_ADD_318_U65 ; P3_SUB_320_U26
g18818 not P3_ADD_318_U67 ; P3_SUB_320_U27
g18819 nand P3_SUB_320_U52 P3_SUB_320_U49 P3_SUB_320_U86 ; P3_SUB_320_U28
g18820 nand P3_SUB_320_U48 P3_SUB_320_U81 P3_SUB_320_U93 ; P3_SUB_320_U29
g18821 nand P3_SUB_320_U47 P3_SUB_320_U79 P3_SUB_320_U94 ; P3_SUB_320_U30
g18822 nand P3_SUB_320_U46 P3_SUB_320_U77 P3_SUB_320_U95 ; P3_SUB_320_U31
g18823 nand P3_SUB_320_U45 P3_SUB_320_U75 P3_SUB_320_U96 ; P3_SUB_320_U32
g18824 nand P3_SUB_320_U44 P3_SUB_320_U73 P3_SUB_320_U97 ; P3_SUB_320_U33
g18825 nand P3_SUB_320_U43 P3_SUB_320_U69 P3_SUB_320_U98 ; P3_SUB_320_U34
g18826 nand P3_SUB_320_U42 P3_SUB_320_U67 P3_SUB_320_U99 ; P3_SUB_320_U35
g18827 nand P3_SUB_320_U41 P3_SUB_320_U65 P3_SUB_320_U100 ; P3_SUB_320_U36
g18828 nand P3_SUB_320_U40 P3_SUB_320_U63 P3_SUB_320_U101 ; P3_SUB_320_U37
g18829 nand P3_SUB_320_U102 P3_SUB_320_U39 ; P3_SUB_320_U38
g18830 not P3_ADD_318_U72 ; P3_SUB_320_U39
g18831 not P3_ADD_318_U73 ; P3_SUB_320_U40
g18832 not P3_ADD_318_U75 ; P3_SUB_320_U41
g18833 not P3_ADD_318_U77 ; P3_SUB_320_U42
g18834 not P3_ADD_318_U79 ; P3_SUB_320_U43
g18835 not P3_ADD_318_U81 ; P3_SUB_320_U44
g18836 not P3_ADD_318_U83 ; P3_SUB_320_U45
g18837 not P3_ADD_318_U85 ; P3_SUB_320_U46
g18838 not P3_ADD_318_U87 ; P3_SUB_320_U47
g18839 not P3_ADD_318_U89 ; P3_SUB_320_U48
g18840 not P3_ADD_318_U91 ; P3_SUB_320_U49
g18841 nand P3_SUB_320_U149 P3_SUB_320_U148 ; P3_SUB_320_U50
g18842 nand P3_SUB_320_U137 P3_SUB_320_U136 ; P3_SUB_320_U51
g18843 not P3_ADD_318_U62 ; P3_SUB_320_U52
g18844 and P3_SUB_320_U129 P3_SUB_320_U128 ; P3_SUB_320_U53
g18845 not P3_ADD_318_U64 ; P3_SUB_320_U54
g18846 and P3_SUB_320_U131 P3_SUB_320_U130 ; P3_SUB_320_U55
g18847 not P3_ADD_318_U66 ; P3_SUB_320_U56
g18848 and P3_SUB_320_U133 P3_SUB_320_U132 ; P3_SUB_320_U57
g18849 not P3_ADD_318_U68 ; P3_SUB_320_U58
g18850 and P3_SUB_320_U135 P3_SUB_320_U134 ; P3_SUB_320_U59
g18851 not P3_ADD_318_U69 ; P3_SUB_320_U60
g18852 not P3_ADD_318_U70 ; P3_SUB_320_U61
g18853 and P3_SUB_320_U139 P3_SUB_320_U138 ; P3_SUB_320_U62
g18854 not P3_ADD_318_U74 ; P3_SUB_320_U63
g18855 and P3_SUB_320_U141 P3_SUB_320_U140 ; P3_SUB_320_U64
g18856 not P3_ADD_318_U76 ; P3_SUB_320_U65
g18857 and P3_SUB_320_U143 P3_SUB_320_U142 ; P3_SUB_320_U66
g18858 not P3_ADD_318_U78 ; P3_SUB_320_U67
g18859 and P3_SUB_320_U145 P3_SUB_320_U144 ; P3_SUB_320_U68
g18860 not P3_ADD_318_U80 ; P3_SUB_320_U69
g18861 and P3_SUB_320_U147 P3_SUB_320_U146 ; P3_SUB_320_U70
g18862 not P3_ADD_318_U4 ; P3_SUB_320_U71
g18863 not P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_320_U72
g18864 not P3_ADD_318_U82 ; P3_SUB_320_U73
g18865 and P3_SUB_320_U151 P3_SUB_320_U150 ; P3_SUB_320_U74
g18866 not P3_ADD_318_U84 ; P3_SUB_320_U75
g18867 and P3_SUB_320_U153 P3_SUB_320_U152 ; P3_SUB_320_U76
g18868 not P3_ADD_318_U86 ; P3_SUB_320_U77
g18869 and P3_SUB_320_U155 P3_SUB_320_U154 ; P3_SUB_320_U78
g18870 not P3_ADD_318_U88 ; P3_SUB_320_U79
g18871 and P3_SUB_320_U157 P3_SUB_320_U156 ; P3_SUB_320_U80
g18872 not P3_ADD_318_U90 ; P3_SUB_320_U81
g18873 and P3_SUB_320_U159 P3_SUB_320_U158 ; P3_SUB_320_U82
g18874 not P3_SUB_320_U21 ; P3_SUB_320_U83
g18875 not P3_SUB_320_U22 ; P3_SUB_320_U84
g18876 not P3_SUB_320_U23 ; P3_SUB_320_U85
g18877 not P3_SUB_320_U24 ; P3_SUB_320_U86
g18878 nand P3_SUB_320_U85 P3_SUB_320_U54 ; P3_SUB_320_U87
g18879 nand P3_ADD_318_U63 P3_SUB_320_U87 ; P3_SUB_320_U88
g18880 nand P3_SUB_320_U84 P3_SUB_320_U56 ; P3_SUB_320_U89
g18881 nand P3_ADD_318_U65 P3_SUB_320_U89 ; P3_SUB_320_U90
g18882 nand P3_SUB_320_U83 P3_SUB_320_U58 ; P3_SUB_320_U91
g18883 nand P3_ADD_318_U67 P3_SUB_320_U91 ; P3_SUB_320_U92
g18884 not P3_SUB_320_U28 ; P3_SUB_320_U93
g18885 not P3_SUB_320_U29 ; P3_SUB_320_U94
g18886 not P3_SUB_320_U30 ; P3_SUB_320_U95
g18887 not P3_SUB_320_U31 ; P3_SUB_320_U96
g18888 not P3_SUB_320_U32 ; P3_SUB_320_U97
g18889 not P3_SUB_320_U33 ; P3_SUB_320_U98
g18890 not P3_SUB_320_U34 ; P3_SUB_320_U99
g18891 not P3_SUB_320_U35 ; P3_SUB_320_U100
g18892 not P3_SUB_320_U36 ; P3_SUB_320_U101
g18893 not P3_SUB_320_U37 ; P3_SUB_320_U102
g18894 not P3_SUB_320_U38 ; P3_SUB_320_U103
g18895 or P3_ADD_318_U4 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_320_U104
g18896 nand P3_ADD_318_U71 P3_SUB_320_U104 ; P3_SUB_320_U105
g18897 nand P3_ADD_318_U72 P3_SUB_320_U37 ; P3_SUB_320_U106
g18898 nand P3_SUB_320_U101 P3_SUB_320_U63 ; P3_SUB_320_U107
g18899 nand P3_ADD_318_U73 P3_SUB_320_U107 ; P3_SUB_320_U108
g18900 nand P3_SUB_320_U100 P3_SUB_320_U65 ; P3_SUB_320_U109
g18901 nand P3_ADD_318_U75 P3_SUB_320_U109 ; P3_SUB_320_U110
g18902 nand P3_SUB_320_U99 P3_SUB_320_U67 ; P3_SUB_320_U111
g18903 nand P3_ADD_318_U77 P3_SUB_320_U111 ; P3_SUB_320_U112
g18904 nand P3_SUB_320_U98 P3_SUB_320_U69 ; P3_SUB_320_U113
g18905 nand P3_ADD_318_U79 P3_SUB_320_U113 ; P3_SUB_320_U114
g18906 nand P3_SUB_320_U97 P3_SUB_320_U73 ; P3_SUB_320_U115
g18907 nand P3_ADD_318_U81 P3_SUB_320_U115 ; P3_SUB_320_U116
g18908 nand P3_SUB_320_U96 P3_SUB_320_U75 ; P3_SUB_320_U117
g18909 nand P3_ADD_318_U83 P3_SUB_320_U117 ; P3_SUB_320_U118
g18910 nand P3_SUB_320_U95 P3_SUB_320_U77 ; P3_SUB_320_U119
g18911 nand P3_ADD_318_U85 P3_SUB_320_U119 ; P3_SUB_320_U120
g18912 nand P3_SUB_320_U94 P3_SUB_320_U79 ; P3_SUB_320_U121
g18913 nand P3_ADD_318_U87 P3_SUB_320_U121 ; P3_SUB_320_U122
g18914 nand P3_SUB_320_U93 P3_SUB_320_U81 ; P3_SUB_320_U123
g18915 nand P3_ADD_318_U89 P3_SUB_320_U123 ; P3_SUB_320_U124
g18916 nand P3_SUB_320_U86 P3_SUB_320_U52 ; P3_SUB_320_U125
g18917 nand P3_ADD_318_U91 P3_SUB_320_U125 ; P3_SUB_320_U126
g18918 nand P3_SUB_320_U103 P3_SUB_320_U61 ; P3_SUB_320_U127
g18919 nand P3_ADD_318_U62 P3_SUB_320_U24 ; P3_SUB_320_U128
g18920 nand P3_SUB_320_U86 P3_SUB_320_U52 ; P3_SUB_320_U129
g18921 nand P3_ADD_318_U64 P3_SUB_320_U23 ; P3_SUB_320_U130
g18922 nand P3_SUB_320_U85 P3_SUB_320_U54 ; P3_SUB_320_U131
g18923 nand P3_ADD_318_U66 P3_SUB_320_U22 ; P3_SUB_320_U132
g18924 nand P3_SUB_320_U84 P3_SUB_320_U56 ; P3_SUB_320_U133
g18925 nand P3_ADD_318_U68 P3_SUB_320_U21 ; P3_SUB_320_U134
g18926 nand P3_SUB_320_U83 P3_SUB_320_U58 ; P3_SUB_320_U135
g18927 nand P3_SUB_320_U127 P3_SUB_320_U60 ; P3_SUB_320_U136
g18928 nand P3_SUB_320_U103 P3_SUB_320_U61 P3_ADD_318_U69 ; P3_SUB_320_U137
g18929 nand P3_ADD_318_U70 P3_SUB_320_U38 ; P3_SUB_320_U138
g18930 nand P3_SUB_320_U103 P3_SUB_320_U61 ; P3_SUB_320_U139
g18931 nand P3_ADD_318_U74 P3_SUB_320_U36 ; P3_SUB_320_U140
g18932 nand P3_SUB_320_U101 P3_SUB_320_U63 ; P3_SUB_320_U141
g18933 nand P3_ADD_318_U76 P3_SUB_320_U35 ; P3_SUB_320_U142
g18934 nand P3_SUB_320_U100 P3_SUB_320_U65 ; P3_SUB_320_U143
g18935 nand P3_ADD_318_U78 P3_SUB_320_U34 ; P3_SUB_320_U144
g18936 nand P3_SUB_320_U99 P3_SUB_320_U67 ; P3_SUB_320_U145
g18937 nand P3_ADD_318_U80 P3_SUB_320_U33 ; P3_SUB_320_U146
g18938 nand P3_SUB_320_U98 P3_SUB_320_U69 ; P3_SUB_320_U147
g18939 nand P3_ADD_318_U4 P3_SUB_320_U72 ; P3_SUB_320_U148
g18940 nand P3_SUB_320_U71 P3_PHYADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_320_U149
g18941 nand P3_ADD_318_U82 P3_SUB_320_U32 ; P3_SUB_320_U150
g18942 nand P3_SUB_320_U97 P3_SUB_320_U73 ; P3_SUB_320_U151
g18943 nand P3_ADD_318_U84 P3_SUB_320_U31 ; P3_SUB_320_U152
g18944 nand P3_SUB_320_U96 P3_SUB_320_U75 ; P3_SUB_320_U153
g18945 nand P3_ADD_318_U86 P3_SUB_320_U30 ; P3_SUB_320_U154
g18946 nand P3_SUB_320_U95 P3_SUB_320_U77 ; P3_SUB_320_U155
g18947 nand P3_ADD_318_U88 P3_SUB_320_U29 ; P3_SUB_320_U156
g18948 nand P3_SUB_320_U94 P3_SUB_320_U79 ; P3_SUB_320_U157
g18949 nand P3_ADD_318_U90 P3_SUB_320_U28 ; P3_SUB_320_U158
g18950 nand P3_SUB_320_U93 P3_SUB_320_U81 ; P3_SUB_320_U159
g18951 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_ADD_505_U5
g18952 and P3_ADD_505_U20 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_505_U6
g18953 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_505_U7
g18954 nand P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_ADD_505_U8
g18955 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_505_U9
g18956 nand P3_ADD_505_U18 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_505_U10
g18957 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_505_U11
g18958 nand P3_ADD_505_U19 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_505_U12
g18959 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_505_U13
g18960 nand P3_ADD_505_U22 P3_ADD_505_U21 ; P3_ADD_505_U14
g18961 nand P3_ADD_505_U24 P3_ADD_505_U23 ; P3_ADD_505_U15
g18962 nand P3_ADD_505_U26 P3_ADD_505_U25 ; P3_ADD_505_U16
g18963 nand P3_ADD_505_U28 P3_ADD_505_U27 ; P3_ADD_505_U17
g18964 not P3_ADD_505_U8 ; P3_ADD_505_U18
g18965 not P3_ADD_505_U10 ; P3_ADD_505_U19
g18966 not P3_ADD_505_U12 ; P3_ADD_505_U20
g18967 nand P3_ADD_505_U12 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_505_U21
g18968 nand P3_ADD_505_U20 P3_ADD_505_U13 ; P3_ADD_505_U22
g18969 nand P3_ADD_505_U10 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_505_U23
g18970 nand P3_ADD_505_U19 P3_ADD_505_U11 ; P3_ADD_505_U24
g18971 nand P3_ADD_505_U8 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_505_U25
g18972 nand P3_ADD_505_U18 P3_ADD_505_U9 ; P3_ADD_505_U26
g18973 nand P3_ADD_505_U5 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_505_U27
g18974 nand P3_ADD_505_U7 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_ADD_505_U28
g18975 nor P3_SUB_485_U6 P3_GTE_485_U7 ; P3_GTE_485_U6
g18976 nor P3_SUB_485_U16 P3_SUB_485_U17 P3_SUB_485_U19 P3_SUB_485_U18 ; P3_GTE_485_U7
g18977 not P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_318_U4
g18978 not P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_318_U5
g18979 nand P3_PHYADDRPOINTER_REG_1__SCAN_IN P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_318_U6
g18980 not P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_318_U7
g18981 nand P3_ADD_318_U94 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_318_U8
g18982 not P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_318_U9
g18983 nand P3_ADD_318_U95 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_318_U10
g18984 not P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_318_U11
g18985 nand P3_ADD_318_U96 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_318_U12
g18986 not P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_318_U13
g18987 nand P3_ADD_318_U97 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_318_U14
g18988 not P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_318_U15
g18989 nand P3_ADD_318_U98 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_318_U16
g18990 not P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_318_U17
g18991 not P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_318_U18
g18992 nand P3_ADD_318_U99 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_318_U19
g18993 nand P3_ADD_318_U100 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_318_U20
g18994 not P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_318_U21
g18995 nand P3_ADD_318_U101 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_318_U22
g18996 not P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_318_U23
g18997 nand P3_ADD_318_U102 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_318_U24
g18998 not P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_318_U25
g18999 nand P3_ADD_318_U103 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_318_U26
g19000 not P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_318_U27
g19001 nand P3_ADD_318_U104 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_318_U28
g19002 not P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_318_U29
g19003 nand P3_ADD_318_U105 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_318_U30
g19004 not P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_318_U31
g19005 nand P3_ADD_318_U106 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_318_U32
g19006 not P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_318_U33
g19007 nand P3_ADD_318_U107 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_318_U34
g19008 not P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_318_U35
g19009 nand P3_ADD_318_U108 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_318_U36
g19010 not P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_318_U37
g19011 nand P3_ADD_318_U109 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_318_U38
g19012 not P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_318_U39
g19013 nand P3_ADD_318_U110 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_318_U40
g19014 not P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_318_U41
g19015 nand P3_ADD_318_U111 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_318_U42
g19016 not P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_318_U43
g19017 nand P3_ADD_318_U112 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_318_U44
g19018 not P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_318_U45
g19019 nand P3_ADD_318_U113 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_318_U46
g19020 not P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_318_U47
g19021 nand P3_ADD_318_U114 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_318_U48
g19022 not P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_318_U49
g19023 nand P3_ADD_318_U115 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_318_U50
g19024 not P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_318_U51
g19025 nand P3_ADD_318_U116 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_318_U52
g19026 not P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_318_U53
g19027 nand P3_ADD_318_U117 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_318_U54
g19028 not P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_318_U55
g19029 nand P3_ADD_318_U118 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_318_U56
g19030 not P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_318_U57
g19031 nand P3_ADD_318_U119 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_318_U58
g19032 not P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_318_U59
g19033 nand P3_ADD_318_U120 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_318_U60
g19034 not P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_318_U61
g19035 nand P3_ADD_318_U124 P3_ADD_318_U123 ; P3_ADD_318_U62
g19036 nand P3_ADD_318_U126 P3_ADD_318_U125 ; P3_ADD_318_U63
g19037 nand P3_ADD_318_U128 P3_ADD_318_U127 ; P3_ADD_318_U64
g19038 nand P3_ADD_318_U130 P3_ADD_318_U129 ; P3_ADD_318_U65
g19039 nand P3_ADD_318_U132 P3_ADD_318_U131 ; P3_ADD_318_U66
g19040 nand P3_ADD_318_U134 P3_ADD_318_U133 ; P3_ADD_318_U67
g19041 nand P3_ADD_318_U136 P3_ADD_318_U135 ; P3_ADD_318_U68
g19042 nand P3_ADD_318_U138 P3_ADD_318_U137 ; P3_ADD_318_U69
g19043 nand P3_ADD_318_U140 P3_ADD_318_U139 ; P3_ADD_318_U70
g19044 nand P3_ADD_318_U142 P3_ADD_318_U141 ; P3_ADD_318_U71
g19045 nand P3_ADD_318_U144 P3_ADD_318_U143 ; P3_ADD_318_U72
g19046 nand P3_ADD_318_U146 P3_ADD_318_U145 ; P3_ADD_318_U73
g19047 nand P3_ADD_318_U148 P3_ADD_318_U147 ; P3_ADD_318_U74
g19048 nand P3_ADD_318_U150 P3_ADD_318_U149 ; P3_ADD_318_U75
g19049 nand P3_ADD_318_U152 P3_ADD_318_U151 ; P3_ADD_318_U76
g19050 nand P3_ADD_318_U154 P3_ADD_318_U153 ; P3_ADD_318_U77
g19051 nand P3_ADD_318_U156 P3_ADD_318_U155 ; P3_ADD_318_U78
g19052 nand P3_ADD_318_U158 P3_ADD_318_U157 ; P3_ADD_318_U79
g19053 nand P3_ADD_318_U160 P3_ADD_318_U159 ; P3_ADD_318_U80
g19054 nand P3_ADD_318_U162 P3_ADD_318_U161 ; P3_ADD_318_U81
g19055 nand P3_ADD_318_U164 P3_ADD_318_U163 ; P3_ADD_318_U82
g19056 nand P3_ADD_318_U166 P3_ADD_318_U165 ; P3_ADD_318_U83
g19057 nand P3_ADD_318_U168 P3_ADD_318_U167 ; P3_ADD_318_U84
g19058 nand P3_ADD_318_U170 P3_ADD_318_U169 ; P3_ADD_318_U85
g19059 nand P3_ADD_318_U172 P3_ADD_318_U171 ; P3_ADD_318_U86
g19060 nand P3_ADD_318_U174 P3_ADD_318_U173 ; P3_ADD_318_U87
g19061 nand P3_ADD_318_U176 P3_ADD_318_U175 ; P3_ADD_318_U88
g19062 nand P3_ADD_318_U178 P3_ADD_318_U177 ; P3_ADD_318_U89
g19063 nand P3_ADD_318_U180 P3_ADD_318_U179 ; P3_ADD_318_U90
g19064 nand P3_ADD_318_U182 P3_ADD_318_U181 ; P3_ADD_318_U91
g19065 not P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_318_U92
g19066 nand P3_ADD_318_U121 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_318_U93
g19067 not P3_ADD_318_U6 ; P3_ADD_318_U94
g19068 not P3_ADD_318_U8 ; P3_ADD_318_U95
g19069 not P3_ADD_318_U10 ; P3_ADD_318_U96
g19070 not P3_ADD_318_U12 ; P3_ADD_318_U97
g19071 not P3_ADD_318_U14 ; P3_ADD_318_U98
g19072 not P3_ADD_318_U16 ; P3_ADD_318_U99
g19073 not P3_ADD_318_U19 ; P3_ADD_318_U100
g19074 not P3_ADD_318_U20 ; P3_ADD_318_U101
g19075 not P3_ADD_318_U22 ; P3_ADD_318_U102
g19076 not P3_ADD_318_U24 ; P3_ADD_318_U103
g19077 not P3_ADD_318_U26 ; P3_ADD_318_U104
g19078 not P3_ADD_318_U28 ; P3_ADD_318_U105
g19079 not P3_ADD_318_U30 ; P3_ADD_318_U106
g19080 not P3_ADD_318_U32 ; P3_ADD_318_U107
g19081 not P3_ADD_318_U34 ; P3_ADD_318_U108
g19082 not P3_ADD_318_U36 ; P3_ADD_318_U109
g19083 not P3_ADD_318_U38 ; P3_ADD_318_U110
g19084 not P3_ADD_318_U40 ; P3_ADD_318_U111
g19085 not P3_ADD_318_U42 ; P3_ADD_318_U112
g19086 not P3_ADD_318_U44 ; P3_ADD_318_U113
g19087 not P3_ADD_318_U46 ; P3_ADD_318_U114
g19088 not P3_ADD_318_U48 ; P3_ADD_318_U115
g19089 not P3_ADD_318_U50 ; P3_ADD_318_U116
g19090 not P3_ADD_318_U52 ; P3_ADD_318_U117
g19091 not P3_ADD_318_U54 ; P3_ADD_318_U118
g19092 not P3_ADD_318_U56 ; P3_ADD_318_U119
g19093 not P3_ADD_318_U58 ; P3_ADD_318_U120
g19094 not P3_ADD_318_U60 ; P3_ADD_318_U121
g19095 not P3_ADD_318_U93 ; P3_ADD_318_U122
g19096 nand P3_ADD_318_U19 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_318_U123
g19097 nand P3_ADD_318_U100 P3_ADD_318_U18 ; P3_ADD_318_U124
g19098 nand P3_ADD_318_U16 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_318_U125
g19099 nand P3_ADD_318_U99 P3_ADD_318_U17 ; P3_ADD_318_U126
g19100 nand P3_ADD_318_U14 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_318_U127
g19101 nand P3_ADD_318_U98 P3_ADD_318_U15 ; P3_ADD_318_U128
g19102 nand P3_ADD_318_U12 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_318_U129
g19103 nand P3_ADD_318_U97 P3_ADD_318_U13 ; P3_ADD_318_U130
g19104 nand P3_ADD_318_U10 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_318_U131
g19105 nand P3_ADD_318_U96 P3_ADD_318_U11 ; P3_ADD_318_U132
g19106 nand P3_ADD_318_U8 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_318_U133
g19107 nand P3_ADD_318_U95 P3_ADD_318_U9 ; P3_ADD_318_U134
g19108 nand P3_ADD_318_U6 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_318_U135
g19109 nand P3_ADD_318_U94 P3_ADD_318_U7 ; P3_ADD_318_U136
g19110 nand P3_ADD_318_U93 P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_318_U137
g19111 nand P3_ADD_318_U122 P3_ADD_318_U92 ; P3_ADD_318_U138
g19112 nand P3_ADD_318_U60 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_318_U139
g19113 nand P3_ADD_318_U121 P3_ADD_318_U61 ; P3_ADD_318_U140
g19114 nand P3_ADD_318_U4 P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_318_U141
g19115 nand P3_ADD_318_U5 P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_318_U142
g19116 nand P3_ADD_318_U58 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_318_U143
g19117 nand P3_ADD_318_U120 P3_ADD_318_U59 ; P3_ADD_318_U144
g19118 nand P3_ADD_318_U56 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_318_U145
g19119 nand P3_ADD_318_U119 P3_ADD_318_U57 ; P3_ADD_318_U146
g19120 nand P3_ADD_318_U54 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_318_U147
g19121 nand P3_ADD_318_U118 P3_ADD_318_U55 ; P3_ADD_318_U148
g19122 nand P3_ADD_318_U52 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_318_U149
g19123 nand P3_ADD_318_U117 P3_ADD_318_U53 ; P3_ADD_318_U150
g19124 nand P3_ADD_318_U50 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_318_U151
g19125 nand P3_ADD_318_U116 P3_ADD_318_U51 ; P3_ADD_318_U152
g19126 nand P3_ADD_318_U48 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_318_U153
g19127 nand P3_ADD_318_U115 P3_ADD_318_U49 ; P3_ADD_318_U154
g19128 nand P3_ADD_318_U46 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_318_U155
g19129 nand P3_ADD_318_U114 P3_ADD_318_U47 ; P3_ADD_318_U156
g19130 nand P3_ADD_318_U44 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_318_U157
g19131 nand P3_ADD_318_U113 P3_ADD_318_U45 ; P3_ADD_318_U158
g19132 nand P3_ADD_318_U42 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_318_U159
g19133 nand P3_ADD_318_U112 P3_ADD_318_U43 ; P3_ADD_318_U160
g19134 nand P3_ADD_318_U40 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_318_U161
g19135 nand P3_ADD_318_U111 P3_ADD_318_U41 ; P3_ADD_318_U162
g19136 nand P3_ADD_318_U38 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_318_U163
g19137 nand P3_ADD_318_U110 P3_ADD_318_U39 ; P3_ADD_318_U164
g19138 nand P3_ADD_318_U36 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_318_U165
g19139 nand P3_ADD_318_U109 P3_ADD_318_U37 ; P3_ADD_318_U166
g19140 nand P3_ADD_318_U34 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_318_U167
g19141 nand P3_ADD_318_U108 P3_ADD_318_U35 ; P3_ADD_318_U168
g19142 nand P3_ADD_318_U32 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_318_U169
g19143 nand P3_ADD_318_U107 P3_ADD_318_U33 ; P3_ADD_318_U170
g19144 nand P3_ADD_318_U30 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_318_U171
g19145 nand P3_ADD_318_U106 P3_ADD_318_U31 ; P3_ADD_318_U172
g19146 nand P3_ADD_318_U28 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_318_U173
g19147 nand P3_ADD_318_U105 P3_ADD_318_U29 ; P3_ADD_318_U174
g19148 nand P3_ADD_318_U26 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_318_U175
g19149 nand P3_ADD_318_U104 P3_ADD_318_U27 ; P3_ADD_318_U176
g19150 nand P3_ADD_318_U24 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_318_U177
g19151 nand P3_ADD_318_U103 P3_ADD_318_U25 ; P3_ADD_318_U178
g19152 nand P3_ADD_318_U22 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_318_U179
g19153 nand P3_ADD_318_U102 P3_ADD_318_U23 ; P3_ADD_318_U180
g19154 nand P3_ADD_318_U20 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_318_U181
g19155 nand P3_ADD_318_U101 P3_ADD_318_U21 ; P3_ADD_318_U182
g19156 nand P3_SUB_370_U45 P3_SUB_370_U44 ; P3_SUB_370_U6
g19157 nand P3_SUB_370_U9 P3_SUB_370_U46 ; P3_SUB_370_U7
g19158 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_370_U8
g19159 nand P3_SUB_370_U18 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_370_U9
g19160 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_370_U10
g19161 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_370_U11
g19162 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_370_U12
g19163 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_370_U13
g19164 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_370_U14
g19165 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_370_U15
g19166 nand P3_SUB_370_U41 P3_SUB_370_U40 ; P3_SUB_370_U16
g19167 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_370_U17
g19168 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_370_U18
g19169 nand P3_SUB_370_U51 P3_SUB_370_U50 ; P3_SUB_370_U19
g19170 nand P3_SUB_370_U56 P3_SUB_370_U55 ; P3_SUB_370_U20
g19171 nand P3_SUB_370_U61 P3_SUB_370_U60 ; P3_SUB_370_U21
g19172 nand P3_SUB_370_U66 P3_SUB_370_U65 ; P3_SUB_370_U22
g19173 nand P3_SUB_370_U48 P3_SUB_370_U47 ; P3_SUB_370_U23
g19174 nand P3_SUB_370_U53 P3_SUB_370_U52 ; P3_SUB_370_U24
g19175 nand P3_SUB_370_U58 P3_SUB_370_U57 ; P3_SUB_370_U25
g19176 nand P3_SUB_370_U63 P3_SUB_370_U62 ; P3_SUB_370_U26
g19177 nand P3_SUB_370_U37 P3_SUB_370_U36 ; P3_SUB_370_U27
g19178 nand P3_SUB_370_U33 P3_SUB_370_U32 ; P3_SUB_370_U28
g19179 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_370_U29
g19180 not P3_SUB_370_U9 ; P3_SUB_370_U30
g19181 nand P3_SUB_370_U30 P3_SUB_370_U10 ; P3_SUB_370_U31
g19182 nand P3_SUB_370_U31 P3_SUB_370_U29 ; P3_SUB_370_U32
g19183 nand P3_SUB_370_U9 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_370_U33
g19184 not P3_SUB_370_U28 ; P3_SUB_370_U34
g19185 nand P3_SUB_370_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_370_U35
g19186 nand P3_SUB_370_U35 P3_SUB_370_U28 ; P3_SUB_370_U36
g19187 nand P3_SUB_370_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_370_U37
g19188 not P3_SUB_370_U27 ; P3_SUB_370_U38
g19189 nand P3_SUB_370_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_370_U39
g19190 nand P3_SUB_370_U39 P3_SUB_370_U27 ; P3_SUB_370_U40
g19191 nand P3_SUB_370_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_370_U41
g19192 not P3_SUB_370_U16 ; P3_SUB_370_U42
g19193 nand P3_SUB_370_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_370_U43
g19194 nand P3_SUB_370_U42 P3_SUB_370_U43 ; P3_SUB_370_U44
g19195 nand P3_SUB_370_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_370_U45
g19196 nand P3_SUB_370_U8 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_370_U46
g19197 nand P3_SUB_370_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_370_U47
g19198 nand P3_SUB_370_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_370_U48
g19199 not P3_SUB_370_U23 ; P3_SUB_370_U49
g19200 nand P3_SUB_370_U49 P3_SUB_370_U42 ; P3_SUB_370_U50
g19201 nand P3_SUB_370_U23 P3_SUB_370_U16 ; P3_SUB_370_U51
g19202 nand P3_SUB_370_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_370_U52
g19203 nand P3_SUB_370_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_370_U53
g19204 not P3_SUB_370_U24 ; P3_SUB_370_U54
g19205 nand P3_SUB_370_U38 P3_SUB_370_U54 ; P3_SUB_370_U55
g19206 nand P3_SUB_370_U24 P3_SUB_370_U27 ; P3_SUB_370_U56
g19207 nand P3_SUB_370_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_370_U57
g19208 nand P3_SUB_370_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_370_U58
g19209 not P3_SUB_370_U25 ; P3_SUB_370_U59
g19210 nand P3_SUB_370_U34 P3_SUB_370_U59 ; P3_SUB_370_U60
g19211 nand P3_SUB_370_U25 P3_SUB_370_U28 ; P3_SUB_370_U61
g19212 nand P3_SUB_370_U10 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_370_U62
g19213 nand P3_SUB_370_U29 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_370_U63
g19214 not P3_SUB_370_U26 ; P3_SUB_370_U64
g19215 nand P3_SUB_370_U64 P3_SUB_370_U30 ; P3_SUB_370_U65
g19216 nand P3_SUB_370_U26 P3_SUB_370_U9 ; P3_SUB_370_U66
g19217 not P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_315_U4
g19218 not P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_315_U5
g19219 nand P3_PHYADDRPOINTER_REG_2__SCAN_IN P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_315_U6
g19220 not P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_315_U7
g19221 nand P3_ADD_315_U91 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_315_U8
g19222 not P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_315_U9
g19223 nand P3_ADD_315_U92 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_315_U10
g19224 not P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_315_U11
g19225 nand P3_ADD_315_U93 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_315_U12
g19226 not P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_315_U13
g19227 nand P3_ADD_315_U94 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_315_U14
g19228 not P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_315_U15
g19229 not P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_315_U16
g19230 nand P3_ADD_315_U95 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_315_U17
g19231 nand P3_ADD_315_U96 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_315_U18
g19232 not P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_315_U19
g19233 nand P3_ADD_315_U97 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_315_U20
g19234 not P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_315_U21
g19235 nand P3_ADD_315_U98 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_315_U22
g19236 not P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_315_U23
g19237 nand P3_ADD_315_U99 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_315_U24
g19238 not P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_315_U25
g19239 nand P3_ADD_315_U100 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_315_U26
g19240 not P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_315_U27
g19241 nand P3_ADD_315_U101 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_315_U28
g19242 not P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_315_U29
g19243 nand P3_ADD_315_U102 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_315_U30
g19244 not P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_315_U31
g19245 nand P3_ADD_315_U103 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_315_U32
g19246 not P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_315_U33
g19247 nand P3_ADD_315_U104 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_315_U34
g19248 not P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_315_U35
g19249 nand P3_ADD_315_U105 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_315_U36
g19250 not P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_315_U37
g19251 nand P3_ADD_315_U106 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_315_U38
g19252 not P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_315_U39
g19253 nand P3_ADD_315_U107 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_315_U40
g19254 not P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_315_U41
g19255 nand P3_ADD_315_U108 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_315_U42
g19256 not P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_315_U43
g19257 nand P3_ADD_315_U109 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_315_U44
g19258 not P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_315_U45
g19259 nand P3_ADD_315_U110 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_315_U46
g19260 not P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_315_U47
g19261 nand P3_ADD_315_U111 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_315_U48
g19262 not P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_315_U49
g19263 nand P3_ADD_315_U112 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_315_U50
g19264 not P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_315_U51
g19265 nand P3_ADD_315_U113 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_315_U52
g19266 not P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_315_U53
g19267 nand P3_ADD_315_U114 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_315_U54
g19268 not P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_315_U55
g19269 nand P3_ADD_315_U115 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_315_U56
g19270 not P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_315_U57
g19271 nand P3_ADD_315_U116 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_315_U58
g19272 not P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_315_U59
g19273 nand P3_ADD_315_U120 P3_ADD_315_U119 ; P3_ADD_315_U60
g19274 nand P3_ADD_315_U122 P3_ADD_315_U121 ; P3_ADD_315_U61
g19275 nand P3_ADD_315_U124 P3_ADD_315_U123 ; P3_ADD_315_U62
g19276 nand P3_ADD_315_U126 P3_ADD_315_U125 ; P3_ADD_315_U63
g19277 nand P3_ADD_315_U128 P3_ADD_315_U127 ; P3_ADD_315_U64
g19278 nand P3_ADD_315_U130 P3_ADD_315_U129 ; P3_ADD_315_U65
g19279 nand P3_ADD_315_U132 P3_ADD_315_U131 ; P3_ADD_315_U66
g19280 nand P3_ADD_315_U134 P3_ADD_315_U133 ; P3_ADD_315_U67
g19281 nand P3_ADD_315_U136 P3_ADD_315_U135 ; P3_ADD_315_U68
g19282 nand P3_ADD_315_U138 P3_ADD_315_U137 ; P3_ADD_315_U69
g19283 nand P3_ADD_315_U140 P3_ADD_315_U139 ; P3_ADD_315_U70
g19284 nand P3_ADD_315_U142 P3_ADD_315_U141 ; P3_ADD_315_U71
g19285 nand P3_ADD_315_U144 P3_ADD_315_U143 ; P3_ADD_315_U72
g19286 nand P3_ADD_315_U146 P3_ADD_315_U145 ; P3_ADD_315_U73
g19287 nand P3_ADD_315_U148 P3_ADD_315_U147 ; P3_ADD_315_U74
g19288 nand P3_ADD_315_U150 P3_ADD_315_U149 ; P3_ADD_315_U75
g19289 nand P3_ADD_315_U152 P3_ADD_315_U151 ; P3_ADD_315_U76
g19290 nand P3_ADD_315_U154 P3_ADD_315_U153 ; P3_ADD_315_U77
g19291 nand P3_ADD_315_U156 P3_ADD_315_U155 ; P3_ADD_315_U78
g19292 nand P3_ADD_315_U158 P3_ADD_315_U157 ; P3_ADD_315_U79
g19293 nand P3_ADD_315_U160 P3_ADD_315_U159 ; P3_ADD_315_U80
g19294 nand P3_ADD_315_U162 P3_ADD_315_U161 ; P3_ADD_315_U81
g19295 nand P3_ADD_315_U164 P3_ADD_315_U163 ; P3_ADD_315_U82
g19296 nand P3_ADD_315_U166 P3_ADD_315_U165 ; P3_ADD_315_U83
g19297 nand P3_ADD_315_U168 P3_ADD_315_U167 ; P3_ADD_315_U84
g19298 nand P3_ADD_315_U170 P3_ADD_315_U169 ; P3_ADD_315_U85
g19299 nand P3_ADD_315_U172 P3_ADD_315_U171 ; P3_ADD_315_U86
g19300 nand P3_ADD_315_U174 P3_ADD_315_U173 ; P3_ADD_315_U87
g19301 nand P3_ADD_315_U176 P3_ADD_315_U175 ; P3_ADD_315_U88
g19302 not P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_315_U89
g19303 nand P3_ADD_315_U117 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_315_U90
g19304 not P3_ADD_315_U6 ; P3_ADD_315_U91
g19305 not P3_ADD_315_U8 ; P3_ADD_315_U92
g19306 not P3_ADD_315_U10 ; P3_ADD_315_U93
g19307 not P3_ADD_315_U12 ; P3_ADD_315_U94
g19308 not P3_ADD_315_U14 ; P3_ADD_315_U95
g19309 not P3_ADD_315_U17 ; P3_ADD_315_U96
g19310 not P3_ADD_315_U18 ; P3_ADD_315_U97
g19311 not P3_ADD_315_U20 ; P3_ADD_315_U98
g19312 not P3_ADD_315_U22 ; P3_ADD_315_U99
g19313 not P3_ADD_315_U24 ; P3_ADD_315_U100
g19314 not P3_ADD_315_U26 ; P3_ADD_315_U101
g19315 not P3_ADD_315_U28 ; P3_ADD_315_U102
g19316 not P3_ADD_315_U30 ; P3_ADD_315_U103
g19317 not P3_ADD_315_U32 ; P3_ADD_315_U104
g19318 not P3_ADD_315_U34 ; P3_ADD_315_U105
g19319 not P3_ADD_315_U36 ; P3_ADD_315_U106
g19320 not P3_ADD_315_U38 ; P3_ADD_315_U107
g19321 not P3_ADD_315_U40 ; P3_ADD_315_U108
g19322 not P3_ADD_315_U42 ; P3_ADD_315_U109
g19323 not P3_ADD_315_U44 ; P3_ADD_315_U110
g19324 not P3_ADD_315_U46 ; P3_ADD_315_U111
g19325 not P3_ADD_315_U48 ; P3_ADD_315_U112
g19326 not P3_ADD_315_U50 ; P3_ADD_315_U113
g19327 not P3_ADD_315_U52 ; P3_ADD_315_U114
g19328 not P3_ADD_315_U54 ; P3_ADD_315_U115
g19329 not P3_ADD_315_U56 ; P3_ADD_315_U116
g19330 not P3_ADD_315_U58 ; P3_ADD_315_U117
g19331 not P3_ADD_315_U90 ; P3_ADD_315_U118
g19332 nand P3_ADD_315_U17 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_315_U119
g19333 nand P3_ADD_315_U96 P3_ADD_315_U16 ; P3_ADD_315_U120
g19334 nand P3_ADD_315_U14 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_315_U121
g19335 nand P3_ADD_315_U95 P3_ADD_315_U15 ; P3_ADD_315_U122
g19336 nand P3_ADD_315_U12 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_315_U123
g19337 nand P3_ADD_315_U94 P3_ADD_315_U13 ; P3_ADD_315_U124
g19338 nand P3_ADD_315_U10 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_315_U125
g19339 nand P3_ADD_315_U93 P3_ADD_315_U11 ; P3_ADD_315_U126
g19340 nand P3_ADD_315_U8 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_315_U127
g19341 nand P3_ADD_315_U92 P3_ADD_315_U9 ; P3_ADD_315_U128
g19342 nand P3_ADD_315_U6 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_315_U129
g19343 nand P3_ADD_315_U91 P3_ADD_315_U7 ; P3_ADD_315_U130
g19344 nand P3_ADD_315_U4 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_315_U131
g19345 nand P3_ADD_315_U5 P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_315_U132
g19346 nand P3_ADD_315_U90 P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_315_U133
g19347 nand P3_ADD_315_U118 P3_ADD_315_U89 ; P3_ADD_315_U134
g19348 nand P3_ADD_315_U58 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_315_U135
g19349 nand P3_ADD_315_U117 P3_ADD_315_U59 ; P3_ADD_315_U136
g19350 nand P3_ADD_315_U56 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_315_U137
g19351 nand P3_ADD_315_U116 P3_ADD_315_U57 ; P3_ADD_315_U138
g19352 nand P3_ADD_315_U54 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_315_U139
g19353 nand P3_ADD_315_U115 P3_ADD_315_U55 ; P3_ADD_315_U140
g19354 nand P3_ADD_315_U52 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_315_U141
g19355 nand P3_ADD_315_U114 P3_ADD_315_U53 ; P3_ADD_315_U142
g19356 nand P3_ADD_315_U50 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_315_U143
g19357 nand P3_ADD_315_U113 P3_ADD_315_U51 ; P3_ADD_315_U144
g19358 nand P3_ADD_315_U48 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_315_U145
g19359 nand P3_ADD_315_U112 P3_ADD_315_U49 ; P3_ADD_315_U146
g19360 nand P3_ADD_315_U46 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_315_U147
g19361 nand P3_ADD_315_U111 P3_ADD_315_U47 ; P3_ADD_315_U148
g19362 nand P3_ADD_315_U44 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_315_U149
g19363 nand P3_ADD_315_U110 P3_ADD_315_U45 ; P3_ADD_315_U150
g19364 nand P3_ADD_315_U42 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_315_U151
g19365 nand P3_ADD_315_U109 P3_ADD_315_U43 ; P3_ADD_315_U152
g19366 nand P3_ADD_315_U40 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_315_U153
g19367 nand P3_ADD_315_U108 P3_ADD_315_U41 ; P3_ADD_315_U154
g19368 nand P3_ADD_315_U38 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_315_U155
g19369 nand P3_ADD_315_U107 P3_ADD_315_U39 ; P3_ADD_315_U156
g19370 nand P3_ADD_315_U36 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_315_U157
g19371 nand P3_ADD_315_U106 P3_ADD_315_U37 ; P3_ADD_315_U158
g19372 nand P3_ADD_315_U34 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_315_U159
g19373 nand P3_ADD_315_U105 P3_ADD_315_U35 ; P3_ADD_315_U160
g19374 nand P3_ADD_315_U32 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_315_U161
g19375 nand P3_ADD_315_U104 P3_ADD_315_U33 ; P3_ADD_315_U162
g19376 nand P3_ADD_315_U30 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_315_U163
g19377 nand P3_ADD_315_U103 P3_ADD_315_U31 ; P3_ADD_315_U164
g19378 nand P3_ADD_315_U28 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_315_U165
g19379 nand P3_ADD_315_U102 P3_ADD_315_U29 ; P3_ADD_315_U166
g19380 nand P3_ADD_315_U26 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_315_U167
g19381 nand P3_ADD_315_U101 P3_ADD_315_U27 ; P3_ADD_315_U168
g19382 nand P3_ADD_315_U24 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_315_U169
g19383 nand P3_ADD_315_U100 P3_ADD_315_U25 ; P3_ADD_315_U170
g19384 nand P3_ADD_315_U22 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_315_U171
g19385 nand P3_ADD_315_U99 P3_ADD_315_U23 ; P3_ADD_315_U172
g19386 nand P3_ADD_315_U20 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_315_U173
g19387 nand P3_ADD_315_U98 P3_ADD_315_U21 ; P3_ADD_315_U174
g19388 nand P3_ADD_315_U18 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_315_U175
g19389 nand P3_ADD_315_U97 P3_ADD_315_U19 ; P3_ADD_315_U176
g19390 nor P3_SUB_355_U6 P3_GTE_355_U8 ; P3_GTE_355_U6
g19391 and P3_SUB_355_U7 P3_SUB_355_U22 ; P3_GTE_355_U7
g19392 nor P3_SUB_355_U19 P3_SUB_355_U20 P3_GTE_355_U7 P3_SUB_355_U21 ; P3_GTE_355_U8
g19393 and P3_ADD_360_1242_U186 P3_ADD_360_1242_U45 ; P3_ADD_360_1242_U4
g19394 and P3_ADD_360_1242_U184 P3_ADD_360_1242_U46 ; P3_ADD_360_1242_U5
g19395 and P3_ADD_360_1242_U182 P3_ADD_360_1242_U76 ; P3_ADD_360_1242_U6
g19396 and P3_ADD_360_1242_U181 P3_ADD_360_1242_U50 ; P3_ADD_360_1242_U7
g19397 and P3_ADD_360_1242_U179 P3_ADD_360_1242_U53 ; P3_ADD_360_1242_U8
g19398 and P3_ADD_360_1242_U177 P3_ADD_360_1242_U56 ; P3_ADD_360_1242_U9
g19399 and P3_ADD_360_1242_U175 P3_ADD_360_1242_U58 ; P3_ADD_360_1242_U10
g19400 and P3_ADD_360_1242_U174 P3_ADD_360_1242_U60 ; P3_ADD_360_1242_U11
g19401 and P3_ADD_360_1242_U173 P3_ADD_360_1242_U63 ; P3_ADD_360_1242_U12
g19402 and P3_ADD_360_1242_U171 P3_ADD_360_1242_U66 ; P3_ADD_360_1242_U13
g19403 and P3_ADD_360_1242_U169 P3_ADD_360_1242_U68 ; P3_ADD_360_1242_U14
g19404 and P3_ADD_360_1242_U168 P3_ADD_360_1242_U71 ; P3_ADD_360_1242_U15
g19405 and P3_ADD_360_1242_U166 P3_ADD_360_1242_U73 ; P3_ADD_360_1242_U16
g19406 and P3_ADD_360_1242_U153 P3_ADD_360_1242_U152 ; P3_ADD_360_1242_U17
g19407 and P3_ADD_360_1242_U151 P3_ADD_360_1242_U149 ; P3_ADD_360_1242_U18
g19408 nand P3_ADD_360_1242_U248 P3_ADD_360_1242_U247 P3_ADD_360_1242_U192 ; P3_ADD_360_1242_U19
g19409 not P3_ADD_360_U19 ; P3_ADD_360_1242_U20
g19410 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_360_1242_U21
g19411 not P3_ADD_360_U20 ; P3_ADD_360_1242_U22
g19412 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_360_1242_U23
g19413 not P3_U2621 ; P3_ADD_360_1242_U24
g19414 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_360_1242_U25
g19415 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_360_1242_U26
g19416 nand P3_U2621 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_360_1242_U27
g19417 not P3_ADD_360_U4 ; P3_ADD_360_1242_U28
g19418 not P3_ADD_360_U21 ; P3_ADD_360_1242_U29
g19419 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_360_1242_U30
g19420 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_360_1242_U31
g19421 not P3_ADD_360_U18 ; P3_ADD_360_1242_U32
g19422 not P3_ADD_360_U17 ; P3_ADD_360_1242_U33
g19423 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_360_1242_U34
g19424 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_360_1242_U35
g19425 not P3_ADD_360_U16 ; P3_ADD_360_1242_U36
g19426 not P3_ADD_360_U5 ; P3_ADD_360_1242_U37
g19427 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_360_1242_U38
g19428 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_360_1242_U39
g19429 nand P3_ADD_360_1242_U131 P3_ADD_360_1242_U130 ; P3_ADD_360_1242_U40
g19430 nand P3_ADD_360_1242_U40 P3_ADD_360_1242_U133 ; P3_ADD_360_1242_U41
g19431 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_360_1242_U42
g19432 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_360_1242_U43
g19433 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_360_1242_U44
g19434 nand P3_ADD_360_1242_U97 P3_ADD_360_1242_U105 ; P3_ADD_360_1242_U45
g19435 nand P3_ADD_360_1242_U98 P3_ADD_360_1242_U119 ; P3_ADD_360_1242_U46
g19436 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_360_1242_U47
g19437 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_360_1242_U48
g19438 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_360_1242_U49
g19439 nand P3_ADD_360_1242_U154 P3_ADD_360_1242_U99 ; P3_ADD_360_1242_U50
g19440 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_360_1242_U51
g19441 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_360_1242_U52
g19442 nand P3_ADD_360_1242_U100 P3_ADD_360_1242_U156 ; P3_ADD_360_1242_U53
g19443 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_360_1242_U54
g19444 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_360_1242_U55
g19445 nand P3_ADD_360_1242_U101 P3_ADD_360_1242_U157 ; P3_ADD_360_1242_U56
g19446 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_360_1242_U57
g19447 nand P3_ADD_360_1242_U158 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_360_1242_U58
g19448 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_360_1242_U59
g19449 nand P3_ADD_360_1242_U159 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_360_1242_U60
g19450 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_360_1242_U61
g19451 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_360_1242_U62
g19452 nand P3_ADD_360_1242_U102 P3_ADD_360_1242_U160 ; P3_ADD_360_1242_U63
g19453 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_360_1242_U64
g19454 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_360_1242_U65
g19455 nand P3_ADD_360_1242_U103 P3_ADD_360_1242_U161 ; P3_ADD_360_1242_U66
g19456 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_360_1242_U67
g19457 nand P3_ADD_360_1242_U162 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_360_1242_U68
g19458 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_360_1242_U69
g19459 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_360_1242_U70
g19460 nand P3_ADD_360_1242_U104 P3_ADD_360_1242_U163 ; P3_ADD_360_1242_U71
g19461 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_360_1242_U72
g19462 nand P3_ADD_360_1242_U164 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_360_1242_U73
g19463 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_360_1242_U74
g19464 nand P3_ADD_360_U4 P3_ADD_360_1242_U124 ; P3_ADD_360_1242_U75
g19465 nand P3_ADD_360_1242_U154 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_360_1242_U76
g19466 nand P3_ADD_360_1242_U230 P3_ADD_360_1242_U229 ; P3_ADD_360_1242_U77
g19467 nand P3_ADD_360_1242_U239 P3_ADD_360_1242_U238 ; P3_ADD_360_1242_U78
g19468 nand P3_ADD_360_1242_U241 P3_ADD_360_1242_U240 ; P3_ADD_360_1242_U79
g19469 nand P3_ADD_360_1242_U243 P3_ADD_360_1242_U242 ; P3_ADD_360_1242_U80
g19470 nand P3_ADD_360_1242_U250 P3_ADD_360_1242_U249 ; P3_ADD_360_1242_U81
g19471 nand P3_ADD_360_1242_U252 P3_ADD_360_1242_U251 ; P3_ADD_360_1242_U82
g19472 nand P3_ADD_360_1242_U254 P3_ADD_360_1242_U253 ; P3_ADD_360_1242_U83
g19473 nand P3_ADD_360_1242_U256 P3_ADD_360_1242_U255 ; P3_ADD_360_1242_U84
g19474 nand P3_ADD_360_1242_U258 P3_ADD_360_1242_U257 ; P3_ADD_360_1242_U85
g19475 nand P3_ADD_360_1242_U201 P3_ADD_360_1242_U200 ; P3_ADD_360_1242_U86
g19476 nand P3_ADD_360_1242_U208 P3_ADD_360_1242_U207 ; P3_ADD_360_1242_U87
g19477 nand P3_ADD_360_1242_U215 P3_ADD_360_1242_U214 ; P3_ADD_360_1242_U88
g19478 nand P3_ADD_360_1242_U222 P3_ADD_360_1242_U221 ; P3_ADD_360_1242_U89
g19479 nand P3_ADD_360_1242_U228 P3_ADD_360_1242_U227 ; P3_ADD_360_1242_U90
g19480 nand P3_ADD_360_1242_U237 P3_ADD_360_1242_U236 ; P3_ADD_360_1242_U91
g19481 and P3_ADD_360_U20 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_360_1242_U92
g19482 and P3_ADD_360_1242_U133 P3_ADD_360_1242_U123 ; P3_ADD_360_1242_U93
g19483 and P3_ADD_360_1242_U190 P3_ADD_360_1242_U125 ; P3_ADD_360_1242_U94
g19484 and P3_ADD_360_1242_U224 P3_ADD_360_1242_U223 P3_ADD_360_1242_U135 ; P3_ADD_360_1242_U95
g19485 and P3_ADD_360_1242_U125 P3_ADD_360_1242_U123 ; P3_ADD_360_1242_U96
g19486 and P3_INSTADDRPOINTER_REG_9__SCAN_IN P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_360_1242_U97
g19487 and P3_INSTADDRPOINTER_REG_11__SCAN_IN P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_360_1242_U98
g19488 and P3_INSTADDRPOINTER_REG_13__SCAN_IN P3_INSTADDRPOINTER_REG_14__SCAN_IN P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_360_1242_U99
g19489 and P3_INSTADDRPOINTER_REG_16__SCAN_IN P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_360_1242_U100
g19490 and P3_INSTADDRPOINTER_REG_18__SCAN_IN P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_360_1242_U101
g19491 and P3_INSTADDRPOINTER_REG_22__SCAN_IN P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_360_1242_U102
g19492 and P3_INSTADDRPOINTER_REG_24__SCAN_IN P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_360_1242_U103
g19493 and P3_INSTADDRPOINTER_REG_27__SCAN_IN P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_360_1242_U104
g19494 nand P3_ADD_360_1242_U147 P3_ADD_360_1242_U146 ; P3_ADD_360_1242_U105
g19495 and P3_ADD_360_1242_U194 P3_ADD_360_1242_U193 ; P3_ADD_360_1242_U106
g19496 and P3_ADD_360_1242_U196 P3_ADD_360_1242_U195 ; P3_ADD_360_1242_U107
g19497 nand P3_ADD_360_1242_U143 P3_ADD_360_1242_U120 P3_ADD_360_1242_U189 ; P3_ADD_360_1242_U108
g19498 and P3_ADD_360_1242_U203 P3_ADD_360_1242_U202 ; P3_ADD_360_1242_U109
g19499 nand P3_ADD_360_1242_U141 P3_ADD_360_1242_U140 ; P3_ADD_360_1242_U110
g19500 and P3_ADD_360_1242_U210 P3_ADD_360_1242_U209 ; P3_ADD_360_1242_U111
g19501 nand P3_ADD_360_1242_U137 P3_ADD_360_1242_U121 P3_ADD_360_1242_U188 ; P3_ADD_360_1242_U112
g19502 and P3_ADD_360_1242_U217 P3_ADD_360_1242_U216 ; P3_ADD_360_1242_U113
g19503 nand P3_ADD_360_1242_U94 P3_ADD_360_1242_U191 ; P3_ADD_360_1242_U114
g19504 and P3_ADD_360_1242_U226 P3_ADD_360_1242_U225 ; P3_ADD_360_1242_U115
g19505 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_360_1242_U116
g19506 and P3_ADD_360_1242_U232 P3_ADD_360_1242_U231 ; P3_ADD_360_1242_U117
g19507 nand P3_ADD_360_1242_U75 P3_ADD_360_1242_U127 ; P3_ADD_360_1242_U118
g19508 not P3_ADD_360_1242_U45 ; P3_ADD_360_1242_U119
g19509 nand P3_ADD_360_1242_U110 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_360_1242_U120
g19510 nand P3_ADD_360_1242_U114 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_360_1242_U121
g19511 not P3_ADD_360_1242_U75 ; P3_ADD_360_1242_U122
g19512 or P3_ADD_360_U19 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_360_1242_U123
g19513 not P3_ADD_360_1242_U27 ; P3_ADD_360_1242_U124
g19514 nand P3_ADD_360_U19 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_360_1242_U125
g19515 nand P3_ADD_360_1242_U28 P3_ADD_360_1242_U27 ; P3_ADD_360_1242_U126
g19516 nand P3_ADD_360_1242_U126 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_360_1242_U127
g19517 not P3_ADD_360_1242_U118 ; P3_ADD_360_1242_U128
g19518 or P3_ADD_360_U21 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_360_1242_U129
g19519 nand P3_ADD_360_1242_U129 P3_ADD_360_1242_U118 ; P3_ADD_360_1242_U130
g19520 nand P3_ADD_360_U21 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_360_1242_U131
g19521 not P3_ADD_360_1242_U40 ; P3_ADD_360_1242_U132
g19522 or P3_ADD_360_U20 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_360_1242_U133
g19523 not P3_ADD_360_1242_U41 ; P3_ADD_360_1242_U134
g19524 nand P3_ADD_360_U20 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_360_1242_U135
g19525 not P3_ADD_360_1242_U114 ; P3_ADD_360_1242_U136
g19526 nand P3_ADD_360_U18 P3_ADD_360_1242_U114 ; P3_ADD_360_1242_U137
g19527 not P3_ADD_360_1242_U112 ; P3_ADD_360_1242_U138
g19528 or P3_ADD_360_U17 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_360_1242_U139
g19529 nand P3_ADD_360_1242_U139 P3_ADD_360_1242_U112 ; P3_ADD_360_1242_U140
g19530 nand P3_ADD_360_U17 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_360_1242_U141
g19531 not P3_ADD_360_1242_U110 ; P3_ADD_360_1242_U142
g19532 nand P3_ADD_360_U16 P3_ADD_360_1242_U110 ; P3_ADD_360_1242_U143
g19533 not P3_ADD_360_1242_U108 ; P3_ADD_360_1242_U144
g19534 or P3_ADD_360_U5 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_360_1242_U145
g19535 nand P3_ADD_360_1242_U145 P3_ADD_360_1242_U108 ; P3_ADD_360_1242_U146
g19536 nand P3_ADD_360_U5 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_360_1242_U147
g19537 not P3_ADD_360_1242_U105 ; P3_ADD_360_1242_U148
g19538 nand P3_ADD_360_1242_U95 P3_ADD_360_1242_U41 ; P3_ADD_360_1242_U149
g19539 nand P3_ADD_360_1242_U135 P3_ADD_360_1242_U41 ; P3_ADD_360_1242_U150
g19540 nand P3_ADD_360_1242_U96 P3_ADD_360_1242_U150 ; P3_ADD_360_1242_U151
g19541 nand P3_ADD_360_1242_U115 P3_ADD_360_1242_U132 ; P3_ADD_360_1242_U152
g19542 nand P3_ADD_360_1242_U134 P3_ADD_360_1242_U135 ; P3_ADD_360_1242_U153
g19543 not P3_ADD_360_1242_U46 ; P3_ADD_360_1242_U154
g19544 not P3_ADD_360_1242_U76 ; P3_ADD_360_1242_U155
g19545 not P3_ADD_360_1242_U50 ; P3_ADD_360_1242_U156
g19546 not P3_ADD_360_1242_U53 ; P3_ADD_360_1242_U157
g19547 not P3_ADD_360_1242_U56 ; P3_ADD_360_1242_U158
g19548 not P3_ADD_360_1242_U58 ; P3_ADD_360_1242_U159
g19549 not P3_ADD_360_1242_U60 ; P3_ADD_360_1242_U160
g19550 not P3_ADD_360_1242_U63 ; P3_ADD_360_1242_U161
g19551 not P3_ADD_360_1242_U66 ; P3_ADD_360_1242_U162
g19552 not P3_ADD_360_1242_U68 ; P3_ADD_360_1242_U163
g19553 not P3_ADD_360_1242_U71 ; P3_ADD_360_1242_U164
g19554 not P3_ADD_360_1242_U73 ; P3_ADD_360_1242_U165
g19555 nand P3_ADD_360_1242_U72 P3_ADD_360_1242_U71 ; P3_ADD_360_1242_U166
g19556 nand P3_ADD_360_1242_U163 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_360_1242_U167
g19557 nand P3_ADD_360_1242_U69 P3_ADD_360_1242_U167 ; P3_ADD_360_1242_U168
g19558 nand P3_ADD_360_1242_U67 P3_ADD_360_1242_U66 ; P3_ADD_360_1242_U169
g19559 nand P3_ADD_360_1242_U161 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_360_1242_U170
g19560 nand P3_ADD_360_1242_U64 P3_ADD_360_1242_U170 ; P3_ADD_360_1242_U171
g19561 nand P3_ADD_360_1242_U160 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_360_1242_U172
g19562 nand P3_ADD_360_1242_U61 P3_ADD_360_1242_U172 ; P3_ADD_360_1242_U173
g19563 nand P3_ADD_360_1242_U59 P3_ADD_360_1242_U58 ; P3_ADD_360_1242_U174
g19564 nand P3_ADD_360_1242_U57 P3_ADD_360_1242_U56 ; P3_ADD_360_1242_U175
g19565 nand P3_ADD_360_1242_U157 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_360_1242_U176
g19566 nand P3_ADD_360_1242_U55 P3_ADD_360_1242_U176 ; P3_ADD_360_1242_U177
g19567 nand P3_ADD_360_1242_U156 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_360_1242_U178
g19568 nand P3_ADD_360_1242_U51 P3_ADD_360_1242_U178 ; P3_ADD_360_1242_U179
g19569 nand P3_ADD_360_1242_U155 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_360_1242_U180
g19570 nand P3_ADD_360_1242_U48 P3_ADD_360_1242_U180 ; P3_ADD_360_1242_U181
g19571 nand P3_ADD_360_1242_U47 P3_ADD_360_1242_U46 ; P3_ADD_360_1242_U182
g19572 nand P3_ADD_360_1242_U119 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_360_1242_U183
g19573 nand P3_ADD_360_1242_U44 P3_ADD_360_1242_U183 ; P3_ADD_360_1242_U184
g19574 nand P3_ADD_360_1242_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_360_1242_U185
g19575 nand P3_ADD_360_1242_U42 P3_ADD_360_1242_U185 ; P3_ADD_360_1242_U186
g19576 nand P3_ADD_360_1242_U165 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_360_1242_U187
g19577 nand P3_ADD_360_U18 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_360_1242_U188
g19578 nand P3_ADD_360_U16 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_360_1242_U189
g19579 nand P3_ADD_360_1242_U92 P3_ADD_360_1242_U123 ; P3_ADD_360_1242_U190
g19580 nand P3_ADD_360_1242_U93 P3_ADD_360_1242_U40 ; P3_ADD_360_1242_U191
g19581 nand P3_ADD_360_1242_U122 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_360_1242_U192
g19582 nand P3_ADD_360_1242_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_360_1242_U193
g19583 nand P3_ADD_360_1242_U148 P3_ADD_360_1242_U39 ; P3_ADD_360_1242_U194
g19584 nand P3_ADD_360_1242_U37 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_360_1242_U195
g19585 nand P3_ADD_360_U5 P3_ADD_360_1242_U38 ; P3_ADD_360_1242_U196
g19586 nand P3_ADD_360_1242_U37 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_360_1242_U197
g19587 nand P3_ADD_360_U5 P3_ADD_360_1242_U38 ; P3_ADD_360_1242_U198
g19588 nand P3_ADD_360_1242_U198 P3_ADD_360_1242_U197 ; P3_ADD_360_1242_U199
g19589 nand P3_ADD_360_1242_U107 P3_ADD_360_1242_U108 ; P3_ADD_360_1242_U200
g19590 nand P3_ADD_360_1242_U144 P3_ADD_360_1242_U199 ; P3_ADD_360_1242_U201
g19591 nand P3_ADD_360_1242_U36 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_360_1242_U202
g19592 nand P3_ADD_360_U16 P3_ADD_360_1242_U35 ; P3_ADD_360_1242_U203
g19593 nand P3_ADD_360_1242_U36 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_360_1242_U204
g19594 nand P3_ADD_360_U16 P3_ADD_360_1242_U35 ; P3_ADD_360_1242_U205
g19595 nand P3_ADD_360_1242_U205 P3_ADD_360_1242_U204 ; P3_ADD_360_1242_U206
g19596 nand P3_ADD_360_1242_U109 P3_ADD_360_1242_U110 ; P3_ADD_360_1242_U207
g19597 nand P3_ADD_360_1242_U142 P3_ADD_360_1242_U206 ; P3_ADD_360_1242_U208
g19598 nand P3_ADD_360_1242_U33 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_360_1242_U209
g19599 nand P3_ADD_360_U17 P3_ADD_360_1242_U34 ; P3_ADD_360_1242_U210
g19600 nand P3_ADD_360_1242_U33 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_360_1242_U211
g19601 nand P3_ADD_360_U17 P3_ADD_360_1242_U34 ; P3_ADD_360_1242_U212
g19602 nand P3_ADD_360_1242_U212 P3_ADD_360_1242_U211 ; P3_ADD_360_1242_U213
g19603 nand P3_ADD_360_1242_U111 P3_ADD_360_1242_U112 ; P3_ADD_360_1242_U214
g19604 nand P3_ADD_360_1242_U138 P3_ADD_360_1242_U213 ; P3_ADD_360_1242_U215
g19605 nand P3_ADD_360_1242_U32 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_360_1242_U216
g19606 nand P3_ADD_360_U18 P3_ADD_360_1242_U31 ; P3_ADD_360_1242_U217
g19607 nand P3_ADD_360_1242_U32 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_360_1242_U218
g19608 nand P3_ADD_360_U18 P3_ADD_360_1242_U31 ; P3_ADD_360_1242_U219
g19609 nand P3_ADD_360_1242_U219 P3_ADD_360_1242_U218 ; P3_ADD_360_1242_U220
g19610 nand P3_ADD_360_1242_U113 P3_ADD_360_1242_U114 ; P3_ADD_360_1242_U221
g19611 nand P3_ADD_360_1242_U136 P3_ADD_360_1242_U220 ; P3_ADD_360_1242_U222
g19612 nand P3_ADD_360_1242_U20 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_360_1242_U223
g19613 nand P3_ADD_360_U19 P3_ADD_360_1242_U21 ; P3_ADD_360_1242_U224
g19614 nand P3_ADD_360_1242_U22 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_360_1242_U225
g19615 nand P3_ADD_360_U20 P3_ADD_360_1242_U23 ; P3_ADD_360_1242_U226
g19616 nand P3_ADD_360_1242_U187 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_360_1242_U227
g19617 nand P3_ADD_360_1242_U165 P3_ADD_360_1242_U116 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_360_1242_U228
g19618 nand P3_ADD_360_1242_U73 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_360_1242_U229
g19619 nand P3_ADD_360_1242_U165 P3_ADD_360_1242_U74 ; P3_ADD_360_1242_U230
g19620 nand P3_ADD_360_1242_U29 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_360_1242_U231
g19621 nand P3_ADD_360_U21 P3_ADD_360_1242_U30 ; P3_ADD_360_1242_U232
g19622 nand P3_ADD_360_1242_U29 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_360_1242_U233
g19623 nand P3_ADD_360_U21 P3_ADD_360_1242_U30 ; P3_ADD_360_1242_U234
g19624 nand P3_ADD_360_1242_U234 P3_ADD_360_1242_U233 ; P3_ADD_360_1242_U235
g19625 nand P3_ADD_360_1242_U117 P3_ADD_360_1242_U118 ; P3_ADD_360_1242_U236
g19626 nand P3_ADD_360_1242_U128 P3_ADD_360_1242_U235 ; P3_ADD_360_1242_U237
g19627 nand P3_ADD_360_1242_U68 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_360_1242_U238
g19628 nand P3_ADD_360_1242_U163 P3_ADD_360_1242_U70 ; P3_ADD_360_1242_U239
g19629 nand P3_ADD_360_1242_U63 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_360_1242_U240
g19630 nand P3_ADD_360_1242_U161 P3_ADD_360_1242_U65 ; P3_ADD_360_1242_U241
g19631 nand P3_ADD_360_1242_U60 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_360_1242_U242
g19632 nand P3_ADD_360_1242_U160 P3_ADD_360_1242_U62 ; P3_ADD_360_1242_U243
g19633 nand P3_ADD_360_1242_U27 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_360_1242_U244
g19634 nand P3_ADD_360_1242_U124 P3_ADD_360_1242_U26 ; P3_ADD_360_1242_U245
g19635 nand P3_ADD_360_1242_U245 P3_ADD_360_1242_U244 ; P3_ADD_360_1242_U246
g19636 nand P3_ADD_360_1242_U27 P3_ADD_360_1242_U26 P3_ADD_360_U4 ; P3_ADD_360_1242_U247
g19637 nand P3_ADD_360_1242_U246 P3_ADD_360_1242_U28 ; P3_ADD_360_1242_U248
g19638 nand P3_ADD_360_1242_U53 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_360_1242_U249
g19639 nand P3_ADD_360_1242_U157 P3_ADD_360_1242_U54 ; P3_ADD_360_1242_U250
g19640 nand P3_ADD_360_1242_U50 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_360_1242_U251
g19641 nand P3_ADD_360_1242_U156 P3_ADD_360_1242_U52 ; P3_ADD_360_1242_U252
g19642 nand P3_ADD_360_1242_U76 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_360_1242_U253
g19643 nand P3_ADD_360_1242_U155 P3_ADD_360_1242_U49 ; P3_ADD_360_1242_U254
g19644 nand P3_ADD_360_1242_U119 P3_ADD_360_1242_U43 ; P3_ADD_360_1242_U255
g19645 nand P3_ADD_360_1242_U45 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_360_1242_U256
g19646 nand P3_ADD_360_1242_U24 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_360_1242_U257
g19647 nand P3_U2621 P3_ADD_360_1242_U25 ; P3_ADD_360_1242_U258
g19648 or P3_LT_563_1260_U7 P3_U3304 ; P3_LT_563_1260_U6
g19649 nor P3_SUB_563_U7 P3_SUB_563_U6 ; P3_LT_563_1260_U7
g19650 not P3_U3301 ; P3_SUB_589_U6
g19651 not P3_U3302 ; P3_SUB_589_U7
g19652 not P3_U2632 ; P3_SUB_589_U8
g19653 not P3_U3300 ; P3_SUB_589_U9
g19654 not P3_REIP_REG_1__SCAN_IN ; P3_ADD_467_U4
g19655 not P3_REIP_REG_2__SCAN_IN ; P3_ADD_467_U5
g19656 nand P3_REIP_REG_1__SCAN_IN P3_REIP_REG_2__SCAN_IN ; P3_ADD_467_U6
g19657 not P3_REIP_REG_3__SCAN_IN ; P3_ADD_467_U7
g19658 nand P3_ADD_467_U94 P3_REIP_REG_3__SCAN_IN ; P3_ADD_467_U8
g19659 not P3_REIP_REG_4__SCAN_IN ; P3_ADD_467_U9
g19660 nand P3_ADD_467_U95 P3_REIP_REG_4__SCAN_IN ; P3_ADD_467_U10
g19661 not P3_REIP_REG_5__SCAN_IN ; P3_ADD_467_U11
g19662 nand P3_ADD_467_U96 P3_REIP_REG_5__SCAN_IN ; P3_ADD_467_U12
g19663 not P3_REIP_REG_6__SCAN_IN ; P3_ADD_467_U13
g19664 nand P3_ADD_467_U97 P3_REIP_REG_6__SCAN_IN ; P3_ADD_467_U14
g19665 not P3_REIP_REG_7__SCAN_IN ; P3_ADD_467_U15
g19666 nand P3_ADD_467_U98 P3_REIP_REG_7__SCAN_IN ; P3_ADD_467_U16
g19667 not P3_REIP_REG_8__SCAN_IN ; P3_ADD_467_U17
g19668 not P3_REIP_REG_9__SCAN_IN ; P3_ADD_467_U18
g19669 nand P3_ADD_467_U99 P3_REIP_REG_8__SCAN_IN ; P3_ADD_467_U19
g19670 nand P3_ADD_467_U100 P3_REIP_REG_9__SCAN_IN ; P3_ADD_467_U20
g19671 not P3_REIP_REG_10__SCAN_IN ; P3_ADD_467_U21
g19672 nand P3_ADD_467_U101 P3_REIP_REG_10__SCAN_IN ; P3_ADD_467_U22
g19673 not P3_REIP_REG_11__SCAN_IN ; P3_ADD_467_U23
g19674 nand P3_ADD_467_U102 P3_REIP_REG_11__SCAN_IN ; P3_ADD_467_U24
g19675 not P3_REIP_REG_12__SCAN_IN ; P3_ADD_467_U25
g19676 nand P3_ADD_467_U103 P3_REIP_REG_12__SCAN_IN ; P3_ADD_467_U26
g19677 not P3_REIP_REG_13__SCAN_IN ; P3_ADD_467_U27
g19678 nand P3_ADD_467_U104 P3_REIP_REG_13__SCAN_IN ; P3_ADD_467_U28
g19679 not P3_REIP_REG_14__SCAN_IN ; P3_ADD_467_U29
g19680 nand P3_ADD_467_U105 P3_REIP_REG_14__SCAN_IN ; P3_ADD_467_U30
g19681 not P3_REIP_REG_15__SCAN_IN ; P3_ADD_467_U31
g19682 nand P3_ADD_467_U106 P3_REIP_REG_15__SCAN_IN ; P3_ADD_467_U32
g19683 not P3_REIP_REG_16__SCAN_IN ; P3_ADD_467_U33
g19684 nand P3_ADD_467_U107 P3_REIP_REG_16__SCAN_IN ; P3_ADD_467_U34
g19685 not P3_REIP_REG_17__SCAN_IN ; P3_ADD_467_U35
g19686 nand P3_ADD_467_U108 P3_REIP_REG_17__SCAN_IN ; P3_ADD_467_U36
g19687 not P3_REIP_REG_18__SCAN_IN ; P3_ADD_467_U37
g19688 nand P3_ADD_467_U109 P3_REIP_REG_18__SCAN_IN ; P3_ADD_467_U38
g19689 not P3_REIP_REG_19__SCAN_IN ; P3_ADD_467_U39
g19690 nand P3_ADD_467_U110 P3_REIP_REG_19__SCAN_IN ; P3_ADD_467_U40
g19691 not P3_REIP_REG_20__SCAN_IN ; P3_ADD_467_U41
g19692 nand P3_ADD_467_U111 P3_REIP_REG_20__SCAN_IN ; P3_ADD_467_U42
g19693 not P3_REIP_REG_21__SCAN_IN ; P3_ADD_467_U43
g19694 nand P3_ADD_467_U112 P3_REIP_REG_21__SCAN_IN ; P3_ADD_467_U44
g19695 not P3_REIP_REG_22__SCAN_IN ; P3_ADD_467_U45
g19696 nand P3_ADD_467_U113 P3_REIP_REG_22__SCAN_IN ; P3_ADD_467_U46
g19697 not P3_REIP_REG_23__SCAN_IN ; P3_ADD_467_U47
g19698 nand P3_ADD_467_U114 P3_REIP_REG_23__SCAN_IN ; P3_ADD_467_U48
g19699 not P3_REIP_REG_24__SCAN_IN ; P3_ADD_467_U49
g19700 nand P3_ADD_467_U115 P3_REIP_REG_24__SCAN_IN ; P3_ADD_467_U50
g19701 not P3_REIP_REG_25__SCAN_IN ; P3_ADD_467_U51
g19702 nand P3_ADD_467_U116 P3_REIP_REG_25__SCAN_IN ; P3_ADD_467_U52
g19703 not P3_REIP_REG_26__SCAN_IN ; P3_ADD_467_U53
g19704 nand P3_ADD_467_U117 P3_REIP_REG_26__SCAN_IN ; P3_ADD_467_U54
g19705 not P3_REIP_REG_27__SCAN_IN ; P3_ADD_467_U55
g19706 nand P3_ADD_467_U118 P3_REIP_REG_27__SCAN_IN ; P3_ADD_467_U56
g19707 not P3_REIP_REG_28__SCAN_IN ; P3_ADD_467_U57
g19708 nand P3_ADD_467_U119 P3_REIP_REG_28__SCAN_IN ; P3_ADD_467_U58
g19709 not P3_REIP_REG_29__SCAN_IN ; P3_ADD_467_U59
g19710 nand P3_ADD_467_U120 P3_REIP_REG_29__SCAN_IN ; P3_ADD_467_U60
g19711 not P3_REIP_REG_30__SCAN_IN ; P3_ADD_467_U61
g19712 nand P3_ADD_467_U124 P3_ADD_467_U123 ; P3_ADD_467_U62
g19713 nand P3_ADD_467_U126 P3_ADD_467_U125 ; P3_ADD_467_U63
g19714 nand P3_ADD_467_U128 P3_ADD_467_U127 ; P3_ADD_467_U64
g19715 nand P3_ADD_467_U130 P3_ADD_467_U129 ; P3_ADD_467_U65
g19716 nand P3_ADD_467_U132 P3_ADD_467_U131 ; P3_ADD_467_U66
g19717 nand P3_ADD_467_U134 P3_ADD_467_U133 ; P3_ADD_467_U67
g19718 nand P3_ADD_467_U136 P3_ADD_467_U135 ; P3_ADD_467_U68
g19719 nand P3_ADD_467_U138 P3_ADD_467_U137 ; P3_ADD_467_U69
g19720 nand P3_ADD_467_U140 P3_ADD_467_U139 ; P3_ADD_467_U70
g19721 nand P3_ADD_467_U142 P3_ADD_467_U141 ; P3_ADD_467_U71
g19722 nand P3_ADD_467_U144 P3_ADD_467_U143 ; P3_ADD_467_U72
g19723 nand P3_ADD_467_U146 P3_ADD_467_U145 ; P3_ADD_467_U73
g19724 nand P3_ADD_467_U148 P3_ADD_467_U147 ; P3_ADD_467_U74
g19725 nand P3_ADD_467_U150 P3_ADD_467_U149 ; P3_ADD_467_U75
g19726 nand P3_ADD_467_U152 P3_ADD_467_U151 ; P3_ADD_467_U76
g19727 nand P3_ADD_467_U154 P3_ADD_467_U153 ; P3_ADD_467_U77
g19728 nand P3_ADD_467_U156 P3_ADD_467_U155 ; P3_ADD_467_U78
g19729 nand P3_ADD_467_U158 P3_ADD_467_U157 ; P3_ADD_467_U79
g19730 nand P3_ADD_467_U160 P3_ADD_467_U159 ; P3_ADD_467_U80
g19731 nand P3_ADD_467_U162 P3_ADD_467_U161 ; P3_ADD_467_U81
g19732 nand P3_ADD_467_U164 P3_ADD_467_U163 ; P3_ADD_467_U82
g19733 nand P3_ADD_467_U166 P3_ADD_467_U165 ; P3_ADD_467_U83
g19734 nand P3_ADD_467_U168 P3_ADD_467_U167 ; P3_ADD_467_U84
g19735 nand P3_ADD_467_U170 P3_ADD_467_U169 ; P3_ADD_467_U85
g19736 nand P3_ADD_467_U172 P3_ADD_467_U171 ; P3_ADD_467_U86
g19737 nand P3_ADD_467_U174 P3_ADD_467_U173 ; P3_ADD_467_U87
g19738 nand P3_ADD_467_U176 P3_ADD_467_U175 ; P3_ADD_467_U88
g19739 nand P3_ADD_467_U178 P3_ADD_467_U177 ; P3_ADD_467_U89
g19740 nand P3_ADD_467_U180 P3_ADD_467_U179 ; P3_ADD_467_U90
g19741 nand P3_ADD_467_U182 P3_ADD_467_U181 ; P3_ADD_467_U91
g19742 not P3_REIP_REG_31__SCAN_IN ; P3_ADD_467_U92
g19743 nand P3_ADD_467_U121 P3_REIP_REG_30__SCAN_IN ; P3_ADD_467_U93
g19744 not P3_ADD_467_U6 ; P3_ADD_467_U94
g19745 not P3_ADD_467_U8 ; P3_ADD_467_U95
g19746 not P3_ADD_467_U10 ; P3_ADD_467_U96
g19747 not P3_ADD_467_U12 ; P3_ADD_467_U97
g19748 not P3_ADD_467_U14 ; P3_ADD_467_U98
g19749 not P3_ADD_467_U16 ; P3_ADD_467_U99
g19750 not P3_ADD_467_U19 ; P3_ADD_467_U100
g19751 not P3_ADD_467_U20 ; P3_ADD_467_U101
g19752 not P3_ADD_467_U22 ; P3_ADD_467_U102
g19753 not P3_ADD_467_U24 ; P3_ADD_467_U103
g19754 not P3_ADD_467_U26 ; P3_ADD_467_U104
g19755 not P3_ADD_467_U28 ; P3_ADD_467_U105
g19756 not P3_ADD_467_U30 ; P3_ADD_467_U106
g19757 not P3_ADD_467_U32 ; P3_ADD_467_U107
g19758 not P3_ADD_467_U34 ; P3_ADD_467_U108
g19759 not P3_ADD_467_U36 ; P3_ADD_467_U109
g19760 not P3_ADD_467_U38 ; P3_ADD_467_U110
g19761 not P3_ADD_467_U40 ; P3_ADD_467_U111
g19762 not P3_ADD_467_U42 ; P3_ADD_467_U112
g19763 not P3_ADD_467_U44 ; P3_ADD_467_U113
g19764 not P3_ADD_467_U46 ; P3_ADD_467_U114
g19765 not P3_ADD_467_U48 ; P3_ADD_467_U115
g19766 not P3_ADD_467_U50 ; P3_ADD_467_U116
g19767 not P3_ADD_467_U52 ; P3_ADD_467_U117
g19768 not P3_ADD_467_U54 ; P3_ADD_467_U118
g19769 not P3_ADD_467_U56 ; P3_ADD_467_U119
g19770 not P3_ADD_467_U58 ; P3_ADD_467_U120
g19771 not P3_ADD_467_U60 ; P3_ADD_467_U121
g19772 not P3_ADD_467_U93 ; P3_ADD_467_U122
g19773 nand P3_ADD_467_U19 P3_REIP_REG_9__SCAN_IN ; P3_ADD_467_U123
g19774 nand P3_ADD_467_U100 P3_ADD_467_U18 ; P3_ADD_467_U124
g19775 nand P3_ADD_467_U16 P3_REIP_REG_8__SCAN_IN ; P3_ADD_467_U125
g19776 nand P3_ADD_467_U99 P3_ADD_467_U17 ; P3_ADD_467_U126
g19777 nand P3_ADD_467_U14 P3_REIP_REG_7__SCAN_IN ; P3_ADD_467_U127
g19778 nand P3_ADD_467_U98 P3_ADD_467_U15 ; P3_ADD_467_U128
g19779 nand P3_ADD_467_U12 P3_REIP_REG_6__SCAN_IN ; P3_ADD_467_U129
g19780 nand P3_ADD_467_U97 P3_ADD_467_U13 ; P3_ADD_467_U130
g19781 nand P3_ADD_467_U10 P3_REIP_REG_5__SCAN_IN ; P3_ADD_467_U131
g19782 nand P3_ADD_467_U96 P3_ADD_467_U11 ; P3_ADD_467_U132
g19783 nand P3_ADD_467_U8 P3_REIP_REG_4__SCAN_IN ; P3_ADD_467_U133
g19784 nand P3_ADD_467_U95 P3_ADD_467_U9 ; P3_ADD_467_U134
g19785 nand P3_ADD_467_U6 P3_REIP_REG_3__SCAN_IN ; P3_ADD_467_U135
g19786 nand P3_ADD_467_U94 P3_ADD_467_U7 ; P3_ADD_467_U136
g19787 nand P3_ADD_467_U93 P3_REIP_REG_31__SCAN_IN ; P3_ADD_467_U137
g19788 nand P3_ADD_467_U122 P3_ADD_467_U92 ; P3_ADD_467_U138
g19789 nand P3_ADD_467_U60 P3_REIP_REG_30__SCAN_IN ; P3_ADD_467_U139
g19790 nand P3_ADD_467_U121 P3_ADD_467_U61 ; P3_ADD_467_U140
g19791 nand P3_ADD_467_U4 P3_REIP_REG_2__SCAN_IN ; P3_ADD_467_U141
g19792 nand P3_ADD_467_U5 P3_REIP_REG_1__SCAN_IN ; P3_ADD_467_U142
g19793 nand P3_ADD_467_U58 P3_REIP_REG_29__SCAN_IN ; P3_ADD_467_U143
g19794 nand P3_ADD_467_U120 P3_ADD_467_U59 ; P3_ADD_467_U144
g19795 nand P3_ADD_467_U56 P3_REIP_REG_28__SCAN_IN ; P3_ADD_467_U145
g19796 nand P3_ADD_467_U119 P3_ADD_467_U57 ; P3_ADD_467_U146
g19797 nand P3_ADD_467_U54 P3_REIP_REG_27__SCAN_IN ; P3_ADD_467_U147
g19798 nand P3_ADD_467_U118 P3_ADD_467_U55 ; P3_ADD_467_U148
g19799 nand P3_ADD_467_U52 P3_REIP_REG_26__SCAN_IN ; P3_ADD_467_U149
g19800 nand P3_ADD_467_U117 P3_ADD_467_U53 ; P3_ADD_467_U150
g19801 nand P3_ADD_467_U50 P3_REIP_REG_25__SCAN_IN ; P3_ADD_467_U151
g19802 nand P3_ADD_467_U116 P3_ADD_467_U51 ; P3_ADD_467_U152
g19803 nand P3_ADD_467_U48 P3_REIP_REG_24__SCAN_IN ; P3_ADD_467_U153
g19804 nand P3_ADD_467_U115 P3_ADD_467_U49 ; P3_ADD_467_U154
g19805 nand P3_ADD_467_U46 P3_REIP_REG_23__SCAN_IN ; P3_ADD_467_U155
g19806 nand P3_ADD_467_U114 P3_ADD_467_U47 ; P3_ADD_467_U156
g19807 nand P3_ADD_467_U44 P3_REIP_REG_22__SCAN_IN ; P3_ADD_467_U157
g19808 nand P3_ADD_467_U113 P3_ADD_467_U45 ; P3_ADD_467_U158
g19809 nand P3_ADD_467_U42 P3_REIP_REG_21__SCAN_IN ; P3_ADD_467_U159
g19810 nand P3_ADD_467_U112 P3_ADD_467_U43 ; P3_ADD_467_U160
g19811 nand P3_ADD_467_U40 P3_REIP_REG_20__SCAN_IN ; P3_ADD_467_U161
g19812 nand P3_ADD_467_U111 P3_ADD_467_U41 ; P3_ADD_467_U162
g19813 nand P3_ADD_467_U38 P3_REIP_REG_19__SCAN_IN ; P3_ADD_467_U163
g19814 nand P3_ADD_467_U110 P3_ADD_467_U39 ; P3_ADD_467_U164
g19815 nand P3_ADD_467_U36 P3_REIP_REG_18__SCAN_IN ; P3_ADD_467_U165
g19816 nand P3_ADD_467_U109 P3_ADD_467_U37 ; P3_ADD_467_U166
g19817 nand P3_ADD_467_U34 P3_REIP_REG_17__SCAN_IN ; P3_ADD_467_U167
g19818 nand P3_ADD_467_U108 P3_ADD_467_U35 ; P3_ADD_467_U168
g19819 nand P3_ADD_467_U32 P3_REIP_REG_16__SCAN_IN ; P3_ADD_467_U169
g19820 nand P3_ADD_467_U107 P3_ADD_467_U33 ; P3_ADD_467_U170
g19821 nand P3_ADD_467_U30 P3_REIP_REG_15__SCAN_IN ; P3_ADD_467_U171
g19822 nand P3_ADD_467_U106 P3_ADD_467_U31 ; P3_ADD_467_U172
g19823 nand P3_ADD_467_U28 P3_REIP_REG_14__SCAN_IN ; P3_ADD_467_U173
g19824 nand P3_ADD_467_U105 P3_ADD_467_U29 ; P3_ADD_467_U174
g19825 nand P3_ADD_467_U26 P3_REIP_REG_13__SCAN_IN ; P3_ADD_467_U175
g19826 nand P3_ADD_467_U104 P3_ADD_467_U27 ; P3_ADD_467_U176
g19827 nand P3_ADD_467_U24 P3_REIP_REG_12__SCAN_IN ; P3_ADD_467_U177
g19828 nand P3_ADD_467_U103 P3_ADD_467_U25 ; P3_ADD_467_U178
g19829 nand P3_ADD_467_U22 P3_REIP_REG_11__SCAN_IN ; P3_ADD_467_U179
g19830 nand P3_ADD_467_U102 P3_ADD_467_U23 ; P3_ADD_467_U180
g19831 nand P3_ADD_467_U20 P3_REIP_REG_10__SCAN_IN ; P3_ADD_467_U181
g19832 nand P3_ADD_467_U101 P3_ADD_467_U21 ; P3_ADD_467_U182
g19833 not P3_REIP_REG_1__SCAN_IN ; P3_ADD_430_U4
g19834 not P3_REIP_REG_2__SCAN_IN ; P3_ADD_430_U5
g19835 nand P3_REIP_REG_1__SCAN_IN P3_REIP_REG_2__SCAN_IN ; P3_ADD_430_U6
g19836 not P3_REIP_REG_3__SCAN_IN ; P3_ADD_430_U7
g19837 nand P3_ADD_430_U94 P3_REIP_REG_3__SCAN_IN ; P3_ADD_430_U8
g19838 not P3_REIP_REG_4__SCAN_IN ; P3_ADD_430_U9
g19839 nand P3_ADD_430_U95 P3_REIP_REG_4__SCAN_IN ; P3_ADD_430_U10
g19840 not P3_REIP_REG_5__SCAN_IN ; P3_ADD_430_U11
g19841 nand P3_ADD_430_U96 P3_REIP_REG_5__SCAN_IN ; P3_ADD_430_U12
g19842 not P3_REIP_REG_6__SCAN_IN ; P3_ADD_430_U13
g19843 nand P3_ADD_430_U97 P3_REIP_REG_6__SCAN_IN ; P3_ADD_430_U14
g19844 not P3_REIP_REG_7__SCAN_IN ; P3_ADD_430_U15
g19845 nand P3_ADD_430_U98 P3_REIP_REG_7__SCAN_IN ; P3_ADD_430_U16
g19846 not P3_REIP_REG_8__SCAN_IN ; P3_ADD_430_U17
g19847 not P3_REIP_REG_9__SCAN_IN ; P3_ADD_430_U18
g19848 nand P3_ADD_430_U99 P3_REIP_REG_8__SCAN_IN ; P3_ADD_430_U19
g19849 nand P3_ADD_430_U100 P3_REIP_REG_9__SCAN_IN ; P3_ADD_430_U20
g19850 not P3_REIP_REG_10__SCAN_IN ; P3_ADD_430_U21
g19851 nand P3_ADD_430_U101 P3_REIP_REG_10__SCAN_IN ; P3_ADD_430_U22
g19852 not P3_REIP_REG_11__SCAN_IN ; P3_ADD_430_U23
g19853 nand P3_ADD_430_U102 P3_REIP_REG_11__SCAN_IN ; P3_ADD_430_U24
g19854 not P3_REIP_REG_12__SCAN_IN ; P3_ADD_430_U25
g19855 nand P3_ADD_430_U103 P3_REIP_REG_12__SCAN_IN ; P3_ADD_430_U26
g19856 not P3_REIP_REG_13__SCAN_IN ; P3_ADD_430_U27
g19857 nand P3_ADD_430_U104 P3_REIP_REG_13__SCAN_IN ; P3_ADD_430_U28
g19858 not P3_REIP_REG_14__SCAN_IN ; P3_ADD_430_U29
g19859 nand P3_ADD_430_U105 P3_REIP_REG_14__SCAN_IN ; P3_ADD_430_U30
g19860 not P3_REIP_REG_15__SCAN_IN ; P3_ADD_430_U31
g19861 nand P3_ADD_430_U106 P3_REIP_REG_15__SCAN_IN ; P3_ADD_430_U32
g19862 not P3_REIP_REG_16__SCAN_IN ; P3_ADD_430_U33
g19863 nand P3_ADD_430_U107 P3_REIP_REG_16__SCAN_IN ; P3_ADD_430_U34
g19864 not P3_REIP_REG_17__SCAN_IN ; P3_ADD_430_U35
g19865 nand P3_ADD_430_U108 P3_REIP_REG_17__SCAN_IN ; P3_ADD_430_U36
g19866 not P3_REIP_REG_18__SCAN_IN ; P3_ADD_430_U37
g19867 nand P3_ADD_430_U109 P3_REIP_REG_18__SCAN_IN ; P3_ADD_430_U38
g19868 not P3_REIP_REG_19__SCAN_IN ; P3_ADD_430_U39
g19869 nand P3_ADD_430_U110 P3_REIP_REG_19__SCAN_IN ; P3_ADD_430_U40
g19870 not P3_REIP_REG_20__SCAN_IN ; P3_ADD_430_U41
g19871 nand P3_ADD_430_U111 P3_REIP_REG_20__SCAN_IN ; P3_ADD_430_U42
g19872 not P3_REIP_REG_21__SCAN_IN ; P3_ADD_430_U43
g19873 nand P3_ADD_430_U112 P3_REIP_REG_21__SCAN_IN ; P3_ADD_430_U44
g19874 not P3_REIP_REG_22__SCAN_IN ; P3_ADD_430_U45
g19875 nand P3_ADD_430_U113 P3_REIP_REG_22__SCAN_IN ; P3_ADD_430_U46
g19876 not P3_REIP_REG_23__SCAN_IN ; P3_ADD_430_U47
g19877 nand P3_ADD_430_U114 P3_REIP_REG_23__SCAN_IN ; P3_ADD_430_U48
g19878 not P3_REIP_REG_24__SCAN_IN ; P3_ADD_430_U49
g19879 nand P3_ADD_430_U115 P3_REIP_REG_24__SCAN_IN ; P3_ADD_430_U50
g19880 not P3_REIP_REG_25__SCAN_IN ; P3_ADD_430_U51
g19881 nand P3_ADD_430_U116 P3_REIP_REG_25__SCAN_IN ; P3_ADD_430_U52
g19882 not P3_REIP_REG_26__SCAN_IN ; P3_ADD_430_U53
g19883 nand P3_ADD_430_U117 P3_REIP_REG_26__SCAN_IN ; P3_ADD_430_U54
g19884 not P3_REIP_REG_27__SCAN_IN ; P3_ADD_430_U55
g19885 nand P3_ADD_430_U118 P3_REIP_REG_27__SCAN_IN ; P3_ADD_430_U56
g19886 not P3_REIP_REG_28__SCAN_IN ; P3_ADD_430_U57
g19887 nand P3_ADD_430_U119 P3_REIP_REG_28__SCAN_IN ; P3_ADD_430_U58
g19888 not P3_REIP_REG_29__SCAN_IN ; P3_ADD_430_U59
g19889 nand P3_ADD_430_U120 P3_REIP_REG_29__SCAN_IN ; P3_ADD_430_U60
g19890 not P3_REIP_REG_30__SCAN_IN ; P3_ADD_430_U61
g19891 nand P3_ADD_430_U124 P3_ADD_430_U123 ; P3_ADD_430_U62
g19892 nand P3_ADD_430_U126 P3_ADD_430_U125 ; P3_ADD_430_U63
g19893 nand P3_ADD_430_U128 P3_ADD_430_U127 ; P3_ADD_430_U64
g19894 nand P3_ADD_430_U130 P3_ADD_430_U129 ; P3_ADD_430_U65
g19895 nand P3_ADD_430_U132 P3_ADD_430_U131 ; P3_ADD_430_U66
g19896 nand P3_ADD_430_U134 P3_ADD_430_U133 ; P3_ADD_430_U67
g19897 nand P3_ADD_430_U136 P3_ADD_430_U135 ; P3_ADD_430_U68
g19898 nand P3_ADD_430_U138 P3_ADD_430_U137 ; P3_ADD_430_U69
g19899 nand P3_ADD_430_U140 P3_ADD_430_U139 ; P3_ADD_430_U70
g19900 nand P3_ADD_430_U142 P3_ADD_430_U141 ; P3_ADD_430_U71
g19901 nand P3_ADD_430_U144 P3_ADD_430_U143 ; P3_ADD_430_U72
g19902 nand P3_ADD_430_U146 P3_ADD_430_U145 ; P3_ADD_430_U73
g19903 nand P3_ADD_430_U148 P3_ADD_430_U147 ; P3_ADD_430_U74
g19904 nand P3_ADD_430_U150 P3_ADD_430_U149 ; P3_ADD_430_U75
g19905 nand P3_ADD_430_U152 P3_ADD_430_U151 ; P3_ADD_430_U76
g19906 nand P3_ADD_430_U154 P3_ADD_430_U153 ; P3_ADD_430_U77
g19907 nand P3_ADD_430_U156 P3_ADD_430_U155 ; P3_ADD_430_U78
g19908 nand P3_ADD_430_U158 P3_ADD_430_U157 ; P3_ADD_430_U79
g19909 nand P3_ADD_430_U160 P3_ADD_430_U159 ; P3_ADD_430_U80
g19910 nand P3_ADD_430_U162 P3_ADD_430_U161 ; P3_ADD_430_U81
g19911 nand P3_ADD_430_U164 P3_ADD_430_U163 ; P3_ADD_430_U82
g19912 nand P3_ADD_430_U166 P3_ADD_430_U165 ; P3_ADD_430_U83
g19913 nand P3_ADD_430_U168 P3_ADD_430_U167 ; P3_ADD_430_U84
g19914 nand P3_ADD_430_U170 P3_ADD_430_U169 ; P3_ADD_430_U85
g19915 nand P3_ADD_430_U172 P3_ADD_430_U171 ; P3_ADD_430_U86
g19916 nand P3_ADD_430_U174 P3_ADD_430_U173 ; P3_ADD_430_U87
g19917 nand P3_ADD_430_U176 P3_ADD_430_U175 ; P3_ADD_430_U88
g19918 nand P3_ADD_430_U178 P3_ADD_430_U177 ; P3_ADD_430_U89
g19919 nand P3_ADD_430_U180 P3_ADD_430_U179 ; P3_ADD_430_U90
g19920 nand P3_ADD_430_U182 P3_ADD_430_U181 ; P3_ADD_430_U91
g19921 not P3_REIP_REG_31__SCAN_IN ; P3_ADD_430_U92
g19922 nand P3_ADD_430_U121 P3_REIP_REG_30__SCAN_IN ; P3_ADD_430_U93
g19923 not P3_ADD_430_U6 ; P3_ADD_430_U94
g19924 not P3_ADD_430_U8 ; P3_ADD_430_U95
g19925 not P3_ADD_430_U10 ; P3_ADD_430_U96
g19926 not P3_ADD_430_U12 ; P3_ADD_430_U97
g19927 not P3_ADD_430_U14 ; P3_ADD_430_U98
g19928 not P3_ADD_430_U16 ; P3_ADD_430_U99
g19929 not P3_ADD_430_U19 ; P3_ADD_430_U100
g19930 not P3_ADD_430_U20 ; P3_ADD_430_U101
g19931 not P3_ADD_430_U22 ; P3_ADD_430_U102
g19932 not P3_ADD_430_U24 ; P3_ADD_430_U103
g19933 not P3_ADD_430_U26 ; P3_ADD_430_U104
g19934 not P3_ADD_430_U28 ; P3_ADD_430_U105
g19935 not P3_ADD_430_U30 ; P3_ADD_430_U106
g19936 not P3_ADD_430_U32 ; P3_ADD_430_U107
g19937 not P3_ADD_430_U34 ; P3_ADD_430_U108
g19938 not P3_ADD_430_U36 ; P3_ADD_430_U109
g19939 not P3_ADD_430_U38 ; P3_ADD_430_U110
g19940 not P3_ADD_430_U40 ; P3_ADD_430_U111
g19941 not P3_ADD_430_U42 ; P3_ADD_430_U112
g19942 not P3_ADD_430_U44 ; P3_ADD_430_U113
g19943 not P3_ADD_430_U46 ; P3_ADD_430_U114
g19944 not P3_ADD_430_U48 ; P3_ADD_430_U115
g19945 not P3_ADD_430_U50 ; P3_ADD_430_U116
g19946 not P3_ADD_430_U52 ; P3_ADD_430_U117
g19947 not P3_ADD_430_U54 ; P3_ADD_430_U118
g19948 not P3_ADD_430_U56 ; P3_ADD_430_U119
g19949 not P3_ADD_430_U58 ; P3_ADD_430_U120
g19950 not P3_ADD_430_U60 ; P3_ADD_430_U121
g19951 not P3_ADD_430_U93 ; P3_ADD_430_U122
g19952 nand P3_ADD_430_U19 P3_REIP_REG_9__SCAN_IN ; P3_ADD_430_U123
g19953 nand P3_ADD_430_U100 P3_ADD_430_U18 ; P3_ADD_430_U124
g19954 nand P3_ADD_430_U16 P3_REIP_REG_8__SCAN_IN ; P3_ADD_430_U125
g19955 nand P3_ADD_430_U99 P3_ADD_430_U17 ; P3_ADD_430_U126
g19956 nand P3_ADD_430_U14 P3_REIP_REG_7__SCAN_IN ; P3_ADD_430_U127
g19957 nand P3_ADD_430_U98 P3_ADD_430_U15 ; P3_ADD_430_U128
g19958 nand P3_ADD_430_U12 P3_REIP_REG_6__SCAN_IN ; P3_ADD_430_U129
g19959 nand P3_ADD_430_U97 P3_ADD_430_U13 ; P3_ADD_430_U130
g19960 nand P3_ADD_430_U10 P3_REIP_REG_5__SCAN_IN ; P3_ADD_430_U131
g19961 nand P3_ADD_430_U96 P3_ADD_430_U11 ; P3_ADD_430_U132
g19962 nand P3_ADD_430_U8 P3_REIP_REG_4__SCAN_IN ; P3_ADD_430_U133
g19963 nand P3_ADD_430_U95 P3_ADD_430_U9 ; P3_ADD_430_U134
g19964 nand P3_ADD_430_U6 P3_REIP_REG_3__SCAN_IN ; P3_ADD_430_U135
g19965 nand P3_ADD_430_U94 P3_ADD_430_U7 ; P3_ADD_430_U136
g19966 nand P3_ADD_430_U93 P3_REIP_REG_31__SCAN_IN ; P3_ADD_430_U137
g19967 nand P3_ADD_430_U122 P3_ADD_430_U92 ; P3_ADD_430_U138
g19968 nand P3_ADD_430_U60 P3_REIP_REG_30__SCAN_IN ; P3_ADD_430_U139
g19969 nand P3_ADD_430_U121 P3_ADD_430_U61 ; P3_ADD_430_U140
g19970 nand P3_ADD_430_U4 P3_REIP_REG_2__SCAN_IN ; P3_ADD_430_U141
g19971 nand P3_ADD_430_U5 P3_REIP_REG_1__SCAN_IN ; P3_ADD_430_U142
g19972 nand P3_ADD_430_U58 P3_REIP_REG_29__SCAN_IN ; P3_ADD_430_U143
g19973 nand P3_ADD_430_U120 P3_ADD_430_U59 ; P3_ADD_430_U144
g19974 nand P3_ADD_430_U56 P3_REIP_REG_28__SCAN_IN ; P3_ADD_430_U145
g19975 nand P3_ADD_430_U119 P3_ADD_430_U57 ; P3_ADD_430_U146
g19976 nand P3_ADD_430_U54 P3_REIP_REG_27__SCAN_IN ; P3_ADD_430_U147
g19977 nand P3_ADD_430_U118 P3_ADD_430_U55 ; P3_ADD_430_U148
g19978 nand P3_ADD_430_U52 P3_REIP_REG_26__SCAN_IN ; P3_ADD_430_U149
g19979 nand P3_ADD_430_U117 P3_ADD_430_U53 ; P3_ADD_430_U150
g19980 nand P3_ADD_430_U50 P3_REIP_REG_25__SCAN_IN ; P3_ADD_430_U151
g19981 nand P3_ADD_430_U116 P3_ADD_430_U51 ; P3_ADD_430_U152
g19982 nand P3_ADD_430_U48 P3_REIP_REG_24__SCAN_IN ; P3_ADD_430_U153
g19983 nand P3_ADD_430_U115 P3_ADD_430_U49 ; P3_ADD_430_U154
g19984 nand P3_ADD_430_U46 P3_REIP_REG_23__SCAN_IN ; P3_ADD_430_U155
g19985 nand P3_ADD_430_U114 P3_ADD_430_U47 ; P3_ADD_430_U156
g19986 nand P3_ADD_430_U44 P3_REIP_REG_22__SCAN_IN ; P3_ADD_430_U157
g19987 nand P3_ADD_430_U113 P3_ADD_430_U45 ; P3_ADD_430_U158
g19988 nand P3_ADD_430_U42 P3_REIP_REG_21__SCAN_IN ; P3_ADD_430_U159
g19989 nand P3_ADD_430_U112 P3_ADD_430_U43 ; P3_ADD_430_U160
g19990 nand P3_ADD_430_U40 P3_REIP_REG_20__SCAN_IN ; P3_ADD_430_U161
g19991 nand P3_ADD_430_U111 P3_ADD_430_U41 ; P3_ADD_430_U162
g19992 nand P3_ADD_430_U38 P3_REIP_REG_19__SCAN_IN ; P3_ADD_430_U163
g19993 nand P3_ADD_430_U110 P3_ADD_430_U39 ; P3_ADD_430_U164
g19994 nand P3_ADD_430_U36 P3_REIP_REG_18__SCAN_IN ; P3_ADD_430_U165
g19995 nand P3_ADD_430_U109 P3_ADD_430_U37 ; P3_ADD_430_U166
g19996 nand P3_ADD_430_U34 P3_REIP_REG_17__SCAN_IN ; P3_ADD_430_U167
g19997 nand P3_ADD_430_U108 P3_ADD_430_U35 ; P3_ADD_430_U168
g19998 nand P3_ADD_430_U32 P3_REIP_REG_16__SCAN_IN ; P3_ADD_430_U169
g19999 nand P3_ADD_430_U107 P3_ADD_430_U33 ; P3_ADD_430_U170
g20000 nand P3_ADD_430_U30 P3_REIP_REG_15__SCAN_IN ; P3_ADD_430_U171
g20001 nand P3_ADD_430_U106 P3_ADD_430_U31 ; P3_ADD_430_U172
g20002 nand P3_ADD_430_U28 P3_REIP_REG_14__SCAN_IN ; P3_ADD_430_U173
g20003 nand P3_ADD_430_U105 P3_ADD_430_U29 ; P3_ADD_430_U174
g20004 nand P3_ADD_430_U26 P3_REIP_REG_13__SCAN_IN ; P3_ADD_430_U175
g20005 nand P3_ADD_430_U104 P3_ADD_430_U27 ; P3_ADD_430_U176
g20006 nand P3_ADD_430_U24 P3_REIP_REG_12__SCAN_IN ; P3_ADD_430_U177
g20007 nand P3_ADD_430_U103 P3_ADD_430_U25 ; P3_ADD_430_U178
g20008 nand P3_ADD_430_U22 P3_REIP_REG_11__SCAN_IN ; P3_ADD_430_U179
g20009 nand P3_ADD_430_U102 P3_ADD_430_U23 ; P3_ADD_430_U180
g20010 nand P3_ADD_430_U20 P3_REIP_REG_10__SCAN_IN ; P3_ADD_430_U181
g20011 nand P3_ADD_430_U101 P3_ADD_430_U21 ; P3_ADD_430_U182
g20012 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_380_U5
g20013 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_380_U6
g20014 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_380_U7
g20015 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_380_U8
g20016 nand P3_ADD_380_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_380_U9
g20017 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_380_U10
g20018 nand P3_ADD_380_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_380_U11
g20019 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_380_U12
g20020 nand P3_ADD_380_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_380_U13
g20021 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_380_U14
g20022 nand P3_ADD_380_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_380_U15
g20023 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_380_U16
g20024 nand P3_ADD_380_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_380_U17
g20025 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_380_U18
g20026 nand P3_ADD_380_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_380_U19
g20027 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_380_U20
g20028 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_380_U21
g20029 nand P3_ADD_380_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_380_U22
g20030 nand P3_ADD_380_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_380_U23
g20031 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_380_U24
g20032 nand P3_ADD_380_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_380_U25
g20033 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_380_U26
g20034 nand P3_ADD_380_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_380_U27
g20035 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_380_U28
g20036 nand P3_ADD_380_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_380_U29
g20037 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_380_U30
g20038 nand P3_ADD_380_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_380_U31
g20039 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_380_U32
g20040 nand P3_ADD_380_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_380_U33
g20041 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_380_U34
g20042 nand P3_ADD_380_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_380_U35
g20043 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_380_U36
g20044 nand P3_ADD_380_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_380_U37
g20045 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_380_U38
g20046 nand P3_ADD_380_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_380_U39
g20047 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_380_U40
g20048 nand P3_ADD_380_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_380_U41
g20049 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_380_U42
g20050 nand P3_ADD_380_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_380_U43
g20051 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_380_U44
g20052 nand P3_ADD_380_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_380_U45
g20053 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_380_U46
g20054 nand P3_ADD_380_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_380_U47
g20055 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_380_U48
g20056 nand P3_ADD_380_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_380_U49
g20057 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_380_U50
g20058 nand P3_ADD_380_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_380_U51
g20059 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_380_U52
g20060 nand P3_ADD_380_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_380_U53
g20061 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_380_U54
g20062 nand P3_ADD_380_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_380_U55
g20063 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_380_U56
g20064 nand P3_ADD_380_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_380_U57
g20065 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_380_U58
g20066 nand P3_ADD_380_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_380_U59
g20067 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_380_U60
g20068 nand P3_ADD_380_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_380_U61
g20069 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_380_U62
g20070 nand P3_ADD_380_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_380_U63
g20071 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_380_U64
g20072 nand P3_ADD_380_U129 P3_ADD_380_U128 ; P3_ADD_380_U65
g20073 nand P3_ADD_380_U131 P3_ADD_380_U130 ; P3_ADD_380_U66
g20074 nand P3_ADD_380_U133 P3_ADD_380_U132 ; P3_ADD_380_U67
g20075 nand P3_ADD_380_U135 P3_ADD_380_U134 ; P3_ADD_380_U68
g20076 nand P3_ADD_380_U137 P3_ADD_380_U136 ; P3_ADD_380_U69
g20077 nand P3_ADD_380_U139 P3_ADD_380_U138 ; P3_ADD_380_U70
g20078 nand P3_ADD_380_U141 P3_ADD_380_U140 ; P3_ADD_380_U71
g20079 nand P3_ADD_380_U143 P3_ADD_380_U142 ; P3_ADD_380_U72
g20080 nand P3_ADD_380_U145 P3_ADD_380_U144 ; P3_ADD_380_U73
g20081 nand P3_ADD_380_U147 P3_ADD_380_U146 ; P3_ADD_380_U74
g20082 nand P3_ADD_380_U149 P3_ADD_380_U148 ; P3_ADD_380_U75
g20083 nand P3_ADD_380_U151 P3_ADD_380_U150 ; P3_ADD_380_U76
g20084 nand P3_ADD_380_U153 P3_ADD_380_U152 ; P3_ADD_380_U77
g20085 nand P3_ADD_380_U155 P3_ADD_380_U154 ; P3_ADD_380_U78
g20086 nand P3_ADD_380_U157 P3_ADD_380_U156 ; P3_ADD_380_U79
g20087 nand P3_ADD_380_U159 P3_ADD_380_U158 ; P3_ADD_380_U80
g20088 nand P3_ADD_380_U161 P3_ADD_380_U160 ; P3_ADD_380_U81
g20089 nand P3_ADD_380_U163 P3_ADD_380_U162 ; P3_ADD_380_U82
g20090 nand P3_ADD_380_U165 P3_ADD_380_U164 ; P3_ADD_380_U83
g20091 nand P3_ADD_380_U167 P3_ADD_380_U166 ; P3_ADD_380_U84
g20092 nand P3_ADD_380_U169 P3_ADD_380_U168 ; P3_ADD_380_U85
g20093 nand P3_ADD_380_U171 P3_ADD_380_U170 ; P3_ADD_380_U86
g20094 nand P3_ADD_380_U173 P3_ADD_380_U172 ; P3_ADD_380_U87
g20095 nand P3_ADD_380_U175 P3_ADD_380_U174 ; P3_ADD_380_U88
g20096 nand P3_ADD_380_U177 P3_ADD_380_U176 ; P3_ADD_380_U89
g20097 nand P3_ADD_380_U179 P3_ADD_380_U178 ; P3_ADD_380_U90
g20098 nand P3_ADD_380_U181 P3_ADD_380_U180 ; P3_ADD_380_U91
g20099 nand P3_ADD_380_U183 P3_ADD_380_U182 ; P3_ADD_380_U92
g20100 nand P3_ADD_380_U185 P3_ADD_380_U184 ; P3_ADD_380_U93
g20101 nand P3_ADD_380_U187 P3_ADD_380_U186 ; P3_ADD_380_U94
g20102 nand P3_ADD_380_U189 P3_ADD_380_U188 ; P3_ADD_380_U95
g20103 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_380_U96
g20104 nand P3_ADD_380_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_380_U97
g20105 not P3_ADD_380_U7 ; P3_ADD_380_U98
g20106 not P3_ADD_380_U9 ; P3_ADD_380_U99
g20107 not P3_ADD_380_U11 ; P3_ADD_380_U100
g20108 not P3_ADD_380_U13 ; P3_ADD_380_U101
g20109 not P3_ADD_380_U15 ; P3_ADD_380_U102
g20110 not P3_ADD_380_U17 ; P3_ADD_380_U103
g20111 not P3_ADD_380_U19 ; P3_ADD_380_U104
g20112 not P3_ADD_380_U22 ; P3_ADD_380_U105
g20113 not P3_ADD_380_U23 ; P3_ADD_380_U106
g20114 not P3_ADD_380_U25 ; P3_ADD_380_U107
g20115 not P3_ADD_380_U27 ; P3_ADD_380_U108
g20116 not P3_ADD_380_U29 ; P3_ADD_380_U109
g20117 not P3_ADD_380_U31 ; P3_ADD_380_U110
g20118 not P3_ADD_380_U33 ; P3_ADD_380_U111
g20119 not P3_ADD_380_U35 ; P3_ADD_380_U112
g20120 not P3_ADD_380_U37 ; P3_ADD_380_U113
g20121 not P3_ADD_380_U39 ; P3_ADD_380_U114
g20122 not P3_ADD_380_U41 ; P3_ADD_380_U115
g20123 not P3_ADD_380_U43 ; P3_ADD_380_U116
g20124 not P3_ADD_380_U45 ; P3_ADD_380_U117
g20125 not P3_ADD_380_U47 ; P3_ADD_380_U118
g20126 not P3_ADD_380_U49 ; P3_ADD_380_U119
g20127 not P3_ADD_380_U51 ; P3_ADD_380_U120
g20128 not P3_ADD_380_U53 ; P3_ADD_380_U121
g20129 not P3_ADD_380_U55 ; P3_ADD_380_U122
g20130 not P3_ADD_380_U57 ; P3_ADD_380_U123
g20131 not P3_ADD_380_U59 ; P3_ADD_380_U124
g20132 not P3_ADD_380_U61 ; P3_ADD_380_U125
g20133 not P3_ADD_380_U63 ; P3_ADD_380_U126
g20134 not P3_ADD_380_U97 ; P3_ADD_380_U127
g20135 nand P3_ADD_380_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_380_U128
g20136 nand P3_ADD_380_U105 P3_ADD_380_U21 ; P3_ADD_380_U129
g20137 nand P3_ADD_380_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_380_U130
g20138 nand P3_ADD_380_U104 P3_ADD_380_U20 ; P3_ADD_380_U131
g20139 nand P3_ADD_380_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_380_U132
g20140 nand P3_ADD_380_U103 P3_ADD_380_U18 ; P3_ADD_380_U133
g20141 nand P3_ADD_380_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_380_U134
g20142 nand P3_ADD_380_U102 P3_ADD_380_U16 ; P3_ADD_380_U135
g20143 nand P3_ADD_380_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_380_U136
g20144 nand P3_ADD_380_U101 P3_ADD_380_U14 ; P3_ADD_380_U137
g20145 nand P3_ADD_380_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_380_U138
g20146 nand P3_ADD_380_U100 P3_ADD_380_U12 ; P3_ADD_380_U139
g20147 nand P3_ADD_380_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_380_U140
g20148 nand P3_ADD_380_U99 P3_ADD_380_U10 ; P3_ADD_380_U141
g20149 nand P3_ADD_380_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_380_U142
g20150 nand P3_ADD_380_U127 P3_ADD_380_U96 ; P3_ADD_380_U143
g20151 nand P3_ADD_380_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_380_U144
g20152 nand P3_ADD_380_U126 P3_ADD_380_U64 ; P3_ADD_380_U145
g20153 nand P3_ADD_380_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_380_U146
g20154 nand P3_ADD_380_U98 P3_ADD_380_U8 ; P3_ADD_380_U147
g20155 nand P3_ADD_380_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_380_U148
g20156 nand P3_ADD_380_U125 P3_ADD_380_U62 ; P3_ADD_380_U149
g20157 nand P3_ADD_380_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_380_U150
g20158 nand P3_ADD_380_U124 P3_ADD_380_U60 ; P3_ADD_380_U151
g20159 nand P3_ADD_380_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_380_U152
g20160 nand P3_ADD_380_U123 P3_ADD_380_U58 ; P3_ADD_380_U153
g20161 nand P3_ADD_380_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_380_U154
g20162 nand P3_ADD_380_U122 P3_ADD_380_U56 ; P3_ADD_380_U155
g20163 nand P3_ADD_380_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_380_U156
g20164 nand P3_ADD_380_U121 P3_ADD_380_U54 ; P3_ADD_380_U157
g20165 nand P3_ADD_380_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_380_U158
g20166 nand P3_ADD_380_U120 P3_ADD_380_U52 ; P3_ADD_380_U159
g20167 nand P3_ADD_380_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_380_U160
g20168 nand P3_ADD_380_U119 P3_ADD_380_U50 ; P3_ADD_380_U161
g20169 nand P3_ADD_380_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_380_U162
g20170 nand P3_ADD_380_U118 P3_ADD_380_U48 ; P3_ADD_380_U163
g20171 nand P3_ADD_380_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_380_U164
g20172 nand P3_ADD_380_U117 P3_ADD_380_U46 ; P3_ADD_380_U165
g20173 nand P3_ADD_380_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_380_U166
g20174 nand P3_ADD_380_U116 P3_ADD_380_U44 ; P3_ADD_380_U167
g20175 nand P3_ADD_380_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_380_U168
g20176 nand P3_ADD_380_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_380_U169
g20177 nand P3_ADD_380_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_380_U170
g20178 nand P3_ADD_380_U115 P3_ADD_380_U42 ; P3_ADD_380_U171
g20179 nand P3_ADD_380_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_380_U172
g20180 nand P3_ADD_380_U114 P3_ADD_380_U40 ; P3_ADD_380_U173
g20181 nand P3_ADD_380_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_380_U174
g20182 nand P3_ADD_380_U113 P3_ADD_380_U38 ; P3_ADD_380_U175
g20183 nand P3_ADD_380_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_380_U176
g20184 nand P3_ADD_380_U112 P3_ADD_380_U36 ; P3_ADD_380_U177
g20185 nand P3_ADD_380_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_380_U178
g20186 nand P3_ADD_380_U111 P3_ADD_380_U34 ; P3_ADD_380_U179
g20187 nand P3_ADD_380_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_380_U180
g20188 nand P3_ADD_380_U110 P3_ADD_380_U32 ; P3_ADD_380_U181
g20189 nand P3_ADD_380_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_380_U182
g20190 nand P3_ADD_380_U109 P3_ADD_380_U30 ; P3_ADD_380_U183
g20191 nand P3_ADD_380_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_380_U184
g20192 nand P3_ADD_380_U108 P3_ADD_380_U28 ; P3_ADD_380_U185
g20193 nand P3_ADD_380_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_380_U186
g20194 nand P3_ADD_380_U107 P3_ADD_380_U26 ; P3_ADD_380_U187
g20195 nand P3_ADD_380_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_380_U188
g20196 nand P3_ADD_380_U106 P3_ADD_380_U24 ; P3_ADD_380_U189
g20197 nor P3_SUB_370_U6 P3_GTE_370_U8 ; P3_GTE_370_U6
g20198 and P3_SUB_370_U21 P3_GTE_370_U9 ; P3_GTE_370_U7
g20199 nor P3_SUB_370_U19 P3_GTE_370_U7 P3_SUB_370_U20 ; P3_GTE_370_U8
g20200 or P3_SUB_370_U7 P3_SUB_370_U22 ; P3_GTE_370_U9
g20201 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_344_U5
g20202 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_344_U6
g20203 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_344_U7
g20204 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_344_U8
g20205 nand P3_ADD_344_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_344_U9
g20206 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_344_U10
g20207 nand P3_ADD_344_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_344_U11
g20208 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_344_U12
g20209 nand P3_ADD_344_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_344_U13
g20210 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_344_U14
g20211 nand P3_ADD_344_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_344_U15
g20212 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_344_U16
g20213 nand P3_ADD_344_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_344_U17
g20214 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_344_U18
g20215 nand P3_ADD_344_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_344_U19
g20216 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_344_U20
g20217 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_344_U21
g20218 nand P3_ADD_344_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_344_U22
g20219 nand P3_ADD_344_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_344_U23
g20220 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_344_U24
g20221 nand P3_ADD_344_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_344_U25
g20222 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_344_U26
g20223 nand P3_ADD_344_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_344_U27
g20224 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_344_U28
g20225 nand P3_ADD_344_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_344_U29
g20226 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_344_U30
g20227 nand P3_ADD_344_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_344_U31
g20228 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_344_U32
g20229 nand P3_ADD_344_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_344_U33
g20230 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_344_U34
g20231 nand P3_ADD_344_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_344_U35
g20232 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_344_U36
g20233 nand P3_ADD_344_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_344_U37
g20234 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_344_U38
g20235 nand P3_ADD_344_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_344_U39
g20236 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_344_U40
g20237 nand P3_ADD_344_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_344_U41
g20238 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_344_U42
g20239 nand P3_ADD_344_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_344_U43
g20240 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_344_U44
g20241 nand P3_ADD_344_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_344_U45
g20242 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_344_U46
g20243 nand P3_ADD_344_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_344_U47
g20244 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_344_U48
g20245 nand P3_ADD_344_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_344_U49
g20246 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_344_U50
g20247 nand P3_ADD_344_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_344_U51
g20248 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_344_U52
g20249 nand P3_ADD_344_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_344_U53
g20250 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_344_U54
g20251 nand P3_ADD_344_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_344_U55
g20252 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_344_U56
g20253 nand P3_ADD_344_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_344_U57
g20254 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_344_U58
g20255 nand P3_ADD_344_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_344_U59
g20256 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_344_U60
g20257 nand P3_ADD_344_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_344_U61
g20258 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_344_U62
g20259 nand P3_ADD_344_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_344_U63
g20260 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_344_U64
g20261 nand P3_ADD_344_U129 P3_ADD_344_U128 ; P3_ADD_344_U65
g20262 nand P3_ADD_344_U131 P3_ADD_344_U130 ; P3_ADD_344_U66
g20263 nand P3_ADD_344_U133 P3_ADD_344_U132 ; P3_ADD_344_U67
g20264 nand P3_ADD_344_U135 P3_ADD_344_U134 ; P3_ADD_344_U68
g20265 nand P3_ADD_344_U137 P3_ADD_344_U136 ; P3_ADD_344_U69
g20266 nand P3_ADD_344_U139 P3_ADD_344_U138 ; P3_ADD_344_U70
g20267 nand P3_ADD_344_U141 P3_ADD_344_U140 ; P3_ADD_344_U71
g20268 nand P3_ADD_344_U143 P3_ADD_344_U142 ; P3_ADD_344_U72
g20269 nand P3_ADD_344_U145 P3_ADD_344_U144 ; P3_ADD_344_U73
g20270 nand P3_ADD_344_U147 P3_ADD_344_U146 ; P3_ADD_344_U74
g20271 nand P3_ADD_344_U149 P3_ADD_344_U148 ; P3_ADD_344_U75
g20272 nand P3_ADD_344_U151 P3_ADD_344_U150 ; P3_ADD_344_U76
g20273 nand P3_ADD_344_U153 P3_ADD_344_U152 ; P3_ADD_344_U77
g20274 nand P3_ADD_344_U155 P3_ADD_344_U154 ; P3_ADD_344_U78
g20275 nand P3_ADD_344_U157 P3_ADD_344_U156 ; P3_ADD_344_U79
g20276 nand P3_ADD_344_U159 P3_ADD_344_U158 ; P3_ADD_344_U80
g20277 nand P3_ADD_344_U161 P3_ADD_344_U160 ; P3_ADD_344_U81
g20278 nand P3_ADD_344_U163 P3_ADD_344_U162 ; P3_ADD_344_U82
g20279 nand P3_ADD_344_U165 P3_ADD_344_U164 ; P3_ADD_344_U83
g20280 nand P3_ADD_344_U167 P3_ADD_344_U166 ; P3_ADD_344_U84
g20281 nand P3_ADD_344_U169 P3_ADD_344_U168 ; P3_ADD_344_U85
g20282 nand P3_ADD_344_U171 P3_ADD_344_U170 ; P3_ADD_344_U86
g20283 nand P3_ADD_344_U173 P3_ADD_344_U172 ; P3_ADD_344_U87
g20284 nand P3_ADD_344_U175 P3_ADD_344_U174 ; P3_ADD_344_U88
g20285 nand P3_ADD_344_U177 P3_ADD_344_U176 ; P3_ADD_344_U89
g20286 nand P3_ADD_344_U179 P3_ADD_344_U178 ; P3_ADD_344_U90
g20287 nand P3_ADD_344_U181 P3_ADD_344_U180 ; P3_ADD_344_U91
g20288 nand P3_ADD_344_U183 P3_ADD_344_U182 ; P3_ADD_344_U92
g20289 nand P3_ADD_344_U185 P3_ADD_344_U184 ; P3_ADD_344_U93
g20290 nand P3_ADD_344_U187 P3_ADD_344_U186 ; P3_ADD_344_U94
g20291 nand P3_ADD_344_U189 P3_ADD_344_U188 ; P3_ADD_344_U95
g20292 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_344_U96
g20293 nand P3_ADD_344_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_344_U97
g20294 not P3_ADD_344_U7 ; P3_ADD_344_U98
g20295 not P3_ADD_344_U9 ; P3_ADD_344_U99
g20296 not P3_ADD_344_U11 ; P3_ADD_344_U100
g20297 not P3_ADD_344_U13 ; P3_ADD_344_U101
g20298 not P3_ADD_344_U15 ; P3_ADD_344_U102
g20299 not P3_ADD_344_U17 ; P3_ADD_344_U103
g20300 not P3_ADD_344_U19 ; P3_ADD_344_U104
g20301 not P3_ADD_344_U22 ; P3_ADD_344_U105
g20302 not P3_ADD_344_U23 ; P3_ADD_344_U106
g20303 not P3_ADD_344_U25 ; P3_ADD_344_U107
g20304 not P3_ADD_344_U27 ; P3_ADD_344_U108
g20305 not P3_ADD_344_U29 ; P3_ADD_344_U109
g20306 not P3_ADD_344_U31 ; P3_ADD_344_U110
g20307 not P3_ADD_344_U33 ; P3_ADD_344_U111
g20308 not P3_ADD_344_U35 ; P3_ADD_344_U112
g20309 not P3_ADD_344_U37 ; P3_ADD_344_U113
g20310 not P3_ADD_344_U39 ; P3_ADD_344_U114
g20311 not P3_ADD_344_U41 ; P3_ADD_344_U115
g20312 not P3_ADD_344_U43 ; P3_ADD_344_U116
g20313 not P3_ADD_344_U45 ; P3_ADD_344_U117
g20314 not P3_ADD_344_U47 ; P3_ADD_344_U118
g20315 not P3_ADD_344_U49 ; P3_ADD_344_U119
g20316 not P3_ADD_344_U51 ; P3_ADD_344_U120
g20317 not P3_ADD_344_U53 ; P3_ADD_344_U121
g20318 not P3_ADD_344_U55 ; P3_ADD_344_U122
g20319 not P3_ADD_344_U57 ; P3_ADD_344_U123
g20320 not P3_ADD_344_U59 ; P3_ADD_344_U124
g20321 not P3_ADD_344_U61 ; P3_ADD_344_U125
g20322 not P3_ADD_344_U63 ; P3_ADD_344_U126
g20323 not P3_ADD_344_U97 ; P3_ADD_344_U127
g20324 nand P3_ADD_344_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_344_U128
g20325 nand P3_ADD_344_U105 P3_ADD_344_U21 ; P3_ADD_344_U129
g20326 nand P3_ADD_344_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_344_U130
g20327 nand P3_ADD_344_U104 P3_ADD_344_U20 ; P3_ADD_344_U131
g20328 nand P3_ADD_344_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_344_U132
g20329 nand P3_ADD_344_U103 P3_ADD_344_U18 ; P3_ADD_344_U133
g20330 nand P3_ADD_344_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_344_U134
g20331 nand P3_ADD_344_U102 P3_ADD_344_U16 ; P3_ADD_344_U135
g20332 nand P3_ADD_344_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_344_U136
g20333 nand P3_ADD_344_U101 P3_ADD_344_U14 ; P3_ADD_344_U137
g20334 nand P3_ADD_344_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_344_U138
g20335 nand P3_ADD_344_U100 P3_ADD_344_U12 ; P3_ADD_344_U139
g20336 nand P3_ADD_344_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_344_U140
g20337 nand P3_ADD_344_U99 P3_ADD_344_U10 ; P3_ADD_344_U141
g20338 nand P3_ADD_344_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_344_U142
g20339 nand P3_ADD_344_U127 P3_ADD_344_U96 ; P3_ADD_344_U143
g20340 nand P3_ADD_344_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_344_U144
g20341 nand P3_ADD_344_U126 P3_ADD_344_U64 ; P3_ADD_344_U145
g20342 nand P3_ADD_344_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_344_U146
g20343 nand P3_ADD_344_U98 P3_ADD_344_U8 ; P3_ADD_344_U147
g20344 nand P3_ADD_344_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_344_U148
g20345 nand P3_ADD_344_U125 P3_ADD_344_U62 ; P3_ADD_344_U149
g20346 nand P3_ADD_344_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_344_U150
g20347 nand P3_ADD_344_U124 P3_ADD_344_U60 ; P3_ADD_344_U151
g20348 nand P3_ADD_344_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_344_U152
g20349 nand P3_ADD_344_U123 P3_ADD_344_U58 ; P3_ADD_344_U153
g20350 nand P3_ADD_344_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_344_U154
g20351 nand P3_ADD_344_U122 P3_ADD_344_U56 ; P3_ADD_344_U155
g20352 nand P3_ADD_344_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_344_U156
g20353 nand P3_ADD_344_U121 P3_ADD_344_U54 ; P3_ADD_344_U157
g20354 nand P3_ADD_344_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_344_U158
g20355 nand P3_ADD_344_U120 P3_ADD_344_U52 ; P3_ADD_344_U159
g20356 nand P3_ADD_344_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_344_U160
g20357 nand P3_ADD_344_U119 P3_ADD_344_U50 ; P3_ADD_344_U161
g20358 nand P3_ADD_344_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_344_U162
g20359 nand P3_ADD_344_U118 P3_ADD_344_U48 ; P3_ADD_344_U163
g20360 nand P3_ADD_344_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_344_U164
g20361 nand P3_ADD_344_U117 P3_ADD_344_U46 ; P3_ADD_344_U165
g20362 nand P3_ADD_344_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_344_U166
g20363 nand P3_ADD_344_U116 P3_ADD_344_U44 ; P3_ADD_344_U167
g20364 nand P3_ADD_344_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_344_U168
g20365 nand P3_ADD_344_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_344_U169
g20366 nand P3_ADD_344_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_344_U170
g20367 nand P3_ADD_344_U115 P3_ADD_344_U42 ; P3_ADD_344_U171
g20368 nand P3_ADD_344_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_344_U172
g20369 nand P3_ADD_344_U114 P3_ADD_344_U40 ; P3_ADD_344_U173
g20370 nand P3_ADD_344_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_344_U174
g20371 nand P3_ADD_344_U113 P3_ADD_344_U38 ; P3_ADD_344_U175
g20372 nand P3_ADD_344_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_344_U176
g20373 nand P3_ADD_344_U112 P3_ADD_344_U36 ; P3_ADD_344_U177
g20374 nand P3_ADD_344_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_344_U178
g20375 nand P3_ADD_344_U111 P3_ADD_344_U34 ; P3_ADD_344_U179
g20376 nand P3_ADD_344_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_344_U180
g20377 nand P3_ADD_344_U110 P3_ADD_344_U32 ; P3_ADD_344_U181
g20378 nand P3_ADD_344_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_344_U182
g20379 nand P3_ADD_344_U109 P3_ADD_344_U30 ; P3_ADD_344_U183
g20380 nand P3_ADD_344_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_344_U184
g20381 nand P3_ADD_344_U108 P3_ADD_344_U28 ; P3_ADD_344_U185
g20382 nand P3_ADD_344_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_344_U186
g20383 nand P3_ADD_344_U107 P3_ADD_344_U26 ; P3_ADD_344_U187
g20384 nand P3_ADD_344_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_344_U188
g20385 nand P3_ADD_344_U106 P3_ADD_344_U24 ; P3_ADD_344_U189
g20386 nand P3_LT_563_U27 P3_LT_563_U28 ; P3_LT_563_U6
g20387 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_LT_563_U7
g20388 nand P3_LT_563_U15 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_LT_563_U8
g20389 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_LT_563_U9
g20390 not P3_U3306 ; P3_LT_563_U10
g20391 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_LT_563_U11
g20392 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_LT_563_U12
g20393 not P3_U3305 ; P3_LT_563_U13
g20394 not P3_U3304 ; P3_LT_563_U14
g20395 not P3_U3308 ; P3_LT_563_U15
g20396 not P3_LT_563_U8 ; P3_LT_563_U16
g20397 nand P3_LT_563_U16 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_LT_563_U17
g20398 nand P3_U3307 P3_LT_563_U17 ; P3_LT_563_U18
g20399 nand P3_LT_563_U8 P3_LT_563_U9 ; P3_LT_563_U19
g20400 nand P3_U3306 P3_LT_563_U11 ; P3_LT_563_U20
g20401 nand P3_LT_563_U19 P3_LT_563_U20 P3_LT_563_U18 ; P3_LT_563_U21
g20402 nand P3_LT_563_U10 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_LT_563_U22
g20403 nand P3_LT_563_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_LT_563_U23
g20404 nand P3_LT_563_U22 P3_LT_563_U23 P3_LT_563_U21 ; P3_LT_563_U24
g20405 nand P3_U3305 P3_LT_563_U12 ; P3_LT_563_U25
g20406 nand P3_U3304 P3_LT_563_U7 ; P3_LT_563_U26
g20407 nand P3_LT_563_U25 P3_LT_563_U26 P3_LT_563_U24 ; P3_LT_563_U27
g20408 nand P3_LT_563_U14 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_LT_563_U28
g20409 not P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_339_U4
g20410 not P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_339_U5
g20411 nand P3_PHYADDRPOINTER_REG_1__SCAN_IN P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_339_U6
g20412 not P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_339_U7
g20413 nand P3_ADD_339_U94 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_339_U8
g20414 not P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_339_U9
g20415 nand P3_ADD_339_U95 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_339_U10
g20416 not P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_339_U11
g20417 nand P3_ADD_339_U96 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_339_U12
g20418 not P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_339_U13
g20419 nand P3_ADD_339_U97 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_339_U14
g20420 not P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_339_U15
g20421 nand P3_ADD_339_U98 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_339_U16
g20422 not P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_339_U17
g20423 not P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_339_U18
g20424 nand P3_ADD_339_U99 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_339_U19
g20425 nand P3_ADD_339_U100 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_339_U20
g20426 not P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_339_U21
g20427 nand P3_ADD_339_U101 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_339_U22
g20428 not P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_339_U23
g20429 nand P3_ADD_339_U102 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_339_U24
g20430 not P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_339_U25
g20431 nand P3_ADD_339_U103 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_339_U26
g20432 not P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_339_U27
g20433 nand P3_ADD_339_U104 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_339_U28
g20434 not P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_339_U29
g20435 nand P3_ADD_339_U105 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_339_U30
g20436 not P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_339_U31
g20437 nand P3_ADD_339_U106 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_339_U32
g20438 not P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_339_U33
g20439 nand P3_ADD_339_U107 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_339_U34
g20440 not P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_339_U35
g20441 nand P3_ADD_339_U108 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_339_U36
g20442 not P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_339_U37
g20443 nand P3_ADD_339_U109 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_339_U38
g20444 not P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_339_U39
g20445 nand P3_ADD_339_U110 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_339_U40
g20446 not P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_339_U41
g20447 nand P3_ADD_339_U111 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_339_U42
g20448 not P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_339_U43
g20449 nand P3_ADD_339_U112 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_339_U44
g20450 not P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_339_U45
g20451 nand P3_ADD_339_U113 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_339_U46
g20452 not P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_339_U47
g20453 nand P3_ADD_339_U114 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_339_U48
g20454 not P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_339_U49
g20455 nand P3_ADD_339_U115 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_339_U50
g20456 not P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_339_U51
g20457 nand P3_ADD_339_U116 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_339_U52
g20458 not P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_339_U53
g20459 nand P3_ADD_339_U117 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_339_U54
g20460 not P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_339_U55
g20461 nand P3_ADD_339_U118 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_339_U56
g20462 not P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_339_U57
g20463 nand P3_ADD_339_U119 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_339_U58
g20464 not P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_339_U59
g20465 nand P3_ADD_339_U120 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_339_U60
g20466 not P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_339_U61
g20467 nand P3_ADD_339_U124 P3_ADD_339_U123 ; P3_ADD_339_U62
g20468 nand P3_ADD_339_U126 P3_ADD_339_U125 ; P3_ADD_339_U63
g20469 nand P3_ADD_339_U128 P3_ADD_339_U127 ; P3_ADD_339_U64
g20470 nand P3_ADD_339_U130 P3_ADD_339_U129 ; P3_ADD_339_U65
g20471 nand P3_ADD_339_U132 P3_ADD_339_U131 ; P3_ADD_339_U66
g20472 nand P3_ADD_339_U134 P3_ADD_339_U133 ; P3_ADD_339_U67
g20473 nand P3_ADD_339_U136 P3_ADD_339_U135 ; P3_ADD_339_U68
g20474 nand P3_ADD_339_U138 P3_ADD_339_U137 ; P3_ADD_339_U69
g20475 nand P3_ADD_339_U140 P3_ADD_339_U139 ; P3_ADD_339_U70
g20476 nand P3_ADD_339_U142 P3_ADD_339_U141 ; P3_ADD_339_U71
g20477 nand P3_ADD_339_U144 P3_ADD_339_U143 ; P3_ADD_339_U72
g20478 nand P3_ADD_339_U146 P3_ADD_339_U145 ; P3_ADD_339_U73
g20479 nand P3_ADD_339_U148 P3_ADD_339_U147 ; P3_ADD_339_U74
g20480 nand P3_ADD_339_U150 P3_ADD_339_U149 ; P3_ADD_339_U75
g20481 nand P3_ADD_339_U152 P3_ADD_339_U151 ; P3_ADD_339_U76
g20482 nand P3_ADD_339_U154 P3_ADD_339_U153 ; P3_ADD_339_U77
g20483 nand P3_ADD_339_U156 P3_ADD_339_U155 ; P3_ADD_339_U78
g20484 nand P3_ADD_339_U158 P3_ADD_339_U157 ; P3_ADD_339_U79
g20485 nand P3_ADD_339_U160 P3_ADD_339_U159 ; P3_ADD_339_U80
g20486 nand P3_ADD_339_U162 P3_ADD_339_U161 ; P3_ADD_339_U81
g20487 nand P3_ADD_339_U164 P3_ADD_339_U163 ; P3_ADD_339_U82
g20488 nand P3_ADD_339_U166 P3_ADD_339_U165 ; P3_ADD_339_U83
g20489 nand P3_ADD_339_U168 P3_ADD_339_U167 ; P3_ADD_339_U84
g20490 nand P3_ADD_339_U170 P3_ADD_339_U169 ; P3_ADD_339_U85
g20491 nand P3_ADD_339_U172 P3_ADD_339_U171 ; P3_ADD_339_U86
g20492 nand P3_ADD_339_U174 P3_ADD_339_U173 ; P3_ADD_339_U87
g20493 nand P3_ADD_339_U176 P3_ADD_339_U175 ; P3_ADD_339_U88
g20494 nand P3_ADD_339_U178 P3_ADD_339_U177 ; P3_ADD_339_U89
g20495 nand P3_ADD_339_U180 P3_ADD_339_U179 ; P3_ADD_339_U90
g20496 nand P3_ADD_339_U182 P3_ADD_339_U181 ; P3_ADD_339_U91
g20497 not P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_339_U92
g20498 nand P3_ADD_339_U121 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_339_U93
g20499 not P3_ADD_339_U6 ; P3_ADD_339_U94
g20500 not P3_ADD_339_U8 ; P3_ADD_339_U95
g20501 not P3_ADD_339_U10 ; P3_ADD_339_U96
g20502 not P3_ADD_339_U12 ; P3_ADD_339_U97
g20503 not P3_ADD_339_U14 ; P3_ADD_339_U98
g20504 not P3_ADD_339_U16 ; P3_ADD_339_U99
g20505 not P3_ADD_339_U19 ; P3_ADD_339_U100
g20506 not P3_ADD_339_U20 ; P3_ADD_339_U101
g20507 not P3_ADD_339_U22 ; P3_ADD_339_U102
g20508 not P3_ADD_339_U24 ; P3_ADD_339_U103
g20509 not P3_ADD_339_U26 ; P3_ADD_339_U104
g20510 not P3_ADD_339_U28 ; P3_ADD_339_U105
g20511 not P3_ADD_339_U30 ; P3_ADD_339_U106
g20512 not P3_ADD_339_U32 ; P3_ADD_339_U107
g20513 not P3_ADD_339_U34 ; P3_ADD_339_U108
g20514 not P3_ADD_339_U36 ; P3_ADD_339_U109
g20515 not P3_ADD_339_U38 ; P3_ADD_339_U110
g20516 not P3_ADD_339_U40 ; P3_ADD_339_U111
g20517 not P3_ADD_339_U42 ; P3_ADD_339_U112
g20518 not P3_ADD_339_U44 ; P3_ADD_339_U113
g20519 not P3_ADD_339_U46 ; P3_ADD_339_U114
g20520 not P3_ADD_339_U48 ; P3_ADD_339_U115
g20521 not P3_ADD_339_U50 ; P3_ADD_339_U116
g20522 not P3_ADD_339_U52 ; P3_ADD_339_U117
g20523 not P3_ADD_339_U54 ; P3_ADD_339_U118
g20524 not P3_ADD_339_U56 ; P3_ADD_339_U119
g20525 not P3_ADD_339_U58 ; P3_ADD_339_U120
g20526 not P3_ADD_339_U60 ; P3_ADD_339_U121
g20527 not P3_ADD_339_U93 ; P3_ADD_339_U122
g20528 nand P3_ADD_339_U19 P3_PHYADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_339_U123
g20529 nand P3_ADD_339_U100 P3_ADD_339_U18 ; P3_ADD_339_U124
g20530 nand P3_ADD_339_U16 P3_PHYADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_339_U125
g20531 nand P3_ADD_339_U99 P3_ADD_339_U17 ; P3_ADD_339_U126
g20532 nand P3_ADD_339_U14 P3_PHYADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_339_U127
g20533 nand P3_ADD_339_U98 P3_ADD_339_U15 ; P3_ADD_339_U128
g20534 nand P3_ADD_339_U12 P3_PHYADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_339_U129
g20535 nand P3_ADD_339_U97 P3_ADD_339_U13 ; P3_ADD_339_U130
g20536 nand P3_ADD_339_U10 P3_PHYADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_339_U131
g20537 nand P3_ADD_339_U96 P3_ADD_339_U11 ; P3_ADD_339_U132
g20538 nand P3_ADD_339_U8 P3_PHYADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_339_U133
g20539 nand P3_ADD_339_U95 P3_ADD_339_U9 ; P3_ADD_339_U134
g20540 nand P3_ADD_339_U6 P3_PHYADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_339_U135
g20541 nand P3_ADD_339_U94 P3_ADD_339_U7 ; P3_ADD_339_U136
g20542 nand P3_ADD_339_U93 P3_PHYADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_339_U137
g20543 nand P3_ADD_339_U122 P3_ADD_339_U92 ; P3_ADD_339_U138
g20544 nand P3_ADD_339_U60 P3_PHYADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_339_U139
g20545 nand P3_ADD_339_U121 P3_ADD_339_U61 ; P3_ADD_339_U140
g20546 nand P3_ADD_339_U4 P3_PHYADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_339_U141
g20547 nand P3_ADD_339_U5 P3_PHYADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_339_U142
g20548 nand P3_ADD_339_U58 P3_PHYADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_339_U143
g20549 nand P3_ADD_339_U120 P3_ADD_339_U59 ; P3_ADD_339_U144
g20550 nand P3_ADD_339_U56 P3_PHYADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_339_U145
g20551 nand P3_ADD_339_U119 P3_ADD_339_U57 ; P3_ADD_339_U146
g20552 nand P3_ADD_339_U54 P3_PHYADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_339_U147
g20553 nand P3_ADD_339_U118 P3_ADD_339_U55 ; P3_ADD_339_U148
g20554 nand P3_ADD_339_U52 P3_PHYADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_339_U149
g20555 nand P3_ADD_339_U117 P3_ADD_339_U53 ; P3_ADD_339_U150
g20556 nand P3_ADD_339_U50 P3_PHYADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_339_U151
g20557 nand P3_ADD_339_U116 P3_ADD_339_U51 ; P3_ADD_339_U152
g20558 nand P3_ADD_339_U48 P3_PHYADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_339_U153
g20559 nand P3_ADD_339_U115 P3_ADD_339_U49 ; P3_ADD_339_U154
g20560 nand P3_ADD_339_U46 P3_PHYADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_339_U155
g20561 nand P3_ADD_339_U114 P3_ADD_339_U47 ; P3_ADD_339_U156
g20562 nand P3_ADD_339_U44 P3_PHYADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_339_U157
g20563 nand P3_ADD_339_U113 P3_ADD_339_U45 ; P3_ADD_339_U158
g20564 nand P3_ADD_339_U42 P3_PHYADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_339_U159
g20565 nand P3_ADD_339_U112 P3_ADD_339_U43 ; P3_ADD_339_U160
g20566 nand P3_ADD_339_U40 P3_PHYADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_339_U161
g20567 nand P3_ADD_339_U111 P3_ADD_339_U41 ; P3_ADD_339_U162
g20568 nand P3_ADD_339_U38 P3_PHYADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_339_U163
g20569 nand P3_ADD_339_U110 P3_ADD_339_U39 ; P3_ADD_339_U164
g20570 nand P3_ADD_339_U36 P3_PHYADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_339_U165
g20571 nand P3_ADD_339_U109 P3_ADD_339_U37 ; P3_ADD_339_U166
g20572 nand P3_ADD_339_U34 P3_PHYADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_339_U167
g20573 nand P3_ADD_339_U108 P3_ADD_339_U35 ; P3_ADD_339_U168
g20574 nand P3_ADD_339_U32 P3_PHYADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_339_U169
g20575 nand P3_ADD_339_U107 P3_ADD_339_U33 ; P3_ADD_339_U170
g20576 nand P3_ADD_339_U30 P3_PHYADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_339_U171
g20577 nand P3_ADD_339_U106 P3_ADD_339_U31 ; P3_ADD_339_U172
g20578 nand P3_ADD_339_U28 P3_PHYADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_339_U173
g20579 nand P3_ADD_339_U105 P3_ADD_339_U29 ; P3_ADD_339_U174
g20580 nand P3_ADD_339_U26 P3_PHYADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_339_U175
g20581 nand P3_ADD_339_U104 P3_ADD_339_U27 ; P3_ADD_339_U176
g20582 nand P3_ADD_339_U24 P3_PHYADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_339_U177
g20583 nand P3_ADD_339_U103 P3_ADD_339_U25 ; P3_ADD_339_U178
g20584 nand P3_ADD_339_U22 P3_PHYADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_339_U179
g20585 nand P3_ADD_339_U102 P3_ADD_339_U23 ; P3_ADD_339_U180
g20586 nand P3_ADD_339_U20 P3_PHYADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_339_U181
g20587 nand P3_ADD_339_U101 P3_ADD_339_U21 ; P3_ADD_339_U182
g20588 not P3_U2622 ; P3_ADD_360_U4
g20589 and P3_ADD_360_U22 P3_ADD_360_U27 ; P3_ADD_360_U5
g20590 not P3_U2623 ; P3_ADD_360_U6
g20591 nand P3_U2623 P3_U2622 ; P3_ADD_360_U7
g20592 not P3_U2624 ; P3_ADD_360_U8
g20593 nand P3_U2624 P3_ADD_360_U24 ; P3_ADD_360_U9
g20594 not P3_U2625 ; P3_ADD_360_U10
g20595 nand P3_U2625 P3_ADD_360_U25 ; P3_ADD_360_U11
g20596 not P3_U2626 ; P3_ADD_360_U12
g20597 nand P3_U2626 P3_ADD_360_U26 ; P3_ADD_360_U13
g20598 not P3_U2628 ; P3_ADD_360_U14
g20599 not P3_U2627 ; P3_ADD_360_U15
g20600 nand P3_ADD_360_U30 P3_ADD_360_U29 ; P3_ADD_360_U16
g20601 nand P3_ADD_360_U32 P3_ADD_360_U31 ; P3_ADD_360_U17
g20602 nand P3_ADD_360_U34 P3_ADD_360_U33 ; P3_ADD_360_U18
g20603 nand P3_ADD_360_U36 P3_ADD_360_U35 ; P3_ADD_360_U19
g20604 nand P3_ADD_360_U38 P3_ADD_360_U37 ; P3_ADD_360_U20
g20605 nand P3_ADD_360_U40 P3_ADD_360_U39 ; P3_ADD_360_U21
g20606 and P3_U2628 P3_U2627 ; P3_ADD_360_U22
g20607 nand P3_U2627 P3_ADD_360_U27 ; P3_ADD_360_U23
g20608 not P3_ADD_360_U7 ; P3_ADD_360_U24
g20609 not P3_ADD_360_U9 ; P3_ADD_360_U25
g20610 not P3_ADD_360_U11 ; P3_ADD_360_U26
g20611 not P3_ADD_360_U13 ; P3_ADD_360_U27
g20612 not P3_ADD_360_U23 ; P3_ADD_360_U28
g20613 nand P3_U2628 P3_ADD_360_U23 ; P3_ADD_360_U29
g20614 nand P3_ADD_360_U28 P3_ADD_360_U14 ; P3_ADD_360_U30
g20615 nand P3_U2627 P3_ADD_360_U13 ; P3_ADD_360_U31
g20616 nand P3_ADD_360_U27 P3_ADD_360_U15 ; P3_ADD_360_U32
g20617 nand P3_U2626 P3_ADD_360_U11 ; P3_ADD_360_U33
g20618 nand P3_ADD_360_U26 P3_ADD_360_U12 ; P3_ADD_360_U34
g20619 nand P3_U2625 P3_ADD_360_U9 ; P3_ADD_360_U35
g20620 nand P3_ADD_360_U25 P3_ADD_360_U10 ; P3_ADD_360_U36
g20621 nand P3_U2624 P3_ADD_360_U7 ; P3_ADD_360_U37
g20622 nand P3_ADD_360_U24 P3_ADD_360_U8 ; P3_ADD_360_U38
g20623 nand P3_U2623 P3_ADD_360_U4 ; P3_ADD_360_U39
g20624 nand P3_U2622 P3_ADD_360_U6 ; P3_ADD_360_U40
g20625 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_LTE_597_U6
g20626 nand P3_SUB_580_U10 P3_SUB_580_U9 ; P3_SUB_580_U6
g20627 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_580_U7
g20628 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_580_U8
g20629 nand P3_SUB_580_U8 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_580_U9
g20630 nand P3_SUB_580_U7 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_580_U10
g20631 or P3_LT_589_U8 P3_U2629 ; P3_LT_589_U6
g20632 and P3_SUB_589_U7 P3_SUB_589_U6 ; P3_LT_589_U7
g20633 nor P3_LT_589_U7 P3_SUB_589_U8 P3_SUB_589_U9 ; P3_LT_589_U8
g20634 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_541_U4
g20635 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_541_U5
g20636 nand P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_541_U6
g20637 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_541_U7
g20638 nand P3_ADD_541_U94 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_541_U8
g20639 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_541_U9
g20640 nand P3_ADD_541_U95 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_541_U10
g20641 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_541_U11
g20642 nand P3_ADD_541_U96 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_541_U12
g20643 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_541_U13
g20644 nand P3_ADD_541_U97 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_541_U14
g20645 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_541_U15
g20646 nand P3_ADD_541_U98 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_541_U16
g20647 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_541_U17
g20648 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_541_U18
g20649 nand P3_ADD_541_U99 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_541_U19
g20650 nand P3_ADD_541_U100 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_541_U20
g20651 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_541_U21
g20652 nand P3_ADD_541_U101 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_541_U22
g20653 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_541_U23
g20654 nand P3_ADD_541_U102 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_541_U24
g20655 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_541_U25
g20656 nand P3_ADD_541_U103 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_541_U26
g20657 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_541_U27
g20658 nand P3_ADD_541_U104 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_541_U28
g20659 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_541_U29
g20660 nand P3_ADD_541_U105 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_541_U30
g20661 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_541_U31
g20662 nand P3_ADD_541_U106 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_541_U32
g20663 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_541_U33
g20664 nand P3_ADD_541_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_541_U34
g20665 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_541_U35
g20666 nand P3_ADD_541_U108 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_541_U36
g20667 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_541_U37
g20668 nand P3_ADD_541_U109 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_541_U38
g20669 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_541_U39
g20670 nand P3_ADD_541_U110 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_541_U40
g20671 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_541_U41
g20672 nand P3_ADD_541_U111 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_541_U42
g20673 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_541_U43
g20674 nand P3_ADD_541_U112 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_541_U44
g20675 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_541_U45
g20676 nand P3_ADD_541_U113 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_541_U46
g20677 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_541_U47
g20678 nand P3_ADD_541_U114 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_541_U48
g20679 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_541_U49
g20680 nand P3_ADD_541_U115 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_541_U50
g20681 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_541_U51
g20682 nand P3_ADD_541_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_541_U52
g20683 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_541_U53
g20684 nand P3_ADD_541_U117 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_541_U54
g20685 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_541_U55
g20686 nand P3_ADD_541_U118 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_541_U56
g20687 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_541_U57
g20688 nand P3_ADD_541_U119 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_541_U58
g20689 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_541_U59
g20690 nand P3_ADD_541_U120 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_541_U60
g20691 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_541_U61
g20692 nand P3_ADD_541_U124 P3_ADD_541_U123 ; P3_ADD_541_U62
g20693 nand P3_ADD_541_U126 P3_ADD_541_U125 ; P3_ADD_541_U63
g20694 nand P3_ADD_541_U128 P3_ADD_541_U127 ; P3_ADD_541_U64
g20695 nand P3_ADD_541_U130 P3_ADD_541_U129 ; P3_ADD_541_U65
g20696 nand P3_ADD_541_U132 P3_ADD_541_U131 ; P3_ADD_541_U66
g20697 nand P3_ADD_541_U134 P3_ADD_541_U133 ; P3_ADD_541_U67
g20698 nand P3_ADD_541_U136 P3_ADD_541_U135 ; P3_ADD_541_U68
g20699 nand P3_ADD_541_U138 P3_ADD_541_U137 ; P3_ADD_541_U69
g20700 nand P3_ADD_541_U140 P3_ADD_541_U139 ; P3_ADD_541_U70
g20701 nand P3_ADD_541_U142 P3_ADD_541_U141 ; P3_ADD_541_U71
g20702 nand P3_ADD_541_U144 P3_ADD_541_U143 ; P3_ADD_541_U72
g20703 nand P3_ADD_541_U146 P3_ADD_541_U145 ; P3_ADD_541_U73
g20704 nand P3_ADD_541_U148 P3_ADD_541_U147 ; P3_ADD_541_U74
g20705 nand P3_ADD_541_U150 P3_ADD_541_U149 ; P3_ADD_541_U75
g20706 nand P3_ADD_541_U152 P3_ADD_541_U151 ; P3_ADD_541_U76
g20707 nand P3_ADD_541_U154 P3_ADD_541_U153 ; P3_ADD_541_U77
g20708 nand P3_ADD_541_U156 P3_ADD_541_U155 ; P3_ADD_541_U78
g20709 nand P3_ADD_541_U158 P3_ADD_541_U157 ; P3_ADD_541_U79
g20710 nand P3_ADD_541_U160 P3_ADD_541_U159 ; P3_ADD_541_U80
g20711 nand P3_ADD_541_U162 P3_ADD_541_U161 ; P3_ADD_541_U81
g20712 nand P3_ADD_541_U164 P3_ADD_541_U163 ; P3_ADD_541_U82
g20713 nand P3_ADD_541_U166 P3_ADD_541_U165 ; P3_ADD_541_U83
g20714 nand P3_ADD_541_U168 P3_ADD_541_U167 ; P3_ADD_541_U84
g20715 nand P3_ADD_541_U170 P3_ADD_541_U169 ; P3_ADD_541_U85
g20716 nand P3_ADD_541_U172 P3_ADD_541_U171 ; P3_ADD_541_U86
g20717 nand P3_ADD_541_U174 P3_ADD_541_U173 ; P3_ADD_541_U87
g20718 nand P3_ADD_541_U176 P3_ADD_541_U175 ; P3_ADD_541_U88
g20719 nand P3_ADD_541_U178 P3_ADD_541_U177 ; P3_ADD_541_U89
g20720 nand P3_ADD_541_U180 P3_ADD_541_U179 ; P3_ADD_541_U90
g20721 nand P3_ADD_541_U182 P3_ADD_541_U181 ; P3_ADD_541_U91
g20722 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_541_U92
g20723 nand P3_ADD_541_U121 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_541_U93
g20724 not P3_ADD_541_U6 ; P3_ADD_541_U94
g20725 not P3_ADD_541_U8 ; P3_ADD_541_U95
g20726 not P3_ADD_541_U10 ; P3_ADD_541_U96
g20727 not P3_ADD_541_U12 ; P3_ADD_541_U97
g20728 not P3_ADD_541_U14 ; P3_ADD_541_U98
g20729 not P3_ADD_541_U16 ; P3_ADD_541_U99
g20730 not P3_ADD_541_U19 ; P3_ADD_541_U100
g20731 not P3_ADD_541_U20 ; P3_ADD_541_U101
g20732 not P3_ADD_541_U22 ; P3_ADD_541_U102
g20733 not P3_ADD_541_U24 ; P3_ADD_541_U103
g20734 not P3_ADD_541_U26 ; P3_ADD_541_U104
g20735 not P3_ADD_541_U28 ; P3_ADD_541_U105
g20736 not P3_ADD_541_U30 ; P3_ADD_541_U106
g20737 not P3_ADD_541_U32 ; P3_ADD_541_U107
g20738 not P3_ADD_541_U34 ; P3_ADD_541_U108
g20739 not P3_ADD_541_U36 ; P3_ADD_541_U109
g20740 not P3_ADD_541_U38 ; P3_ADD_541_U110
g20741 not P3_ADD_541_U40 ; P3_ADD_541_U111
g20742 not P3_ADD_541_U42 ; P3_ADD_541_U112
g20743 not P3_ADD_541_U44 ; P3_ADD_541_U113
g20744 not P3_ADD_541_U46 ; P3_ADD_541_U114
g20745 not P3_ADD_541_U48 ; P3_ADD_541_U115
g20746 not P3_ADD_541_U50 ; P3_ADD_541_U116
g20747 not P3_ADD_541_U52 ; P3_ADD_541_U117
g20748 not P3_ADD_541_U54 ; P3_ADD_541_U118
g20749 not P3_ADD_541_U56 ; P3_ADD_541_U119
g20750 not P3_ADD_541_U58 ; P3_ADD_541_U120
g20751 not P3_ADD_541_U60 ; P3_ADD_541_U121
g20752 not P3_ADD_541_U93 ; P3_ADD_541_U122
g20753 nand P3_ADD_541_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_541_U123
g20754 nand P3_ADD_541_U100 P3_ADD_541_U18 ; P3_ADD_541_U124
g20755 nand P3_ADD_541_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_541_U125
g20756 nand P3_ADD_541_U99 P3_ADD_541_U17 ; P3_ADD_541_U126
g20757 nand P3_ADD_541_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_541_U127
g20758 nand P3_ADD_541_U98 P3_ADD_541_U15 ; P3_ADD_541_U128
g20759 nand P3_ADD_541_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_541_U129
g20760 nand P3_ADD_541_U97 P3_ADD_541_U13 ; P3_ADD_541_U130
g20761 nand P3_ADD_541_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_541_U131
g20762 nand P3_ADD_541_U96 P3_ADD_541_U11 ; P3_ADD_541_U132
g20763 nand P3_ADD_541_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_541_U133
g20764 nand P3_ADD_541_U95 P3_ADD_541_U9 ; P3_ADD_541_U134
g20765 nand P3_ADD_541_U6 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_541_U135
g20766 nand P3_ADD_541_U94 P3_ADD_541_U7 ; P3_ADD_541_U136
g20767 nand P3_ADD_541_U93 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_541_U137
g20768 nand P3_ADD_541_U122 P3_ADD_541_U92 ; P3_ADD_541_U138
g20769 nand P3_ADD_541_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_541_U139
g20770 nand P3_ADD_541_U121 P3_ADD_541_U61 ; P3_ADD_541_U140
g20771 nand P3_ADD_541_U4 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_541_U141
g20772 nand P3_ADD_541_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_541_U142
g20773 nand P3_ADD_541_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_541_U143
g20774 nand P3_ADD_541_U120 P3_ADD_541_U59 ; P3_ADD_541_U144
g20775 nand P3_ADD_541_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_541_U145
g20776 nand P3_ADD_541_U119 P3_ADD_541_U57 ; P3_ADD_541_U146
g20777 nand P3_ADD_541_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_541_U147
g20778 nand P3_ADD_541_U118 P3_ADD_541_U55 ; P3_ADD_541_U148
g20779 nand P3_ADD_541_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_541_U149
g20780 nand P3_ADD_541_U117 P3_ADD_541_U53 ; P3_ADD_541_U150
g20781 nand P3_ADD_541_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_541_U151
g20782 nand P3_ADD_541_U116 P3_ADD_541_U51 ; P3_ADD_541_U152
g20783 nand P3_ADD_541_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_541_U153
g20784 nand P3_ADD_541_U115 P3_ADD_541_U49 ; P3_ADD_541_U154
g20785 nand P3_ADD_541_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_541_U155
g20786 nand P3_ADD_541_U114 P3_ADD_541_U47 ; P3_ADD_541_U156
g20787 nand P3_ADD_541_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_541_U157
g20788 nand P3_ADD_541_U113 P3_ADD_541_U45 ; P3_ADD_541_U158
g20789 nand P3_ADD_541_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_541_U159
g20790 nand P3_ADD_541_U112 P3_ADD_541_U43 ; P3_ADD_541_U160
g20791 nand P3_ADD_541_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_541_U161
g20792 nand P3_ADD_541_U111 P3_ADD_541_U41 ; P3_ADD_541_U162
g20793 nand P3_ADD_541_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_541_U163
g20794 nand P3_ADD_541_U110 P3_ADD_541_U39 ; P3_ADD_541_U164
g20795 nand P3_ADD_541_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_541_U165
g20796 nand P3_ADD_541_U109 P3_ADD_541_U37 ; P3_ADD_541_U166
g20797 nand P3_ADD_541_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_541_U167
g20798 nand P3_ADD_541_U108 P3_ADD_541_U35 ; P3_ADD_541_U168
g20799 nand P3_ADD_541_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_541_U169
g20800 nand P3_ADD_541_U107 P3_ADD_541_U33 ; P3_ADD_541_U170
g20801 nand P3_ADD_541_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_541_U171
g20802 nand P3_ADD_541_U106 P3_ADD_541_U31 ; P3_ADD_541_U172
g20803 nand P3_ADD_541_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_541_U173
g20804 nand P3_ADD_541_U105 P3_ADD_541_U29 ; P3_ADD_541_U174
g20805 nand P3_ADD_541_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_541_U175
g20806 nand P3_ADD_541_U104 P3_ADD_541_U27 ; P3_ADD_541_U176
g20807 nand P3_ADD_541_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_541_U177
g20808 nand P3_ADD_541_U103 P3_ADD_541_U25 ; P3_ADD_541_U178
g20809 nand P3_ADD_541_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_541_U179
g20810 nand P3_ADD_541_U102 P3_ADD_541_U23 ; P3_ADD_541_U180
g20811 nand P3_ADD_541_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_541_U181
g20812 nand P3_ADD_541_U101 P3_ADD_541_U21 ; P3_ADD_541_U182
g20813 nand P3_SUB_355_U45 P3_SUB_355_U44 ; P3_SUB_355_U6
g20814 nand P3_SUB_355_U9 P3_SUB_355_U46 ; P3_SUB_355_U7
g20815 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_355_U8
g20816 nand P3_SUB_355_U18 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_355_U9
g20817 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_355_U10
g20818 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_355_U11
g20819 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_355_U12
g20820 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_355_U13
g20821 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_355_U14
g20822 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_355_U15
g20823 nand P3_SUB_355_U41 P3_SUB_355_U40 ; P3_SUB_355_U16
g20824 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_355_U17
g20825 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_355_U18
g20826 nand P3_SUB_355_U51 P3_SUB_355_U50 ; P3_SUB_355_U19
g20827 nand P3_SUB_355_U56 P3_SUB_355_U55 ; P3_SUB_355_U20
g20828 nand P3_SUB_355_U61 P3_SUB_355_U60 ; P3_SUB_355_U21
g20829 nand P3_SUB_355_U66 P3_SUB_355_U65 ; P3_SUB_355_U22
g20830 nand P3_SUB_355_U48 P3_SUB_355_U47 ; P3_SUB_355_U23
g20831 nand P3_SUB_355_U53 P3_SUB_355_U52 ; P3_SUB_355_U24
g20832 nand P3_SUB_355_U58 P3_SUB_355_U57 ; P3_SUB_355_U25
g20833 nand P3_SUB_355_U63 P3_SUB_355_U62 ; P3_SUB_355_U26
g20834 nand P3_SUB_355_U37 P3_SUB_355_U36 ; P3_SUB_355_U27
g20835 nand P3_SUB_355_U33 P3_SUB_355_U32 ; P3_SUB_355_U28
g20836 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_355_U29
g20837 not P3_SUB_355_U9 ; P3_SUB_355_U30
g20838 nand P3_SUB_355_U30 P3_SUB_355_U10 ; P3_SUB_355_U31
g20839 nand P3_SUB_355_U31 P3_SUB_355_U29 ; P3_SUB_355_U32
g20840 nand P3_SUB_355_U9 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_355_U33
g20841 not P3_SUB_355_U28 ; P3_SUB_355_U34
g20842 nand P3_SUB_355_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_355_U35
g20843 nand P3_SUB_355_U35 P3_SUB_355_U28 ; P3_SUB_355_U36
g20844 nand P3_SUB_355_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_355_U37
g20845 not P3_SUB_355_U27 ; P3_SUB_355_U38
g20846 nand P3_SUB_355_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_355_U39
g20847 nand P3_SUB_355_U39 P3_SUB_355_U27 ; P3_SUB_355_U40
g20848 nand P3_SUB_355_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_355_U41
g20849 not P3_SUB_355_U16 ; P3_SUB_355_U42
g20850 nand P3_SUB_355_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_355_U43
g20851 nand P3_SUB_355_U42 P3_SUB_355_U43 ; P3_SUB_355_U44
g20852 nand P3_SUB_355_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_355_U45
g20853 nand P3_SUB_355_U8 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_355_U46
g20854 nand P3_SUB_355_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_355_U47
g20855 nand P3_SUB_355_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_355_U48
g20856 not P3_SUB_355_U23 ; P3_SUB_355_U49
g20857 nand P3_SUB_355_U49 P3_SUB_355_U42 ; P3_SUB_355_U50
g20858 nand P3_SUB_355_U23 P3_SUB_355_U16 ; P3_SUB_355_U51
g20859 nand P3_SUB_355_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_355_U52
g20860 nand P3_SUB_355_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_355_U53
g20861 not P3_SUB_355_U24 ; P3_SUB_355_U54
g20862 nand P3_SUB_355_U38 P3_SUB_355_U54 ; P3_SUB_355_U55
g20863 nand P3_SUB_355_U24 P3_SUB_355_U27 ; P3_SUB_355_U56
g20864 nand P3_SUB_355_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_355_U57
g20865 nand P3_SUB_355_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_355_U58
g20866 not P3_SUB_355_U25 ; P3_SUB_355_U59
g20867 nand P3_SUB_355_U34 P3_SUB_355_U59 ; P3_SUB_355_U60
g20868 nand P3_SUB_355_U25 P3_SUB_355_U28 ; P3_SUB_355_U61
g20869 nand P3_SUB_355_U10 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_355_U62
g20870 nand P3_SUB_355_U29 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_355_U63
g20871 not P3_SUB_355_U26 ; P3_SUB_355_U64
g20872 nand P3_SUB_355_U64 P3_SUB_355_U30 ; P3_SUB_355_U65
g20873 nand P3_SUB_355_U26 P3_SUB_355_U9 ; P3_SUB_355_U66
g20874 nand P3_SUB_450_U43 P3_SUB_450_U42 ; P3_SUB_450_U6
g20875 nand P3_SUB_450_U27 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_450_U7
g20876 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_450_U8
g20877 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_450_U9
g20878 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_450_U10
g20879 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_450_U11
g20880 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_450_U12
g20881 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_450_U13
g20882 nand P3_SUB_450_U39 P3_SUB_450_U38 ; P3_SUB_450_U14
g20883 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_450_U15
g20884 nand P3_SUB_450_U48 P3_SUB_450_U47 ; P3_SUB_450_U16
g20885 nand P3_SUB_450_U53 P3_SUB_450_U52 ; P3_SUB_450_U17
g20886 nand P3_SUB_450_U58 P3_SUB_450_U57 ; P3_SUB_450_U18
g20887 nand P3_SUB_450_U63 P3_SUB_450_U62 ; P3_SUB_450_U19
g20888 nand P3_SUB_450_U45 P3_SUB_450_U44 ; P3_SUB_450_U20
g20889 nand P3_SUB_450_U50 P3_SUB_450_U49 ; P3_SUB_450_U21
g20890 nand P3_SUB_450_U55 P3_SUB_450_U54 ; P3_SUB_450_U22
g20891 nand P3_SUB_450_U60 P3_SUB_450_U59 ; P3_SUB_450_U23
g20892 nand P3_SUB_450_U35 P3_SUB_450_U34 ; P3_SUB_450_U24
g20893 nand P3_SUB_450_U31 P3_SUB_450_U30 ; P3_SUB_450_U25
g20894 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_450_U26
g20895 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_450_U27
g20896 not P3_SUB_450_U7 ; P3_SUB_450_U28
g20897 nand P3_SUB_450_U28 P3_SUB_450_U8 ; P3_SUB_450_U29
g20898 nand P3_SUB_450_U29 P3_SUB_450_U26 ; P3_SUB_450_U30
g20899 nand P3_SUB_450_U7 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_450_U31
g20900 not P3_SUB_450_U25 ; P3_SUB_450_U32
g20901 nand P3_SUB_450_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_450_U33
g20902 nand P3_SUB_450_U33 P3_SUB_450_U25 ; P3_SUB_450_U34
g20903 nand P3_SUB_450_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_450_U35
g20904 not P3_SUB_450_U24 ; P3_SUB_450_U36
g20905 nand P3_SUB_450_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_450_U37
g20906 nand P3_SUB_450_U37 P3_SUB_450_U24 ; P3_SUB_450_U38
g20907 nand P3_SUB_450_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_450_U39
g20908 not P3_SUB_450_U14 ; P3_SUB_450_U40
g20909 nand P3_SUB_450_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_450_U41
g20910 nand P3_SUB_450_U40 P3_SUB_450_U41 ; P3_SUB_450_U42
g20911 nand P3_SUB_450_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_450_U43
g20912 nand P3_SUB_450_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_450_U44
g20913 nand P3_SUB_450_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_450_U45
g20914 not P3_SUB_450_U20 ; P3_SUB_450_U46
g20915 nand P3_SUB_450_U46 P3_SUB_450_U40 ; P3_SUB_450_U47
g20916 nand P3_SUB_450_U20 P3_SUB_450_U14 ; P3_SUB_450_U48
g20917 nand P3_SUB_450_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_450_U49
g20918 nand P3_SUB_450_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_450_U50
g20919 not P3_SUB_450_U21 ; P3_SUB_450_U51
g20920 nand P3_SUB_450_U36 P3_SUB_450_U51 ; P3_SUB_450_U52
g20921 nand P3_SUB_450_U21 P3_SUB_450_U24 ; P3_SUB_450_U53
g20922 nand P3_SUB_450_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_450_U54
g20923 nand P3_SUB_450_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_450_U55
g20924 not P3_SUB_450_U22 ; P3_SUB_450_U56
g20925 nand P3_SUB_450_U32 P3_SUB_450_U56 ; P3_SUB_450_U57
g20926 nand P3_SUB_450_U22 P3_SUB_450_U25 ; P3_SUB_450_U58
g20927 nand P3_SUB_450_U8 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_450_U59
g20928 nand P3_SUB_450_U26 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_450_U60
g20929 not P3_SUB_450_U23 ; P3_SUB_450_U61
g20930 nand P3_SUB_450_U61 P3_SUB_450_U28 ; P3_SUB_450_U62
g20931 nand P3_SUB_450_U23 P3_SUB_450_U7 ; P3_SUB_450_U63
g20932 and P3_INSTADDRPOINTER_REG_27__SCAN_IN P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_SUB_357_1258_U4
g20933 and P3_SUB_357_1258_U188 P3_SUB_357_1258_U186 ; P3_SUB_357_1258_U5
g20934 and P3_SUB_357_1258_U187 P3_SUB_357_1258_U178 ; P3_SUB_357_1258_U6
g20935 and P3_SUB_357_1258_U6 P3_SUB_357_1258_U189 ; P3_SUB_357_1258_U7
g20936 and P3_SUB_357_1258_U5 P3_SUB_357_1258_U190 ; P3_SUB_357_1258_U8
g20937 and P3_SUB_357_1258_U209 P3_SUB_357_1258_U204 ; P3_SUB_357_1258_U9
g20938 and P3_SUB_357_1258_U210 P3_SUB_357_1258_U205 P3_SUB_357_1258_U206 P3_SUB_357_1258_U156 ; P3_SUB_357_1258_U10
g20939 and P3_SUB_357_1258_U9 P3_SUB_357_1258_U211 ; P3_SUB_357_1258_U11
g20940 and P3_SUB_357_1258_U10 P3_SUB_357_1258_U212 ; P3_SUB_357_1258_U12
g20941 and P3_SUB_357_1258_U11 P3_SUB_357_1258_U213 ; P3_SUB_357_1258_U13
g20942 and P3_SUB_357_1258_U12 P3_SUB_357_1258_U214 ; P3_SUB_357_1258_U14
g20943 and P3_SUB_357_1258_U255 P3_SUB_357_1258_U252 ; P3_SUB_357_1258_U15
g20944 and P3_SUB_357_1258_U249 P3_SUB_357_1258_U248 ; P3_SUB_357_1258_U16
g20945 and P3_SUB_357_1258_U244 P3_SUB_357_1258_U241 ; P3_SUB_357_1258_U17
g20946 and P3_SUB_357_1258_U233 P3_SUB_357_1258_U230 ; P3_SUB_357_1258_U18
g20947 and P3_SUB_357_1258_U227 P3_SUB_357_1258_U303 ; P3_SUB_357_1258_U19
g20948 and P3_SUB_357_1258_U225 P3_SUB_357_1258_U296 ; P3_SUB_357_1258_U20
g20949 nand P3_SUB_357_1258_U426 P3_SUB_357_1258_U425 P3_SUB_357_1258_U307 ; P3_SUB_357_1258_U21
g20950 not P3_ADD_357_U9 ; P3_SUB_357_1258_U22
g20951 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_SUB_357_1258_U23
g20952 not P3_ADD_357_U8 ; P3_SUB_357_1258_U24
g20953 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_SUB_357_1258_U25
g20954 not P3_ADD_357_U19 ; P3_SUB_357_1258_U26
g20955 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_SUB_357_1258_U27
g20956 not P3_ADD_357_U10 ; P3_SUB_357_1258_U28
g20957 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_357_1258_U29
g20958 nand P3_ADD_357_U10 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_357_1258_U30
g20959 not P3_SUB_357_U7 ; P3_SUB_357_1258_U31
g20960 not P3_ADD_357_U13 ; P3_SUB_357_1258_U32
g20961 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_SUB_357_1258_U33
g20962 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_357_1258_U34
g20963 not P3_ADD_357_U7 ; P3_SUB_357_1258_U35
g20964 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_SUB_357_1258_U36
g20965 not P3_ADD_357_U17 ; P3_SUB_357_1258_U37
g20966 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_SUB_357_1258_U38
g20967 not P3_ADD_357_U6 ; P3_SUB_357_1258_U39
g20968 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_SUB_357_1258_U40
g20969 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_SUB_357_1258_U41
g20970 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_SUB_357_1258_U42
g20971 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_SUB_357_1258_U43
g20972 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_SUB_357_1258_U44
g20973 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_SUB_357_1258_U45
g20974 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_SUB_357_1258_U46
g20975 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_SUB_357_1258_U47
g20976 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_SUB_357_1258_U48
g20977 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_SUB_357_1258_U49
g20978 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_SUB_357_1258_U50
g20979 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_SUB_357_1258_U51
g20980 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_SUB_357_1258_U52
g20981 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_SUB_357_1258_U53
g20982 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_SUB_357_1258_U54
g20983 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_SUB_357_1258_U55
g20984 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_SUB_357_1258_U56
g20985 nand P3_INSTADDRPOINTER_REG_19__SCAN_IN P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_SUB_357_1258_U57
g20986 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_SUB_357_1258_U58
g20987 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_SUB_357_1258_U59
g20988 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_SUB_357_1258_U60
g20989 nand P3_SUB_357_1258_U222 P3_SUB_357_1258_U151 P3_SUB_357_1258_U269 ; P3_SUB_357_1258_U61
g20990 nand P3_SUB_357_1258_U105 P3_SUB_357_1258_U218 ; P3_SUB_357_1258_U62
g20991 nand P3_SUB_357_1258_U104 P3_SUB_357_1258_U284 ; P3_SUB_357_1258_U63
g20992 nand P3_SUB_357_1258_U276 P3_SUB_357_1258_U205 ; P3_SUB_357_1258_U64
g20993 nand P3_SUB_357_1258_U277 P3_SUB_357_1258_U47 ; P3_SUB_357_1258_U65
g20994 nand P3_SUB_357_U7 P3_SUB_357_1258_U161 ; P3_SUB_357_1258_U66
g20995 nand P3_SUB_357_1258_U102 P3_SUB_357_1258_U198 ; P3_SUB_357_1258_U67
g20996 nand P3_SUB_357_1258_U290 P3_SUB_357_1258_U8 ; P3_SUB_357_1258_U68
g20997 nand P3_SUB_357_1258_U484 P3_SUB_357_1258_U483 ; P3_SUB_357_1258_U69
g20998 nand P3_SUB_357_1258_U312 P3_SUB_357_1258_U311 ; P3_SUB_357_1258_U70
g20999 nand P3_SUB_357_1258_U319 P3_SUB_357_1258_U318 ; P3_SUB_357_1258_U71
g21000 nand P3_SUB_357_1258_U326 P3_SUB_357_1258_U325 ; P3_SUB_357_1258_U72
g21001 nand P3_SUB_357_1258_U333 P3_SUB_357_1258_U332 ; P3_SUB_357_1258_U73
g21002 nand P3_SUB_357_1258_U340 P3_SUB_357_1258_U339 ; P3_SUB_357_1258_U74
g21003 nand P3_SUB_357_1258_U345 P3_SUB_357_1258_U344 ; P3_SUB_357_1258_U75
g21004 nand P3_SUB_357_1258_U350 P3_SUB_357_1258_U349 ; P3_SUB_357_1258_U76
g21005 nand P3_SUB_357_1258_U361 P3_SUB_357_1258_U360 ; P3_SUB_357_1258_U77
g21006 nand P3_SUB_357_1258_U366 P3_SUB_357_1258_U365 ; P3_SUB_357_1258_U78
g21007 nand P3_SUB_357_1258_U373 P3_SUB_357_1258_U372 ; P3_SUB_357_1258_U79
g21008 nand P3_SUB_357_1258_U384 P3_SUB_357_1258_U383 ; P3_SUB_357_1258_U80
g21009 nand P3_SUB_357_1258_U391 P3_SUB_357_1258_U390 ; P3_SUB_357_1258_U81
g21010 nand P3_SUB_357_1258_U398 P3_SUB_357_1258_U397 ; P3_SUB_357_1258_U82
g21011 nand P3_SUB_357_1258_U405 P3_SUB_357_1258_U404 ; P3_SUB_357_1258_U83
g21012 nand P3_SUB_357_1258_U412 P3_SUB_357_1258_U411 ; P3_SUB_357_1258_U84
g21013 nand P3_SUB_357_1258_U419 P3_SUB_357_1258_U418 ; P3_SUB_357_1258_U85
g21014 nand P3_SUB_357_1258_U431 P3_SUB_357_1258_U430 ; P3_SUB_357_1258_U86
g21015 nand P3_SUB_357_1258_U438 P3_SUB_357_1258_U437 ; P3_SUB_357_1258_U87
g21016 nand P3_SUB_357_1258_U449 P3_SUB_357_1258_U448 ; P3_SUB_357_1258_U88
g21017 nand P3_SUB_357_1258_U456 P3_SUB_357_1258_U455 ; P3_SUB_357_1258_U89
g21018 nand P3_SUB_357_1258_U463 P3_SUB_357_1258_U462 ; P3_SUB_357_1258_U90
g21019 nand P3_SUB_357_1258_U470 P3_SUB_357_1258_U469 ; P3_SUB_357_1258_U91
g21020 nand P3_SUB_357_1258_U477 P3_SUB_357_1258_U476 ; P3_SUB_357_1258_U92
g21021 nand P3_SUB_357_1258_U482 P3_SUB_357_1258_U481 ; P3_SUB_357_1258_U93
g21022 and P3_SUB_357_1258_U163 P3_SUB_357_1258_U164 P3_SUB_357_1258_U160 ; P3_SUB_357_1258_U94
g21023 and P3_ADD_357_U7 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_SUB_357_1258_U95
g21024 and P3_SUB_357_1258_U168 P3_SUB_357_1258_U162 ; P3_SUB_357_1258_U96
g21025 and P3_SUB_357_1258_U164 P3_SUB_357_1258_U163 ; P3_SUB_357_1258_U97
g21026 and P3_SUB_357_1258_U7 P3_SUB_357_1258_U154 ; P3_SUB_357_1258_U98
g21027 and P3_SUB_357_1258_U192 P3_SUB_357_1258_U155 ; P3_SUB_357_1258_U99
g21028 and P3_SUB_357_1258_U99 P3_SUB_357_1258_U8 ; P3_SUB_357_1258_U100
g21029 and P3_INSTADDRPOINTER_REG_16__SCAN_IN P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_SUB_357_1258_U101
g21030 and P3_SUB_357_1258_U199 P3_SUB_357_1258_U56 ; P3_SUB_357_1258_U102
g21031 and P3_SUB_357_1258_U215 P3_SUB_357_1258_U13 ; P3_SUB_357_1258_U103
g21032 and P3_SUB_357_1258_U14 P3_SUB_357_1258_U216 ; P3_SUB_357_1258_U104
g21033 and P3_SUB_357_1258_U157 P3_SUB_357_1258_U58 P3_SUB_357_1258_U219 ; P3_SUB_357_1258_U105
g21034 and P3_SUB_357_1258_U219 P3_SUB_357_1258_U157 ; P3_SUB_357_1258_U106
g21035 and P3_SUB_357_1258_U60 P3_SUB_357_1258_U269 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_SUB_357_1258_U107
g21036 and P3_INSTADDRPOINTER_REG_30__SCAN_IN P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_SUB_357_1258_U108
g21037 and P3_SUB_357_1258_U386 P3_SUB_357_1258_U385 P3_SUB_357_1258_U157 ; P3_SUB_357_1258_U109
g21038 and P3_SUB_357_1258_U232 P3_SUB_357_1258_U153 ; P3_SUB_357_1258_U110
g21039 and P3_SUB_357_1258_U237 P3_SUB_357_1258_U156 ; P3_SUB_357_1258_U111
g21040 and P3_SUB_357_1258_U243 P3_SUB_357_1258_U156 ; P3_SUB_357_1258_U112
g21041 and P3_SUB_357_1258_U465 P3_SUB_357_1258_U464 P3_SUB_357_1258_U155 ; P3_SUB_357_1258_U113
g21042 and P3_SUB_357_1258_U254 P3_SUB_357_1258_U154 ; P3_SUB_357_1258_U114
g21043 nand P3_SUB_357_1258_U176 P3_SUB_357_1258_U152 P3_SUB_357_1258_U268 ; P3_SUB_357_1258_U115
g21044 and P3_SUB_357_1258_U314 P3_SUB_357_1258_U313 ; P3_SUB_357_1258_U116
g21045 nand P3_SUB_357_1258_U300 P3_SUB_357_1258_U267 ; P3_SUB_357_1258_U117
g21046 and P3_SUB_357_1258_U321 P3_SUB_357_1258_U320 ; P3_SUB_357_1258_U118
g21047 nand P3_SUB_357_1258_U173 P3_SUB_357_1258_U172 ; P3_SUB_357_1258_U119
g21048 and P3_SUB_357_1258_U328 P3_SUB_357_1258_U327 ; P3_SUB_357_1258_U120
g21049 nand P3_SUB_357_1258_U298 P3_SUB_357_1258_U266 ; P3_SUB_357_1258_U121
g21050 and P3_SUB_357_1258_U335 P3_SUB_357_1258_U334 ; P3_SUB_357_1258_U122
g21051 nand P3_SUB_357_1258_U96 P3_SUB_357_1258_U167 ; P3_SUB_357_1258_U123
g21052 nand P3_SUB_357_1258_U181 P3_SUB_357_1258_U180 ; P3_SUB_357_1258_U124
g21053 nand P3_SUB_357_1258_U159 P3_SUB_357_1258_U183 ; P3_SUB_357_1258_U125
g21054 and P3_SUB_357_1258_U356 P3_SUB_357_1258_U355 ; P3_SUB_357_1258_U126
g21055 nand P3_SUB_357_1258_U270 P3_SUB_357_1258_U66 P3_SUB_357_1258_U271 ; P3_SUB_357_1258_U127
g21056 and P3_SUB_357_1258_U368 P3_SUB_357_1258_U367 ; P3_SUB_357_1258_U128
g21057 nand P3_SUB_357_1258_U275 P3_SUB_357_1258_U274 P3_SUB_357_1258_U304 ; P3_SUB_357_1258_U129
g21058 and P3_SUB_357_1258_U379 P3_SUB_357_1258_U378 ; P3_SUB_357_1258_U130
g21059 nand P3_SUB_357_1258_U106 P3_SUB_357_1258_U218 ; P3_SUB_357_1258_U131
g21060 and P3_SUB_357_1258_U393 P3_SUB_357_1258_U392 ; P3_SUB_357_1258_U132
g21061 nand P3_SUB_357_1258_U282 P3_SUB_357_1258_U14 ; P3_SUB_357_1258_U133
g21062 and P3_SUB_357_1258_U400 P3_SUB_357_1258_U399 ; P3_SUB_357_1258_U134
g21063 nand P3_SUB_357_1258_U280 P3_SUB_357_1258_U12 ; P3_SUB_357_1258_U135
g21064 and P3_SUB_357_1258_U407 P3_SUB_357_1258_U406 ; P3_SUB_357_1258_U136
g21065 nand P3_SUB_357_1258_U278 P3_SUB_357_1258_U10 ; P3_SUB_357_1258_U137
g21066 and P3_SUB_357_1258_U414 P3_SUB_357_1258_U413 ; P3_SUB_357_1258_U138
g21067 nand P3_SUB_357_1258_U111 P3_SUB_357_1258_U236 ; P3_SUB_357_1258_U139
g21068 and P3_SUB_357_1258_U433 P3_SUB_357_1258_U432 ; P3_SUB_357_1258_U140
g21069 nand P3_SUB_357_1258_U272 P3_SUB_357_1258_U201 P3_SUB_357_1258_U273 ; P3_SUB_357_1258_U141
g21070 and P3_SUB_357_1258_U444 P3_SUB_357_1258_U443 ; P3_SUB_357_1258_U142
g21071 nand P3_SUB_357_1258_U199 P3_SUB_357_1258_U198 ; P3_SUB_357_1258_U143
g21072 and P3_SUB_357_1258_U451 P3_SUB_357_1258_U450 ; P3_SUB_357_1258_U144
g21073 nand P3_SUB_357_1258_U195 P3_SUB_357_1258_U194 ; P3_SUB_357_1258_U145
g21074 and P3_SUB_357_1258_U458 P3_SUB_357_1258_U457 ; P3_SUB_357_1258_U146
g21075 nand P3_SUB_357_1258_U100 P3_SUB_357_1258_U292 ; P3_SUB_357_1258_U147
g21076 and P3_SUB_357_1258_U472 P3_SUB_357_1258_U471 ; P3_SUB_357_1258_U148
g21077 nand P3_SUB_357_1258_U288 P3_SUB_357_1258_U5 ; P3_SUB_357_1258_U149
g21078 nand P3_SUB_357_1258_U286 P3_SUB_357_1258_U186 ; P3_SUB_357_1258_U150
g21079 nand P3_ADD_357_U6 P3_SUB_357_1258_U129 ; P3_SUB_357_1258_U151
g21080 nand P3_ADD_357_U6 P3_SUB_357_1258_U117 ; P3_SUB_357_1258_U152
g21081 nand P3_SUB_357_1258_U217 P3_SUB_357_1258_U39 ; P3_SUB_357_1258_U153
g21082 nand P3_SUB_357_1258_U191 P3_SUB_357_1258_U39 ; P3_SUB_357_1258_U154
g21083 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_SUB_357_1258_U155
g21084 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_SUB_357_1258_U156
g21085 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_SUB_357_1258_U157
g21086 not P3_SUB_357_1258_U66 ; P3_SUB_357_1258_U158
g21087 nand P3_ADD_357_U13 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_SUB_357_1258_U159
g21088 or P3_ADD_357_U19 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_SUB_357_1258_U160
g21089 not P3_SUB_357_1258_U30 ; P3_SUB_357_1258_U161
g21090 nand P3_ADD_357_U19 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_SUB_357_1258_U162
g21091 or P3_ADD_357_U7 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_SUB_357_1258_U163
g21092 or P3_ADD_357_U13 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_SUB_357_1258_U164
g21093 not P3_SUB_357_1258_U127 ; P3_SUB_357_1258_U165
g21094 nand P3_SUB_357_1258_U271 P3_SUB_357_1258_U270 P3_SUB_357_1258_U159 P3_SUB_357_1258_U66 ; P3_SUB_357_1258_U166
g21095 nand P3_SUB_357_1258_U94 P3_SUB_357_1258_U166 ; P3_SUB_357_1258_U167
g21096 nand P3_SUB_357_1258_U95 P3_SUB_357_1258_U160 ; P3_SUB_357_1258_U168
g21097 not P3_SUB_357_1258_U123 ; P3_SUB_357_1258_U169
g21098 or P3_ADD_357_U8 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_SUB_357_1258_U170
g21099 or P3_ADD_357_U17 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_SUB_357_1258_U171
g21100 nand P3_SUB_357_1258_U171 P3_SUB_357_1258_U121 ; P3_SUB_357_1258_U172
g21101 nand P3_ADD_357_U17 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_SUB_357_1258_U173
g21102 not P3_SUB_357_1258_U119 ; P3_SUB_357_1258_U174
g21103 or P3_ADD_357_U9 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_SUB_357_1258_U175
g21104 nand P3_SUB_357_1258_U117 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_SUB_357_1258_U176
g21105 not P3_SUB_357_1258_U115 ; P3_SUB_357_1258_U177
g21106 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_SUB_357_1258_U178
g21107 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_SUB_357_1258_U179
g21108 nand P3_SUB_357_1258_U97 P3_SUB_357_1258_U166 ; P3_SUB_357_1258_U180
g21109 nand P3_ADD_357_U7 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_SUB_357_1258_U181
g21110 not P3_SUB_357_1258_U124 ; P3_SUB_357_1258_U182
g21111 nand P3_SUB_357_1258_U127 P3_SUB_357_1258_U164 ; P3_SUB_357_1258_U183
g21112 not P3_SUB_357_1258_U125 ; P3_SUB_357_1258_U184
g21113 nand P3_ADD_357_U7 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_SUB_357_1258_U185
g21114 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_SUB_357_1258_U186
g21115 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_SUB_357_1258_U187
g21116 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_SUB_357_1258_U188
g21117 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_SUB_357_1258_U189
g21118 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_SUB_357_1258_U190
g21119 nand P3_INSTADDRPOINTER_REG_12__SCAN_IN P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_SUB_357_1258_U191
g21120 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_SUB_357_1258_U192
g21121 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_SUB_357_1258_U193
g21122 nand P3_SUB_357_1258_U193 P3_SUB_357_1258_U147 ; P3_SUB_357_1258_U194
g21123 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_SUB_357_1258_U195
g21124 not P3_SUB_357_1258_U145 ; P3_SUB_357_1258_U196
g21125 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_SUB_357_1258_U197
g21126 nand P3_SUB_357_1258_U197 P3_SUB_357_1258_U145 ; P3_SUB_357_1258_U198
g21127 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_SUB_357_1258_U199
g21128 not P3_SUB_357_1258_U143 ; P3_SUB_357_1258_U200
g21129 nand P3_SUB_357_1258_U101 P3_SUB_357_1258_U143 ; P3_SUB_357_1258_U201
g21130 not P3_SUB_357_1258_U67 ; P3_SUB_357_1258_U202
g21131 not P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U203
g21132 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_SUB_357_1258_U204
g21133 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_SUB_357_1258_U205
g21134 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_SUB_357_1258_U206
g21135 not P3_SUB_357_1258_U57 ; P3_SUB_357_1258_U207
g21136 nand P3_SUB_357_1258_U207 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_SUB_357_1258_U208
g21137 nand P3_SUB_357_1258_U39 P3_SUB_357_1258_U208 ; P3_SUB_357_1258_U209
g21138 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_SUB_357_1258_U210
g21139 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_SUB_357_1258_U211
g21140 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_SUB_357_1258_U212
g21141 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_SUB_357_1258_U213
g21142 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_SUB_357_1258_U214
g21143 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_SUB_357_1258_U215
g21144 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_SUB_357_1258_U216
g21145 nand P3_INSTADDRPOINTER_REG_25__SCAN_IN P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_SUB_357_1258_U217
g21146 nand P3_SUB_357_1258_U63 P3_SUB_357_1258_U153 ; P3_SUB_357_1258_U218
g21147 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_SUB_357_1258_U219
g21148 not P3_SUB_357_1258_U131 ; P3_SUB_357_1258_U220
g21149 not P3_SUB_357_1258_U62 ; P3_SUB_357_1258_U221
g21150 nand P3_SUB_357_1258_U129 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_SUB_357_1258_U222
g21151 not P3_SUB_357_1258_U61 ; P3_SUB_357_1258_U223
g21152 nand P3_SUB_357_1258_U151 P3_SUB_357_1258_U107 ; P3_SUB_357_1258_U224
g21153 nand P3_SUB_357_1258_U354 P3_SUB_357_1258_U353 P3_SUB_357_1258_U294 ; P3_SUB_357_1258_U225
g21154 nand P3_SUB_357_1258_U221 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_SUB_357_1258_U226
g21155 nand P3_SUB_357_1258_U377 P3_SUB_357_1258_U376 P3_SUB_357_1258_U62 ; P3_SUB_357_1258_U227
g21156 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_SUB_357_1258_U228
g21157 nand P3_SUB_357_1258_U228 P3_SUB_357_1258_U63 ; P3_SUB_357_1258_U229
g21158 nand P3_SUB_357_1258_U109 P3_SUB_357_1258_U229 ; P3_SUB_357_1258_U230
g21159 nand P3_SUB_357_1258_U285 P3_SUB_357_1258_U157 ; P3_SUB_357_1258_U231
g21160 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_SUB_357_1258_U232
g21161 nand P3_SUB_357_1258_U110 P3_SUB_357_1258_U231 ; P3_SUB_357_1258_U233
g21162 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_SUB_357_1258_U234
g21163 not P3_SUB_357_1258_U65 ; P3_SUB_357_1258_U235
g21164 nand P3_ADD_357_U6 P3_SUB_357_1258_U65 ; P3_SUB_357_1258_U236
g21165 nand P3_SUB_357_1258_U207 P3_SUB_357_1258_U64 ; P3_SUB_357_1258_U237
g21166 not P3_SUB_357_1258_U139 ; P3_SUB_357_1258_U238
g21167 nand P3_SUB_357_1258_U235 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_SUB_357_1258_U239
g21168 nand P3_SUB_357_1258_U64 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_SUB_357_1258_U240
g21169 nand P3_SUB_357_1258_U421 P3_SUB_357_1258_U420 P3_SUB_357_1258_U240 ; P3_SUB_357_1258_U241
g21170 nand P3_SUB_357_1258_U277 P3_SUB_357_1258_U206 ; P3_SUB_357_1258_U242
g21171 nand P3_SUB_357_1258_U57 P3_SUB_357_1258_U39 ; P3_SUB_357_1258_U243
g21172 nand P3_SUB_357_1258_U112 P3_SUB_357_1258_U242 ; P3_SUB_357_1258_U244
g21173 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_SUB_357_1258_U245
g21174 nand P3_SUB_357_1258_U202 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_SUB_357_1258_U246
g21175 nand P3_SUB_357_1258_U143 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_SUB_357_1258_U247
g21176 nand P3_SUB_357_1258_U440 P3_SUB_357_1258_U439 P3_SUB_357_1258_U247 ; P3_SUB_357_1258_U248
g21177 nand P3_SUB_357_1258_U442 P3_SUB_357_1258_U441 P3_SUB_357_1258_U67 ; P3_SUB_357_1258_U249
g21178 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_SUB_357_1258_U250
g21179 nand P3_SUB_357_1258_U250 P3_SUB_357_1258_U68 ; P3_SUB_357_1258_U251
g21180 nand P3_SUB_357_1258_U113 P3_SUB_357_1258_U251 ; P3_SUB_357_1258_U252
g21181 nand P3_SUB_357_1258_U291 P3_SUB_357_1258_U155 ; P3_SUB_357_1258_U253
g21182 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_SUB_357_1258_U254
g21183 nand P3_SUB_357_1258_U114 P3_SUB_357_1258_U253 ; P3_SUB_357_1258_U255
g21184 or P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_SUB_357_1258_U256
g21185 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_SUB_357_1258_U257
g21186 nand P3_SUB_357_1258_U179 P3_SUB_357_1258_U178 ; P3_SUB_357_1258_U258
g21187 nand P3_SUB_357_1258_U162 P3_SUB_357_1258_U160 ; P3_SUB_357_1258_U259
g21188 nand P3_SUB_357_1258_U185 P3_SUB_357_1258_U163 ; P3_SUB_357_1258_U260
g21189 nand P3_SUB_357_1258_U164 P3_SUB_357_1258_U159 ; P3_SUB_357_1258_U261
g21190 nand P3_SUB_357_1258_U234 P3_SUB_357_1258_U157 ; P3_SUB_357_1258_U262
g21191 nand P3_SUB_357_1258_U245 P3_SUB_357_1258_U206 ; P3_SUB_357_1258_U263
g21192 nand P3_SUB_357_1258_U256 P3_SUB_357_1258_U155 ; P3_SUB_357_1258_U264
g21193 nand P3_SUB_357_1258_U257 P3_SUB_357_1258_U187 ; P3_SUB_357_1258_U265
g21194 nand P3_ADD_357_U8 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_SUB_357_1258_U266
g21195 nand P3_ADD_357_U9 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_SUB_357_1258_U267
g21196 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_SUB_357_1258_U268
g21197 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_SUB_357_1258_U269
g21198 nand P3_SUB_357_1258_U161 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_357_1258_U270
g21199 nand P3_SUB_357_U7 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_357_1258_U271
g21200 nand P3_ADD_357_U6 P3_SUB_357_1258_U67 ; P3_SUB_357_1258_U272
g21201 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_SUB_357_1258_U273
g21202 nand P3_ADD_357_U6 P3_SUB_357_1258_U62 ; P3_SUB_357_1258_U274
g21203 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_SUB_357_1258_U275
g21204 nand P3_SUB_357_1258_U204 P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U276
g21205 not P3_SUB_357_1258_U64 ; P3_SUB_357_1258_U277
g21206 nand P3_SUB_357_1258_U9 P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U278
g21207 not P3_SUB_357_1258_U137 ; P3_SUB_357_1258_U279
g21208 nand P3_SUB_357_1258_U11 P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U280
g21209 not P3_SUB_357_1258_U135 ; P3_SUB_357_1258_U281
g21210 nand P3_SUB_357_1258_U13 P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U282
g21211 not P3_SUB_357_1258_U133 ; P3_SUB_357_1258_U283
g21212 nand P3_SUB_357_1258_U103 P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U284
g21213 not P3_SUB_357_1258_U63 ; P3_SUB_357_1258_U285
g21214 nand P3_SUB_357_1258_U178 P3_SUB_357_1258_U115 ; P3_SUB_357_1258_U286
g21215 not P3_SUB_357_1258_U150 ; P3_SUB_357_1258_U287
g21216 nand P3_SUB_357_1258_U6 P3_SUB_357_1258_U115 ; P3_SUB_357_1258_U288
g21217 not P3_SUB_357_1258_U149 ; P3_SUB_357_1258_U289
g21218 nand P3_SUB_357_1258_U7 P3_SUB_357_1258_U115 ; P3_SUB_357_1258_U290
g21219 not P3_SUB_357_1258_U68 ; P3_SUB_357_1258_U291
g21220 nand P3_SUB_357_1258_U98 P3_SUB_357_1258_U115 ; P3_SUB_357_1258_U292
g21221 not P3_SUB_357_1258_U147 ; P3_SUB_357_1258_U293
g21222 nand P3_SUB_357_1258_U223 P3_SUB_357_1258_U60 ; P3_SUB_357_1258_U294
g21223 nand P3_SUB_357_1258_U61 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_SUB_357_1258_U295
g21224 nand P3_SUB_357_1258_U352 P3_SUB_357_1258_U351 P3_SUB_357_1258_U295 ; P3_SUB_357_1258_U296
g21225 nand P3_SUB_357_1258_U108 P3_SUB_357_1258_U61 ; P3_SUB_357_1258_U297
g21226 nand P3_SUB_357_1258_U170 P3_SUB_357_1258_U123 ; P3_SUB_357_1258_U298
g21227 not P3_SUB_357_1258_U121 ; P3_SUB_357_1258_U299
g21228 nand P3_SUB_357_1258_U175 P3_SUB_357_1258_U119 ; P3_SUB_357_1258_U300
g21229 not P3_SUB_357_1258_U117 ; P3_SUB_357_1258_U301
g21230 nand P3_SUB_357_1258_U131 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_SUB_357_1258_U302
g21231 nand P3_SUB_357_1258_U375 P3_SUB_357_1258_U374 P3_SUB_357_1258_U302 ; P3_SUB_357_1258_U303
g21232 nand P3_SUB_357_1258_U4 P3_SUB_357_1258_U131 ; P3_SUB_357_1258_U304
g21233 not P3_SUB_357_1258_U129 ; P3_SUB_357_1258_U305
g21234 nand P3_SUB_357_1258_U4 P3_SUB_357_1258_U131 ; P3_SUB_357_1258_U306
g21235 nand P3_SUB_357_1258_U158 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_357_1258_U307
g21236 nand P3_ADD_357_U6 P3_SUB_357_1258_U41 ; P3_SUB_357_1258_U308
g21237 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_SUB_357_1258_U309
g21238 nand P3_SUB_357_1258_U309 P3_SUB_357_1258_U308 ; P3_SUB_357_1258_U310
g21239 nand P3_SUB_357_1258_U258 P3_SUB_357_1258_U115 ; P3_SUB_357_1258_U311
g21240 nand P3_SUB_357_1258_U177 P3_SUB_357_1258_U310 ; P3_SUB_357_1258_U312
g21241 nand P3_ADD_357_U6 P3_SUB_357_1258_U40 ; P3_SUB_357_1258_U313
g21242 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_SUB_357_1258_U314
g21243 nand P3_ADD_357_U6 P3_SUB_357_1258_U40 ; P3_SUB_357_1258_U315
g21244 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_SUB_357_1258_U316
g21245 nand P3_SUB_357_1258_U316 P3_SUB_357_1258_U315 ; P3_SUB_357_1258_U317
g21246 nand P3_SUB_357_1258_U116 P3_SUB_357_1258_U117 ; P3_SUB_357_1258_U318
g21247 nand P3_SUB_357_1258_U301 P3_SUB_357_1258_U317 ; P3_SUB_357_1258_U319
g21248 nand P3_SUB_357_1258_U22 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_SUB_357_1258_U320
g21249 nand P3_ADD_357_U9 P3_SUB_357_1258_U23 ; P3_SUB_357_1258_U321
g21250 nand P3_SUB_357_1258_U22 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_SUB_357_1258_U322
g21251 nand P3_ADD_357_U9 P3_SUB_357_1258_U23 ; P3_SUB_357_1258_U323
g21252 nand P3_SUB_357_1258_U323 P3_SUB_357_1258_U322 ; P3_SUB_357_1258_U324
g21253 nand P3_SUB_357_1258_U118 P3_SUB_357_1258_U119 ; P3_SUB_357_1258_U325
g21254 nand P3_SUB_357_1258_U174 P3_SUB_357_1258_U324 ; P3_SUB_357_1258_U326
g21255 nand P3_SUB_357_1258_U37 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_SUB_357_1258_U327
g21256 nand P3_ADD_357_U17 P3_SUB_357_1258_U38 ; P3_SUB_357_1258_U328
g21257 nand P3_SUB_357_1258_U37 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_SUB_357_1258_U329
g21258 nand P3_ADD_357_U17 P3_SUB_357_1258_U38 ; P3_SUB_357_1258_U330
g21259 nand P3_SUB_357_1258_U330 P3_SUB_357_1258_U329 ; P3_SUB_357_1258_U331
g21260 nand P3_SUB_357_1258_U120 P3_SUB_357_1258_U121 ; P3_SUB_357_1258_U332
g21261 nand P3_SUB_357_1258_U299 P3_SUB_357_1258_U331 ; P3_SUB_357_1258_U333
g21262 nand P3_SUB_357_1258_U24 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_SUB_357_1258_U334
g21263 nand P3_ADD_357_U8 P3_SUB_357_1258_U25 ; P3_SUB_357_1258_U335
g21264 nand P3_SUB_357_1258_U24 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_SUB_357_1258_U336
g21265 nand P3_ADD_357_U8 P3_SUB_357_1258_U25 ; P3_SUB_357_1258_U337
g21266 nand P3_SUB_357_1258_U337 P3_SUB_357_1258_U336 ; P3_SUB_357_1258_U338
g21267 nand P3_SUB_357_1258_U122 P3_SUB_357_1258_U123 ; P3_SUB_357_1258_U339
g21268 nand P3_SUB_357_1258_U169 P3_SUB_357_1258_U338 ; P3_SUB_357_1258_U340
g21269 nand P3_SUB_357_1258_U26 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_SUB_357_1258_U341
g21270 nand P3_ADD_357_U19 P3_SUB_357_1258_U27 ; P3_SUB_357_1258_U342
g21271 nand P3_SUB_357_1258_U342 P3_SUB_357_1258_U341 ; P3_SUB_357_1258_U343
g21272 nand P3_SUB_357_1258_U259 P3_SUB_357_1258_U124 ; P3_SUB_357_1258_U344
g21273 nand P3_SUB_357_1258_U182 P3_SUB_357_1258_U343 ; P3_SUB_357_1258_U345
g21274 nand P3_SUB_357_1258_U35 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_SUB_357_1258_U346
g21275 nand P3_ADD_357_U7 P3_SUB_357_1258_U36 ; P3_SUB_357_1258_U347
g21276 nand P3_SUB_357_1258_U347 P3_SUB_357_1258_U346 ; P3_SUB_357_1258_U348
g21277 nand P3_SUB_357_1258_U260 P3_SUB_357_1258_U125 ; P3_SUB_357_1258_U349
g21278 nand P3_SUB_357_1258_U184 P3_SUB_357_1258_U348 ; P3_SUB_357_1258_U350
g21279 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_SUB_357_1258_U351
g21280 nand P3_ADD_357_U6 P3_SUB_357_1258_U224 ; P3_SUB_357_1258_U352
g21281 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_SUB_357_1258_U353
g21282 nand P3_SUB_357_1258_U297 P3_SUB_357_1258_U39 ; P3_SUB_357_1258_U354
g21283 nand P3_ADD_357_U6 P3_SUB_357_1258_U60 ; P3_SUB_357_1258_U355
g21284 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_SUB_357_1258_U356
g21285 nand P3_ADD_357_U6 P3_SUB_357_1258_U60 ; P3_SUB_357_1258_U357
g21286 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_SUB_357_1258_U358
g21287 nand P3_SUB_357_1258_U358 P3_SUB_357_1258_U357 ; P3_SUB_357_1258_U359
g21288 nand P3_SUB_357_1258_U126 P3_SUB_357_1258_U61 ; P3_SUB_357_1258_U360
g21289 nand P3_SUB_357_1258_U359 P3_SUB_357_1258_U223 ; P3_SUB_357_1258_U361
g21290 nand P3_SUB_357_1258_U32 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_SUB_357_1258_U362
g21291 nand P3_ADD_357_U13 P3_SUB_357_1258_U33 ; P3_SUB_357_1258_U363
g21292 nand P3_SUB_357_1258_U363 P3_SUB_357_1258_U362 ; P3_SUB_357_1258_U364
g21293 nand P3_SUB_357_1258_U261 P3_SUB_357_1258_U127 ; P3_SUB_357_1258_U365
g21294 nand P3_SUB_357_1258_U165 P3_SUB_357_1258_U364 ; P3_SUB_357_1258_U366
g21295 nand P3_ADD_357_U6 P3_SUB_357_1258_U59 ; P3_SUB_357_1258_U367
g21296 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_SUB_357_1258_U368
g21297 nand P3_ADD_357_U6 P3_SUB_357_1258_U59 ; P3_SUB_357_1258_U369
g21298 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_SUB_357_1258_U370
g21299 nand P3_SUB_357_1258_U370 P3_SUB_357_1258_U369 ; P3_SUB_357_1258_U371
g21300 nand P3_SUB_357_1258_U128 P3_SUB_357_1258_U129 ; P3_SUB_357_1258_U372
g21301 nand P3_SUB_357_1258_U305 P3_SUB_357_1258_U371 ; P3_SUB_357_1258_U373
g21302 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_SUB_357_1258_U374
g21303 nand P3_ADD_357_U6 P3_SUB_357_1258_U226 ; P3_SUB_357_1258_U375
g21304 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_SUB_357_1258_U376
g21305 nand P3_SUB_357_1258_U306 P3_SUB_357_1258_U39 ; P3_SUB_357_1258_U377
g21306 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_SUB_357_1258_U378
g21307 nand P3_ADD_357_U6 P3_SUB_357_1258_U58 ; P3_SUB_357_1258_U379
g21308 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_SUB_357_1258_U380
g21309 nand P3_ADD_357_U6 P3_SUB_357_1258_U58 ; P3_SUB_357_1258_U381
g21310 nand P3_SUB_357_1258_U381 P3_SUB_357_1258_U380 ; P3_SUB_357_1258_U382
g21311 nand P3_SUB_357_1258_U130 P3_SUB_357_1258_U131 ; P3_SUB_357_1258_U383
g21312 nand P3_SUB_357_1258_U220 P3_SUB_357_1258_U382 ; P3_SUB_357_1258_U384
g21313 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_SUB_357_1258_U385
g21314 nand P3_ADD_357_U6 P3_SUB_357_1258_U43 ; P3_SUB_357_1258_U386
g21315 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_SUB_357_1258_U387
g21316 nand P3_ADD_357_U6 P3_SUB_357_1258_U42 ; P3_SUB_357_1258_U388
g21317 nand P3_SUB_357_1258_U388 P3_SUB_357_1258_U387 ; P3_SUB_357_1258_U389
g21318 nand P3_SUB_357_1258_U63 P3_SUB_357_1258_U262 ; P3_SUB_357_1258_U390
g21319 nand P3_SUB_357_1258_U389 P3_SUB_357_1258_U285 ; P3_SUB_357_1258_U391
g21320 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_SUB_357_1258_U392
g21321 nand P3_ADD_357_U6 P3_SUB_357_1258_U44 ; P3_SUB_357_1258_U393
g21322 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_SUB_357_1258_U394
g21323 nand P3_ADD_357_U6 P3_SUB_357_1258_U44 ; P3_SUB_357_1258_U395
g21324 nand P3_SUB_357_1258_U395 P3_SUB_357_1258_U394 ; P3_SUB_357_1258_U396
g21325 nand P3_SUB_357_1258_U132 P3_SUB_357_1258_U133 ; P3_SUB_357_1258_U397
g21326 nand P3_SUB_357_1258_U283 P3_SUB_357_1258_U396 ; P3_SUB_357_1258_U398
g21327 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_SUB_357_1258_U399
g21328 nand P3_ADD_357_U6 P3_SUB_357_1258_U45 ; P3_SUB_357_1258_U400
g21329 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_SUB_357_1258_U401
g21330 nand P3_ADD_357_U6 P3_SUB_357_1258_U45 ; P3_SUB_357_1258_U402
g21331 nand P3_SUB_357_1258_U402 P3_SUB_357_1258_U401 ; P3_SUB_357_1258_U403
g21332 nand P3_SUB_357_1258_U134 P3_SUB_357_1258_U135 ; P3_SUB_357_1258_U404
g21333 nand P3_SUB_357_1258_U281 P3_SUB_357_1258_U403 ; P3_SUB_357_1258_U405
g21334 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_SUB_357_1258_U406
g21335 nand P3_ADD_357_U6 P3_SUB_357_1258_U46 ; P3_SUB_357_1258_U407
g21336 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_SUB_357_1258_U408
g21337 nand P3_ADD_357_U6 P3_SUB_357_1258_U46 ; P3_SUB_357_1258_U409
g21338 nand P3_SUB_357_1258_U409 P3_SUB_357_1258_U408 ; P3_SUB_357_1258_U410
g21339 nand P3_SUB_357_1258_U136 P3_SUB_357_1258_U137 ; P3_SUB_357_1258_U411
g21340 nand P3_SUB_357_1258_U279 P3_SUB_357_1258_U410 ; P3_SUB_357_1258_U412
g21341 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_SUB_357_1258_U413
g21342 nand P3_ADD_357_U6 P3_SUB_357_1258_U48 ; P3_SUB_357_1258_U414
g21343 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_SUB_357_1258_U415
g21344 nand P3_ADD_357_U6 P3_SUB_357_1258_U48 ; P3_SUB_357_1258_U416
g21345 nand P3_SUB_357_1258_U416 P3_SUB_357_1258_U415 ; P3_SUB_357_1258_U417
g21346 nand P3_SUB_357_1258_U138 P3_SUB_357_1258_U139 ; P3_SUB_357_1258_U418
g21347 nand P3_SUB_357_1258_U238 P3_SUB_357_1258_U417 ; P3_SUB_357_1258_U419
g21348 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_SUB_357_1258_U420
g21349 nand P3_ADD_357_U6 P3_SUB_357_1258_U239 ; P3_SUB_357_1258_U421
g21350 nand P3_SUB_357_1258_U30 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_SUB_357_1258_U422
g21351 nand P3_SUB_357_1258_U161 P3_SUB_357_1258_U34 ; P3_SUB_357_1258_U423
g21352 nand P3_SUB_357_1258_U423 P3_SUB_357_1258_U422 ; P3_SUB_357_1258_U424
g21353 nand P3_SUB_357_1258_U30 P3_SUB_357_1258_U34 P3_SUB_357_U7 ; P3_SUB_357_1258_U425
g21354 nand P3_SUB_357_1258_U424 P3_SUB_357_1258_U31 ; P3_SUB_357_1258_U426
g21355 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_SUB_357_1258_U427
g21356 nand P3_ADD_357_U6 P3_SUB_357_1258_U47 ; P3_SUB_357_1258_U428
g21357 nand P3_SUB_357_1258_U428 P3_SUB_357_1258_U427 ; P3_SUB_357_1258_U429
g21358 nand P3_SUB_357_1258_U64 P3_SUB_357_1258_U263 ; P3_SUB_357_1258_U430
g21359 nand P3_SUB_357_1258_U429 P3_SUB_357_1258_U277 ; P3_SUB_357_1258_U431
g21360 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_SUB_357_1258_U432
g21361 nand P3_ADD_357_U6 P3_SUB_357_1258_U49 ; P3_SUB_357_1258_U433
g21362 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_SUB_357_1258_U434
g21363 nand P3_ADD_357_U6 P3_SUB_357_1258_U49 ; P3_SUB_357_1258_U435
g21364 nand P3_SUB_357_1258_U435 P3_SUB_357_1258_U434 ; P3_SUB_357_1258_U436
g21365 nand P3_SUB_357_1258_U140 P3_SUB_357_1258_U141 ; P3_SUB_357_1258_U437
g21366 nand P3_SUB_357_1258_U203 P3_SUB_357_1258_U436 ; P3_SUB_357_1258_U438
g21367 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_SUB_357_1258_U439
g21368 nand P3_ADD_357_U6 P3_SUB_357_1258_U246 ; P3_SUB_357_1258_U440
g21369 nand P3_ADD_357_U6 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_SUB_357_1258_U441
g21370 nand P3_SUB_357_1258_U201 P3_SUB_357_1258_U39 ; P3_SUB_357_1258_U442
g21371 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_SUB_357_1258_U443
g21372 nand P3_ADD_357_U6 P3_SUB_357_1258_U56 ; P3_SUB_357_1258_U444
g21373 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_SUB_357_1258_U445
g21374 nand P3_ADD_357_U6 P3_SUB_357_1258_U56 ; P3_SUB_357_1258_U446
g21375 nand P3_SUB_357_1258_U446 P3_SUB_357_1258_U445 ; P3_SUB_357_1258_U447
g21376 nand P3_SUB_357_1258_U142 P3_SUB_357_1258_U143 ; P3_SUB_357_1258_U448
g21377 nand P3_SUB_357_1258_U200 P3_SUB_357_1258_U447 ; P3_SUB_357_1258_U449
g21378 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_SUB_357_1258_U450
g21379 nand P3_ADD_357_U6 P3_SUB_357_1258_U55 ; P3_SUB_357_1258_U451
g21380 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_SUB_357_1258_U452
g21381 nand P3_ADD_357_U6 P3_SUB_357_1258_U55 ; P3_SUB_357_1258_U453
g21382 nand P3_SUB_357_1258_U453 P3_SUB_357_1258_U452 ; P3_SUB_357_1258_U454
g21383 nand P3_SUB_357_1258_U144 P3_SUB_357_1258_U145 ; P3_SUB_357_1258_U455
g21384 nand P3_SUB_357_1258_U196 P3_SUB_357_1258_U454 ; P3_SUB_357_1258_U456
g21385 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_SUB_357_1258_U457
g21386 nand P3_ADD_357_U6 P3_SUB_357_1258_U54 ; P3_SUB_357_1258_U458
g21387 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_SUB_357_1258_U459
g21388 nand P3_ADD_357_U6 P3_SUB_357_1258_U54 ; P3_SUB_357_1258_U460
g21389 nand P3_SUB_357_1258_U460 P3_SUB_357_1258_U459 ; P3_SUB_357_1258_U461
g21390 nand P3_SUB_357_1258_U146 P3_SUB_357_1258_U147 ; P3_SUB_357_1258_U462
g21391 nand P3_SUB_357_1258_U293 P3_SUB_357_1258_U461 ; P3_SUB_357_1258_U463
g21392 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_SUB_357_1258_U464
g21393 nand P3_ADD_357_U6 P3_SUB_357_1258_U51 ; P3_SUB_357_1258_U465
g21394 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_SUB_357_1258_U466
g21395 nand P3_ADD_357_U6 P3_SUB_357_1258_U50 ; P3_SUB_357_1258_U467
g21396 nand P3_SUB_357_1258_U467 P3_SUB_357_1258_U466 ; P3_SUB_357_1258_U468
g21397 nand P3_SUB_357_1258_U68 P3_SUB_357_1258_U264 ; P3_SUB_357_1258_U469
g21398 nand P3_SUB_357_1258_U468 P3_SUB_357_1258_U291 ; P3_SUB_357_1258_U470
g21399 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_SUB_357_1258_U471
g21400 nand P3_ADD_357_U6 P3_SUB_357_1258_U52 ; P3_SUB_357_1258_U472
g21401 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_SUB_357_1258_U473
g21402 nand P3_ADD_357_U6 P3_SUB_357_1258_U52 ; P3_SUB_357_1258_U474
g21403 nand P3_SUB_357_1258_U474 P3_SUB_357_1258_U473 ; P3_SUB_357_1258_U475
g21404 nand P3_SUB_357_1258_U148 P3_SUB_357_1258_U149 ; P3_SUB_357_1258_U476
g21405 nand P3_SUB_357_1258_U289 P3_SUB_357_1258_U475 ; P3_SUB_357_1258_U477
g21406 nand P3_SUB_357_1258_U39 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_SUB_357_1258_U478
g21407 nand P3_ADD_357_U6 P3_SUB_357_1258_U53 ; P3_SUB_357_1258_U479
g21408 nand P3_SUB_357_1258_U479 P3_SUB_357_1258_U478 ; P3_SUB_357_1258_U480
g21409 nand P3_SUB_357_1258_U150 P3_SUB_357_1258_U265 ; P3_SUB_357_1258_U481
g21410 nand P3_SUB_357_1258_U287 P3_SUB_357_1258_U480 ; P3_SUB_357_1258_U482
g21411 nand P3_SUB_357_1258_U28 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_SUB_357_1258_U483
g21412 nand P3_ADD_357_U10 P3_SUB_357_1258_U29 ; P3_SUB_357_1258_U484
g21413 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_ADD_486_U5
g21414 and P3_ADD_486_U20 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_486_U6
g21415 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_486_U7
g21416 nand P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_ADD_486_U8
g21417 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_486_U9
g21418 nand P3_ADD_486_U18 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_486_U10
g21419 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_486_U11
g21420 nand P3_ADD_486_U19 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_486_U12
g21421 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_486_U13
g21422 nand P3_ADD_486_U22 P3_ADD_486_U21 ; P3_ADD_486_U14
g21423 nand P3_ADD_486_U24 P3_ADD_486_U23 ; P3_ADD_486_U15
g21424 nand P3_ADD_486_U26 P3_ADD_486_U25 ; P3_ADD_486_U16
g21425 nand P3_ADD_486_U28 P3_ADD_486_U27 ; P3_ADD_486_U17
g21426 not P3_ADD_486_U8 ; P3_ADD_486_U18
g21427 not P3_ADD_486_U10 ; P3_ADD_486_U19
g21428 not P3_ADD_486_U12 ; P3_ADD_486_U20
g21429 nand P3_ADD_486_U12 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_486_U21
g21430 nand P3_ADD_486_U20 P3_ADD_486_U13 ; P3_ADD_486_U22
g21431 nand P3_ADD_486_U10 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_486_U23
g21432 nand P3_ADD_486_U19 P3_ADD_486_U11 ; P3_ADD_486_U24
g21433 nand P3_ADD_486_U8 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_486_U25
g21434 nand P3_ADD_486_U18 P3_ADD_486_U9 ; P3_ADD_486_U26
g21435 nand P3_ADD_486_U5 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_486_U27
g21436 nand P3_ADD_486_U7 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_ADD_486_U28
g21437 nand P3_SUB_485_U43 P3_SUB_485_U42 ; P3_SUB_485_U6
g21438 nand P3_SUB_485_U27 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_485_U7
g21439 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_485_U8
g21440 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_485_U9
g21441 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_485_U10
g21442 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_485_U11
g21443 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_485_U12
g21444 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_485_U13
g21445 nand P3_SUB_485_U39 P3_SUB_485_U38 ; P3_SUB_485_U14
g21446 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_485_U15
g21447 nand P3_SUB_485_U48 P3_SUB_485_U47 ; P3_SUB_485_U16
g21448 nand P3_SUB_485_U53 P3_SUB_485_U52 ; P3_SUB_485_U17
g21449 nand P3_SUB_485_U58 P3_SUB_485_U57 ; P3_SUB_485_U18
g21450 nand P3_SUB_485_U63 P3_SUB_485_U62 ; P3_SUB_485_U19
g21451 nand P3_SUB_485_U45 P3_SUB_485_U44 ; P3_SUB_485_U20
g21452 nand P3_SUB_485_U50 P3_SUB_485_U49 ; P3_SUB_485_U21
g21453 nand P3_SUB_485_U55 P3_SUB_485_U54 ; P3_SUB_485_U22
g21454 nand P3_SUB_485_U60 P3_SUB_485_U59 ; P3_SUB_485_U23
g21455 nand P3_SUB_485_U35 P3_SUB_485_U34 ; P3_SUB_485_U24
g21456 nand P3_SUB_485_U31 P3_SUB_485_U30 ; P3_SUB_485_U25
g21457 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_485_U26
g21458 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_485_U27
g21459 not P3_SUB_485_U7 ; P3_SUB_485_U28
g21460 nand P3_SUB_485_U28 P3_SUB_485_U8 ; P3_SUB_485_U29
g21461 nand P3_SUB_485_U29 P3_SUB_485_U26 ; P3_SUB_485_U30
g21462 nand P3_SUB_485_U7 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_485_U31
g21463 not P3_SUB_485_U25 ; P3_SUB_485_U32
g21464 nand P3_SUB_485_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_485_U33
g21465 nand P3_SUB_485_U33 P3_SUB_485_U25 ; P3_SUB_485_U34
g21466 nand P3_SUB_485_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_485_U35
g21467 not P3_SUB_485_U24 ; P3_SUB_485_U36
g21468 nand P3_SUB_485_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_485_U37
g21469 nand P3_SUB_485_U37 P3_SUB_485_U24 ; P3_SUB_485_U38
g21470 nand P3_SUB_485_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_485_U39
g21471 not P3_SUB_485_U14 ; P3_SUB_485_U40
g21472 nand P3_SUB_485_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_485_U41
g21473 nand P3_SUB_485_U40 P3_SUB_485_U41 ; P3_SUB_485_U42
g21474 nand P3_SUB_485_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_485_U43
g21475 nand P3_SUB_485_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_485_U44
g21476 nand P3_SUB_485_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_485_U45
g21477 not P3_SUB_485_U20 ; P3_SUB_485_U46
g21478 nand P3_SUB_485_U46 P3_SUB_485_U40 ; P3_SUB_485_U47
g21479 nand P3_SUB_485_U20 P3_SUB_485_U14 ; P3_SUB_485_U48
g21480 nand P3_SUB_485_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_485_U49
g21481 nand P3_SUB_485_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_485_U50
g21482 not P3_SUB_485_U21 ; P3_SUB_485_U51
g21483 nand P3_SUB_485_U36 P3_SUB_485_U51 ; P3_SUB_485_U52
g21484 nand P3_SUB_485_U21 P3_SUB_485_U24 ; P3_SUB_485_U53
g21485 nand P3_SUB_485_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_485_U54
g21486 nand P3_SUB_485_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_485_U55
g21487 not P3_SUB_485_U22 ; P3_SUB_485_U56
g21488 nand P3_SUB_485_U32 P3_SUB_485_U56 ; P3_SUB_485_U57
g21489 nand P3_SUB_485_U22 P3_SUB_485_U25 ; P3_SUB_485_U58
g21490 nand P3_SUB_485_U8 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_485_U59
g21491 nand P3_SUB_485_U26 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_485_U60
g21492 not P3_SUB_485_U23 ; P3_SUB_485_U61
g21493 nand P3_SUB_485_U61 P3_SUB_485_U28 ; P3_SUB_485_U62
g21494 nand P3_SUB_485_U23 P3_SUB_485_U7 ; P3_SUB_485_U63
g21495 not P3_U3305 ; P3_SUB_563_U6
g21496 not P3_U3306 ; P3_SUB_563_U7
g21497 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_515_U4
g21498 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_515_U5
g21499 nand P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_515_U6
g21500 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_515_U7
g21501 nand P3_ADD_515_U94 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_515_U8
g21502 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_515_U9
g21503 nand P3_ADD_515_U95 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_515_U10
g21504 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_515_U11
g21505 nand P3_ADD_515_U96 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_515_U12
g21506 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_515_U13
g21507 nand P3_ADD_515_U97 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_515_U14
g21508 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_515_U15
g21509 nand P3_ADD_515_U98 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_515_U16
g21510 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_515_U17
g21511 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_515_U18
g21512 nand P3_ADD_515_U99 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_515_U19
g21513 nand P3_ADD_515_U100 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_515_U20
g21514 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_515_U21
g21515 nand P3_ADD_515_U101 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_515_U22
g21516 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_515_U23
g21517 nand P3_ADD_515_U102 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_515_U24
g21518 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_515_U25
g21519 nand P3_ADD_515_U103 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_515_U26
g21520 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_515_U27
g21521 nand P3_ADD_515_U104 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_515_U28
g21522 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_515_U29
g21523 nand P3_ADD_515_U105 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_515_U30
g21524 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_515_U31
g21525 nand P3_ADD_515_U106 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_515_U32
g21526 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_515_U33
g21527 nand P3_ADD_515_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_515_U34
g21528 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_515_U35
g21529 nand P3_ADD_515_U108 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_515_U36
g21530 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_515_U37
g21531 nand P3_ADD_515_U109 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_515_U38
g21532 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_515_U39
g21533 nand P3_ADD_515_U110 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_515_U40
g21534 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_515_U41
g21535 nand P3_ADD_515_U111 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_515_U42
g21536 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_515_U43
g21537 nand P3_ADD_515_U112 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_515_U44
g21538 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_515_U45
g21539 nand P3_ADD_515_U113 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_515_U46
g21540 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_515_U47
g21541 nand P3_ADD_515_U114 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_515_U48
g21542 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_515_U49
g21543 nand P3_ADD_515_U115 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_515_U50
g21544 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_515_U51
g21545 nand P3_ADD_515_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_515_U52
g21546 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_515_U53
g21547 nand P3_ADD_515_U117 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_515_U54
g21548 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_515_U55
g21549 nand P3_ADD_515_U118 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_515_U56
g21550 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_515_U57
g21551 nand P3_ADD_515_U119 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_515_U58
g21552 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_515_U59
g21553 nand P3_ADD_515_U120 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_515_U60
g21554 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_515_U61
g21555 nand P3_ADD_515_U124 P3_ADD_515_U123 ; P3_ADD_515_U62
g21556 nand P3_ADD_515_U126 P3_ADD_515_U125 ; P3_ADD_515_U63
g21557 nand P3_ADD_515_U128 P3_ADD_515_U127 ; P3_ADD_515_U64
g21558 nand P3_ADD_515_U130 P3_ADD_515_U129 ; P3_ADD_515_U65
g21559 nand P3_ADD_515_U132 P3_ADD_515_U131 ; P3_ADD_515_U66
g21560 nand P3_ADD_515_U134 P3_ADD_515_U133 ; P3_ADD_515_U67
g21561 nand P3_ADD_515_U136 P3_ADD_515_U135 ; P3_ADD_515_U68
g21562 nand P3_ADD_515_U138 P3_ADD_515_U137 ; P3_ADD_515_U69
g21563 nand P3_ADD_515_U140 P3_ADD_515_U139 ; P3_ADD_515_U70
g21564 nand P3_ADD_515_U142 P3_ADD_515_U141 ; P3_ADD_515_U71
g21565 nand P3_ADD_515_U144 P3_ADD_515_U143 ; P3_ADD_515_U72
g21566 nand P3_ADD_515_U146 P3_ADD_515_U145 ; P3_ADD_515_U73
g21567 nand P3_ADD_515_U148 P3_ADD_515_U147 ; P3_ADD_515_U74
g21568 nand P3_ADD_515_U150 P3_ADD_515_U149 ; P3_ADD_515_U75
g21569 nand P3_ADD_515_U152 P3_ADD_515_U151 ; P3_ADD_515_U76
g21570 nand P3_ADD_515_U154 P3_ADD_515_U153 ; P3_ADD_515_U77
g21571 nand P3_ADD_515_U156 P3_ADD_515_U155 ; P3_ADD_515_U78
g21572 nand P3_ADD_515_U158 P3_ADD_515_U157 ; P3_ADD_515_U79
g21573 nand P3_ADD_515_U160 P3_ADD_515_U159 ; P3_ADD_515_U80
g21574 nand P3_ADD_515_U162 P3_ADD_515_U161 ; P3_ADD_515_U81
g21575 nand P3_ADD_515_U164 P3_ADD_515_U163 ; P3_ADD_515_U82
g21576 nand P3_ADD_515_U166 P3_ADD_515_U165 ; P3_ADD_515_U83
g21577 nand P3_ADD_515_U168 P3_ADD_515_U167 ; P3_ADD_515_U84
g21578 nand P3_ADD_515_U170 P3_ADD_515_U169 ; P3_ADD_515_U85
g21579 nand P3_ADD_515_U172 P3_ADD_515_U171 ; P3_ADD_515_U86
g21580 nand P3_ADD_515_U174 P3_ADD_515_U173 ; P3_ADD_515_U87
g21581 nand P3_ADD_515_U176 P3_ADD_515_U175 ; P3_ADD_515_U88
g21582 nand P3_ADD_515_U178 P3_ADD_515_U177 ; P3_ADD_515_U89
g21583 nand P3_ADD_515_U180 P3_ADD_515_U179 ; P3_ADD_515_U90
g21584 nand P3_ADD_515_U182 P3_ADD_515_U181 ; P3_ADD_515_U91
g21585 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_515_U92
g21586 nand P3_ADD_515_U121 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_515_U93
g21587 not P3_ADD_515_U6 ; P3_ADD_515_U94
g21588 not P3_ADD_515_U8 ; P3_ADD_515_U95
g21589 not P3_ADD_515_U10 ; P3_ADD_515_U96
g21590 not P3_ADD_515_U12 ; P3_ADD_515_U97
g21591 not P3_ADD_515_U14 ; P3_ADD_515_U98
g21592 not P3_ADD_515_U16 ; P3_ADD_515_U99
g21593 not P3_ADD_515_U19 ; P3_ADD_515_U100
g21594 not P3_ADD_515_U20 ; P3_ADD_515_U101
g21595 not P3_ADD_515_U22 ; P3_ADD_515_U102
g21596 not P3_ADD_515_U24 ; P3_ADD_515_U103
g21597 not P3_ADD_515_U26 ; P3_ADD_515_U104
g21598 not P3_ADD_515_U28 ; P3_ADD_515_U105
g21599 not P3_ADD_515_U30 ; P3_ADD_515_U106
g21600 not P3_ADD_515_U32 ; P3_ADD_515_U107
g21601 not P3_ADD_515_U34 ; P3_ADD_515_U108
g21602 not P3_ADD_515_U36 ; P3_ADD_515_U109
g21603 not P3_ADD_515_U38 ; P3_ADD_515_U110
g21604 not P3_ADD_515_U40 ; P3_ADD_515_U111
g21605 not P3_ADD_515_U42 ; P3_ADD_515_U112
g21606 not P3_ADD_515_U44 ; P3_ADD_515_U113
g21607 not P3_ADD_515_U46 ; P3_ADD_515_U114
g21608 not P3_ADD_515_U48 ; P3_ADD_515_U115
g21609 not P3_ADD_515_U50 ; P3_ADD_515_U116
g21610 not P3_ADD_515_U52 ; P3_ADD_515_U117
g21611 not P3_ADD_515_U54 ; P3_ADD_515_U118
g21612 not P3_ADD_515_U56 ; P3_ADD_515_U119
g21613 not P3_ADD_515_U58 ; P3_ADD_515_U120
g21614 not P3_ADD_515_U60 ; P3_ADD_515_U121
g21615 not P3_ADD_515_U93 ; P3_ADD_515_U122
g21616 nand P3_ADD_515_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_515_U123
g21617 nand P3_ADD_515_U100 P3_ADD_515_U18 ; P3_ADD_515_U124
g21618 nand P3_ADD_515_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_515_U125
g21619 nand P3_ADD_515_U99 P3_ADD_515_U17 ; P3_ADD_515_U126
g21620 nand P3_ADD_515_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_515_U127
g21621 nand P3_ADD_515_U98 P3_ADD_515_U15 ; P3_ADD_515_U128
g21622 nand P3_ADD_515_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_515_U129
g21623 nand P3_ADD_515_U97 P3_ADD_515_U13 ; P3_ADD_515_U130
g21624 nand P3_ADD_515_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_515_U131
g21625 nand P3_ADD_515_U96 P3_ADD_515_U11 ; P3_ADD_515_U132
g21626 nand P3_ADD_515_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_515_U133
g21627 nand P3_ADD_515_U95 P3_ADD_515_U9 ; P3_ADD_515_U134
g21628 nand P3_ADD_515_U6 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_515_U135
g21629 nand P3_ADD_515_U94 P3_ADD_515_U7 ; P3_ADD_515_U136
g21630 nand P3_ADD_515_U93 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_515_U137
g21631 nand P3_ADD_515_U122 P3_ADD_515_U92 ; P3_ADD_515_U138
g21632 nand P3_ADD_515_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_515_U139
g21633 nand P3_ADD_515_U121 P3_ADD_515_U61 ; P3_ADD_515_U140
g21634 nand P3_ADD_515_U4 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_515_U141
g21635 nand P3_ADD_515_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_515_U142
g21636 nand P3_ADD_515_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_515_U143
g21637 nand P3_ADD_515_U120 P3_ADD_515_U59 ; P3_ADD_515_U144
g21638 nand P3_ADD_515_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_515_U145
g21639 nand P3_ADD_515_U119 P3_ADD_515_U57 ; P3_ADD_515_U146
g21640 nand P3_ADD_515_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_515_U147
g21641 nand P3_ADD_515_U118 P3_ADD_515_U55 ; P3_ADD_515_U148
g21642 nand P3_ADD_515_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_515_U149
g21643 nand P3_ADD_515_U117 P3_ADD_515_U53 ; P3_ADD_515_U150
g21644 nand P3_ADD_515_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_515_U151
g21645 nand P3_ADD_515_U116 P3_ADD_515_U51 ; P3_ADD_515_U152
g21646 nand P3_ADD_515_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_515_U153
g21647 nand P3_ADD_515_U115 P3_ADD_515_U49 ; P3_ADD_515_U154
g21648 nand P3_ADD_515_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_515_U155
g21649 nand P3_ADD_515_U114 P3_ADD_515_U47 ; P3_ADD_515_U156
g21650 nand P3_ADD_515_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_515_U157
g21651 nand P3_ADD_515_U113 P3_ADD_515_U45 ; P3_ADD_515_U158
g21652 nand P3_ADD_515_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_515_U159
g21653 nand P3_ADD_515_U112 P3_ADD_515_U43 ; P3_ADD_515_U160
g21654 nand P3_ADD_515_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_515_U161
g21655 nand P3_ADD_515_U111 P3_ADD_515_U41 ; P3_ADD_515_U162
g21656 nand P3_ADD_515_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_515_U163
g21657 nand P3_ADD_515_U110 P3_ADD_515_U39 ; P3_ADD_515_U164
g21658 nand P3_ADD_515_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_515_U165
g21659 nand P3_ADD_515_U109 P3_ADD_515_U37 ; P3_ADD_515_U166
g21660 nand P3_ADD_515_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_515_U167
g21661 nand P3_ADD_515_U108 P3_ADD_515_U35 ; P3_ADD_515_U168
g21662 nand P3_ADD_515_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_515_U169
g21663 nand P3_ADD_515_U107 P3_ADD_515_U33 ; P3_ADD_515_U170
g21664 nand P3_ADD_515_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_515_U171
g21665 nand P3_ADD_515_U106 P3_ADD_515_U31 ; P3_ADD_515_U172
g21666 nand P3_ADD_515_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_515_U173
g21667 nand P3_ADD_515_U105 P3_ADD_515_U29 ; P3_ADD_515_U174
g21668 nand P3_ADD_515_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_515_U175
g21669 nand P3_ADD_515_U104 P3_ADD_515_U27 ; P3_ADD_515_U176
g21670 nand P3_ADD_515_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_515_U177
g21671 nand P3_ADD_515_U103 P3_ADD_515_U25 ; P3_ADD_515_U178
g21672 nand P3_ADD_515_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_515_U179
g21673 nand P3_ADD_515_U102 P3_ADD_515_U23 ; P3_ADD_515_U180
g21674 nand P3_ADD_515_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_515_U181
g21675 nand P3_ADD_515_U101 P3_ADD_515_U21 ; P3_ADD_515_U182
g21676 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_394_U4
g21677 nand P3_ADD_394_U92 P3_ADD_394_U126 ; P3_ADD_394_U5
g21678 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_394_U6
g21679 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_394_U7
g21680 nand P3_ADD_394_U92 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_394_U8
g21681 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_394_U9
g21682 nand P3_ADD_394_U98 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_394_U10
g21683 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_394_U11
g21684 nand P3_ADD_394_U99 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_394_U12
g21685 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_394_U13
g21686 nand P3_ADD_394_U100 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_394_U14
g21687 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_394_U15
g21688 nand P3_ADD_394_U101 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_394_U16
g21689 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_394_U17
g21690 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_394_U18
g21691 nand P3_ADD_394_U102 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_394_U19
g21692 nand P3_ADD_394_U103 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_394_U20
g21693 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_394_U21
g21694 nand P3_ADD_394_U104 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_394_U22
g21695 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_394_U23
g21696 nand P3_ADD_394_U105 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_394_U24
g21697 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_394_U25
g21698 nand P3_ADD_394_U106 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_394_U26
g21699 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_394_U27
g21700 nand P3_ADD_394_U107 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_394_U28
g21701 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_394_U29
g21702 nand P3_ADD_394_U108 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_394_U30
g21703 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_394_U31
g21704 nand P3_ADD_394_U109 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_394_U32
g21705 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_394_U33
g21706 nand P3_ADD_394_U110 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_394_U34
g21707 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_394_U35
g21708 nand P3_ADD_394_U111 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_394_U36
g21709 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_394_U37
g21710 nand P3_ADD_394_U112 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_394_U38
g21711 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_394_U39
g21712 nand P3_ADD_394_U113 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_394_U40
g21713 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_394_U41
g21714 nand P3_ADD_394_U114 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_394_U42
g21715 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_394_U43
g21716 nand P3_ADD_394_U115 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_394_U44
g21717 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_394_U45
g21718 nand P3_ADD_394_U116 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_394_U46
g21719 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_394_U47
g21720 nand P3_ADD_394_U117 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_394_U48
g21721 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_394_U49
g21722 nand P3_ADD_394_U118 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_394_U50
g21723 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_394_U51
g21724 nand P3_ADD_394_U119 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_394_U52
g21725 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_394_U53
g21726 nand P3_ADD_394_U120 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_394_U54
g21727 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_394_U55
g21728 nand P3_ADD_394_U121 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_394_U56
g21729 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_394_U57
g21730 nand P3_ADD_394_U122 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_394_U58
g21731 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_394_U59
g21732 nand P3_ADD_394_U123 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_394_U60
g21733 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_394_U61
g21734 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_394_U62
g21735 nand P3_ADD_394_U128 P3_ADD_394_U127 ; P3_ADD_394_U63
g21736 nand P3_ADD_394_U130 P3_ADD_394_U129 ; P3_ADD_394_U64
g21737 nand P3_ADD_394_U132 P3_ADD_394_U131 ; P3_ADD_394_U65
g21738 nand P3_ADD_394_U134 P3_ADD_394_U133 ; P3_ADD_394_U66
g21739 nand P3_ADD_394_U136 P3_ADD_394_U135 ; P3_ADD_394_U67
g21740 nand P3_ADD_394_U138 P3_ADD_394_U137 ; P3_ADD_394_U68
g21741 nand P3_ADD_394_U142 P3_ADD_394_U141 ; P3_ADD_394_U69
g21742 nand P3_ADD_394_U144 P3_ADD_394_U143 ; P3_ADD_394_U70
g21743 nand P3_ADD_394_U146 P3_ADD_394_U145 ; P3_ADD_394_U71
g21744 nand P3_ADD_394_U148 P3_ADD_394_U147 ; P3_ADD_394_U72
g21745 nand P3_ADD_394_U150 P3_ADD_394_U149 ; P3_ADD_394_U73
g21746 nand P3_ADD_394_U152 P3_ADD_394_U151 ; P3_ADD_394_U74
g21747 nand P3_ADD_394_U154 P3_ADD_394_U153 ; P3_ADD_394_U75
g21748 nand P3_ADD_394_U156 P3_ADD_394_U155 ; P3_ADD_394_U76
g21749 nand P3_ADD_394_U158 P3_ADD_394_U157 ; P3_ADD_394_U77
g21750 nand P3_ADD_394_U160 P3_ADD_394_U159 ; P3_ADD_394_U78
g21751 nand P3_ADD_394_U162 P3_ADD_394_U161 ; P3_ADD_394_U79
g21752 nand P3_ADD_394_U164 P3_ADD_394_U163 ; P3_ADD_394_U80
g21753 nand P3_ADD_394_U166 P3_ADD_394_U165 ; P3_ADD_394_U81
g21754 nand P3_ADD_394_U168 P3_ADD_394_U167 ; P3_ADD_394_U82
g21755 nand P3_ADD_394_U170 P3_ADD_394_U169 ; P3_ADD_394_U83
g21756 nand P3_ADD_394_U172 P3_ADD_394_U171 ; P3_ADD_394_U84
g21757 nand P3_ADD_394_U174 P3_ADD_394_U173 ; P3_ADD_394_U85
g21758 nand P3_ADD_394_U176 P3_ADD_394_U175 ; P3_ADD_394_U86
g21759 nand P3_ADD_394_U178 P3_ADD_394_U177 ; P3_ADD_394_U87
g21760 nand P3_ADD_394_U180 P3_ADD_394_U179 ; P3_ADD_394_U88
g21761 nand P3_ADD_394_U182 P3_ADD_394_U181 ; P3_ADD_394_U89
g21762 nand P3_ADD_394_U184 P3_ADD_394_U183 ; P3_ADD_394_U90
g21763 nand P3_ADD_394_U186 P3_ADD_394_U185 ; P3_ADD_394_U91
g21764 nand P3_ADD_394_U62 P3_ADD_394_U96 ; P3_ADD_394_U92
g21765 and P3_ADD_394_U140 P3_ADD_394_U139 ; P3_ADD_394_U93
g21766 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_394_U94
g21767 nand P3_ADD_394_U124 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_394_U95
g21768 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_394_U96
g21769 not P3_ADD_394_U92 ; P3_ADD_394_U97
g21770 not P3_ADD_394_U8 ; P3_ADD_394_U98
g21771 not P3_ADD_394_U10 ; P3_ADD_394_U99
g21772 not P3_ADD_394_U12 ; P3_ADD_394_U100
g21773 not P3_ADD_394_U14 ; P3_ADD_394_U101
g21774 not P3_ADD_394_U16 ; P3_ADD_394_U102
g21775 not P3_ADD_394_U19 ; P3_ADD_394_U103
g21776 not P3_ADD_394_U20 ; P3_ADD_394_U104
g21777 not P3_ADD_394_U22 ; P3_ADD_394_U105
g21778 not P3_ADD_394_U24 ; P3_ADD_394_U106
g21779 not P3_ADD_394_U26 ; P3_ADD_394_U107
g21780 not P3_ADD_394_U28 ; P3_ADD_394_U108
g21781 not P3_ADD_394_U30 ; P3_ADD_394_U109
g21782 not P3_ADD_394_U32 ; P3_ADD_394_U110
g21783 not P3_ADD_394_U34 ; P3_ADD_394_U111
g21784 not P3_ADD_394_U36 ; P3_ADD_394_U112
g21785 not P3_ADD_394_U38 ; P3_ADD_394_U113
g21786 not P3_ADD_394_U40 ; P3_ADD_394_U114
g21787 not P3_ADD_394_U42 ; P3_ADD_394_U115
g21788 not P3_ADD_394_U44 ; P3_ADD_394_U116
g21789 not P3_ADD_394_U46 ; P3_ADD_394_U117
g21790 not P3_ADD_394_U48 ; P3_ADD_394_U118
g21791 not P3_ADD_394_U50 ; P3_ADD_394_U119
g21792 not P3_ADD_394_U52 ; P3_ADD_394_U120
g21793 not P3_ADD_394_U54 ; P3_ADD_394_U121
g21794 not P3_ADD_394_U56 ; P3_ADD_394_U122
g21795 not P3_ADD_394_U58 ; P3_ADD_394_U123
g21796 not P3_ADD_394_U60 ; P3_ADD_394_U124
g21797 not P3_ADD_394_U95 ; P3_ADD_394_U125
g21798 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_394_U126
g21799 nand P3_ADD_394_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_394_U127
g21800 nand P3_ADD_394_U103 P3_ADD_394_U18 ; P3_ADD_394_U128
g21801 nand P3_ADD_394_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_394_U129
g21802 nand P3_ADD_394_U102 P3_ADD_394_U17 ; P3_ADD_394_U130
g21803 nand P3_ADD_394_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_394_U131
g21804 nand P3_ADD_394_U101 P3_ADD_394_U15 ; P3_ADD_394_U132
g21805 nand P3_ADD_394_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_394_U133
g21806 nand P3_ADD_394_U100 P3_ADD_394_U13 ; P3_ADD_394_U134
g21807 nand P3_ADD_394_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_394_U135
g21808 nand P3_ADD_394_U99 P3_ADD_394_U11 ; P3_ADD_394_U136
g21809 nand P3_ADD_394_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_394_U137
g21810 nand P3_ADD_394_U98 P3_ADD_394_U9 ; P3_ADD_394_U138
g21811 nand P3_ADD_394_U92 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_394_U139
g21812 nand P3_ADD_394_U97 P3_ADD_394_U7 ; P3_ADD_394_U140
g21813 nand P3_ADD_394_U95 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_394_U141
g21814 nand P3_ADD_394_U125 P3_ADD_394_U94 ; P3_ADD_394_U142
g21815 nand P3_ADD_394_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_394_U143
g21816 nand P3_ADD_394_U124 P3_ADD_394_U61 ; P3_ADD_394_U144
g21817 nand P3_ADD_394_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_394_U145
g21818 nand P3_ADD_394_U123 P3_ADD_394_U59 ; P3_ADD_394_U146
g21819 nand P3_ADD_394_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_394_U147
g21820 nand P3_ADD_394_U122 P3_ADD_394_U57 ; P3_ADD_394_U148
g21821 nand P3_ADD_394_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_394_U149
g21822 nand P3_ADD_394_U121 P3_ADD_394_U55 ; P3_ADD_394_U150
g21823 nand P3_ADD_394_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_394_U151
g21824 nand P3_ADD_394_U120 P3_ADD_394_U53 ; P3_ADD_394_U152
g21825 nand P3_ADD_394_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_394_U153
g21826 nand P3_ADD_394_U119 P3_ADD_394_U51 ; P3_ADD_394_U154
g21827 nand P3_ADD_394_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_394_U155
g21828 nand P3_ADD_394_U118 P3_ADD_394_U49 ; P3_ADD_394_U156
g21829 nand P3_ADD_394_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_394_U157
g21830 nand P3_ADD_394_U117 P3_ADD_394_U47 ; P3_ADD_394_U158
g21831 nand P3_ADD_394_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_394_U159
g21832 nand P3_ADD_394_U116 P3_ADD_394_U45 ; P3_ADD_394_U160
g21833 nand P3_ADD_394_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_394_U161
g21834 nand P3_ADD_394_U115 P3_ADD_394_U43 ; P3_ADD_394_U162
g21835 nand P3_ADD_394_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_394_U163
g21836 nand P3_ADD_394_U114 P3_ADD_394_U41 ; P3_ADD_394_U164
g21837 nand P3_ADD_394_U4 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_394_U165
g21838 nand P3_ADD_394_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_394_U166
g21839 nand P3_ADD_394_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_394_U167
g21840 nand P3_ADD_394_U113 P3_ADD_394_U39 ; P3_ADD_394_U168
g21841 nand P3_ADD_394_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_394_U169
g21842 nand P3_ADD_394_U112 P3_ADD_394_U37 ; P3_ADD_394_U170
g21843 nand P3_ADD_394_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_394_U171
g21844 nand P3_ADD_394_U111 P3_ADD_394_U35 ; P3_ADD_394_U172
g21845 nand P3_ADD_394_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_394_U173
g21846 nand P3_ADD_394_U110 P3_ADD_394_U33 ; P3_ADD_394_U174
g21847 nand P3_ADD_394_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_394_U175
g21848 nand P3_ADD_394_U109 P3_ADD_394_U31 ; P3_ADD_394_U176
g21849 nand P3_ADD_394_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_394_U177
g21850 nand P3_ADD_394_U108 P3_ADD_394_U29 ; P3_ADD_394_U178
g21851 nand P3_ADD_394_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_394_U179
g21852 nand P3_ADD_394_U107 P3_ADD_394_U27 ; P3_ADD_394_U180
g21853 nand P3_ADD_394_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_394_U181
g21854 nand P3_ADD_394_U106 P3_ADD_394_U25 ; P3_ADD_394_U182
g21855 nand P3_ADD_394_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_394_U183
g21856 nand P3_ADD_394_U105 P3_ADD_394_U23 ; P3_ADD_394_U184
g21857 nand P3_ADD_394_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_394_U185
g21858 nand P3_ADD_394_U104 P3_ADD_394_U21 ; P3_ADD_394_U186
g21859 nor P3_SUB_450_U6 P3_GTE_450_U7 ; P3_GTE_450_U6
g21860 nor P3_SUB_450_U16 P3_SUB_450_U17 P3_SUB_450_U19 P3_SUB_450_U18 ; P3_GTE_450_U7
g21861 and P3_SUB_414_U126 P3_SUB_414_U28 ; P3_SUB_414_U6
g21862 and P3_SUB_414_U124 P3_SUB_414_U29 ; P3_SUB_414_U7
g21863 and P3_SUB_414_U122 P3_SUB_414_U30 ; P3_SUB_414_U8
g21864 and P3_SUB_414_U120 P3_SUB_414_U31 ; P3_SUB_414_U9
g21865 and P3_SUB_414_U118 P3_SUB_414_U32 ; P3_SUB_414_U10
g21866 and P3_SUB_414_U116 P3_SUB_414_U33 ; P3_SUB_414_U11
g21867 and P3_SUB_414_U114 P3_SUB_414_U34 ; P3_SUB_414_U12
g21868 and P3_SUB_414_U112 P3_SUB_414_U35 ; P3_SUB_414_U13
g21869 and P3_SUB_414_U110 P3_SUB_414_U36 ; P3_SUB_414_U14
g21870 and P3_SUB_414_U108 P3_SUB_414_U37 ; P3_SUB_414_U15
g21871 and P3_SUB_414_U106 P3_SUB_414_U38 ; P3_SUB_414_U16
g21872 and P3_SUB_414_U105 P3_SUB_414_U21 ; P3_SUB_414_U17
g21873 and P3_SUB_414_U92 P3_SUB_414_U22 ; P3_SUB_414_U18
g21874 and P3_SUB_414_U90 P3_SUB_414_U23 ; P3_SUB_414_U19
g21875 and P3_SUB_414_U88 P3_SUB_414_U24 ; P3_SUB_414_U20
g21876 or P3_EBX_REG_0__SCAN_IN P3_EBX_REG_1__SCAN_IN P3_EBX_REG_2__SCAN_IN ; P3_SUB_414_U21
g21877 nand P3_SUB_414_U27 P3_SUB_414_U58 P3_SUB_414_U83 ; P3_SUB_414_U22
g21878 nand P3_SUB_414_U26 P3_SUB_414_U56 P3_SUB_414_U84 ; P3_SUB_414_U23
g21879 nand P3_SUB_414_U25 P3_SUB_414_U54 P3_SUB_414_U85 ; P3_SUB_414_U24
g21880 not P3_EBX_REG_8__SCAN_IN ; P3_SUB_414_U25
g21881 not P3_EBX_REG_6__SCAN_IN ; P3_SUB_414_U26
g21882 not P3_EBX_REG_4__SCAN_IN ; P3_SUB_414_U27
g21883 nand P3_SUB_414_U52 P3_SUB_414_U49 P3_SUB_414_U86 ; P3_SUB_414_U28
g21884 nand P3_SUB_414_U48 P3_SUB_414_U81 P3_SUB_414_U93 ; P3_SUB_414_U29
g21885 nand P3_SUB_414_U47 P3_SUB_414_U79 P3_SUB_414_U94 ; P3_SUB_414_U30
g21886 nand P3_SUB_414_U46 P3_SUB_414_U77 P3_SUB_414_U95 ; P3_SUB_414_U31
g21887 nand P3_SUB_414_U45 P3_SUB_414_U75 P3_SUB_414_U96 ; P3_SUB_414_U32
g21888 nand P3_SUB_414_U44 P3_SUB_414_U73 P3_SUB_414_U97 ; P3_SUB_414_U33
g21889 nand P3_SUB_414_U43 P3_SUB_414_U69 P3_SUB_414_U98 ; P3_SUB_414_U34
g21890 nand P3_SUB_414_U42 P3_SUB_414_U67 P3_SUB_414_U99 ; P3_SUB_414_U35
g21891 nand P3_SUB_414_U41 P3_SUB_414_U65 P3_SUB_414_U100 ; P3_SUB_414_U36
g21892 nand P3_SUB_414_U40 P3_SUB_414_U63 P3_SUB_414_U101 ; P3_SUB_414_U37
g21893 nand P3_SUB_414_U102 P3_SUB_414_U39 ; P3_SUB_414_U38
g21894 not P3_EBX_REG_29__SCAN_IN ; P3_SUB_414_U39
g21895 not P3_EBX_REG_28__SCAN_IN ; P3_SUB_414_U40
g21896 not P3_EBX_REG_26__SCAN_IN ; P3_SUB_414_U41
g21897 not P3_EBX_REG_24__SCAN_IN ; P3_SUB_414_U42
g21898 not P3_EBX_REG_22__SCAN_IN ; P3_SUB_414_U43
g21899 not P3_EBX_REG_20__SCAN_IN ; P3_SUB_414_U44
g21900 not P3_EBX_REG_18__SCAN_IN ; P3_SUB_414_U45
g21901 not P3_EBX_REG_16__SCAN_IN ; P3_SUB_414_U46
g21902 not P3_EBX_REG_14__SCAN_IN ; P3_SUB_414_U47
g21903 not P3_EBX_REG_12__SCAN_IN ; P3_SUB_414_U48
g21904 not P3_EBX_REG_10__SCAN_IN ; P3_SUB_414_U49
g21905 nand P3_SUB_414_U149 P3_SUB_414_U148 ; P3_SUB_414_U50
g21906 nand P3_SUB_414_U137 P3_SUB_414_U136 ; P3_SUB_414_U51
g21907 not P3_EBX_REG_9__SCAN_IN ; P3_SUB_414_U52
g21908 and P3_SUB_414_U129 P3_SUB_414_U128 ; P3_SUB_414_U53
g21909 not P3_EBX_REG_7__SCAN_IN ; P3_SUB_414_U54
g21910 and P3_SUB_414_U131 P3_SUB_414_U130 ; P3_SUB_414_U55
g21911 not P3_EBX_REG_5__SCAN_IN ; P3_SUB_414_U56
g21912 and P3_SUB_414_U133 P3_SUB_414_U132 ; P3_SUB_414_U57
g21913 not P3_EBX_REG_3__SCAN_IN ; P3_SUB_414_U58
g21914 and P3_SUB_414_U135 P3_SUB_414_U134 ; P3_SUB_414_U59
g21915 not P3_EBX_REG_31__SCAN_IN ; P3_SUB_414_U60
g21916 not P3_EBX_REG_30__SCAN_IN ; P3_SUB_414_U61
g21917 and P3_SUB_414_U139 P3_SUB_414_U138 ; P3_SUB_414_U62
g21918 not P3_EBX_REG_27__SCAN_IN ; P3_SUB_414_U63
g21919 and P3_SUB_414_U141 P3_SUB_414_U140 ; P3_SUB_414_U64
g21920 not P3_EBX_REG_25__SCAN_IN ; P3_SUB_414_U65
g21921 and P3_SUB_414_U143 P3_SUB_414_U142 ; P3_SUB_414_U66
g21922 not P3_EBX_REG_23__SCAN_IN ; P3_SUB_414_U67
g21923 and P3_SUB_414_U145 P3_SUB_414_U144 ; P3_SUB_414_U68
g21924 not P3_EBX_REG_21__SCAN_IN ; P3_SUB_414_U69
g21925 and P3_SUB_414_U147 P3_SUB_414_U146 ; P3_SUB_414_U70
g21926 not P3_EBX_REG_1__SCAN_IN ; P3_SUB_414_U71
g21927 not P3_EBX_REG_0__SCAN_IN ; P3_SUB_414_U72
g21928 not P3_EBX_REG_19__SCAN_IN ; P3_SUB_414_U73
g21929 and P3_SUB_414_U151 P3_SUB_414_U150 ; P3_SUB_414_U74
g21930 not P3_EBX_REG_17__SCAN_IN ; P3_SUB_414_U75
g21931 and P3_SUB_414_U153 P3_SUB_414_U152 ; P3_SUB_414_U76
g21932 not P3_EBX_REG_15__SCAN_IN ; P3_SUB_414_U77
g21933 and P3_SUB_414_U155 P3_SUB_414_U154 ; P3_SUB_414_U78
g21934 not P3_EBX_REG_13__SCAN_IN ; P3_SUB_414_U79
g21935 and P3_SUB_414_U157 P3_SUB_414_U156 ; P3_SUB_414_U80
g21936 not P3_EBX_REG_11__SCAN_IN ; P3_SUB_414_U81
g21937 and P3_SUB_414_U159 P3_SUB_414_U158 ; P3_SUB_414_U82
g21938 not P3_SUB_414_U21 ; P3_SUB_414_U83
g21939 not P3_SUB_414_U22 ; P3_SUB_414_U84
g21940 not P3_SUB_414_U23 ; P3_SUB_414_U85
g21941 not P3_SUB_414_U24 ; P3_SUB_414_U86
g21942 nand P3_SUB_414_U85 P3_SUB_414_U54 ; P3_SUB_414_U87
g21943 nand P3_SUB_414_U87 P3_EBX_REG_8__SCAN_IN ; P3_SUB_414_U88
g21944 nand P3_SUB_414_U84 P3_SUB_414_U56 ; P3_SUB_414_U89
g21945 nand P3_SUB_414_U89 P3_EBX_REG_6__SCAN_IN ; P3_SUB_414_U90
g21946 nand P3_SUB_414_U83 P3_SUB_414_U58 ; P3_SUB_414_U91
g21947 nand P3_SUB_414_U91 P3_EBX_REG_4__SCAN_IN ; P3_SUB_414_U92
g21948 not P3_SUB_414_U28 ; P3_SUB_414_U93
g21949 not P3_SUB_414_U29 ; P3_SUB_414_U94
g21950 not P3_SUB_414_U30 ; P3_SUB_414_U95
g21951 not P3_SUB_414_U31 ; P3_SUB_414_U96
g21952 not P3_SUB_414_U32 ; P3_SUB_414_U97
g21953 not P3_SUB_414_U33 ; P3_SUB_414_U98
g21954 not P3_SUB_414_U34 ; P3_SUB_414_U99
g21955 not P3_SUB_414_U35 ; P3_SUB_414_U100
g21956 not P3_SUB_414_U36 ; P3_SUB_414_U101
g21957 not P3_SUB_414_U37 ; P3_SUB_414_U102
g21958 not P3_SUB_414_U38 ; P3_SUB_414_U103
g21959 or P3_EBX_REG_0__SCAN_IN P3_EBX_REG_1__SCAN_IN ; P3_SUB_414_U104
g21960 nand P3_SUB_414_U104 P3_EBX_REG_2__SCAN_IN ; P3_SUB_414_U105
g21961 nand P3_SUB_414_U37 P3_EBX_REG_29__SCAN_IN ; P3_SUB_414_U106
g21962 nand P3_SUB_414_U101 P3_SUB_414_U63 ; P3_SUB_414_U107
g21963 nand P3_SUB_414_U107 P3_EBX_REG_28__SCAN_IN ; P3_SUB_414_U108
g21964 nand P3_SUB_414_U100 P3_SUB_414_U65 ; P3_SUB_414_U109
g21965 nand P3_SUB_414_U109 P3_EBX_REG_26__SCAN_IN ; P3_SUB_414_U110
g21966 nand P3_SUB_414_U99 P3_SUB_414_U67 ; P3_SUB_414_U111
g21967 nand P3_SUB_414_U111 P3_EBX_REG_24__SCAN_IN ; P3_SUB_414_U112
g21968 nand P3_SUB_414_U98 P3_SUB_414_U69 ; P3_SUB_414_U113
g21969 nand P3_SUB_414_U113 P3_EBX_REG_22__SCAN_IN ; P3_SUB_414_U114
g21970 nand P3_SUB_414_U97 P3_SUB_414_U73 ; P3_SUB_414_U115
g21971 nand P3_SUB_414_U115 P3_EBX_REG_20__SCAN_IN ; P3_SUB_414_U116
g21972 nand P3_SUB_414_U96 P3_SUB_414_U75 ; P3_SUB_414_U117
g21973 nand P3_SUB_414_U117 P3_EBX_REG_18__SCAN_IN ; P3_SUB_414_U118
g21974 nand P3_SUB_414_U95 P3_SUB_414_U77 ; P3_SUB_414_U119
g21975 nand P3_SUB_414_U119 P3_EBX_REG_16__SCAN_IN ; P3_SUB_414_U120
g21976 nand P3_SUB_414_U94 P3_SUB_414_U79 ; P3_SUB_414_U121
g21977 nand P3_SUB_414_U121 P3_EBX_REG_14__SCAN_IN ; P3_SUB_414_U122
g21978 nand P3_SUB_414_U93 P3_SUB_414_U81 ; P3_SUB_414_U123
g21979 nand P3_SUB_414_U123 P3_EBX_REG_12__SCAN_IN ; P3_SUB_414_U124
g21980 nand P3_SUB_414_U86 P3_SUB_414_U52 ; P3_SUB_414_U125
g21981 nand P3_SUB_414_U125 P3_EBX_REG_10__SCAN_IN ; P3_SUB_414_U126
g21982 nand P3_SUB_414_U103 P3_SUB_414_U61 ; P3_SUB_414_U127
g21983 nand P3_SUB_414_U24 P3_EBX_REG_9__SCAN_IN ; P3_SUB_414_U128
g21984 nand P3_SUB_414_U86 P3_SUB_414_U52 ; P3_SUB_414_U129
g21985 nand P3_SUB_414_U23 P3_EBX_REG_7__SCAN_IN ; P3_SUB_414_U130
g21986 nand P3_SUB_414_U85 P3_SUB_414_U54 ; P3_SUB_414_U131
g21987 nand P3_SUB_414_U22 P3_EBX_REG_5__SCAN_IN ; P3_SUB_414_U132
g21988 nand P3_SUB_414_U84 P3_SUB_414_U56 ; P3_SUB_414_U133
g21989 nand P3_SUB_414_U21 P3_EBX_REG_3__SCAN_IN ; P3_SUB_414_U134
g21990 nand P3_SUB_414_U83 P3_SUB_414_U58 ; P3_SUB_414_U135
g21991 nand P3_SUB_414_U127 P3_SUB_414_U60 ; P3_SUB_414_U136
g21992 nand P3_SUB_414_U103 P3_SUB_414_U61 P3_EBX_REG_31__SCAN_IN ; P3_SUB_414_U137
g21993 nand P3_SUB_414_U38 P3_EBX_REG_30__SCAN_IN ; P3_SUB_414_U138
g21994 nand P3_SUB_414_U103 P3_SUB_414_U61 ; P3_SUB_414_U139
g21995 nand P3_SUB_414_U36 P3_EBX_REG_27__SCAN_IN ; P3_SUB_414_U140
g21996 nand P3_SUB_414_U101 P3_SUB_414_U63 ; P3_SUB_414_U141
g21997 nand P3_SUB_414_U35 P3_EBX_REG_25__SCAN_IN ; P3_SUB_414_U142
g21998 nand P3_SUB_414_U100 P3_SUB_414_U65 ; P3_SUB_414_U143
g21999 nand P3_SUB_414_U34 P3_EBX_REG_23__SCAN_IN ; P3_SUB_414_U144
g22000 nand P3_SUB_414_U99 P3_SUB_414_U67 ; P3_SUB_414_U145
g22001 nand P3_SUB_414_U33 P3_EBX_REG_21__SCAN_IN ; P3_SUB_414_U146
g22002 nand P3_SUB_414_U98 P3_SUB_414_U69 ; P3_SUB_414_U147
g22003 nand P3_SUB_414_U72 P3_EBX_REG_1__SCAN_IN ; P3_SUB_414_U148
g22004 nand P3_SUB_414_U71 P3_EBX_REG_0__SCAN_IN ; P3_SUB_414_U149
g22005 nand P3_SUB_414_U32 P3_EBX_REG_19__SCAN_IN ; P3_SUB_414_U150
g22006 nand P3_SUB_414_U97 P3_SUB_414_U73 ; P3_SUB_414_U151
g22007 nand P3_SUB_414_U31 P3_EBX_REG_17__SCAN_IN ; P3_SUB_414_U152
g22008 nand P3_SUB_414_U96 P3_SUB_414_U75 ; P3_SUB_414_U153
g22009 nand P3_SUB_414_U30 P3_EBX_REG_15__SCAN_IN ; P3_SUB_414_U154
g22010 nand P3_SUB_414_U95 P3_SUB_414_U77 ; P3_SUB_414_U155
g22011 nand P3_SUB_414_U29 P3_EBX_REG_13__SCAN_IN ; P3_SUB_414_U156
g22012 nand P3_SUB_414_U94 P3_SUB_414_U79 ; P3_SUB_414_U157
g22013 nand P3_SUB_414_U28 P3_EBX_REG_11__SCAN_IN ; P3_SUB_414_U158
g22014 nand P3_SUB_414_U93 P3_SUB_414_U81 ; P3_SUB_414_U159
g22015 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_441_U4
g22016 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_441_U5
g22017 nand P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_441_U6
g22018 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_441_U7
g22019 nand P3_ADD_441_U94 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_441_U8
g22020 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_441_U9
g22021 nand P3_ADD_441_U95 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_441_U10
g22022 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_441_U11
g22023 nand P3_ADD_441_U96 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_441_U12
g22024 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_441_U13
g22025 nand P3_ADD_441_U97 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_441_U14
g22026 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_441_U15
g22027 nand P3_ADD_441_U98 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_441_U16
g22028 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_441_U17
g22029 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_441_U18
g22030 nand P3_ADD_441_U99 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_441_U19
g22031 nand P3_ADD_441_U100 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_441_U20
g22032 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_441_U21
g22033 nand P3_ADD_441_U101 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_441_U22
g22034 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_441_U23
g22035 nand P3_ADD_441_U102 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_441_U24
g22036 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_441_U25
g22037 nand P3_ADD_441_U103 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_441_U26
g22038 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_441_U27
g22039 nand P3_ADD_441_U104 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_441_U28
g22040 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_441_U29
g22041 nand P3_ADD_441_U105 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_441_U30
g22042 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_441_U31
g22043 nand P3_ADD_441_U106 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_441_U32
g22044 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_441_U33
g22045 nand P3_ADD_441_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_441_U34
g22046 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_441_U35
g22047 nand P3_ADD_441_U108 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_441_U36
g22048 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_441_U37
g22049 nand P3_ADD_441_U109 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_441_U38
g22050 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_441_U39
g22051 nand P3_ADD_441_U110 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_441_U40
g22052 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_441_U41
g22053 nand P3_ADD_441_U111 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_441_U42
g22054 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_441_U43
g22055 nand P3_ADD_441_U112 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_441_U44
g22056 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_441_U45
g22057 nand P3_ADD_441_U113 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_441_U46
g22058 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_441_U47
g22059 nand P3_ADD_441_U114 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_441_U48
g22060 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_441_U49
g22061 nand P3_ADD_441_U115 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_441_U50
g22062 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_441_U51
g22063 nand P3_ADD_441_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_441_U52
g22064 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_441_U53
g22065 nand P3_ADD_441_U117 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_441_U54
g22066 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_441_U55
g22067 nand P3_ADD_441_U118 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_441_U56
g22068 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_441_U57
g22069 nand P3_ADD_441_U119 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_441_U58
g22070 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_441_U59
g22071 nand P3_ADD_441_U120 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_441_U60
g22072 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_441_U61
g22073 nand P3_ADD_441_U124 P3_ADD_441_U123 ; P3_ADD_441_U62
g22074 nand P3_ADD_441_U126 P3_ADD_441_U125 ; P3_ADD_441_U63
g22075 nand P3_ADD_441_U128 P3_ADD_441_U127 ; P3_ADD_441_U64
g22076 nand P3_ADD_441_U130 P3_ADD_441_U129 ; P3_ADD_441_U65
g22077 nand P3_ADD_441_U132 P3_ADD_441_U131 ; P3_ADD_441_U66
g22078 nand P3_ADD_441_U134 P3_ADD_441_U133 ; P3_ADD_441_U67
g22079 nand P3_ADD_441_U136 P3_ADD_441_U135 ; P3_ADD_441_U68
g22080 nand P3_ADD_441_U138 P3_ADD_441_U137 ; P3_ADD_441_U69
g22081 nand P3_ADD_441_U140 P3_ADD_441_U139 ; P3_ADD_441_U70
g22082 nand P3_ADD_441_U142 P3_ADD_441_U141 ; P3_ADD_441_U71
g22083 nand P3_ADD_441_U144 P3_ADD_441_U143 ; P3_ADD_441_U72
g22084 nand P3_ADD_441_U146 P3_ADD_441_U145 ; P3_ADD_441_U73
g22085 nand P3_ADD_441_U148 P3_ADD_441_U147 ; P3_ADD_441_U74
g22086 nand P3_ADD_441_U150 P3_ADD_441_U149 ; P3_ADD_441_U75
g22087 nand P3_ADD_441_U152 P3_ADD_441_U151 ; P3_ADD_441_U76
g22088 nand P3_ADD_441_U154 P3_ADD_441_U153 ; P3_ADD_441_U77
g22089 nand P3_ADD_441_U156 P3_ADD_441_U155 ; P3_ADD_441_U78
g22090 nand P3_ADD_441_U158 P3_ADD_441_U157 ; P3_ADD_441_U79
g22091 nand P3_ADD_441_U160 P3_ADD_441_U159 ; P3_ADD_441_U80
g22092 nand P3_ADD_441_U162 P3_ADD_441_U161 ; P3_ADD_441_U81
g22093 nand P3_ADD_441_U164 P3_ADD_441_U163 ; P3_ADD_441_U82
g22094 nand P3_ADD_441_U166 P3_ADD_441_U165 ; P3_ADD_441_U83
g22095 nand P3_ADD_441_U168 P3_ADD_441_U167 ; P3_ADD_441_U84
g22096 nand P3_ADD_441_U170 P3_ADD_441_U169 ; P3_ADD_441_U85
g22097 nand P3_ADD_441_U172 P3_ADD_441_U171 ; P3_ADD_441_U86
g22098 nand P3_ADD_441_U174 P3_ADD_441_U173 ; P3_ADD_441_U87
g22099 nand P3_ADD_441_U176 P3_ADD_441_U175 ; P3_ADD_441_U88
g22100 nand P3_ADD_441_U178 P3_ADD_441_U177 ; P3_ADD_441_U89
g22101 nand P3_ADD_441_U180 P3_ADD_441_U179 ; P3_ADD_441_U90
g22102 nand P3_ADD_441_U182 P3_ADD_441_U181 ; P3_ADD_441_U91
g22103 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_441_U92
g22104 nand P3_ADD_441_U121 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_441_U93
g22105 not P3_ADD_441_U6 ; P3_ADD_441_U94
g22106 not P3_ADD_441_U8 ; P3_ADD_441_U95
g22107 not P3_ADD_441_U10 ; P3_ADD_441_U96
g22108 not P3_ADD_441_U12 ; P3_ADD_441_U97
g22109 not P3_ADD_441_U14 ; P3_ADD_441_U98
g22110 not P3_ADD_441_U16 ; P3_ADD_441_U99
g22111 not P3_ADD_441_U19 ; P3_ADD_441_U100
g22112 not P3_ADD_441_U20 ; P3_ADD_441_U101
g22113 not P3_ADD_441_U22 ; P3_ADD_441_U102
g22114 not P3_ADD_441_U24 ; P3_ADD_441_U103
g22115 not P3_ADD_441_U26 ; P3_ADD_441_U104
g22116 not P3_ADD_441_U28 ; P3_ADD_441_U105
g22117 not P3_ADD_441_U30 ; P3_ADD_441_U106
g22118 not P3_ADD_441_U32 ; P3_ADD_441_U107
g22119 not P3_ADD_441_U34 ; P3_ADD_441_U108
g22120 not P3_ADD_441_U36 ; P3_ADD_441_U109
g22121 not P3_ADD_441_U38 ; P3_ADD_441_U110
g22122 not P3_ADD_441_U40 ; P3_ADD_441_U111
g22123 not P3_ADD_441_U42 ; P3_ADD_441_U112
g22124 not P3_ADD_441_U44 ; P3_ADD_441_U113
g22125 not P3_ADD_441_U46 ; P3_ADD_441_U114
g22126 not P3_ADD_441_U48 ; P3_ADD_441_U115
g22127 not P3_ADD_441_U50 ; P3_ADD_441_U116
g22128 not P3_ADD_441_U52 ; P3_ADD_441_U117
g22129 not P3_ADD_441_U54 ; P3_ADD_441_U118
g22130 not P3_ADD_441_U56 ; P3_ADD_441_U119
g22131 not P3_ADD_441_U58 ; P3_ADD_441_U120
g22132 not P3_ADD_441_U60 ; P3_ADD_441_U121
g22133 not P3_ADD_441_U93 ; P3_ADD_441_U122
g22134 nand P3_ADD_441_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_441_U123
g22135 nand P3_ADD_441_U100 P3_ADD_441_U18 ; P3_ADD_441_U124
g22136 nand P3_ADD_441_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_441_U125
g22137 nand P3_ADD_441_U99 P3_ADD_441_U17 ; P3_ADD_441_U126
g22138 nand P3_ADD_441_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_441_U127
g22139 nand P3_ADD_441_U98 P3_ADD_441_U15 ; P3_ADD_441_U128
g22140 nand P3_ADD_441_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_441_U129
g22141 nand P3_ADD_441_U97 P3_ADD_441_U13 ; P3_ADD_441_U130
g22142 nand P3_ADD_441_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_441_U131
g22143 nand P3_ADD_441_U96 P3_ADD_441_U11 ; P3_ADD_441_U132
g22144 nand P3_ADD_441_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_441_U133
g22145 nand P3_ADD_441_U95 P3_ADD_441_U9 ; P3_ADD_441_U134
g22146 nand P3_ADD_441_U6 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_441_U135
g22147 nand P3_ADD_441_U94 P3_ADD_441_U7 ; P3_ADD_441_U136
g22148 nand P3_ADD_441_U93 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_441_U137
g22149 nand P3_ADD_441_U122 P3_ADD_441_U92 ; P3_ADD_441_U138
g22150 nand P3_ADD_441_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_441_U139
g22151 nand P3_ADD_441_U121 P3_ADD_441_U61 ; P3_ADD_441_U140
g22152 nand P3_ADD_441_U4 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_441_U141
g22153 nand P3_ADD_441_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_441_U142
g22154 nand P3_ADD_441_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_441_U143
g22155 nand P3_ADD_441_U120 P3_ADD_441_U59 ; P3_ADD_441_U144
g22156 nand P3_ADD_441_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_441_U145
g22157 nand P3_ADD_441_U119 P3_ADD_441_U57 ; P3_ADD_441_U146
g22158 nand P3_ADD_441_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_441_U147
g22159 nand P3_ADD_441_U118 P3_ADD_441_U55 ; P3_ADD_441_U148
g22160 nand P3_ADD_441_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_441_U149
g22161 nand P3_ADD_441_U117 P3_ADD_441_U53 ; P3_ADD_441_U150
g22162 nand P3_ADD_441_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_441_U151
g22163 nand P3_ADD_441_U116 P3_ADD_441_U51 ; P3_ADD_441_U152
g22164 nand P3_ADD_441_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_441_U153
g22165 nand P3_ADD_441_U115 P3_ADD_441_U49 ; P3_ADD_441_U154
g22166 nand P3_ADD_441_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_441_U155
g22167 nand P3_ADD_441_U114 P3_ADD_441_U47 ; P3_ADD_441_U156
g22168 nand P3_ADD_441_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_441_U157
g22169 nand P3_ADD_441_U113 P3_ADD_441_U45 ; P3_ADD_441_U158
g22170 nand P3_ADD_441_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_441_U159
g22171 nand P3_ADD_441_U112 P3_ADD_441_U43 ; P3_ADD_441_U160
g22172 nand P3_ADD_441_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_441_U161
g22173 nand P3_ADD_441_U111 P3_ADD_441_U41 ; P3_ADD_441_U162
g22174 nand P3_ADD_441_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_441_U163
g22175 nand P3_ADD_441_U110 P3_ADD_441_U39 ; P3_ADD_441_U164
g22176 nand P3_ADD_441_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_441_U165
g22177 nand P3_ADD_441_U109 P3_ADD_441_U37 ; P3_ADD_441_U166
g22178 nand P3_ADD_441_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_441_U167
g22179 nand P3_ADD_441_U108 P3_ADD_441_U35 ; P3_ADD_441_U168
g22180 nand P3_ADD_441_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_441_U169
g22181 nand P3_ADD_441_U107 P3_ADD_441_U33 ; P3_ADD_441_U170
g22182 nand P3_ADD_441_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_441_U171
g22183 nand P3_ADD_441_U106 P3_ADD_441_U31 ; P3_ADD_441_U172
g22184 nand P3_ADD_441_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_441_U173
g22185 nand P3_ADD_441_U105 P3_ADD_441_U29 ; P3_ADD_441_U174
g22186 nand P3_ADD_441_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_441_U175
g22187 nand P3_ADD_441_U104 P3_ADD_441_U27 ; P3_ADD_441_U176
g22188 nand P3_ADD_441_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_441_U177
g22189 nand P3_ADD_441_U103 P3_ADD_441_U25 ; P3_ADD_441_U178
g22190 nand P3_ADD_441_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_441_U179
g22191 nand P3_ADD_441_U102 P3_ADD_441_U23 ; P3_ADD_441_U180
g22192 nand P3_ADD_441_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_441_U181
g22193 nand P3_ADD_441_U101 P3_ADD_441_U21 ; P3_ADD_441_U182
g22194 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_349_U5
g22195 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_349_U6
g22196 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_349_U7
g22197 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_349_U8
g22198 nand P3_ADD_349_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_349_U9
g22199 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_349_U10
g22200 nand P3_ADD_349_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_349_U11
g22201 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_349_U12
g22202 nand P3_ADD_349_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_349_U13
g22203 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_349_U14
g22204 nand P3_ADD_349_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_349_U15
g22205 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_349_U16
g22206 nand P3_ADD_349_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_349_U17
g22207 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_349_U18
g22208 nand P3_ADD_349_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_349_U19
g22209 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_349_U20
g22210 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_349_U21
g22211 nand P3_ADD_349_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_349_U22
g22212 nand P3_ADD_349_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_349_U23
g22213 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_349_U24
g22214 nand P3_ADD_349_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_349_U25
g22215 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_349_U26
g22216 nand P3_ADD_349_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_349_U27
g22217 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_349_U28
g22218 nand P3_ADD_349_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_349_U29
g22219 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_349_U30
g22220 nand P3_ADD_349_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_349_U31
g22221 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_349_U32
g22222 nand P3_ADD_349_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_349_U33
g22223 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_349_U34
g22224 nand P3_ADD_349_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_349_U35
g22225 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_349_U36
g22226 nand P3_ADD_349_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_349_U37
g22227 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_349_U38
g22228 nand P3_ADD_349_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_349_U39
g22229 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_349_U40
g22230 nand P3_ADD_349_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_349_U41
g22231 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_349_U42
g22232 nand P3_ADD_349_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_349_U43
g22233 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_349_U44
g22234 nand P3_ADD_349_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_349_U45
g22235 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_349_U46
g22236 nand P3_ADD_349_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_349_U47
g22237 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_349_U48
g22238 nand P3_ADD_349_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_349_U49
g22239 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_349_U50
g22240 nand P3_ADD_349_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_349_U51
g22241 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_349_U52
g22242 nand P3_ADD_349_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_349_U53
g22243 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_349_U54
g22244 nand P3_ADD_349_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_349_U55
g22245 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_349_U56
g22246 nand P3_ADD_349_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_349_U57
g22247 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_349_U58
g22248 nand P3_ADD_349_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_349_U59
g22249 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_349_U60
g22250 nand P3_ADD_349_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_349_U61
g22251 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_349_U62
g22252 nand P3_ADD_349_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_349_U63
g22253 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_349_U64
g22254 nand P3_ADD_349_U129 P3_ADD_349_U128 ; P3_ADD_349_U65
g22255 nand P3_ADD_349_U131 P3_ADD_349_U130 ; P3_ADD_349_U66
g22256 nand P3_ADD_349_U133 P3_ADD_349_U132 ; P3_ADD_349_U67
g22257 nand P3_ADD_349_U135 P3_ADD_349_U134 ; P3_ADD_349_U68
g22258 nand P3_ADD_349_U137 P3_ADD_349_U136 ; P3_ADD_349_U69
g22259 nand P3_ADD_349_U139 P3_ADD_349_U138 ; P3_ADD_349_U70
g22260 nand P3_ADD_349_U141 P3_ADD_349_U140 ; P3_ADD_349_U71
g22261 nand P3_ADD_349_U143 P3_ADD_349_U142 ; P3_ADD_349_U72
g22262 nand P3_ADD_349_U145 P3_ADD_349_U144 ; P3_ADD_349_U73
g22263 nand P3_ADD_349_U147 P3_ADD_349_U146 ; P3_ADD_349_U74
g22264 nand P3_ADD_349_U149 P3_ADD_349_U148 ; P3_ADD_349_U75
g22265 nand P3_ADD_349_U151 P3_ADD_349_U150 ; P3_ADD_349_U76
g22266 nand P3_ADD_349_U153 P3_ADD_349_U152 ; P3_ADD_349_U77
g22267 nand P3_ADD_349_U155 P3_ADD_349_U154 ; P3_ADD_349_U78
g22268 nand P3_ADD_349_U157 P3_ADD_349_U156 ; P3_ADD_349_U79
g22269 nand P3_ADD_349_U159 P3_ADD_349_U158 ; P3_ADD_349_U80
g22270 nand P3_ADD_349_U161 P3_ADD_349_U160 ; P3_ADD_349_U81
g22271 nand P3_ADD_349_U163 P3_ADD_349_U162 ; P3_ADD_349_U82
g22272 nand P3_ADD_349_U165 P3_ADD_349_U164 ; P3_ADD_349_U83
g22273 nand P3_ADD_349_U167 P3_ADD_349_U166 ; P3_ADD_349_U84
g22274 nand P3_ADD_349_U169 P3_ADD_349_U168 ; P3_ADD_349_U85
g22275 nand P3_ADD_349_U171 P3_ADD_349_U170 ; P3_ADD_349_U86
g22276 nand P3_ADD_349_U173 P3_ADD_349_U172 ; P3_ADD_349_U87
g22277 nand P3_ADD_349_U175 P3_ADD_349_U174 ; P3_ADD_349_U88
g22278 nand P3_ADD_349_U177 P3_ADD_349_U176 ; P3_ADD_349_U89
g22279 nand P3_ADD_349_U179 P3_ADD_349_U178 ; P3_ADD_349_U90
g22280 nand P3_ADD_349_U181 P3_ADD_349_U180 ; P3_ADD_349_U91
g22281 nand P3_ADD_349_U183 P3_ADD_349_U182 ; P3_ADD_349_U92
g22282 nand P3_ADD_349_U185 P3_ADD_349_U184 ; P3_ADD_349_U93
g22283 nand P3_ADD_349_U187 P3_ADD_349_U186 ; P3_ADD_349_U94
g22284 nand P3_ADD_349_U189 P3_ADD_349_U188 ; P3_ADD_349_U95
g22285 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_349_U96
g22286 nand P3_ADD_349_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_349_U97
g22287 not P3_ADD_349_U7 ; P3_ADD_349_U98
g22288 not P3_ADD_349_U9 ; P3_ADD_349_U99
g22289 not P3_ADD_349_U11 ; P3_ADD_349_U100
g22290 not P3_ADD_349_U13 ; P3_ADD_349_U101
g22291 not P3_ADD_349_U15 ; P3_ADD_349_U102
g22292 not P3_ADD_349_U17 ; P3_ADD_349_U103
g22293 not P3_ADD_349_U19 ; P3_ADD_349_U104
g22294 not P3_ADD_349_U22 ; P3_ADD_349_U105
g22295 not P3_ADD_349_U23 ; P3_ADD_349_U106
g22296 not P3_ADD_349_U25 ; P3_ADD_349_U107
g22297 not P3_ADD_349_U27 ; P3_ADD_349_U108
g22298 not P3_ADD_349_U29 ; P3_ADD_349_U109
g22299 not P3_ADD_349_U31 ; P3_ADD_349_U110
g22300 not P3_ADD_349_U33 ; P3_ADD_349_U111
g22301 not P3_ADD_349_U35 ; P3_ADD_349_U112
g22302 not P3_ADD_349_U37 ; P3_ADD_349_U113
g22303 not P3_ADD_349_U39 ; P3_ADD_349_U114
g22304 not P3_ADD_349_U41 ; P3_ADD_349_U115
g22305 not P3_ADD_349_U43 ; P3_ADD_349_U116
g22306 not P3_ADD_349_U45 ; P3_ADD_349_U117
g22307 not P3_ADD_349_U47 ; P3_ADD_349_U118
g22308 not P3_ADD_349_U49 ; P3_ADD_349_U119
g22309 not P3_ADD_349_U51 ; P3_ADD_349_U120
g22310 not P3_ADD_349_U53 ; P3_ADD_349_U121
g22311 not P3_ADD_349_U55 ; P3_ADD_349_U122
g22312 not P3_ADD_349_U57 ; P3_ADD_349_U123
g22313 not P3_ADD_349_U59 ; P3_ADD_349_U124
g22314 not P3_ADD_349_U61 ; P3_ADD_349_U125
g22315 not P3_ADD_349_U63 ; P3_ADD_349_U126
g22316 not P3_ADD_349_U97 ; P3_ADD_349_U127
g22317 nand P3_ADD_349_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_349_U128
g22318 nand P3_ADD_349_U105 P3_ADD_349_U21 ; P3_ADD_349_U129
g22319 nand P3_ADD_349_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_349_U130
g22320 nand P3_ADD_349_U104 P3_ADD_349_U20 ; P3_ADD_349_U131
g22321 nand P3_ADD_349_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_349_U132
g22322 nand P3_ADD_349_U103 P3_ADD_349_U18 ; P3_ADD_349_U133
g22323 nand P3_ADD_349_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_349_U134
g22324 nand P3_ADD_349_U102 P3_ADD_349_U16 ; P3_ADD_349_U135
g22325 nand P3_ADD_349_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_349_U136
g22326 nand P3_ADD_349_U101 P3_ADD_349_U14 ; P3_ADD_349_U137
g22327 nand P3_ADD_349_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_349_U138
g22328 nand P3_ADD_349_U100 P3_ADD_349_U12 ; P3_ADD_349_U139
g22329 nand P3_ADD_349_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_349_U140
g22330 nand P3_ADD_349_U99 P3_ADD_349_U10 ; P3_ADD_349_U141
g22331 nand P3_ADD_349_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_349_U142
g22332 nand P3_ADD_349_U127 P3_ADD_349_U96 ; P3_ADD_349_U143
g22333 nand P3_ADD_349_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_349_U144
g22334 nand P3_ADD_349_U126 P3_ADD_349_U64 ; P3_ADD_349_U145
g22335 nand P3_ADD_349_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_349_U146
g22336 nand P3_ADD_349_U98 P3_ADD_349_U8 ; P3_ADD_349_U147
g22337 nand P3_ADD_349_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_349_U148
g22338 nand P3_ADD_349_U125 P3_ADD_349_U62 ; P3_ADD_349_U149
g22339 nand P3_ADD_349_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_349_U150
g22340 nand P3_ADD_349_U124 P3_ADD_349_U60 ; P3_ADD_349_U151
g22341 nand P3_ADD_349_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_349_U152
g22342 nand P3_ADD_349_U123 P3_ADD_349_U58 ; P3_ADD_349_U153
g22343 nand P3_ADD_349_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_349_U154
g22344 nand P3_ADD_349_U122 P3_ADD_349_U56 ; P3_ADD_349_U155
g22345 nand P3_ADD_349_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_349_U156
g22346 nand P3_ADD_349_U121 P3_ADD_349_U54 ; P3_ADD_349_U157
g22347 nand P3_ADD_349_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_349_U158
g22348 nand P3_ADD_349_U120 P3_ADD_349_U52 ; P3_ADD_349_U159
g22349 nand P3_ADD_349_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_349_U160
g22350 nand P3_ADD_349_U119 P3_ADD_349_U50 ; P3_ADD_349_U161
g22351 nand P3_ADD_349_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_349_U162
g22352 nand P3_ADD_349_U118 P3_ADD_349_U48 ; P3_ADD_349_U163
g22353 nand P3_ADD_349_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_349_U164
g22354 nand P3_ADD_349_U117 P3_ADD_349_U46 ; P3_ADD_349_U165
g22355 nand P3_ADD_349_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_349_U166
g22356 nand P3_ADD_349_U116 P3_ADD_349_U44 ; P3_ADD_349_U167
g22357 nand P3_ADD_349_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_349_U168
g22358 nand P3_ADD_349_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_349_U169
g22359 nand P3_ADD_349_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_349_U170
g22360 nand P3_ADD_349_U115 P3_ADD_349_U42 ; P3_ADD_349_U171
g22361 nand P3_ADD_349_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_349_U172
g22362 nand P3_ADD_349_U114 P3_ADD_349_U40 ; P3_ADD_349_U173
g22363 nand P3_ADD_349_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_349_U174
g22364 nand P3_ADD_349_U113 P3_ADD_349_U38 ; P3_ADD_349_U175
g22365 nand P3_ADD_349_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_349_U176
g22366 nand P3_ADD_349_U112 P3_ADD_349_U36 ; P3_ADD_349_U177
g22367 nand P3_ADD_349_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_349_U178
g22368 nand P3_ADD_349_U111 P3_ADD_349_U34 ; P3_ADD_349_U179
g22369 nand P3_ADD_349_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_349_U180
g22370 nand P3_ADD_349_U110 P3_ADD_349_U32 ; P3_ADD_349_U181
g22371 nand P3_ADD_349_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_349_U182
g22372 nand P3_ADD_349_U109 P3_ADD_349_U30 ; P3_ADD_349_U183
g22373 nand P3_ADD_349_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_349_U184
g22374 nand P3_ADD_349_U108 P3_ADD_349_U28 ; P3_ADD_349_U185
g22375 nand P3_ADD_349_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_349_U186
g22376 nand P3_ADD_349_U107 P3_ADD_349_U26 ; P3_ADD_349_U187
g22377 nand P3_ADD_349_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_349_U188
g22378 nand P3_ADD_349_U106 P3_ADD_349_U24 ; P3_ADD_349_U189
g22379 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_405_U4
g22380 nand P3_ADD_405_U92 P3_ADD_405_U126 ; P3_ADD_405_U5
g22381 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_405_U6
g22382 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_405_U7
g22383 nand P3_ADD_405_U92 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_405_U8
g22384 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_405_U9
g22385 nand P3_ADD_405_U98 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_405_U10
g22386 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_405_U11
g22387 nand P3_ADD_405_U99 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_405_U12
g22388 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_405_U13
g22389 nand P3_ADD_405_U100 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_405_U14
g22390 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_405_U15
g22391 nand P3_ADD_405_U101 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_405_U16
g22392 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_405_U17
g22393 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_405_U18
g22394 nand P3_ADD_405_U102 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_405_U19
g22395 nand P3_ADD_405_U103 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_405_U20
g22396 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_405_U21
g22397 nand P3_ADD_405_U104 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_405_U22
g22398 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_405_U23
g22399 nand P3_ADD_405_U105 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_405_U24
g22400 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_405_U25
g22401 nand P3_ADD_405_U106 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_405_U26
g22402 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_405_U27
g22403 nand P3_ADD_405_U107 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_405_U28
g22404 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_405_U29
g22405 nand P3_ADD_405_U108 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_405_U30
g22406 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_405_U31
g22407 nand P3_ADD_405_U109 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_405_U32
g22408 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_405_U33
g22409 nand P3_ADD_405_U110 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_405_U34
g22410 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_405_U35
g22411 nand P3_ADD_405_U111 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_405_U36
g22412 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_405_U37
g22413 nand P3_ADD_405_U112 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_405_U38
g22414 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_405_U39
g22415 nand P3_ADD_405_U113 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_405_U40
g22416 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_405_U41
g22417 nand P3_ADD_405_U114 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_405_U42
g22418 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_405_U43
g22419 nand P3_ADD_405_U115 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_405_U44
g22420 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_405_U45
g22421 nand P3_ADD_405_U116 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_405_U46
g22422 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_405_U47
g22423 nand P3_ADD_405_U117 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_405_U48
g22424 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_405_U49
g22425 nand P3_ADD_405_U118 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_405_U50
g22426 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_405_U51
g22427 nand P3_ADD_405_U119 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_405_U52
g22428 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_405_U53
g22429 nand P3_ADD_405_U120 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_405_U54
g22430 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_405_U55
g22431 nand P3_ADD_405_U121 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_405_U56
g22432 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_405_U57
g22433 nand P3_ADD_405_U122 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_405_U58
g22434 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_405_U59
g22435 nand P3_ADD_405_U123 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_405_U60
g22436 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_405_U61
g22437 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_405_U62
g22438 nand P3_ADD_405_U128 P3_ADD_405_U127 ; P3_ADD_405_U63
g22439 nand P3_ADD_405_U130 P3_ADD_405_U129 ; P3_ADD_405_U64
g22440 nand P3_ADD_405_U132 P3_ADD_405_U131 ; P3_ADD_405_U65
g22441 nand P3_ADD_405_U134 P3_ADD_405_U133 ; P3_ADD_405_U66
g22442 nand P3_ADD_405_U136 P3_ADD_405_U135 ; P3_ADD_405_U67
g22443 nand P3_ADD_405_U138 P3_ADD_405_U137 ; P3_ADD_405_U68
g22444 nand P3_ADD_405_U142 P3_ADD_405_U141 ; P3_ADD_405_U69
g22445 nand P3_ADD_405_U144 P3_ADD_405_U143 ; P3_ADD_405_U70
g22446 nand P3_ADD_405_U146 P3_ADD_405_U145 ; P3_ADD_405_U71
g22447 nand P3_ADD_405_U148 P3_ADD_405_U147 ; P3_ADD_405_U72
g22448 nand P3_ADD_405_U150 P3_ADD_405_U149 ; P3_ADD_405_U73
g22449 nand P3_ADD_405_U152 P3_ADD_405_U151 ; P3_ADD_405_U74
g22450 nand P3_ADD_405_U154 P3_ADD_405_U153 ; P3_ADD_405_U75
g22451 nand P3_ADD_405_U156 P3_ADD_405_U155 ; P3_ADD_405_U76
g22452 nand P3_ADD_405_U158 P3_ADD_405_U157 ; P3_ADD_405_U77
g22453 nand P3_ADD_405_U160 P3_ADD_405_U159 ; P3_ADD_405_U78
g22454 nand P3_ADD_405_U162 P3_ADD_405_U161 ; P3_ADD_405_U79
g22455 nand P3_ADD_405_U164 P3_ADD_405_U163 ; P3_ADD_405_U80
g22456 nand P3_ADD_405_U166 P3_ADD_405_U165 ; P3_ADD_405_U81
g22457 nand P3_ADD_405_U168 P3_ADD_405_U167 ; P3_ADD_405_U82
g22458 nand P3_ADD_405_U170 P3_ADD_405_U169 ; P3_ADD_405_U83
g22459 nand P3_ADD_405_U172 P3_ADD_405_U171 ; P3_ADD_405_U84
g22460 nand P3_ADD_405_U174 P3_ADD_405_U173 ; P3_ADD_405_U85
g22461 nand P3_ADD_405_U176 P3_ADD_405_U175 ; P3_ADD_405_U86
g22462 nand P3_ADD_405_U178 P3_ADD_405_U177 ; P3_ADD_405_U87
g22463 nand P3_ADD_405_U180 P3_ADD_405_U179 ; P3_ADD_405_U88
g22464 nand P3_ADD_405_U182 P3_ADD_405_U181 ; P3_ADD_405_U89
g22465 nand P3_ADD_405_U184 P3_ADD_405_U183 ; P3_ADD_405_U90
g22466 nand P3_ADD_405_U186 P3_ADD_405_U185 ; P3_ADD_405_U91
g22467 nand P3_ADD_405_U62 P3_ADD_405_U96 ; P3_ADD_405_U92
g22468 and P3_ADD_405_U140 P3_ADD_405_U139 ; P3_ADD_405_U93
g22469 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_405_U94
g22470 nand P3_ADD_405_U124 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_405_U95
g22471 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_405_U96
g22472 not P3_ADD_405_U92 ; P3_ADD_405_U97
g22473 not P3_ADD_405_U8 ; P3_ADD_405_U98
g22474 not P3_ADD_405_U10 ; P3_ADD_405_U99
g22475 not P3_ADD_405_U12 ; P3_ADD_405_U100
g22476 not P3_ADD_405_U14 ; P3_ADD_405_U101
g22477 not P3_ADD_405_U16 ; P3_ADD_405_U102
g22478 not P3_ADD_405_U19 ; P3_ADD_405_U103
g22479 not P3_ADD_405_U20 ; P3_ADD_405_U104
g22480 not P3_ADD_405_U22 ; P3_ADD_405_U105
g22481 not P3_ADD_405_U24 ; P3_ADD_405_U106
g22482 not P3_ADD_405_U26 ; P3_ADD_405_U107
g22483 not P3_ADD_405_U28 ; P3_ADD_405_U108
g22484 not P3_ADD_405_U30 ; P3_ADD_405_U109
g22485 not P3_ADD_405_U32 ; P3_ADD_405_U110
g22486 not P3_ADD_405_U34 ; P3_ADD_405_U111
g22487 not P3_ADD_405_U36 ; P3_ADD_405_U112
g22488 not P3_ADD_405_U38 ; P3_ADD_405_U113
g22489 not P3_ADD_405_U40 ; P3_ADD_405_U114
g22490 not P3_ADD_405_U42 ; P3_ADD_405_U115
g22491 not P3_ADD_405_U44 ; P3_ADD_405_U116
g22492 not P3_ADD_405_U46 ; P3_ADD_405_U117
g22493 not P3_ADD_405_U48 ; P3_ADD_405_U118
g22494 not P3_ADD_405_U50 ; P3_ADD_405_U119
g22495 not P3_ADD_405_U52 ; P3_ADD_405_U120
g22496 not P3_ADD_405_U54 ; P3_ADD_405_U121
g22497 not P3_ADD_405_U56 ; P3_ADD_405_U122
g22498 not P3_ADD_405_U58 ; P3_ADD_405_U123
g22499 not P3_ADD_405_U60 ; P3_ADD_405_U124
g22500 not P3_ADD_405_U95 ; P3_ADD_405_U125
g22501 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_405_U126
g22502 nand P3_ADD_405_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_405_U127
g22503 nand P3_ADD_405_U103 P3_ADD_405_U18 ; P3_ADD_405_U128
g22504 nand P3_ADD_405_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_405_U129
g22505 nand P3_ADD_405_U102 P3_ADD_405_U17 ; P3_ADD_405_U130
g22506 nand P3_ADD_405_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_405_U131
g22507 nand P3_ADD_405_U101 P3_ADD_405_U15 ; P3_ADD_405_U132
g22508 nand P3_ADD_405_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_405_U133
g22509 nand P3_ADD_405_U100 P3_ADD_405_U13 ; P3_ADD_405_U134
g22510 nand P3_ADD_405_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_405_U135
g22511 nand P3_ADD_405_U99 P3_ADD_405_U11 ; P3_ADD_405_U136
g22512 nand P3_ADD_405_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_405_U137
g22513 nand P3_ADD_405_U98 P3_ADD_405_U9 ; P3_ADD_405_U138
g22514 nand P3_ADD_405_U92 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_405_U139
g22515 nand P3_ADD_405_U97 P3_ADD_405_U7 ; P3_ADD_405_U140
g22516 nand P3_ADD_405_U95 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_405_U141
g22517 nand P3_ADD_405_U125 P3_ADD_405_U94 ; P3_ADD_405_U142
g22518 nand P3_ADD_405_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_405_U143
g22519 nand P3_ADD_405_U124 P3_ADD_405_U61 ; P3_ADD_405_U144
g22520 nand P3_ADD_405_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_405_U145
g22521 nand P3_ADD_405_U123 P3_ADD_405_U59 ; P3_ADD_405_U146
g22522 nand P3_ADD_405_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_405_U147
g22523 nand P3_ADD_405_U122 P3_ADD_405_U57 ; P3_ADD_405_U148
g22524 nand P3_ADD_405_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_405_U149
g22525 nand P3_ADD_405_U121 P3_ADD_405_U55 ; P3_ADD_405_U150
g22526 nand P3_ADD_405_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_405_U151
g22527 nand P3_ADD_405_U120 P3_ADD_405_U53 ; P3_ADD_405_U152
g22528 nand P3_ADD_405_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_405_U153
g22529 nand P3_ADD_405_U119 P3_ADD_405_U51 ; P3_ADD_405_U154
g22530 nand P3_ADD_405_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_405_U155
g22531 nand P3_ADD_405_U118 P3_ADD_405_U49 ; P3_ADD_405_U156
g22532 nand P3_ADD_405_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_405_U157
g22533 nand P3_ADD_405_U117 P3_ADD_405_U47 ; P3_ADD_405_U158
g22534 nand P3_ADD_405_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_405_U159
g22535 nand P3_ADD_405_U116 P3_ADD_405_U45 ; P3_ADD_405_U160
g22536 nand P3_ADD_405_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_405_U161
g22537 nand P3_ADD_405_U115 P3_ADD_405_U43 ; P3_ADD_405_U162
g22538 nand P3_ADD_405_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_405_U163
g22539 nand P3_ADD_405_U114 P3_ADD_405_U41 ; P3_ADD_405_U164
g22540 nand P3_ADD_405_U4 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_405_U165
g22541 nand P3_ADD_405_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_405_U166
g22542 nand P3_ADD_405_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_405_U167
g22543 nand P3_ADD_405_U113 P3_ADD_405_U39 ; P3_ADD_405_U168
g22544 nand P3_ADD_405_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_405_U169
g22545 nand P3_ADD_405_U112 P3_ADD_405_U37 ; P3_ADD_405_U170
g22546 nand P3_ADD_405_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_405_U171
g22547 nand P3_ADD_405_U111 P3_ADD_405_U35 ; P3_ADD_405_U172
g22548 nand P3_ADD_405_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_405_U173
g22549 nand P3_ADD_405_U110 P3_ADD_405_U33 ; P3_ADD_405_U174
g22550 nand P3_ADD_405_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_405_U175
g22551 nand P3_ADD_405_U109 P3_ADD_405_U31 ; P3_ADD_405_U176
g22552 nand P3_ADD_405_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_405_U177
g22553 nand P3_ADD_405_U108 P3_ADD_405_U29 ; P3_ADD_405_U178
g22554 nand P3_ADD_405_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_405_U179
g22555 nand P3_ADD_405_U107 P3_ADD_405_U27 ; P3_ADD_405_U180
g22556 nand P3_ADD_405_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_405_U181
g22557 nand P3_ADD_405_U106 P3_ADD_405_U25 ; P3_ADD_405_U182
g22558 nand P3_ADD_405_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_405_U183
g22559 nand P3_ADD_405_U105 P3_ADD_405_U23 ; P3_ADD_405_U184
g22560 nand P3_ADD_405_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_405_U185
g22561 nand P3_ADD_405_U104 P3_ADD_405_U21 ; P3_ADD_405_U186
g22562 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_553_U5
g22563 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_553_U6
g22564 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_553_U7
g22565 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_553_U8
g22566 nand P3_ADD_553_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_553_U9
g22567 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_553_U10
g22568 nand P3_ADD_553_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_553_U11
g22569 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_553_U12
g22570 nand P3_ADD_553_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_553_U13
g22571 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_553_U14
g22572 nand P3_ADD_553_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_553_U15
g22573 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_553_U16
g22574 nand P3_ADD_553_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_553_U17
g22575 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_553_U18
g22576 nand P3_ADD_553_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_553_U19
g22577 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_553_U20
g22578 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_553_U21
g22579 nand P3_ADD_553_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_553_U22
g22580 nand P3_ADD_553_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_553_U23
g22581 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_553_U24
g22582 nand P3_ADD_553_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_553_U25
g22583 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_553_U26
g22584 nand P3_ADD_553_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_553_U27
g22585 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_553_U28
g22586 nand P3_ADD_553_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_553_U29
g22587 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_553_U30
g22588 nand P3_ADD_553_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_553_U31
g22589 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_553_U32
g22590 nand P3_ADD_553_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_553_U33
g22591 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_553_U34
g22592 nand P3_ADD_553_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_553_U35
g22593 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_553_U36
g22594 nand P3_ADD_553_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_553_U37
g22595 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_553_U38
g22596 nand P3_ADD_553_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_553_U39
g22597 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_553_U40
g22598 nand P3_ADD_553_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_553_U41
g22599 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_553_U42
g22600 nand P3_ADD_553_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_553_U43
g22601 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_553_U44
g22602 nand P3_ADD_553_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_553_U45
g22603 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_553_U46
g22604 nand P3_ADD_553_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_553_U47
g22605 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_553_U48
g22606 nand P3_ADD_553_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_553_U49
g22607 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_553_U50
g22608 nand P3_ADD_553_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_553_U51
g22609 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_553_U52
g22610 nand P3_ADD_553_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_553_U53
g22611 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_553_U54
g22612 nand P3_ADD_553_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_553_U55
g22613 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_553_U56
g22614 nand P3_ADD_553_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_553_U57
g22615 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_553_U58
g22616 nand P3_ADD_553_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_553_U59
g22617 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_553_U60
g22618 nand P3_ADD_553_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_553_U61
g22619 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_553_U62
g22620 nand P3_ADD_553_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_553_U63
g22621 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_553_U64
g22622 nand P3_ADD_553_U129 P3_ADD_553_U128 ; P3_ADD_553_U65
g22623 nand P3_ADD_553_U131 P3_ADD_553_U130 ; P3_ADD_553_U66
g22624 nand P3_ADD_553_U133 P3_ADD_553_U132 ; P3_ADD_553_U67
g22625 nand P3_ADD_553_U135 P3_ADD_553_U134 ; P3_ADD_553_U68
g22626 nand P3_ADD_553_U137 P3_ADD_553_U136 ; P3_ADD_553_U69
g22627 nand P3_ADD_553_U139 P3_ADD_553_U138 ; P3_ADD_553_U70
g22628 nand P3_ADD_553_U141 P3_ADD_553_U140 ; P3_ADD_553_U71
g22629 nand P3_ADD_553_U143 P3_ADD_553_U142 ; P3_ADD_553_U72
g22630 nand P3_ADD_553_U145 P3_ADD_553_U144 ; P3_ADD_553_U73
g22631 nand P3_ADD_553_U147 P3_ADD_553_U146 ; P3_ADD_553_U74
g22632 nand P3_ADD_553_U149 P3_ADD_553_U148 ; P3_ADD_553_U75
g22633 nand P3_ADD_553_U151 P3_ADD_553_U150 ; P3_ADD_553_U76
g22634 nand P3_ADD_553_U153 P3_ADD_553_U152 ; P3_ADD_553_U77
g22635 nand P3_ADD_553_U155 P3_ADD_553_U154 ; P3_ADD_553_U78
g22636 nand P3_ADD_553_U157 P3_ADD_553_U156 ; P3_ADD_553_U79
g22637 nand P3_ADD_553_U159 P3_ADD_553_U158 ; P3_ADD_553_U80
g22638 nand P3_ADD_553_U161 P3_ADD_553_U160 ; P3_ADD_553_U81
g22639 nand P3_ADD_553_U163 P3_ADD_553_U162 ; P3_ADD_553_U82
g22640 nand P3_ADD_553_U165 P3_ADD_553_U164 ; P3_ADD_553_U83
g22641 nand P3_ADD_553_U167 P3_ADD_553_U166 ; P3_ADD_553_U84
g22642 nand P3_ADD_553_U169 P3_ADD_553_U168 ; P3_ADD_553_U85
g22643 nand P3_ADD_553_U171 P3_ADD_553_U170 ; P3_ADD_553_U86
g22644 nand P3_ADD_553_U173 P3_ADD_553_U172 ; P3_ADD_553_U87
g22645 nand P3_ADD_553_U175 P3_ADD_553_U174 ; P3_ADD_553_U88
g22646 nand P3_ADD_553_U177 P3_ADD_553_U176 ; P3_ADD_553_U89
g22647 nand P3_ADD_553_U179 P3_ADD_553_U178 ; P3_ADD_553_U90
g22648 nand P3_ADD_553_U181 P3_ADD_553_U180 ; P3_ADD_553_U91
g22649 nand P3_ADD_553_U183 P3_ADD_553_U182 ; P3_ADD_553_U92
g22650 nand P3_ADD_553_U185 P3_ADD_553_U184 ; P3_ADD_553_U93
g22651 nand P3_ADD_553_U187 P3_ADD_553_U186 ; P3_ADD_553_U94
g22652 nand P3_ADD_553_U189 P3_ADD_553_U188 ; P3_ADD_553_U95
g22653 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_553_U96
g22654 nand P3_ADD_553_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_553_U97
g22655 not P3_ADD_553_U7 ; P3_ADD_553_U98
g22656 not P3_ADD_553_U9 ; P3_ADD_553_U99
g22657 not P3_ADD_553_U11 ; P3_ADD_553_U100
g22658 not P3_ADD_553_U13 ; P3_ADD_553_U101
g22659 not P3_ADD_553_U15 ; P3_ADD_553_U102
g22660 not P3_ADD_553_U17 ; P3_ADD_553_U103
g22661 not P3_ADD_553_U19 ; P3_ADD_553_U104
g22662 not P3_ADD_553_U22 ; P3_ADD_553_U105
g22663 not P3_ADD_553_U23 ; P3_ADD_553_U106
g22664 not P3_ADD_553_U25 ; P3_ADD_553_U107
g22665 not P3_ADD_553_U27 ; P3_ADD_553_U108
g22666 not P3_ADD_553_U29 ; P3_ADD_553_U109
g22667 not P3_ADD_553_U31 ; P3_ADD_553_U110
g22668 not P3_ADD_553_U33 ; P3_ADD_553_U111
g22669 not P3_ADD_553_U35 ; P3_ADD_553_U112
g22670 not P3_ADD_553_U37 ; P3_ADD_553_U113
g22671 not P3_ADD_553_U39 ; P3_ADD_553_U114
g22672 not P3_ADD_553_U41 ; P3_ADD_553_U115
g22673 not P3_ADD_553_U43 ; P3_ADD_553_U116
g22674 not P3_ADD_553_U45 ; P3_ADD_553_U117
g22675 not P3_ADD_553_U47 ; P3_ADD_553_U118
g22676 not P3_ADD_553_U49 ; P3_ADD_553_U119
g22677 not P3_ADD_553_U51 ; P3_ADD_553_U120
g22678 not P3_ADD_553_U53 ; P3_ADD_553_U121
g22679 not P3_ADD_553_U55 ; P3_ADD_553_U122
g22680 not P3_ADD_553_U57 ; P3_ADD_553_U123
g22681 not P3_ADD_553_U59 ; P3_ADD_553_U124
g22682 not P3_ADD_553_U61 ; P3_ADD_553_U125
g22683 not P3_ADD_553_U63 ; P3_ADD_553_U126
g22684 not P3_ADD_553_U97 ; P3_ADD_553_U127
g22685 nand P3_ADD_553_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_553_U128
g22686 nand P3_ADD_553_U105 P3_ADD_553_U21 ; P3_ADD_553_U129
g22687 nand P3_ADD_553_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_553_U130
g22688 nand P3_ADD_553_U104 P3_ADD_553_U20 ; P3_ADD_553_U131
g22689 nand P3_ADD_553_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_553_U132
g22690 nand P3_ADD_553_U103 P3_ADD_553_U18 ; P3_ADD_553_U133
g22691 nand P3_ADD_553_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_553_U134
g22692 nand P3_ADD_553_U102 P3_ADD_553_U16 ; P3_ADD_553_U135
g22693 nand P3_ADD_553_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_553_U136
g22694 nand P3_ADD_553_U101 P3_ADD_553_U14 ; P3_ADD_553_U137
g22695 nand P3_ADD_553_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_553_U138
g22696 nand P3_ADD_553_U100 P3_ADD_553_U12 ; P3_ADD_553_U139
g22697 nand P3_ADD_553_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_553_U140
g22698 nand P3_ADD_553_U99 P3_ADD_553_U10 ; P3_ADD_553_U141
g22699 nand P3_ADD_553_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_553_U142
g22700 nand P3_ADD_553_U127 P3_ADD_553_U96 ; P3_ADD_553_U143
g22701 nand P3_ADD_553_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_553_U144
g22702 nand P3_ADD_553_U126 P3_ADD_553_U64 ; P3_ADD_553_U145
g22703 nand P3_ADD_553_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_553_U146
g22704 nand P3_ADD_553_U98 P3_ADD_553_U8 ; P3_ADD_553_U147
g22705 nand P3_ADD_553_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_553_U148
g22706 nand P3_ADD_553_U125 P3_ADD_553_U62 ; P3_ADD_553_U149
g22707 nand P3_ADD_553_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_553_U150
g22708 nand P3_ADD_553_U124 P3_ADD_553_U60 ; P3_ADD_553_U151
g22709 nand P3_ADD_553_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_553_U152
g22710 nand P3_ADD_553_U123 P3_ADD_553_U58 ; P3_ADD_553_U153
g22711 nand P3_ADD_553_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_553_U154
g22712 nand P3_ADD_553_U122 P3_ADD_553_U56 ; P3_ADD_553_U155
g22713 nand P3_ADD_553_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_553_U156
g22714 nand P3_ADD_553_U121 P3_ADD_553_U54 ; P3_ADD_553_U157
g22715 nand P3_ADD_553_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_553_U158
g22716 nand P3_ADD_553_U120 P3_ADD_553_U52 ; P3_ADD_553_U159
g22717 nand P3_ADD_553_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_553_U160
g22718 nand P3_ADD_553_U119 P3_ADD_553_U50 ; P3_ADD_553_U161
g22719 nand P3_ADD_553_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_553_U162
g22720 nand P3_ADD_553_U118 P3_ADD_553_U48 ; P3_ADD_553_U163
g22721 nand P3_ADD_553_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_553_U164
g22722 nand P3_ADD_553_U117 P3_ADD_553_U46 ; P3_ADD_553_U165
g22723 nand P3_ADD_553_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_553_U166
g22724 nand P3_ADD_553_U116 P3_ADD_553_U44 ; P3_ADD_553_U167
g22725 nand P3_ADD_553_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_553_U168
g22726 nand P3_ADD_553_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_553_U169
g22727 nand P3_ADD_553_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_553_U170
g22728 nand P3_ADD_553_U115 P3_ADD_553_U42 ; P3_ADD_553_U171
g22729 nand P3_ADD_553_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_553_U172
g22730 nand P3_ADD_553_U114 P3_ADD_553_U40 ; P3_ADD_553_U173
g22731 nand P3_ADD_553_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_553_U174
g22732 nand P3_ADD_553_U113 P3_ADD_553_U38 ; P3_ADD_553_U175
g22733 nand P3_ADD_553_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_553_U176
g22734 nand P3_ADD_553_U112 P3_ADD_553_U36 ; P3_ADD_553_U177
g22735 nand P3_ADD_553_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_553_U178
g22736 nand P3_ADD_553_U111 P3_ADD_553_U34 ; P3_ADD_553_U179
g22737 nand P3_ADD_553_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_553_U180
g22738 nand P3_ADD_553_U110 P3_ADD_553_U32 ; P3_ADD_553_U181
g22739 nand P3_ADD_553_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_553_U182
g22740 nand P3_ADD_553_U109 P3_ADD_553_U30 ; P3_ADD_553_U183
g22741 nand P3_ADD_553_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_553_U184
g22742 nand P3_ADD_553_U108 P3_ADD_553_U28 ; P3_ADD_553_U185
g22743 nand P3_ADD_553_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_553_U186
g22744 nand P3_ADD_553_U107 P3_ADD_553_U26 ; P3_ADD_553_U187
g22745 nand P3_ADD_553_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_553_U188
g22746 nand P3_ADD_553_U106 P3_ADD_553_U24 ; P3_ADD_553_U189
g22747 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_558_U5
g22748 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_558_U6
g22749 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_558_U7
g22750 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_558_U8
g22751 nand P3_ADD_558_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_558_U9
g22752 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_558_U10
g22753 nand P3_ADD_558_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_558_U11
g22754 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_558_U12
g22755 nand P3_ADD_558_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_558_U13
g22756 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_558_U14
g22757 nand P3_ADD_558_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_558_U15
g22758 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_558_U16
g22759 nand P3_ADD_558_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_558_U17
g22760 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_558_U18
g22761 nand P3_ADD_558_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_558_U19
g22762 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_558_U20
g22763 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_558_U21
g22764 nand P3_ADD_558_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_558_U22
g22765 nand P3_ADD_558_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_558_U23
g22766 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_558_U24
g22767 nand P3_ADD_558_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_558_U25
g22768 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_558_U26
g22769 nand P3_ADD_558_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_558_U27
g22770 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_558_U28
g22771 nand P3_ADD_558_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_558_U29
g22772 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_558_U30
g22773 nand P3_ADD_558_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_558_U31
g22774 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_558_U32
g22775 nand P3_ADD_558_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_558_U33
g22776 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_558_U34
g22777 nand P3_ADD_558_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_558_U35
g22778 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_558_U36
g22779 nand P3_ADD_558_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_558_U37
g22780 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_558_U38
g22781 nand P3_ADD_558_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_558_U39
g22782 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_558_U40
g22783 nand P3_ADD_558_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_558_U41
g22784 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_558_U42
g22785 nand P3_ADD_558_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_558_U43
g22786 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_558_U44
g22787 nand P3_ADD_558_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_558_U45
g22788 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_558_U46
g22789 nand P3_ADD_558_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_558_U47
g22790 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_558_U48
g22791 nand P3_ADD_558_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_558_U49
g22792 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_558_U50
g22793 nand P3_ADD_558_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_558_U51
g22794 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_558_U52
g22795 nand P3_ADD_558_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_558_U53
g22796 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_558_U54
g22797 nand P3_ADD_558_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_558_U55
g22798 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_558_U56
g22799 nand P3_ADD_558_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_558_U57
g22800 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_558_U58
g22801 nand P3_ADD_558_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_558_U59
g22802 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_558_U60
g22803 nand P3_ADD_558_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_558_U61
g22804 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_558_U62
g22805 nand P3_ADD_558_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_558_U63
g22806 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_558_U64
g22807 nand P3_ADD_558_U129 P3_ADD_558_U128 ; P3_ADD_558_U65
g22808 nand P3_ADD_558_U131 P3_ADD_558_U130 ; P3_ADD_558_U66
g22809 nand P3_ADD_558_U133 P3_ADD_558_U132 ; P3_ADD_558_U67
g22810 nand P3_ADD_558_U135 P3_ADD_558_U134 ; P3_ADD_558_U68
g22811 nand P3_ADD_558_U137 P3_ADD_558_U136 ; P3_ADD_558_U69
g22812 nand P3_ADD_558_U139 P3_ADD_558_U138 ; P3_ADD_558_U70
g22813 nand P3_ADD_558_U141 P3_ADD_558_U140 ; P3_ADD_558_U71
g22814 nand P3_ADD_558_U143 P3_ADD_558_U142 ; P3_ADD_558_U72
g22815 nand P3_ADD_558_U145 P3_ADD_558_U144 ; P3_ADD_558_U73
g22816 nand P3_ADD_558_U147 P3_ADD_558_U146 ; P3_ADD_558_U74
g22817 nand P3_ADD_558_U149 P3_ADD_558_U148 ; P3_ADD_558_U75
g22818 nand P3_ADD_558_U151 P3_ADD_558_U150 ; P3_ADD_558_U76
g22819 nand P3_ADD_558_U153 P3_ADD_558_U152 ; P3_ADD_558_U77
g22820 nand P3_ADD_558_U155 P3_ADD_558_U154 ; P3_ADD_558_U78
g22821 nand P3_ADD_558_U157 P3_ADD_558_U156 ; P3_ADD_558_U79
g22822 nand P3_ADD_558_U159 P3_ADD_558_U158 ; P3_ADD_558_U80
g22823 nand P3_ADD_558_U161 P3_ADD_558_U160 ; P3_ADD_558_U81
g22824 nand P3_ADD_558_U163 P3_ADD_558_U162 ; P3_ADD_558_U82
g22825 nand P3_ADD_558_U165 P3_ADD_558_U164 ; P3_ADD_558_U83
g22826 nand P3_ADD_558_U167 P3_ADD_558_U166 ; P3_ADD_558_U84
g22827 nand P3_ADD_558_U169 P3_ADD_558_U168 ; P3_ADD_558_U85
g22828 nand P3_ADD_558_U171 P3_ADD_558_U170 ; P3_ADD_558_U86
g22829 nand P3_ADD_558_U173 P3_ADD_558_U172 ; P3_ADD_558_U87
g22830 nand P3_ADD_558_U175 P3_ADD_558_U174 ; P3_ADD_558_U88
g22831 nand P3_ADD_558_U177 P3_ADD_558_U176 ; P3_ADD_558_U89
g22832 nand P3_ADD_558_U179 P3_ADD_558_U178 ; P3_ADD_558_U90
g22833 nand P3_ADD_558_U181 P3_ADD_558_U180 ; P3_ADD_558_U91
g22834 nand P3_ADD_558_U183 P3_ADD_558_U182 ; P3_ADD_558_U92
g22835 nand P3_ADD_558_U185 P3_ADD_558_U184 ; P3_ADD_558_U93
g22836 nand P3_ADD_558_U187 P3_ADD_558_U186 ; P3_ADD_558_U94
g22837 nand P3_ADD_558_U189 P3_ADD_558_U188 ; P3_ADD_558_U95
g22838 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_558_U96
g22839 nand P3_ADD_558_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_558_U97
g22840 not P3_ADD_558_U7 ; P3_ADD_558_U98
g22841 not P3_ADD_558_U9 ; P3_ADD_558_U99
g22842 not P3_ADD_558_U11 ; P3_ADD_558_U100
g22843 not P3_ADD_558_U13 ; P3_ADD_558_U101
g22844 not P3_ADD_558_U15 ; P3_ADD_558_U102
g22845 not P3_ADD_558_U17 ; P3_ADD_558_U103
g22846 not P3_ADD_558_U19 ; P3_ADD_558_U104
g22847 not P3_ADD_558_U22 ; P3_ADD_558_U105
g22848 not P3_ADD_558_U23 ; P3_ADD_558_U106
g22849 not P3_ADD_558_U25 ; P3_ADD_558_U107
g22850 not P3_ADD_558_U27 ; P3_ADD_558_U108
g22851 not P3_ADD_558_U29 ; P3_ADD_558_U109
g22852 not P3_ADD_558_U31 ; P3_ADD_558_U110
g22853 not P3_ADD_558_U33 ; P3_ADD_558_U111
g22854 not P3_ADD_558_U35 ; P3_ADD_558_U112
g22855 not P3_ADD_558_U37 ; P3_ADD_558_U113
g22856 not P3_ADD_558_U39 ; P3_ADD_558_U114
g22857 not P3_ADD_558_U41 ; P3_ADD_558_U115
g22858 not P3_ADD_558_U43 ; P3_ADD_558_U116
g22859 not P3_ADD_558_U45 ; P3_ADD_558_U117
g22860 not P3_ADD_558_U47 ; P3_ADD_558_U118
g22861 not P3_ADD_558_U49 ; P3_ADD_558_U119
g22862 not P3_ADD_558_U51 ; P3_ADD_558_U120
g22863 not P3_ADD_558_U53 ; P3_ADD_558_U121
g22864 not P3_ADD_558_U55 ; P3_ADD_558_U122
g22865 not P3_ADD_558_U57 ; P3_ADD_558_U123
g22866 not P3_ADD_558_U59 ; P3_ADD_558_U124
g22867 not P3_ADD_558_U61 ; P3_ADD_558_U125
g22868 not P3_ADD_558_U63 ; P3_ADD_558_U126
g22869 not P3_ADD_558_U97 ; P3_ADD_558_U127
g22870 nand P3_ADD_558_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_558_U128
g22871 nand P3_ADD_558_U105 P3_ADD_558_U21 ; P3_ADD_558_U129
g22872 nand P3_ADD_558_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_558_U130
g22873 nand P3_ADD_558_U104 P3_ADD_558_U20 ; P3_ADD_558_U131
g22874 nand P3_ADD_558_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_558_U132
g22875 nand P3_ADD_558_U103 P3_ADD_558_U18 ; P3_ADD_558_U133
g22876 nand P3_ADD_558_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_558_U134
g22877 nand P3_ADD_558_U102 P3_ADD_558_U16 ; P3_ADD_558_U135
g22878 nand P3_ADD_558_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_558_U136
g22879 nand P3_ADD_558_U101 P3_ADD_558_U14 ; P3_ADD_558_U137
g22880 nand P3_ADD_558_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_558_U138
g22881 nand P3_ADD_558_U100 P3_ADD_558_U12 ; P3_ADD_558_U139
g22882 nand P3_ADD_558_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_558_U140
g22883 nand P3_ADD_558_U99 P3_ADD_558_U10 ; P3_ADD_558_U141
g22884 nand P3_ADD_558_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_558_U142
g22885 nand P3_ADD_558_U127 P3_ADD_558_U96 ; P3_ADD_558_U143
g22886 nand P3_ADD_558_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_558_U144
g22887 nand P3_ADD_558_U126 P3_ADD_558_U64 ; P3_ADD_558_U145
g22888 nand P3_ADD_558_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_558_U146
g22889 nand P3_ADD_558_U98 P3_ADD_558_U8 ; P3_ADD_558_U147
g22890 nand P3_ADD_558_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_558_U148
g22891 nand P3_ADD_558_U125 P3_ADD_558_U62 ; P3_ADD_558_U149
g22892 nand P3_ADD_558_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_558_U150
g22893 nand P3_ADD_558_U124 P3_ADD_558_U60 ; P3_ADD_558_U151
g22894 nand P3_ADD_558_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_558_U152
g22895 nand P3_ADD_558_U123 P3_ADD_558_U58 ; P3_ADD_558_U153
g22896 nand P3_ADD_558_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_558_U154
g22897 nand P3_ADD_558_U122 P3_ADD_558_U56 ; P3_ADD_558_U155
g22898 nand P3_ADD_558_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_558_U156
g22899 nand P3_ADD_558_U121 P3_ADD_558_U54 ; P3_ADD_558_U157
g22900 nand P3_ADD_558_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_558_U158
g22901 nand P3_ADD_558_U120 P3_ADD_558_U52 ; P3_ADD_558_U159
g22902 nand P3_ADD_558_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_558_U160
g22903 nand P3_ADD_558_U119 P3_ADD_558_U50 ; P3_ADD_558_U161
g22904 nand P3_ADD_558_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_558_U162
g22905 nand P3_ADD_558_U118 P3_ADD_558_U48 ; P3_ADD_558_U163
g22906 nand P3_ADD_558_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_558_U164
g22907 nand P3_ADD_558_U117 P3_ADD_558_U46 ; P3_ADD_558_U165
g22908 nand P3_ADD_558_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_558_U166
g22909 nand P3_ADD_558_U116 P3_ADD_558_U44 ; P3_ADD_558_U167
g22910 nand P3_ADD_558_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_558_U168
g22911 nand P3_ADD_558_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_558_U169
g22912 nand P3_ADD_558_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_558_U170
g22913 nand P3_ADD_558_U115 P3_ADD_558_U42 ; P3_ADD_558_U171
g22914 nand P3_ADD_558_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_558_U172
g22915 nand P3_ADD_558_U114 P3_ADD_558_U40 ; P3_ADD_558_U173
g22916 nand P3_ADD_558_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_558_U174
g22917 nand P3_ADD_558_U113 P3_ADD_558_U38 ; P3_ADD_558_U175
g22918 nand P3_ADD_558_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_558_U176
g22919 nand P3_ADD_558_U112 P3_ADD_558_U36 ; P3_ADD_558_U177
g22920 nand P3_ADD_558_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_558_U178
g22921 nand P3_ADD_558_U111 P3_ADD_558_U34 ; P3_ADD_558_U179
g22922 nand P3_ADD_558_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_558_U180
g22923 nand P3_ADD_558_U110 P3_ADD_558_U32 ; P3_ADD_558_U181
g22924 nand P3_ADD_558_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_558_U182
g22925 nand P3_ADD_558_U109 P3_ADD_558_U30 ; P3_ADD_558_U183
g22926 nand P3_ADD_558_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_558_U184
g22927 nand P3_ADD_558_U108 P3_ADD_558_U28 ; P3_ADD_558_U185
g22928 nand P3_ADD_558_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_558_U186
g22929 nand P3_ADD_558_U107 P3_ADD_558_U26 ; P3_ADD_558_U187
g22930 nand P3_ADD_558_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_558_U188
g22931 nand P3_ADD_558_U106 P3_ADD_558_U24 ; P3_ADD_558_U189
g22932 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_385_U5
g22933 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_385_U6
g22934 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_385_U7
g22935 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_385_U8
g22936 nand P3_ADD_385_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_385_U9
g22937 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_385_U10
g22938 nand P3_ADD_385_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_385_U11
g22939 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_385_U12
g22940 nand P3_ADD_385_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_385_U13
g22941 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_385_U14
g22942 nand P3_ADD_385_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_385_U15
g22943 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_385_U16
g22944 nand P3_ADD_385_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_385_U17
g22945 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_385_U18
g22946 nand P3_ADD_385_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_385_U19
g22947 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_385_U20
g22948 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_385_U21
g22949 nand P3_ADD_385_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_385_U22
g22950 nand P3_ADD_385_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_385_U23
g22951 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_385_U24
g22952 nand P3_ADD_385_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_385_U25
g22953 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_385_U26
g22954 nand P3_ADD_385_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_385_U27
g22955 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_385_U28
g22956 nand P3_ADD_385_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_385_U29
g22957 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_385_U30
g22958 nand P3_ADD_385_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_385_U31
g22959 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_385_U32
g22960 nand P3_ADD_385_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_385_U33
g22961 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_385_U34
g22962 nand P3_ADD_385_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_385_U35
g22963 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_385_U36
g22964 nand P3_ADD_385_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_385_U37
g22965 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_385_U38
g22966 nand P3_ADD_385_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_385_U39
g22967 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_385_U40
g22968 nand P3_ADD_385_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_385_U41
g22969 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_385_U42
g22970 nand P3_ADD_385_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_385_U43
g22971 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_385_U44
g22972 nand P3_ADD_385_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_385_U45
g22973 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_385_U46
g22974 nand P3_ADD_385_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_385_U47
g22975 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_385_U48
g22976 nand P3_ADD_385_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_385_U49
g22977 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_385_U50
g22978 nand P3_ADD_385_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_385_U51
g22979 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_385_U52
g22980 nand P3_ADD_385_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_385_U53
g22981 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_385_U54
g22982 nand P3_ADD_385_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_385_U55
g22983 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_385_U56
g22984 nand P3_ADD_385_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_385_U57
g22985 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_385_U58
g22986 nand P3_ADD_385_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_385_U59
g22987 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_385_U60
g22988 nand P3_ADD_385_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_385_U61
g22989 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_385_U62
g22990 nand P3_ADD_385_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_385_U63
g22991 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_385_U64
g22992 nand P3_ADD_385_U129 P3_ADD_385_U128 ; P3_ADD_385_U65
g22993 nand P3_ADD_385_U131 P3_ADD_385_U130 ; P3_ADD_385_U66
g22994 nand P3_ADD_385_U133 P3_ADD_385_U132 ; P3_ADD_385_U67
g22995 nand P3_ADD_385_U135 P3_ADD_385_U134 ; P3_ADD_385_U68
g22996 nand P3_ADD_385_U137 P3_ADD_385_U136 ; P3_ADD_385_U69
g22997 nand P3_ADD_385_U139 P3_ADD_385_U138 ; P3_ADD_385_U70
g22998 nand P3_ADD_385_U141 P3_ADD_385_U140 ; P3_ADD_385_U71
g22999 nand P3_ADD_385_U143 P3_ADD_385_U142 ; P3_ADD_385_U72
g23000 nand P3_ADD_385_U145 P3_ADD_385_U144 ; P3_ADD_385_U73
g23001 nand P3_ADD_385_U147 P3_ADD_385_U146 ; P3_ADD_385_U74
g23002 nand P3_ADD_385_U149 P3_ADD_385_U148 ; P3_ADD_385_U75
g23003 nand P3_ADD_385_U151 P3_ADD_385_U150 ; P3_ADD_385_U76
g23004 nand P3_ADD_385_U153 P3_ADD_385_U152 ; P3_ADD_385_U77
g23005 nand P3_ADD_385_U155 P3_ADD_385_U154 ; P3_ADD_385_U78
g23006 nand P3_ADD_385_U157 P3_ADD_385_U156 ; P3_ADD_385_U79
g23007 nand P3_ADD_385_U159 P3_ADD_385_U158 ; P3_ADD_385_U80
g23008 nand P3_ADD_385_U161 P3_ADD_385_U160 ; P3_ADD_385_U81
g23009 nand P3_ADD_385_U163 P3_ADD_385_U162 ; P3_ADD_385_U82
g23010 nand P3_ADD_385_U165 P3_ADD_385_U164 ; P3_ADD_385_U83
g23011 nand P3_ADD_385_U167 P3_ADD_385_U166 ; P3_ADD_385_U84
g23012 nand P3_ADD_385_U169 P3_ADD_385_U168 ; P3_ADD_385_U85
g23013 nand P3_ADD_385_U171 P3_ADD_385_U170 ; P3_ADD_385_U86
g23014 nand P3_ADD_385_U173 P3_ADD_385_U172 ; P3_ADD_385_U87
g23015 nand P3_ADD_385_U175 P3_ADD_385_U174 ; P3_ADD_385_U88
g23016 nand P3_ADD_385_U177 P3_ADD_385_U176 ; P3_ADD_385_U89
g23017 nand P3_ADD_385_U179 P3_ADD_385_U178 ; P3_ADD_385_U90
g23018 nand P3_ADD_385_U181 P3_ADD_385_U180 ; P3_ADD_385_U91
g23019 nand P3_ADD_385_U183 P3_ADD_385_U182 ; P3_ADD_385_U92
g23020 nand P3_ADD_385_U185 P3_ADD_385_U184 ; P3_ADD_385_U93
g23021 nand P3_ADD_385_U187 P3_ADD_385_U186 ; P3_ADD_385_U94
g23022 nand P3_ADD_385_U189 P3_ADD_385_U188 ; P3_ADD_385_U95
g23023 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_385_U96
g23024 nand P3_ADD_385_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_385_U97
g23025 not P3_ADD_385_U7 ; P3_ADD_385_U98
g23026 not P3_ADD_385_U9 ; P3_ADD_385_U99
g23027 not P3_ADD_385_U11 ; P3_ADD_385_U100
g23028 not P3_ADD_385_U13 ; P3_ADD_385_U101
g23029 not P3_ADD_385_U15 ; P3_ADD_385_U102
g23030 not P3_ADD_385_U17 ; P3_ADD_385_U103
g23031 not P3_ADD_385_U19 ; P3_ADD_385_U104
g23032 not P3_ADD_385_U22 ; P3_ADD_385_U105
g23033 not P3_ADD_385_U23 ; P3_ADD_385_U106
g23034 not P3_ADD_385_U25 ; P3_ADD_385_U107
g23035 not P3_ADD_385_U27 ; P3_ADD_385_U108
g23036 not P3_ADD_385_U29 ; P3_ADD_385_U109
g23037 not P3_ADD_385_U31 ; P3_ADD_385_U110
g23038 not P3_ADD_385_U33 ; P3_ADD_385_U111
g23039 not P3_ADD_385_U35 ; P3_ADD_385_U112
g23040 not P3_ADD_385_U37 ; P3_ADD_385_U113
g23041 not P3_ADD_385_U39 ; P3_ADD_385_U114
g23042 not P3_ADD_385_U41 ; P3_ADD_385_U115
g23043 not P3_ADD_385_U43 ; P3_ADD_385_U116
g23044 not P3_ADD_385_U45 ; P3_ADD_385_U117
g23045 not P3_ADD_385_U47 ; P3_ADD_385_U118
g23046 not P3_ADD_385_U49 ; P3_ADD_385_U119
g23047 not P3_ADD_385_U51 ; P3_ADD_385_U120
g23048 not P3_ADD_385_U53 ; P3_ADD_385_U121
g23049 not P3_ADD_385_U55 ; P3_ADD_385_U122
g23050 not P3_ADD_385_U57 ; P3_ADD_385_U123
g23051 not P3_ADD_385_U59 ; P3_ADD_385_U124
g23052 not P3_ADD_385_U61 ; P3_ADD_385_U125
g23053 not P3_ADD_385_U63 ; P3_ADD_385_U126
g23054 not P3_ADD_385_U97 ; P3_ADD_385_U127
g23055 nand P3_ADD_385_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_385_U128
g23056 nand P3_ADD_385_U105 P3_ADD_385_U21 ; P3_ADD_385_U129
g23057 nand P3_ADD_385_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_385_U130
g23058 nand P3_ADD_385_U104 P3_ADD_385_U20 ; P3_ADD_385_U131
g23059 nand P3_ADD_385_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_385_U132
g23060 nand P3_ADD_385_U103 P3_ADD_385_U18 ; P3_ADD_385_U133
g23061 nand P3_ADD_385_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_385_U134
g23062 nand P3_ADD_385_U102 P3_ADD_385_U16 ; P3_ADD_385_U135
g23063 nand P3_ADD_385_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_385_U136
g23064 nand P3_ADD_385_U101 P3_ADD_385_U14 ; P3_ADD_385_U137
g23065 nand P3_ADD_385_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_385_U138
g23066 nand P3_ADD_385_U100 P3_ADD_385_U12 ; P3_ADD_385_U139
g23067 nand P3_ADD_385_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_385_U140
g23068 nand P3_ADD_385_U99 P3_ADD_385_U10 ; P3_ADD_385_U141
g23069 nand P3_ADD_385_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_385_U142
g23070 nand P3_ADD_385_U127 P3_ADD_385_U96 ; P3_ADD_385_U143
g23071 nand P3_ADD_385_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_385_U144
g23072 nand P3_ADD_385_U126 P3_ADD_385_U64 ; P3_ADD_385_U145
g23073 nand P3_ADD_385_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_385_U146
g23074 nand P3_ADD_385_U98 P3_ADD_385_U8 ; P3_ADD_385_U147
g23075 nand P3_ADD_385_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_385_U148
g23076 nand P3_ADD_385_U125 P3_ADD_385_U62 ; P3_ADD_385_U149
g23077 nand P3_ADD_385_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_385_U150
g23078 nand P3_ADD_385_U124 P3_ADD_385_U60 ; P3_ADD_385_U151
g23079 nand P3_ADD_385_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_385_U152
g23080 nand P3_ADD_385_U123 P3_ADD_385_U58 ; P3_ADD_385_U153
g23081 nand P3_ADD_385_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_385_U154
g23082 nand P3_ADD_385_U122 P3_ADD_385_U56 ; P3_ADD_385_U155
g23083 nand P3_ADD_385_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_385_U156
g23084 nand P3_ADD_385_U121 P3_ADD_385_U54 ; P3_ADD_385_U157
g23085 nand P3_ADD_385_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_385_U158
g23086 nand P3_ADD_385_U120 P3_ADD_385_U52 ; P3_ADD_385_U159
g23087 nand P3_ADD_385_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_385_U160
g23088 nand P3_ADD_385_U119 P3_ADD_385_U50 ; P3_ADD_385_U161
g23089 nand P3_ADD_385_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_385_U162
g23090 nand P3_ADD_385_U118 P3_ADD_385_U48 ; P3_ADD_385_U163
g23091 nand P3_ADD_385_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_385_U164
g23092 nand P3_ADD_385_U117 P3_ADD_385_U46 ; P3_ADD_385_U165
g23093 nand P3_ADD_385_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_385_U166
g23094 nand P3_ADD_385_U116 P3_ADD_385_U44 ; P3_ADD_385_U167
g23095 nand P3_ADD_385_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_385_U168
g23096 nand P3_ADD_385_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_385_U169
g23097 nand P3_ADD_385_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_385_U170
g23098 nand P3_ADD_385_U115 P3_ADD_385_U42 ; P3_ADD_385_U171
g23099 nand P3_ADD_385_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_385_U172
g23100 nand P3_ADD_385_U114 P3_ADD_385_U40 ; P3_ADD_385_U173
g23101 nand P3_ADD_385_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_385_U174
g23102 nand P3_ADD_385_U113 P3_ADD_385_U38 ; P3_ADD_385_U175
g23103 nand P3_ADD_385_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_385_U176
g23104 nand P3_ADD_385_U112 P3_ADD_385_U36 ; P3_ADD_385_U177
g23105 nand P3_ADD_385_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_385_U178
g23106 nand P3_ADD_385_U111 P3_ADD_385_U34 ; P3_ADD_385_U179
g23107 nand P3_ADD_385_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_385_U180
g23108 nand P3_ADD_385_U110 P3_ADD_385_U32 ; P3_ADD_385_U181
g23109 nand P3_ADD_385_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_385_U182
g23110 nand P3_ADD_385_U109 P3_ADD_385_U30 ; P3_ADD_385_U183
g23111 nand P3_ADD_385_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_385_U184
g23112 nand P3_ADD_385_U108 P3_ADD_385_U28 ; P3_ADD_385_U185
g23113 nand P3_ADD_385_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_385_U186
g23114 nand P3_ADD_385_U107 P3_ADD_385_U26 ; P3_ADD_385_U187
g23115 nand P3_ADD_385_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_385_U188
g23116 nand P3_ADD_385_U106 P3_ADD_385_U24 ; P3_ADD_385_U189
g23117 nand P3_ADD_357_U15 P3_ADD_357_U23 ; P3_ADD_357_U6
g23118 and P3_ADD_357_U29 P3_ADD_357_U11 ; P3_ADD_357_U7
g23119 and P3_ADD_357_U27 P3_ADD_357_U12 ; P3_ADD_357_U8
g23120 and P3_ADD_357_U25 P3_ADD_357_U6 ; P3_ADD_357_U9
g23121 not P3_SUB_357_U10 ; P3_ADD_357_U10
g23122 or P3_SUB_357_U7 P3_SUB_357_U12 P3_SUB_357_U11 ; P3_ADD_357_U11
g23123 nand P3_ADD_357_U14 P3_ADD_357_U22 ; P3_ADD_357_U12
g23124 nand P3_ADD_357_U35 P3_ADD_357_U34 ; P3_ADD_357_U13
g23125 nor P3_SUB_357_U13 P3_SUB_357_U9 ; P3_ADD_357_U14
g23126 nor P3_SUB_357_U6 P3_SUB_357_U8 ; P3_ADD_357_U15
g23127 not P3_SUB_357_U6 ; P3_ADD_357_U16
g23128 and P3_ADD_357_U31 P3_ADD_357_U30 ; P3_ADD_357_U17
g23129 not P3_SUB_357_U13 ; P3_ADD_357_U18
g23130 and P3_ADD_357_U33 P3_ADD_357_U32 ; P3_ADD_357_U19
g23131 not P3_SUB_357_U7 ; P3_ADD_357_U20
g23132 not P3_SUB_357_U12 ; P3_ADD_357_U21
g23133 not P3_ADD_357_U11 ; P3_ADD_357_U22
g23134 not P3_ADD_357_U12 ; P3_ADD_357_U23
g23135 nand P3_ADD_357_U23 P3_ADD_357_U16 ; P3_ADD_357_U24
g23136 nand P3_SUB_357_U8 P3_ADD_357_U24 ; P3_ADD_357_U25
g23137 nand P3_ADD_357_U22 P3_ADD_357_U18 ; P3_ADD_357_U26
g23138 nand P3_SUB_357_U9 P3_ADD_357_U26 ; P3_ADD_357_U27
g23139 or P3_SUB_357_U7 P3_SUB_357_U12 ; P3_ADD_357_U28
g23140 nand P3_SUB_357_U11 P3_ADD_357_U28 ; P3_ADD_357_U29
g23141 nand P3_SUB_357_U6 P3_ADD_357_U12 ; P3_ADD_357_U30
g23142 nand P3_ADD_357_U23 P3_ADD_357_U16 ; P3_ADD_357_U31
g23143 nand P3_SUB_357_U13 P3_ADD_357_U11 ; P3_ADD_357_U32
g23144 nand P3_ADD_357_U22 P3_ADD_357_U18 ; P3_ADD_357_U33
g23145 nand P3_SUB_357_U7 P3_ADD_357_U21 ; P3_ADD_357_U34
g23146 nand P3_SUB_357_U12 P3_ADD_357_U20 ; P3_ADD_357_U35
g23147 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_547_U5
g23148 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_547_U6
g23149 nand P3_INSTADDRPOINTER_REG_0__SCAN_IN P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_547_U7
g23150 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_547_U8
g23151 nand P3_ADD_547_U98 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_547_U9
g23152 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_547_U10
g23153 nand P3_ADD_547_U99 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_547_U11
g23154 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_547_U12
g23155 nand P3_ADD_547_U100 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_547_U13
g23156 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_547_U14
g23157 nand P3_ADD_547_U101 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_547_U15
g23158 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_547_U16
g23159 nand P3_ADD_547_U102 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_547_U17
g23160 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_547_U18
g23161 nand P3_ADD_547_U103 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_547_U19
g23162 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_547_U20
g23163 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_547_U21
g23164 nand P3_ADD_547_U104 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_547_U22
g23165 nand P3_ADD_547_U105 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_547_U23
g23166 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_547_U24
g23167 nand P3_ADD_547_U106 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_547_U25
g23168 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_547_U26
g23169 nand P3_ADD_547_U107 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_547_U27
g23170 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_547_U28
g23171 nand P3_ADD_547_U108 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_547_U29
g23172 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_547_U30
g23173 nand P3_ADD_547_U109 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_547_U31
g23174 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_547_U32
g23175 nand P3_ADD_547_U110 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_547_U33
g23176 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_547_U34
g23177 nand P3_ADD_547_U111 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_547_U35
g23178 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_547_U36
g23179 nand P3_ADD_547_U112 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_547_U37
g23180 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_547_U38
g23181 nand P3_ADD_547_U113 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_547_U39
g23182 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_547_U40
g23183 nand P3_ADD_547_U114 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_547_U41
g23184 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_547_U42
g23185 nand P3_ADD_547_U115 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_547_U43
g23186 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_547_U44
g23187 nand P3_ADD_547_U116 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_547_U45
g23188 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_547_U46
g23189 nand P3_ADD_547_U117 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_547_U47
g23190 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_547_U48
g23191 nand P3_ADD_547_U118 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_547_U49
g23192 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_547_U50
g23193 nand P3_ADD_547_U119 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_547_U51
g23194 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_547_U52
g23195 nand P3_ADD_547_U120 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_547_U53
g23196 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_547_U54
g23197 nand P3_ADD_547_U121 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_547_U55
g23198 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_547_U56
g23199 nand P3_ADD_547_U122 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_547_U57
g23200 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_547_U58
g23201 nand P3_ADD_547_U123 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_547_U59
g23202 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_547_U60
g23203 nand P3_ADD_547_U124 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_547_U61
g23204 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_547_U62
g23205 nand P3_ADD_547_U125 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_547_U63
g23206 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_547_U64
g23207 nand P3_ADD_547_U129 P3_ADD_547_U128 ; P3_ADD_547_U65
g23208 nand P3_ADD_547_U131 P3_ADD_547_U130 ; P3_ADD_547_U66
g23209 nand P3_ADD_547_U133 P3_ADD_547_U132 ; P3_ADD_547_U67
g23210 nand P3_ADD_547_U135 P3_ADD_547_U134 ; P3_ADD_547_U68
g23211 nand P3_ADD_547_U137 P3_ADD_547_U136 ; P3_ADD_547_U69
g23212 nand P3_ADD_547_U139 P3_ADD_547_U138 ; P3_ADD_547_U70
g23213 nand P3_ADD_547_U141 P3_ADD_547_U140 ; P3_ADD_547_U71
g23214 nand P3_ADD_547_U143 P3_ADD_547_U142 ; P3_ADD_547_U72
g23215 nand P3_ADD_547_U145 P3_ADD_547_U144 ; P3_ADD_547_U73
g23216 nand P3_ADD_547_U147 P3_ADD_547_U146 ; P3_ADD_547_U74
g23217 nand P3_ADD_547_U149 P3_ADD_547_U148 ; P3_ADD_547_U75
g23218 nand P3_ADD_547_U151 P3_ADD_547_U150 ; P3_ADD_547_U76
g23219 nand P3_ADD_547_U153 P3_ADD_547_U152 ; P3_ADD_547_U77
g23220 nand P3_ADD_547_U155 P3_ADD_547_U154 ; P3_ADD_547_U78
g23221 nand P3_ADD_547_U157 P3_ADD_547_U156 ; P3_ADD_547_U79
g23222 nand P3_ADD_547_U159 P3_ADD_547_U158 ; P3_ADD_547_U80
g23223 nand P3_ADD_547_U161 P3_ADD_547_U160 ; P3_ADD_547_U81
g23224 nand P3_ADD_547_U163 P3_ADD_547_U162 ; P3_ADD_547_U82
g23225 nand P3_ADD_547_U165 P3_ADD_547_U164 ; P3_ADD_547_U83
g23226 nand P3_ADD_547_U167 P3_ADD_547_U166 ; P3_ADD_547_U84
g23227 nand P3_ADD_547_U169 P3_ADD_547_U168 ; P3_ADD_547_U85
g23228 nand P3_ADD_547_U171 P3_ADD_547_U170 ; P3_ADD_547_U86
g23229 nand P3_ADD_547_U173 P3_ADD_547_U172 ; P3_ADD_547_U87
g23230 nand P3_ADD_547_U175 P3_ADD_547_U174 ; P3_ADD_547_U88
g23231 nand P3_ADD_547_U177 P3_ADD_547_U176 ; P3_ADD_547_U89
g23232 nand P3_ADD_547_U179 P3_ADD_547_U178 ; P3_ADD_547_U90
g23233 nand P3_ADD_547_U181 P3_ADD_547_U180 ; P3_ADD_547_U91
g23234 nand P3_ADD_547_U183 P3_ADD_547_U182 ; P3_ADD_547_U92
g23235 nand P3_ADD_547_U185 P3_ADD_547_U184 ; P3_ADD_547_U93
g23236 nand P3_ADD_547_U187 P3_ADD_547_U186 ; P3_ADD_547_U94
g23237 nand P3_ADD_547_U189 P3_ADD_547_U188 ; P3_ADD_547_U95
g23238 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_547_U96
g23239 nand P3_ADD_547_U126 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_547_U97
g23240 not P3_ADD_547_U7 ; P3_ADD_547_U98
g23241 not P3_ADD_547_U9 ; P3_ADD_547_U99
g23242 not P3_ADD_547_U11 ; P3_ADD_547_U100
g23243 not P3_ADD_547_U13 ; P3_ADD_547_U101
g23244 not P3_ADD_547_U15 ; P3_ADD_547_U102
g23245 not P3_ADD_547_U17 ; P3_ADD_547_U103
g23246 not P3_ADD_547_U19 ; P3_ADD_547_U104
g23247 not P3_ADD_547_U22 ; P3_ADD_547_U105
g23248 not P3_ADD_547_U23 ; P3_ADD_547_U106
g23249 not P3_ADD_547_U25 ; P3_ADD_547_U107
g23250 not P3_ADD_547_U27 ; P3_ADD_547_U108
g23251 not P3_ADD_547_U29 ; P3_ADD_547_U109
g23252 not P3_ADD_547_U31 ; P3_ADD_547_U110
g23253 not P3_ADD_547_U33 ; P3_ADD_547_U111
g23254 not P3_ADD_547_U35 ; P3_ADD_547_U112
g23255 not P3_ADD_547_U37 ; P3_ADD_547_U113
g23256 not P3_ADD_547_U39 ; P3_ADD_547_U114
g23257 not P3_ADD_547_U41 ; P3_ADD_547_U115
g23258 not P3_ADD_547_U43 ; P3_ADD_547_U116
g23259 not P3_ADD_547_U45 ; P3_ADD_547_U117
g23260 not P3_ADD_547_U47 ; P3_ADD_547_U118
g23261 not P3_ADD_547_U49 ; P3_ADD_547_U119
g23262 not P3_ADD_547_U51 ; P3_ADD_547_U120
g23263 not P3_ADD_547_U53 ; P3_ADD_547_U121
g23264 not P3_ADD_547_U55 ; P3_ADD_547_U122
g23265 not P3_ADD_547_U57 ; P3_ADD_547_U123
g23266 not P3_ADD_547_U59 ; P3_ADD_547_U124
g23267 not P3_ADD_547_U61 ; P3_ADD_547_U125
g23268 not P3_ADD_547_U63 ; P3_ADD_547_U126
g23269 not P3_ADD_547_U97 ; P3_ADD_547_U127
g23270 nand P3_ADD_547_U22 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_547_U128
g23271 nand P3_ADD_547_U105 P3_ADD_547_U21 ; P3_ADD_547_U129
g23272 nand P3_ADD_547_U19 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_547_U130
g23273 nand P3_ADD_547_U104 P3_ADD_547_U20 ; P3_ADD_547_U131
g23274 nand P3_ADD_547_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_547_U132
g23275 nand P3_ADD_547_U103 P3_ADD_547_U18 ; P3_ADD_547_U133
g23276 nand P3_ADD_547_U15 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_547_U134
g23277 nand P3_ADD_547_U102 P3_ADD_547_U16 ; P3_ADD_547_U135
g23278 nand P3_ADD_547_U13 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_547_U136
g23279 nand P3_ADD_547_U101 P3_ADD_547_U14 ; P3_ADD_547_U137
g23280 nand P3_ADD_547_U11 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_547_U138
g23281 nand P3_ADD_547_U100 P3_ADD_547_U12 ; P3_ADD_547_U139
g23282 nand P3_ADD_547_U9 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_547_U140
g23283 nand P3_ADD_547_U99 P3_ADD_547_U10 ; P3_ADD_547_U141
g23284 nand P3_ADD_547_U97 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_547_U142
g23285 nand P3_ADD_547_U127 P3_ADD_547_U96 ; P3_ADD_547_U143
g23286 nand P3_ADD_547_U63 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_547_U144
g23287 nand P3_ADD_547_U126 P3_ADD_547_U64 ; P3_ADD_547_U145
g23288 nand P3_ADD_547_U7 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_547_U146
g23289 nand P3_ADD_547_U98 P3_ADD_547_U8 ; P3_ADD_547_U147
g23290 nand P3_ADD_547_U61 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_547_U148
g23291 nand P3_ADD_547_U125 P3_ADD_547_U62 ; P3_ADD_547_U149
g23292 nand P3_ADD_547_U59 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_547_U150
g23293 nand P3_ADD_547_U124 P3_ADD_547_U60 ; P3_ADD_547_U151
g23294 nand P3_ADD_547_U57 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_547_U152
g23295 nand P3_ADD_547_U123 P3_ADD_547_U58 ; P3_ADD_547_U153
g23296 nand P3_ADD_547_U55 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_547_U154
g23297 nand P3_ADD_547_U122 P3_ADD_547_U56 ; P3_ADD_547_U155
g23298 nand P3_ADD_547_U53 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_547_U156
g23299 nand P3_ADD_547_U121 P3_ADD_547_U54 ; P3_ADD_547_U157
g23300 nand P3_ADD_547_U51 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_547_U158
g23301 nand P3_ADD_547_U120 P3_ADD_547_U52 ; P3_ADD_547_U159
g23302 nand P3_ADD_547_U49 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_547_U160
g23303 nand P3_ADD_547_U119 P3_ADD_547_U50 ; P3_ADD_547_U161
g23304 nand P3_ADD_547_U47 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_547_U162
g23305 nand P3_ADD_547_U118 P3_ADD_547_U48 ; P3_ADD_547_U163
g23306 nand P3_ADD_547_U45 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_547_U164
g23307 nand P3_ADD_547_U117 P3_ADD_547_U46 ; P3_ADD_547_U165
g23308 nand P3_ADD_547_U43 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_547_U166
g23309 nand P3_ADD_547_U116 P3_ADD_547_U44 ; P3_ADD_547_U167
g23310 nand P3_ADD_547_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_547_U168
g23311 nand P3_ADD_547_U6 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_547_U169
g23312 nand P3_ADD_547_U41 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_547_U170
g23313 nand P3_ADD_547_U115 P3_ADD_547_U42 ; P3_ADD_547_U171
g23314 nand P3_ADD_547_U39 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_547_U172
g23315 nand P3_ADD_547_U114 P3_ADD_547_U40 ; P3_ADD_547_U173
g23316 nand P3_ADD_547_U37 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_547_U174
g23317 nand P3_ADD_547_U113 P3_ADD_547_U38 ; P3_ADD_547_U175
g23318 nand P3_ADD_547_U35 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_547_U176
g23319 nand P3_ADD_547_U112 P3_ADD_547_U36 ; P3_ADD_547_U177
g23320 nand P3_ADD_547_U33 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_547_U178
g23321 nand P3_ADD_547_U111 P3_ADD_547_U34 ; P3_ADD_547_U179
g23322 nand P3_ADD_547_U31 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_547_U180
g23323 nand P3_ADD_547_U110 P3_ADD_547_U32 ; P3_ADD_547_U181
g23324 nand P3_ADD_547_U29 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_547_U182
g23325 nand P3_ADD_547_U109 P3_ADD_547_U30 ; P3_ADD_547_U183
g23326 nand P3_ADD_547_U27 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_547_U184
g23327 nand P3_ADD_547_U108 P3_ADD_547_U28 ; P3_ADD_547_U185
g23328 nand P3_ADD_547_U25 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_547_U186
g23329 nand P3_ADD_547_U107 P3_ADD_547_U26 ; P3_ADD_547_U187
g23330 nand P3_ADD_547_U23 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_547_U188
g23331 nand P3_ADD_547_U106 P3_ADD_547_U24 ; P3_ADD_547_U189
g23332 nand P3_SUB_412_U43 P3_SUB_412_U42 ; P3_SUB_412_U6
g23333 nand P3_SUB_412_U27 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_412_U7
g23334 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_412_U8
g23335 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_412_U9
g23336 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_412_U10
g23337 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_412_U11
g23338 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_412_U12
g23339 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_412_U13
g23340 nand P3_SUB_412_U39 P3_SUB_412_U38 ; P3_SUB_412_U14
g23341 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_412_U15
g23342 nand P3_SUB_412_U48 P3_SUB_412_U47 ; P3_SUB_412_U16
g23343 nand P3_SUB_412_U53 P3_SUB_412_U52 ; P3_SUB_412_U17
g23344 nand P3_SUB_412_U58 P3_SUB_412_U57 ; P3_SUB_412_U18
g23345 nand P3_SUB_412_U63 P3_SUB_412_U62 ; P3_SUB_412_U19
g23346 nand P3_SUB_412_U45 P3_SUB_412_U44 ; P3_SUB_412_U20
g23347 nand P3_SUB_412_U50 P3_SUB_412_U49 ; P3_SUB_412_U21
g23348 nand P3_SUB_412_U55 P3_SUB_412_U54 ; P3_SUB_412_U22
g23349 nand P3_SUB_412_U60 P3_SUB_412_U59 ; P3_SUB_412_U23
g23350 nand P3_SUB_412_U35 P3_SUB_412_U34 ; P3_SUB_412_U24
g23351 nand P3_SUB_412_U31 P3_SUB_412_U30 ; P3_SUB_412_U25
g23352 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_412_U26
g23353 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_412_U27
g23354 not P3_SUB_412_U7 ; P3_SUB_412_U28
g23355 nand P3_SUB_412_U28 P3_SUB_412_U8 ; P3_SUB_412_U29
g23356 nand P3_SUB_412_U29 P3_SUB_412_U26 ; P3_SUB_412_U30
g23357 nand P3_SUB_412_U7 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_412_U31
g23358 not P3_SUB_412_U25 ; P3_SUB_412_U32
g23359 nand P3_SUB_412_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_412_U33
g23360 nand P3_SUB_412_U33 P3_SUB_412_U25 ; P3_SUB_412_U34
g23361 nand P3_SUB_412_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_412_U35
g23362 not P3_SUB_412_U24 ; P3_SUB_412_U36
g23363 nand P3_SUB_412_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_412_U37
g23364 nand P3_SUB_412_U37 P3_SUB_412_U24 ; P3_SUB_412_U38
g23365 nand P3_SUB_412_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_412_U39
g23366 not P3_SUB_412_U14 ; P3_SUB_412_U40
g23367 nand P3_SUB_412_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_412_U41
g23368 nand P3_SUB_412_U40 P3_SUB_412_U41 ; P3_SUB_412_U42
g23369 nand P3_SUB_412_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_412_U43
g23370 nand P3_SUB_412_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_412_U44
g23371 nand P3_SUB_412_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_412_U45
g23372 not P3_SUB_412_U20 ; P3_SUB_412_U46
g23373 nand P3_SUB_412_U46 P3_SUB_412_U40 ; P3_SUB_412_U47
g23374 nand P3_SUB_412_U20 P3_SUB_412_U14 ; P3_SUB_412_U48
g23375 nand P3_SUB_412_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_412_U49
g23376 nand P3_SUB_412_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_412_U50
g23377 not P3_SUB_412_U21 ; P3_SUB_412_U51
g23378 nand P3_SUB_412_U36 P3_SUB_412_U51 ; P3_SUB_412_U52
g23379 nand P3_SUB_412_U21 P3_SUB_412_U24 ; P3_SUB_412_U53
g23380 nand P3_SUB_412_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_412_U54
g23381 nand P3_SUB_412_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_412_U55
g23382 not P3_SUB_412_U22 ; P3_SUB_412_U56
g23383 nand P3_SUB_412_U32 P3_SUB_412_U56 ; P3_SUB_412_U57
g23384 nand P3_SUB_412_U22 P3_SUB_412_U25 ; P3_SUB_412_U58
g23385 nand P3_SUB_412_U8 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_412_U59
g23386 nand P3_SUB_412_U26 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_412_U60
g23387 not P3_SUB_412_U23 ; P3_SUB_412_U61
g23388 nand P3_SUB_412_U61 P3_SUB_412_U28 ; P3_SUB_412_U62
g23389 nand P3_SUB_412_U23 P3_SUB_412_U7 ; P3_SUB_412_U63
g23390 and P3_ADD_371_1212_U133 P3_ADD_371_1212_U132 ; P3_ADD_371_1212_U4
g23391 and P3_ADD_371_1212_U196 P3_ADD_371_1212_U48 ; P3_ADD_371_1212_U5
g23392 and P3_ADD_371_1212_U194 P3_ADD_371_1212_U49 ; P3_ADD_371_1212_U6
g23393 and P3_ADD_371_1212_U192 P3_ADD_371_1212_U78 ; P3_ADD_371_1212_U7
g23394 and P3_ADD_371_1212_U191 P3_ADD_371_1212_U53 ; P3_ADD_371_1212_U8
g23395 and P3_ADD_371_1212_U189 P3_ADD_371_1212_U56 ; P3_ADD_371_1212_U9
g23396 and P3_ADD_371_1212_U187 P3_ADD_371_1212_U59 ; P3_ADD_371_1212_U10
g23397 and P3_ADD_371_1212_U185 P3_ADD_371_1212_U168 ; P3_ADD_371_1212_U11
g23398 and P3_ADD_371_1212_U184 P3_ADD_371_1212_U62 ; P3_ADD_371_1212_U12
g23399 and P3_ADD_371_1212_U183 P3_ADD_371_1212_U65 ; P3_ADD_371_1212_U13
g23400 and P3_ADD_371_1212_U181 P3_ADD_371_1212_U68 ; P3_ADD_371_1212_U14
g23401 and P3_ADD_371_1212_U179 P3_ADD_371_1212_U70 ; P3_ADD_371_1212_U15
g23402 and P3_ADD_371_1212_U178 P3_ADD_371_1212_U73 ; P3_ADD_371_1212_U16
g23403 and P3_ADD_371_1212_U176 P3_ADD_371_1212_U75 ; P3_ADD_371_1212_U17
g23404 and P3_ADD_371_1212_U162 P3_ADD_371_1212_U159 ; P3_ADD_371_1212_U18
g23405 and P3_ADD_371_1212_U155 P3_ADD_371_1212_U152 ; P3_ADD_371_1212_U19
g23406 nand P3_ADD_371_1212_U255 P3_ADD_371_1212_U254 P3_ADD_371_1212_U203 ; P3_ADD_371_1212_U20
g23407 not P3_ADD_371_U20 ; P3_ADD_371_1212_U21
g23408 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_371_1212_U22
g23409 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_371_1212_U23
g23410 nand P3_ADD_371_U20 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_371_1212_U24
g23411 not P3_ADD_371_U19 ; P3_ADD_371_1212_U25
g23412 not P3_ADD_371_U5 ; P3_ADD_371_1212_U26
g23413 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_371_1212_U27
g23414 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_371_1212_U28
g23415 nand P3_ADD_371_U5 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_371_1212_U29
g23416 not P3_ADD_371_U25 ; P3_ADD_371_1212_U30
g23417 not P3_ADD_371_U4 ; P3_ADD_371_1212_U31
g23418 not P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_371_1212_U32
g23419 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_371_1212_U33
g23420 nand P3_ADD_371_U4 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_371_1212_U34
g23421 not P3_ADD_371_U21 ; P3_ADD_371_1212_U35
g23422 not P3_ADD_371_U18 ; P3_ADD_371_1212_U36
g23423 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_371_1212_U37
g23424 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_371_1212_U38
g23425 not P3_ADD_371_U17 ; P3_ADD_371_1212_U39
g23426 not P3_ADD_371_U6 ; P3_ADD_371_1212_U40
g23427 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_371_1212_U41
g23428 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_371_1212_U42
g23429 nand P3_ADD_371_1212_U94 P3_ADD_371_1212_U130 ; P3_ADD_371_1212_U43
g23430 nand P3_ADD_371_1212_U77 P3_ADD_371_1212_U123 ; P3_ADD_371_1212_U44
g23431 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_371_1212_U45
g23432 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_371_1212_U46
g23433 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_371_1212_U47
g23434 nand P3_ADD_371_1212_U99 P3_ADD_371_1212_U108 ; P3_ADD_371_1212_U48
g23435 nand P3_ADD_371_1212_U100 P3_ADD_371_1212_U117 ; P3_ADD_371_1212_U49
g23436 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_371_1212_U50
g23437 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_371_1212_U51
g23438 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_371_1212_U52
g23439 nand P3_ADD_371_1212_U163 P3_ADD_371_1212_U101 ; P3_ADD_371_1212_U53
g23440 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_371_1212_U54
g23441 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_371_1212_U55
g23442 nand P3_ADD_371_1212_U102 P3_ADD_371_1212_U165 ; P3_ADD_371_1212_U56
g23443 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_371_1212_U57
g23444 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_371_1212_U58
g23445 nand P3_ADD_371_1212_U103 P3_ADD_371_1212_U166 ; P3_ADD_371_1212_U59
g23446 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_371_1212_U60
g23447 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_371_1212_U61
g23448 nand P3_ADD_371_1212_U104 P3_ADD_371_1212_U167 ; P3_ADD_371_1212_U62
g23449 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_371_1212_U63
g23450 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_371_1212_U64
g23451 nand P3_ADD_371_1212_U105 P3_ADD_371_1212_U169 ; P3_ADD_371_1212_U65
g23452 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_371_1212_U66
g23453 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_371_1212_U67
g23454 nand P3_ADD_371_1212_U106 P3_ADD_371_1212_U170 ; P3_ADD_371_1212_U68
g23455 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_371_1212_U69
g23456 nand P3_ADD_371_1212_U171 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_371_1212_U70
g23457 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_371_1212_U71
g23458 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_371_1212_U72
g23459 nand P3_ADD_371_1212_U107 P3_ADD_371_1212_U172 ; P3_ADD_371_1212_U73
g23460 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_371_1212_U74
g23461 nand P3_ADD_371_1212_U173 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_371_1212_U75
g23462 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_371_1212_U76
g23463 nand P3_ADD_371_U21 P3_ADD_371_1212_U121 ; P3_ADD_371_1212_U77
g23464 nand P3_ADD_371_1212_U163 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_371_1212_U78
g23465 nand P3_ADD_371_1212_U239 P3_ADD_371_1212_U238 ; P3_ADD_371_1212_U79
g23466 nand P3_ADD_371_1212_U246 P3_ADD_371_1212_U245 ; P3_ADD_371_1212_U80
g23467 nand P3_ADD_371_1212_U248 P3_ADD_371_1212_U247 ; P3_ADD_371_1212_U81
g23468 nand P3_ADD_371_1212_U250 P3_ADD_371_1212_U249 ; P3_ADD_371_1212_U82
g23469 nand P3_ADD_371_1212_U257 P3_ADD_371_1212_U256 ; P3_ADD_371_1212_U83
g23470 nand P3_ADD_371_1212_U259 P3_ADD_371_1212_U258 ; P3_ADD_371_1212_U84
g23471 nand P3_ADD_371_1212_U261 P3_ADD_371_1212_U260 ; P3_ADD_371_1212_U85
g23472 nand P3_ADD_371_1212_U263 P3_ADD_371_1212_U262 ; P3_ADD_371_1212_U86
g23473 nand P3_ADD_371_1212_U265 P3_ADD_371_1212_U264 ; P3_ADD_371_1212_U87
g23474 nand P3_ADD_371_1212_U212 P3_ADD_371_1212_U211 ; P3_ADD_371_1212_U88
g23475 nand P3_ADD_371_1212_U219 P3_ADD_371_1212_U218 ; P3_ADD_371_1212_U89
g23476 nand P3_ADD_371_1212_U226 P3_ADD_371_1212_U225 ; P3_ADD_371_1212_U90
g23477 nand P3_ADD_371_1212_U233 P3_ADD_371_1212_U232 ; P3_ADD_371_1212_U91
g23478 nand P3_ADD_371_1212_U237 P3_ADD_371_1212_U236 ; P3_ADD_371_1212_U92
g23479 nand P3_ADD_371_1212_U244 P3_ADD_371_1212_U243 ; P3_ADD_371_1212_U93
g23480 and P3_ADD_371_1212_U129 P3_ADD_371_1212_U128 ; P3_ADD_371_1212_U94
g23481 and P3_ADD_371_1212_U137 P3_ADD_371_1212_U136 ; P3_ADD_371_1212_U95
g23482 and P3_ADD_371_1212_U228 P3_ADD_371_1212_U227 P3_ADD_371_1212_U24 ; P3_ADD_371_1212_U96
g23483 and P3_ADD_371_1212_U154 P3_ADD_371_1212_U4 ; P3_ADD_371_1212_U97
g23484 and P3_ADD_371_1212_U235 P3_ADD_371_1212_U234 P3_ADD_371_1212_U29 ; P3_ADD_371_1212_U98
g23485 and P3_INSTADDRPOINTER_REG_9__SCAN_IN P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_371_1212_U99
g23486 and P3_INSTADDRPOINTER_REG_11__SCAN_IN P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_371_1212_U100
g23487 and P3_INSTADDRPOINTER_REG_13__SCAN_IN P3_INSTADDRPOINTER_REG_14__SCAN_IN P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_371_1212_U101
g23488 and P3_INSTADDRPOINTER_REG_16__SCAN_IN P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_371_1212_U102
g23489 and P3_INSTADDRPOINTER_REG_18__SCAN_IN P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_371_1212_U103
g23490 and P3_INSTADDRPOINTER_REG_20__SCAN_IN P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_371_1212_U104
g23491 and P3_INSTADDRPOINTER_REG_22__SCAN_IN P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_371_1212_U105
g23492 and P3_INSTADDRPOINTER_REG_24__SCAN_IN P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_371_1212_U106
g23493 and P3_INSTADDRPOINTER_REG_27__SCAN_IN P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_371_1212_U107
g23494 nand P3_ADD_371_1212_U148 P3_ADD_371_1212_U147 ; P3_ADD_371_1212_U108
g23495 and P3_ADD_371_1212_U205 P3_ADD_371_1212_U204 ; P3_ADD_371_1212_U109
g23496 and P3_ADD_371_1212_U207 P3_ADD_371_1212_U206 ; P3_ADD_371_1212_U110
g23497 nand P3_ADD_371_1212_U144 P3_ADD_371_1212_U118 P3_ADD_371_1212_U200 ; P3_ADD_371_1212_U111
g23498 and P3_ADD_371_1212_U214 P3_ADD_371_1212_U213 ; P3_ADD_371_1212_U112
g23499 nand P3_ADD_371_1212_U142 P3_ADD_371_1212_U141 ; P3_ADD_371_1212_U113
g23500 and P3_ADD_371_1212_U221 P3_ADD_371_1212_U220 ; P3_ADD_371_1212_U114
g23501 nand P3_ADD_371_1212_U95 P3_ADD_371_1212_U138 ; P3_ADD_371_1212_U115
g23502 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_371_1212_U116
g23503 not P3_ADD_371_1212_U48 ; P3_ADD_371_1212_U117
g23504 nand P3_ADD_371_1212_U113 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_371_1212_U118
g23505 nand P3_ADD_371_1212_U202 P3_ADD_371_1212_U201 ; P3_ADD_371_1212_U119
g23506 not P3_ADD_371_1212_U77 ; P3_ADD_371_1212_U120
g23507 not P3_ADD_371_1212_U34 ; P3_ADD_371_1212_U121
g23508 nand P3_ADD_371_1212_U35 P3_ADD_371_1212_U34 ; P3_ADD_371_1212_U122
g23509 nand P3_ADD_371_1212_U122 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_371_1212_U123
g23510 not P3_ADD_371_1212_U44 ; P3_ADD_371_1212_U124
g23511 or P3_ADD_371_U5 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_371_1212_U125
g23512 not P3_ADD_371_1212_U29 ; P3_ADD_371_1212_U126
g23513 nand P3_ADD_371_1212_U30 P3_ADD_371_1212_U29 ; P3_ADD_371_1212_U127
g23514 nand P3_ADD_371_1212_U127 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_371_1212_U128
g23515 nand P3_ADD_371_U25 P3_ADD_371_1212_U126 ; P3_ADD_371_1212_U129
g23516 nand P3_ADD_371_1212_U44 P3_ADD_371_1212_U119 ; P3_ADD_371_1212_U130
g23517 not P3_ADD_371_1212_U43 ; P3_ADD_371_1212_U131
g23518 or P3_ADD_371_U19 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_371_1212_U132
g23519 or P3_ADD_371_U20 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_371_1212_U133
g23520 not P3_ADD_371_1212_U24 ; P3_ADD_371_1212_U134
g23521 nand P3_ADD_371_1212_U25 P3_ADD_371_1212_U24 ; P3_ADD_371_1212_U135
g23522 nand P3_ADD_371_1212_U135 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_371_1212_U136
g23523 nand P3_ADD_371_U19 P3_ADD_371_1212_U134 ; P3_ADD_371_1212_U137
g23524 nand P3_ADD_371_1212_U4 P3_ADD_371_1212_U43 ; P3_ADD_371_1212_U138
g23525 not P3_ADD_371_1212_U115 ; P3_ADD_371_1212_U139
g23526 or P3_ADD_371_U18 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_371_1212_U140
g23527 nand P3_ADD_371_1212_U140 P3_ADD_371_1212_U115 ; P3_ADD_371_1212_U141
g23528 nand P3_ADD_371_U18 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_371_1212_U142
g23529 not P3_ADD_371_1212_U113 ; P3_ADD_371_1212_U143
g23530 nand P3_ADD_371_U17 P3_ADD_371_1212_U113 ; P3_ADD_371_1212_U144
g23531 not P3_ADD_371_1212_U111 ; P3_ADD_371_1212_U145
g23532 or P3_ADD_371_U6 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_371_1212_U146
g23533 nand P3_ADD_371_1212_U146 P3_ADD_371_1212_U111 ; P3_ADD_371_1212_U147
g23534 nand P3_ADD_371_U6 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_371_1212_U148
g23535 not P3_ADD_371_1212_U108 ; P3_ADD_371_1212_U149
g23536 or P3_ADD_371_U20 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_371_1212_U150
g23537 nand P3_ADD_371_1212_U150 P3_ADD_371_1212_U43 ; P3_ADD_371_1212_U151
g23538 nand P3_ADD_371_1212_U96 P3_ADD_371_1212_U151 ; P3_ADD_371_1212_U152
g23539 nand P3_ADD_371_1212_U131 P3_ADD_371_1212_U24 ; P3_ADD_371_1212_U153
g23540 nand P3_ADD_371_U19 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_371_1212_U154
g23541 nand P3_ADD_371_1212_U97 P3_ADD_371_1212_U153 ; P3_ADD_371_1212_U155
g23542 or P3_ADD_371_U20 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_371_1212_U156
g23543 or P3_ADD_371_U5 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_371_1212_U157
g23544 nand P3_ADD_371_1212_U157 P3_ADD_371_1212_U44 ; P3_ADD_371_1212_U158
g23545 nand P3_ADD_371_1212_U98 P3_ADD_371_1212_U158 ; P3_ADD_371_1212_U159
g23546 nand P3_ADD_371_1212_U124 P3_ADD_371_1212_U29 ; P3_ADD_371_1212_U160
g23547 nand P3_ADD_371_U25 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_371_1212_U161
g23548 nand P3_ADD_371_1212_U160 P3_ADD_371_1212_U161 P3_ADD_371_1212_U119 ; P3_ADD_371_1212_U162
g23549 not P3_ADD_371_1212_U49 ; P3_ADD_371_1212_U163
g23550 not P3_ADD_371_1212_U78 ; P3_ADD_371_1212_U164
g23551 not P3_ADD_371_1212_U53 ; P3_ADD_371_1212_U165
g23552 not P3_ADD_371_1212_U56 ; P3_ADD_371_1212_U166
g23553 not P3_ADD_371_1212_U59 ; P3_ADD_371_1212_U167
g23554 nand P3_ADD_371_1212_U167 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_371_1212_U168
g23555 not P3_ADD_371_1212_U62 ; P3_ADD_371_1212_U169
g23556 not P3_ADD_371_1212_U65 ; P3_ADD_371_1212_U170
g23557 not P3_ADD_371_1212_U68 ; P3_ADD_371_1212_U171
g23558 not P3_ADD_371_1212_U70 ; P3_ADD_371_1212_U172
g23559 not P3_ADD_371_1212_U73 ; P3_ADD_371_1212_U173
g23560 not P3_ADD_371_1212_U75 ; P3_ADD_371_1212_U174
g23561 or P3_ADD_371_U5 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_371_1212_U175
g23562 nand P3_ADD_371_1212_U74 P3_ADD_371_1212_U73 ; P3_ADD_371_1212_U176
g23563 nand P3_ADD_371_1212_U172 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_371_1212_U177
g23564 nand P3_ADD_371_1212_U71 P3_ADD_371_1212_U177 ; P3_ADD_371_1212_U178
g23565 nand P3_ADD_371_1212_U69 P3_ADD_371_1212_U68 ; P3_ADD_371_1212_U179
g23566 nand P3_ADD_371_1212_U170 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_371_1212_U180
g23567 nand P3_ADD_371_1212_U66 P3_ADD_371_1212_U180 ; P3_ADD_371_1212_U181
g23568 nand P3_ADD_371_1212_U169 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_371_1212_U182
g23569 nand P3_ADD_371_1212_U63 P3_ADD_371_1212_U182 ; P3_ADD_371_1212_U183
g23570 nand P3_ADD_371_1212_U61 P3_ADD_371_1212_U168 ; P3_ADD_371_1212_U184
g23571 nand P3_ADD_371_1212_U60 P3_ADD_371_1212_U59 ; P3_ADD_371_1212_U185
g23572 nand P3_ADD_371_1212_U166 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_371_1212_U186
g23573 nand P3_ADD_371_1212_U58 P3_ADD_371_1212_U186 ; P3_ADD_371_1212_U187
g23574 nand P3_ADD_371_1212_U165 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_371_1212_U188
g23575 nand P3_ADD_371_1212_U54 P3_ADD_371_1212_U188 ; P3_ADD_371_1212_U189
g23576 nand P3_ADD_371_1212_U164 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_371_1212_U190
g23577 nand P3_ADD_371_1212_U51 P3_ADD_371_1212_U190 ; P3_ADD_371_1212_U191
g23578 nand P3_ADD_371_1212_U50 P3_ADD_371_1212_U49 ; P3_ADD_371_1212_U192
g23579 nand P3_ADD_371_1212_U117 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_371_1212_U193
g23580 nand P3_ADD_371_1212_U47 P3_ADD_371_1212_U193 ; P3_ADD_371_1212_U194
g23581 nand P3_ADD_371_1212_U108 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_371_1212_U195
g23582 nand P3_ADD_371_1212_U45 P3_ADD_371_1212_U195 ; P3_ADD_371_1212_U196
g23583 nand P3_ADD_371_1212_U156 P3_ADD_371_1212_U24 ; P3_ADD_371_1212_U197
g23584 nand P3_ADD_371_1212_U174 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_371_1212_U198
g23585 nand P3_ADD_371_1212_U175 P3_ADD_371_1212_U29 ; P3_ADD_371_1212_U199
g23586 nand P3_ADD_371_U17 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_371_1212_U200
g23587 nand P3_ADD_371_1212_U125 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_371_1212_U201
g23588 nand P3_ADD_371_U25 P3_ADD_371_1212_U125 ; P3_ADD_371_1212_U202
g23589 nand P3_ADD_371_1212_U120 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_371_1212_U203
g23590 nand P3_ADD_371_1212_U108 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_371_1212_U204
g23591 nand P3_ADD_371_1212_U149 P3_ADD_371_1212_U42 ; P3_ADD_371_1212_U205
g23592 nand P3_ADD_371_1212_U40 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_371_1212_U206
g23593 nand P3_ADD_371_U6 P3_ADD_371_1212_U41 ; P3_ADD_371_1212_U207
g23594 nand P3_ADD_371_1212_U40 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_371_1212_U208
g23595 nand P3_ADD_371_U6 P3_ADD_371_1212_U41 ; P3_ADD_371_1212_U209
g23596 nand P3_ADD_371_1212_U209 P3_ADD_371_1212_U208 ; P3_ADD_371_1212_U210
g23597 nand P3_ADD_371_1212_U110 P3_ADD_371_1212_U111 ; P3_ADD_371_1212_U211
g23598 nand P3_ADD_371_1212_U145 P3_ADD_371_1212_U210 ; P3_ADD_371_1212_U212
g23599 nand P3_ADD_371_1212_U39 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_371_1212_U213
g23600 nand P3_ADD_371_U17 P3_ADD_371_1212_U38 ; P3_ADD_371_1212_U214
g23601 nand P3_ADD_371_1212_U39 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_371_1212_U215
g23602 nand P3_ADD_371_U17 P3_ADD_371_1212_U38 ; P3_ADD_371_1212_U216
g23603 nand P3_ADD_371_1212_U216 P3_ADD_371_1212_U215 ; P3_ADD_371_1212_U217
g23604 nand P3_ADD_371_1212_U112 P3_ADD_371_1212_U113 ; P3_ADD_371_1212_U218
g23605 nand P3_ADD_371_1212_U143 P3_ADD_371_1212_U217 ; P3_ADD_371_1212_U219
g23606 nand P3_ADD_371_1212_U36 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_371_1212_U220
g23607 nand P3_ADD_371_U18 P3_ADD_371_1212_U37 ; P3_ADD_371_1212_U221
g23608 nand P3_ADD_371_1212_U36 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_371_1212_U222
g23609 nand P3_ADD_371_U18 P3_ADD_371_1212_U37 ; P3_ADD_371_1212_U223
g23610 nand P3_ADD_371_1212_U223 P3_ADD_371_1212_U222 ; P3_ADD_371_1212_U224
g23611 nand P3_ADD_371_1212_U114 P3_ADD_371_1212_U115 ; P3_ADD_371_1212_U225
g23612 nand P3_ADD_371_1212_U139 P3_ADD_371_1212_U224 ; P3_ADD_371_1212_U226
g23613 nand P3_ADD_371_1212_U25 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_371_1212_U227
g23614 nand P3_ADD_371_U19 P3_ADD_371_1212_U23 ; P3_ADD_371_1212_U228
g23615 nand P3_ADD_371_1212_U21 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_371_1212_U229
g23616 nand P3_ADD_371_U20 P3_ADD_371_1212_U22 ; P3_ADD_371_1212_U230
g23617 nand P3_ADD_371_1212_U230 P3_ADD_371_1212_U229 ; P3_ADD_371_1212_U231
g23618 nand P3_ADD_371_1212_U197 P3_ADD_371_1212_U43 ; P3_ADD_371_1212_U232
g23619 nand P3_ADD_371_1212_U231 P3_ADD_371_1212_U131 ; P3_ADD_371_1212_U233
g23620 nand P3_ADD_371_1212_U30 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_371_1212_U234
g23621 nand P3_ADD_371_U25 P3_ADD_371_1212_U28 ; P3_ADD_371_1212_U235
g23622 nand P3_ADD_371_1212_U198 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_371_1212_U236
g23623 nand P3_ADD_371_1212_U174 P3_ADD_371_1212_U116 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_371_1212_U237
g23624 nand P3_ADD_371_1212_U75 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_371_1212_U238
g23625 nand P3_ADD_371_1212_U174 P3_ADD_371_1212_U76 ; P3_ADD_371_1212_U239
g23626 nand P3_ADD_371_1212_U26 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_371_1212_U240
g23627 nand P3_ADD_371_U5 P3_ADD_371_1212_U27 ; P3_ADD_371_1212_U241
g23628 nand P3_ADD_371_1212_U241 P3_ADD_371_1212_U240 ; P3_ADD_371_1212_U242
g23629 nand P3_ADD_371_1212_U199 P3_ADD_371_1212_U44 ; P3_ADD_371_1212_U243
g23630 nand P3_ADD_371_1212_U242 P3_ADD_371_1212_U124 ; P3_ADD_371_1212_U244
g23631 nand P3_ADD_371_1212_U70 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_371_1212_U245
g23632 nand P3_ADD_371_1212_U172 P3_ADD_371_1212_U72 ; P3_ADD_371_1212_U246
g23633 nand P3_ADD_371_1212_U65 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_371_1212_U247
g23634 nand P3_ADD_371_1212_U170 P3_ADD_371_1212_U67 ; P3_ADD_371_1212_U248
g23635 nand P3_ADD_371_1212_U62 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_371_1212_U249
g23636 nand P3_ADD_371_1212_U169 P3_ADD_371_1212_U64 ; P3_ADD_371_1212_U250
g23637 nand P3_ADD_371_1212_U34 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_371_1212_U251
g23638 nand P3_ADD_371_1212_U121 P3_ADD_371_1212_U33 ; P3_ADD_371_1212_U252
g23639 nand P3_ADD_371_1212_U252 P3_ADD_371_1212_U251 ; P3_ADD_371_1212_U253
g23640 nand P3_ADD_371_1212_U34 P3_ADD_371_1212_U33 P3_ADD_371_U21 ; P3_ADD_371_1212_U254
g23641 nand P3_ADD_371_1212_U253 P3_ADD_371_1212_U35 ; P3_ADD_371_1212_U255
g23642 nand P3_ADD_371_1212_U56 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_371_1212_U256
g23643 nand P3_ADD_371_1212_U166 P3_ADD_371_1212_U57 ; P3_ADD_371_1212_U257
g23644 nand P3_ADD_371_1212_U53 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_371_1212_U258
g23645 nand P3_ADD_371_1212_U165 P3_ADD_371_1212_U55 ; P3_ADD_371_1212_U259
g23646 nand P3_ADD_371_1212_U78 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_371_1212_U260
g23647 nand P3_ADD_371_1212_U164 P3_ADD_371_1212_U52 ; P3_ADD_371_1212_U261
g23648 nand P3_ADD_371_1212_U117 P3_ADD_371_1212_U46 ; P3_ADD_371_1212_U262
g23649 nand P3_ADD_371_1212_U48 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_371_1212_U263
g23650 nand P3_ADD_371_1212_U31 P3_INSTADDRPOINTER_REG_0__SCAN_IN ; P3_ADD_371_1212_U264
g23651 nand P3_ADD_371_U4 P3_ADD_371_1212_U32 ; P3_ADD_371_1212_U265
g23652 nand P3_SUB_504_U43 P3_SUB_504_U42 ; P3_SUB_504_U6
g23653 nand P3_SUB_504_U27 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_504_U7
g23654 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_504_U8
g23655 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_504_U9
g23656 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_504_U10
g23657 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_504_U11
g23658 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_504_U12
g23659 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_504_U13
g23660 nand P3_SUB_504_U39 P3_SUB_504_U38 ; P3_SUB_504_U14
g23661 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_504_U15
g23662 nand P3_SUB_504_U48 P3_SUB_504_U47 ; P3_SUB_504_U16
g23663 nand P3_SUB_504_U53 P3_SUB_504_U52 ; P3_SUB_504_U17
g23664 nand P3_SUB_504_U58 P3_SUB_504_U57 ; P3_SUB_504_U18
g23665 nand P3_SUB_504_U63 P3_SUB_504_U62 ; P3_SUB_504_U19
g23666 nand P3_SUB_504_U45 P3_SUB_504_U44 ; P3_SUB_504_U20
g23667 nand P3_SUB_504_U50 P3_SUB_504_U49 ; P3_SUB_504_U21
g23668 nand P3_SUB_504_U55 P3_SUB_504_U54 ; P3_SUB_504_U22
g23669 nand P3_SUB_504_U60 P3_SUB_504_U59 ; P3_SUB_504_U23
g23670 nand P3_SUB_504_U35 P3_SUB_504_U34 ; P3_SUB_504_U24
g23671 nand P3_SUB_504_U31 P3_SUB_504_U30 ; P3_SUB_504_U25
g23672 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_504_U26
g23673 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_504_U27
g23674 not P3_SUB_504_U7 ; P3_SUB_504_U28
g23675 nand P3_SUB_504_U28 P3_SUB_504_U8 ; P3_SUB_504_U29
g23676 nand P3_SUB_504_U29 P3_SUB_504_U26 ; P3_SUB_504_U30
g23677 nand P3_SUB_504_U7 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_504_U31
g23678 not P3_SUB_504_U25 ; P3_SUB_504_U32
g23679 nand P3_SUB_504_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_504_U33
g23680 nand P3_SUB_504_U33 P3_SUB_504_U25 ; P3_SUB_504_U34
g23681 nand P3_SUB_504_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_504_U35
g23682 not P3_SUB_504_U24 ; P3_SUB_504_U36
g23683 nand P3_SUB_504_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_504_U37
g23684 nand P3_SUB_504_U37 P3_SUB_504_U24 ; P3_SUB_504_U38
g23685 nand P3_SUB_504_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_504_U39
g23686 not P3_SUB_504_U14 ; P3_SUB_504_U40
g23687 nand P3_SUB_504_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_504_U41
g23688 nand P3_SUB_504_U40 P3_SUB_504_U41 ; P3_SUB_504_U42
g23689 nand P3_SUB_504_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_504_U43
g23690 nand P3_SUB_504_U13 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_504_U44
g23691 nand P3_SUB_504_U15 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_504_U45
g23692 not P3_SUB_504_U20 ; P3_SUB_504_U46
g23693 nand P3_SUB_504_U46 P3_SUB_504_U40 ; P3_SUB_504_U47
g23694 nand P3_SUB_504_U20 P3_SUB_504_U14 ; P3_SUB_504_U48
g23695 nand P3_SUB_504_U12 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_504_U49
g23696 nand P3_SUB_504_U11 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_504_U50
g23697 not P3_SUB_504_U21 ; P3_SUB_504_U51
g23698 nand P3_SUB_504_U36 P3_SUB_504_U51 ; P3_SUB_504_U52
g23699 nand P3_SUB_504_U21 P3_SUB_504_U24 ; P3_SUB_504_U53
g23700 nand P3_SUB_504_U10 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_504_U54
g23701 nand P3_SUB_504_U9 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_504_U55
g23702 not P3_SUB_504_U22 ; P3_SUB_504_U56
g23703 nand P3_SUB_504_U32 P3_SUB_504_U56 ; P3_SUB_504_U57
g23704 nand P3_SUB_504_U22 P3_SUB_504_U25 ; P3_SUB_504_U58
g23705 nand P3_SUB_504_U8 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_504_U59
g23706 nand P3_SUB_504_U26 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_504_U60
g23707 not P3_SUB_504_U23 ; P3_SUB_504_U61
g23708 nand P3_SUB_504_U61 P3_SUB_504_U28 ; P3_SUB_504_U62
g23709 nand P3_SUB_504_U23 P3_SUB_504_U7 ; P3_SUB_504_U63
g23710 nand P3_SUB_401_U45 P3_SUB_401_U44 ; P3_SUB_401_U6
g23711 nand P3_SUB_401_U9 P3_SUB_401_U46 ; P3_SUB_401_U7
g23712 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_401_U8
g23713 nand P3_SUB_401_U18 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_401_U9
g23714 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_401_U10
g23715 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_401_U11
g23716 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_401_U12
g23717 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_401_U13
g23718 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_401_U14
g23719 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_401_U15
g23720 nand P3_SUB_401_U41 P3_SUB_401_U40 ; P3_SUB_401_U16
g23721 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_401_U17
g23722 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_401_U18
g23723 nand P3_SUB_401_U51 P3_SUB_401_U50 ; P3_SUB_401_U19
g23724 nand P3_SUB_401_U56 P3_SUB_401_U55 ; P3_SUB_401_U20
g23725 nand P3_SUB_401_U61 P3_SUB_401_U60 ; P3_SUB_401_U21
g23726 nand P3_SUB_401_U66 P3_SUB_401_U65 ; P3_SUB_401_U22
g23727 nand P3_SUB_401_U48 P3_SUB_401_U47 ; P3_SUB_401_U23
g23728 nand P3_SUB_401_U53 P3_SUB_401_U52 ; P3_SUB_401_U24
g23729 nand P3_SUB_401_U58 P3_SUB_401_U57 ; P3_SUB_401_U25
g23730 nand P3_SUB_401_U63 P3_SUB_401_U62 ; P3_SUB_401_U26
g23731 nand P3_SUB_401_U37 P3_SUB_401_U36 ; P3_SUB_401_U27
g23732 nand P3_SUB_401_U33 P3_SUB_401_U32 ; P3_SUB_401_U28
g23733 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_401_U29
g23734 not P3_SUB_401_U9 ; P3_SUB_401_U30
g23735 nand P3_SUB_401_U30 P3_SUB_401_U10 ; P3_SUB_401_U31
g23736 nand P3_SUB_401_U31 P3_SUB_401_U29 ; P3_SUB_401_U32
g23737 nand P3_SUB_401_U9 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_401_U33
g23738 not P3_SUB_401_U28 ; P3_SUB_401_U34
g23739 nand P3_SUB_401_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_401_U35
g23740 nand P3_SUB_401_U35 P3_SUB_401_U28 ; P3_SUB_401_U36
g23741 nand P3_SUB_401_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_401_U37
g23742 not P3_SUB_401_U27 ; P3_SUB_401_U38
g23743 nand P3_SUB_401_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_401_U39
g23744 nand P3_SUB_401_U39 P3_SUB_401_U27 ; P3_SUB_401_U40
g23745 nand P3_SUB_401_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_401_U41
g23746 not P3_SUB_401_U16 ; P3_SUB_401_U42
g23747 nand P3_SUB_401_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_401_U43
g23748 nand P3_SUB_401_U42 P3_SUB_401_U43 ; P3_SUB_401_U44
g23749 nand P3_SUB_401_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_401_U45
g23750 nand P3_SUB_401_U8 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_401_U46
g23751 nand P3_SUB_401_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_401_U47
g23752 nand P3_SUB_401_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_401_U48
g23753 not P3_SUB_401_U23 ; P3_SUB_401_U49
g23754 nand P3_SUB_401_U49 P3_SUB_401_U42 ; P3_SUB_401_U50
g23755 nand P3_SUB_401_U23 P3_SUB_401_U16 ; P3_SUB_401_U51
g23756 nand P3_SUB_401_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_401_U52
g23757 nand P3_SUB_401_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_401_U53
g23758 not P3_SUB_401_U24 ; P3_SUB_401_U54
g23759 nand P3_SUB_401_U38 P3_SUB_401_U54 ; P3_SUB_401_U55
g23760 nand P3_SUB_401_U24 P3_SUB_401_U27 ; P3_SUB_401_U56
g23761 nand P3_SUB_401_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_401_U57
g23762 nand P3_SUB_401_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_401_U58
g23763 not P3_SUB_401_U25 ; P3_SUB_401_U59
g23764 nand P3_SUB_401_U34 P3_SUB_401_U59 ; P3_SUB_401_U60
g23765 nand P3_SUB_401_U25 P3_SUB_401_U28 ; P3_SUB_401_U61
g23766 nand P3_SUB_401_U10 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_401_U62
g23767 nand P3_SUB_401_U29 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_401_U63
g23768 not P3_SUB_401_U26 ; P3_SUB_401_U64
g23769 nand P3_SUB_401_U64 P3_SUB_401_U30 ; P3_SUB_401_U65
g23770 nand P3_SUB_401_U26 P3_SUB_401_U9 ; P3_SUB_401_U66
g23771 not P3_U2621 ; P3_ADD_371_U4
g23772 nand P3_ADD_371_U24 P3_ADD_371_U32 ; P3_ADD_371_U5
g23773 and P3_ADD_371_U22 P3_ADD_371_U30 ; P3_ADD_371_U6
g23774 not P3_U2622 ; P3_ADD_371_U7
g23775 not P3_U2624 ; P3_ADD_371_U8
g23776 nand P3_U2624 P3_ADD_371_U24 ; P3_ADD_371_U9
g23777 not P3_U2625 ; P3_ADD_371_U10
g23778 nand P3_U2625 P3_ADD_371_U28 ; P3_ADD_371_U11
g23779 not P3_U2626 ; P3_ADD_371_U12
g23780 nand P3_U2626 P3_ADD_371_U29 ; P3_ADD_371_U13
g23781 not P3_U2628 ; P3_ADD_371_U14
g23782 not P3_U2627 ; P3_ADD_371_U15
g23783 not P3_U2623 ; P3_ADD_371_U16
g23784 nand P3_ADD_371_U34 P3_ADD_371_U33 ; P3_ADD_371_U17
g23785 nand P3_ADD_371_U36 P3_ADD_371_U35 ; P3_ADD_371_U18
g23786 nand P3_ADD_371_U38 P3_ADD_371_U37 ; P3_ADD_371_U19
g23787 nand P3_ADD_371_U40 P3_ADD_371_U39 ; P3_ADD_371_U20
g23788 nand P3_ADD_371_U44 P3_ADD_371_U43 ; P3_ADD_371_U21
g23789 and P3_U2628 P3_U2627 ; P3_ADD_371_U22
g23790 nand P3_U2627 P3_ADD_371_U30 ; P3_ADD_371_U23
g23791 nand P3_ADD_371_U16 P3_ADD_371_U26 ; P3_ADD_371_U24
g23792 and P3_ADD_371_U42 P3_ADD_371_U41 ; P3_ADD_371_U25
g23793 nand P3_U2622 P3_U2621 ; P3_ADD_371_U26
g23794 not P3_ADD_371_U24 ; P3_ADD_371_U27
g23795 not P3_ADD_371_U9 ; P3_ADD_371_U28
g23796 not P3_ADD_371_U11 ; P3_ADD_371_U29
g23797 not P3_ADD_371_U13 ; P3_ADD_371_U30
g23798 not P3_ADD_371_U23 ; P3_ADD_371_U31
g23799 nand P3_U2622 P3_U2621 P3_U2623 ; P3_ADD_371_U32
g23800 nand P3_U2628 P3_ADD_371_U23 ; P3_ADD_371_U33
g23801 nand P3_ADD_371_U31 P3_ADD_371_U14 ; P3_ADD_371_U34
g23802 nand P3_U2627 P3_ADD_371_U13 ; P3_ADD_371_U35
g23803 nand P3_ADD_371_U30 P3_ADD_371_U15 ; P3_ADD_371_U36
g23804 nand P3_U2626 P3_ADD_371_U11 ; P3_ADD_371_U37
g23805 nand P3_ADD_371_U29 P3_ADD_371_U12 ; P3_ADD_371_U38
g23806 nand P3_U2625 P3_ADD_371_U9 ; P3_ADD_371_U39
g23807 nand P3_ADD_371_U28 P3_ADD_371_U10 ; P3_ADD_371_U40
g23808 nand P3_U2624 P3_ADD_371_U24 ; P3_ADD_371_U41
g23809 nand P3_ADD_371_U27 P3_ADD_371_U8 ; P3_ADD_371_U42
g23810 nand P3_U2622 P3_ADD_371_U4 ; P3_ADD_371_U43
g23811 nand P3_U2621 P3_ADD_371_U7 ; P3_ADD_371_U44
g23812 nand P3_SUB_390_U45 P3_SUB_390_U44 ; P3_SUB_390_U6
g23813 nand P3_SUB_390_U9 P3_SUB_390_U46 ; P3_SUB_390_U7
g23814 not P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_390_U8
g23815 nand P3_SUB_390_U18 P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P3_SUB_390_U9
g23816 not P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_390_U10
g23817 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_390_U11
g23818 not P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_390_U12
g23819 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_390_U13
g23820 not P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_390_U14
g23821 not P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_390_U15
g23822 nand P3_SUB_390_U41 P3_SUB_390_U40 ; P3_SUB_390_U16
g23823 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_390_U17
g23824 not P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_390_U18
g23825 nand P3_SUB_390_U51 P3_SUB_390_U50 ; P3_SUB_390_U19
g23826 nand P3_SUB_390_U56 P3_SUB_390_U55 ; P3_SUB_390_U20
g23827 nand P3_SUB_390_U61 P3_SUB_390_U60 ; P3_SUB_390_U21
g23828 nand P3_SUB_390_U66 P3_SUB_390_U65 ; P3_SUB_390_U22
g23829 nand P3_SUB_390_U48 P3_SUB_390_U47 ; P3_SUB_390_U23
g23830 nand P3_SUB_390_U53 P3_SUB_390_U52 ; P3_SUB_390_U24
g23831 nand P3_SUB_390_U58 P3_SUB_390_U57 ; P3_SUB_390_U25
g23832 nand P3_SUB_390_U63 P3_SUB_390_U62 ; P3_SUB_390_U26
g23833 nand P3_SUB_390_U37 P3_SUB_390_U36 ; P3_SUB_390_U27
g23834 nand P3_SUB_390_U33 P3_SUB_390_U32 ; P3_SUB_390_U28
g23835 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_390_U29
g23836 not P3_SUB_390_U9 ; P3_SUB_390_U30
g23837 nand P3_SUB_390_U30 P3_SUB_390_U10 ; P3_SUB_390_U31
g23838 nand P3_SUB_390_U31 P3_SUB_390_U29 ; P3_SUB_390_U32
g23839 nand P3_SUB_390_U9 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_390_U33
g23840 not P3_SUB_390_U28 ; P3_SUB_390_U34
g23841 nand P3_SUB_390_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_390_U35
g23842 nand P3_SUB_390_U35 P3_SUB_390_U28 ; P3_SUB_390_U36
g23843 nand P3_SUB_390_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_390_U37
g23844 not P3_SUB_390_U27 ; P3_SUB_390_U38
g23845 nand P3_SUB_390_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_390_U39
g23846 nand P3_SUB_390_U39 P3_SUB_390_U27 ; P3_SUB_390_U40
g23847 nand P3_SUB_390_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_390_U41
g23848 not P3_SUB_390_U16 ; P3_SUB_390_U42
g23849 nand P3_SUB_390_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_390_U43
g23850 nand P3_SUB_390_U42 P3_SUB_390_U43 ; P3_SUB_390_U44
g23851 nand P3_SUB_390_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_390_U45
g23852 nand P3_SUB_390_U8 P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P3_SUB_390_U46
g23853 nand P3_SUB_390_U15 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_SUB_390_U47
g23854 nand P3_SUB_390_U17 P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P3_SUB_390_U48
g23855 not P3_SUB_390_U23 ; P3_SUB_390_U49
g23856 nand P3_SUB_390_U49 P3_SUB_390_U42 ; P3_SUB_390_U50
g23857 nand P3_SUB_390_U23 P3_SUB_390_U16 ; P3_SUB_390_U51
g23858 nand P3_SUB_390_U14 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_SUB_390_U52
g23859 nand P3_SUB_390_U13 P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P3_SUB_390_U53
g23860 not P3_SUB_390_U24 ; P3_SUB_390_U54
g23861 nand P3_SUB_390_U38 P3_SUB_390_U54 ; P3_SUB_390_U55
g23862 nand P3_SUB_390_U24 P3_SUB_390_U27 ; P3_SUB_390_U56
g23863 nand P3_SUB_390_U12 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_SUB_390_U57
g23864 nand P3_SUB_390_U11 P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P3_SUB_390_U58
g23865 not P3_SUB_390_U25 ; P3_SUB_390_U59
g23866 nand P3_SUB_390_U34 P3_SUB_390_U59 ; P3_SUB_390_U60
g23867 nand P3_SUB_390_U25 P3_SUB_390_U28 ; P3_SUB_390_U61
g23868 nand P3_SUB_390_U10 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_SUB_390_U62
g23869 nand P3_SUB_390_U29 P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P3_SUB_390_U63
g23870 not P3_SUB_390_U26 ; P3_SUB_390_U64
g23871 nand P3_SUB_390_U64 P3_SUB_390_U30 ; P3_SUB_390_U65
g23872 nand P3_SUB_390_U26 P3_SUB_390_U9 ; P3_SUB_390_U66
g23873 not P3_U2627 ; P3_SUB_357_U6
g23874 not P3_U2622 ; P3_SUB_357_U7
g23875 not P3_U2628 ; P3_SUB_357_U8
g23876 not P3_U2626 ; P3_SUB_357_U9
g23877 not P3_U2621 ; P3_SUB_357_U10
g23878 not P3_U2624 ; P3_SUB_357_U11
g23879 not P3_U2623 ; P3_SUB_357_U12
g23880 not P3_U2625 ; P3_SUB_357_U13
g23881 not P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_495_U4
g23882 not P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_495_U5
g23883 nand P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_495_U6
g23884 not P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_495_U7
g23885 nand P3_ADD_495_U16 P3_ADD_495_U15 ; P3_ADD_495_U8
g23886 nand P3_ADD_495_U18 P3_ADD_495_U17 ; P3_ADD_495_U9
g23887 nand P3_ADD_495_U20 P3_ADD_495_U19 ; P3_ADD_495_U10
g23888 not P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_495_U11
g23889 nand P3_ADD_495_U13 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_495_U12
g23890 not P3_ADD_495_U6 ; P3_ADD_495_U13
g23891 not P3_ADD_495_U12 ; P3_ADD_495_U14
g23892 nand P3_ADD_495_U12 P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P3_ADD_495_U15
g23893 nand P3_ADD_495_U14 P3_ADD_495_U11 ; P3_ADD_495_U16
g23894 nand P3_ADD_495_U6 P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P3_ADD_495_U17
g23895 nand P3_ADD_495_U13 P3_ADD_495_U7 ; P3_ADD_495_U18
g23896 nand P3_ADD_495_U4 P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P3_ADD_495_U19
g23897 nand P3_ADD_495_U5 P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P3_ADD_495_U20
g23898 nor P3_SUB_412_U6 P3_GTE_412_U7 ; P3_GTE_412_U6
g23899 nor P3_SUB_412_U16 P3_SUB_412_U17 P3_SUB_412_U19 P3_SUB_412_U18 ; P3_GTE_412_U7
g23900 nor P3_SUB_504_U6 P3_GTE_504_U7 ; P3_GTE_504_U6
g23901 nor P3_SUB_504_U16 P3_SUB_504_U17 P3_SUB_504_U19 P3_SUB_504_U18 ; P3_GTE_504_U7
g23902 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_494_U4
g23903 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_494_U5
g23904 nand P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_494_U6
g23905 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_494_U7
g23906 nand P3_ADD_494_U94 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_494_U8
g23907 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_494_U9
g23908 nand P3_ADD_494_U95 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_494_U10
g23909 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_494_U11
g23910 nand P3_ADD_494_U96 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_494_U12
g23911 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_494_U13
g23912 nand P3_ADD_494_U97 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_494_U14
g23913 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_494_U15
g23914 nand P3_ADD_494_U98 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_494_U16
g23915 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_494_U17
g23916 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_494_U18
g23917 nand P3_ADD_494_U99 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_494_U19
g23918 nand P3_ADD_494_U100 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_494_U20
g23919 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_494_U21
g23920 nand P3_ADD_494_U101 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_494_U22
g23921 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_494_U23
g23922 nand P3_ADD_494_U102 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_494_U24
g23923 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_494_U25
g23924 nand P3_ADD_494_U103 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_494_U26
g23925 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_494_U27
g23926 nand P3_ADD_494_U104 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_494_U28
g23927 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_494_U29
g23928 nand P3_ADD_494_U105 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_494_U30
g23929 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_494_U31
g23930 nand P3_ADD_494_U106 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_494_U32
g23931 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_494_U33
g23932 nand P3_ADD_494_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_494_U34
g23933 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_494_U35
g23934 nand P3_ADD_494_U108 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_494_U36
g23935 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_494_U37
g23936 nand P3_ADD_494_U109 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_494_U38
g23937 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_494_U39
g23938 nand P3_ADD_494_U110 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_494_U40
g23939 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_494_U41
g23940 nand P3_ADD_494_U111 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_494_U42
g23941 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_494_U43
g23942 nand P3_ADD_494_U112 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_494_U44
g23943 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_494_U45
g23944 nand P3_ADD_494_U113 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_494_U46
g23945 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_494_U47
g23946 nand P3_ADD_494_U114 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_494_U48
g23947 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_494_U49
g23948 nand P3_ADD_494_U115 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_494_U50
g23949 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_494_U51
g23950 nand P3_ADD_494_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_494_U52
g23951 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_494_U53
g23952 nand P3_ADD_494_U117 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_494_U54
g23953 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_494_U55
g23954 nand P3_ADD_494_U118 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_494_U56
g23955 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_494_U57
g23956 nand P3_ADD_494_U119 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_494_U58
g23957 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_494_U59
g23958 nand P3_ADD_494_U120 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_494_U60
g23959 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_494_U61
g23960 nand P3_ADD_494_U124 P3_ADD_494_U123 ; P3_ADD_494_U62
g23961 nand P3_ADD_494_U126 P3_ADD_494_U125 ; P3_ADD_494_U63
g23962 nand P3_ADD_494_U128 P3_ADD_494_U127 ; P3_ADD_494_U64
g23963 nand P3_ADD_494_U130 P3_ADD_494_U129 ; P3_ADD_494_U65
g23964 nand P3_ADD_494_U132 P3_ADD_494_U131 ; P3_ADD_494_U66
g23965 nand P3_ADD_494_U134 P3_ADD_494_U133 ; P3_ADD_494_U67
g23966 nand P3_ADD_494_U136 P3_ADD_494_U135 ; P3_ADD_494_U68
g23967 nand P3_ADD_494_U138 P3_ADD_494_U137 ; P3_ADD_494_U69
g23968 nand P3_ADD_494_U140 P3_ADD_494_U139 ; P3_ADD_494_U70
g23969 nand P3_ADD_494_U142 P3_ADD_494_U141 ; P3_ADD_494_U71
g23970 nand P3_ADD_494_U144 P3_ADD_494_U143 ; P3_ADD_494_U72
g23971 nand P3_ADD_494_U146 P3_ADD_494_U145 ; P3_ADD_494_U73
g23972 nand P3_ADD_494_U148 P3_ADD_494_U147 ; P3_ADD_494_U74
g23973 nand P3_ADD_494_U150 P3_ADD_494_U149 ; P3_ADD_494_U75
g23974 nand P3_ADD_494_U152 P3_ADD_494_U151 ; P3_ADD_494_U76
g23975 nand P3_ADD_494_U154 P3_ADD_494_U153 ; P3_ADD_494_U77
g23976 nand P3_ADD_494_U156 P3_ADD_494_U155 ; P3_ADD_494_U78
g23977 nand P3_ADD_494_U158 P3_ADD_494_U157 ; P3_ADD_494_U79
g23978 nand P3_ADD_494_U160 P3_ADD_494_U159 ; P3_ADD_494_U80
g23979 nand P3_ADD_494_U162 P3_ADD_494_U161 ; P3_ADD_494_U81
g23980 nand P3_ADD_494_U164 P3_ADD_494_U163 ; P3_ADD_494_U82
g23981 nand P3_ADD_494_U166 P3_ADD_494_U165 ; P3_ADD_494_U83
g23982 nand P3_ADD_494_U168 P3_ADD_494_U167 ; P3_ADD_494_U84
g23983 nand P3_ADD_494_U170 P3_ADD_494_U169 ; P3_ADD_494_U85
g23984 nand P3_ADD_494_U172 P3_ADD_494_U171 ; P3_ADD_494_U86
g23985 nand P3_ADD_494_U174 P3_ADD_494_U173 ; P3_ADD_494_U87
g23986 nand P3_ADD_494_U176 P3_ADD_494_U175 ; P3_ADD_494_U88
g23987 nand P3_ADD_494_U178 P3_ADD_494_U177 ; P3_ADD_494_U89
g23988 nand P3_ADD_494_U180 P3_ADD_494_U179 ; P3_ADD_494_U90
g23989 nand P3_ADD_494_U182 P3_ADD_494_U181 ; P3_ADD_494_U91
g23990 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_494_U92
g23991 nand P3_ADD_494_U121 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_494_U93
g23992 not P3_ADD_494_U6 ; P3_ADD_494_U94
g23993 not P3_ADD_494_U8 ; P3_ADD_494_U95
g23994 not P3_ADD_494_U10 ; P3_ADD_494_U96
g23995 not P3_ADD_494_U12 ; P3_ADD_494_U97
g23996 not P3_ADD_494_U14 ; P3_ADD_494_U98
g23997 not P3_ADD_494_U16 ; P3_ADD_494_U99
g23998 not P3_ADD_494_U19 ; P3_ADD_494_U100
g23999 not P3_ADD_494_U20 ; P3_ADD_494_U101
g24000 not P3_ADD_494_U22 ; P3_ADD_494_U102
g24001 not P3_ADD_494_U24 ; P3_ADD_494_U103
g24002 not P3_ADD_494_U26 ; P3_ADD_494_U104
g24003 not P3_ADD_494_U28 ; P3_ADD_494_U105
g24004 not P3_ADD_494_U30 ; P3_ADD_494_U106
g24005 not P3_ADD_494_U32 ; P3_ADD_494_U107
g24006 not P3_ADD_494_U34 ; P3_ADD_494_U108
g24007 not P3_ADD_494_U36 ; P3_ADD_494_U109
g24008 not P3_ADD_494_U38 ; P3_ADD_494_U110
g24009 not P3_ADD_494_U40 ; P3_ADD_494_U111
g24010 not P3_ADD_494_U42 ; P3_ADD_494_U112
g24011 not P3_ADD_494_U44 ; P3_ADD_494_U113
g24012 not P3_ADD_494_U46 ; P3_ADD_494_U114
g24013 not P3_ADD_494_U48 ; P3_ADD_494_U115
g24014 not P3_ADD_494_U50 ; P3_ADD_494_U116
g24015 not P3_ADD_494_U52 ; P3_ADD_494_U117
g24016 not P3_ADD_494_U54 ; P3_ADD_494_U118
g24017 not P3_ADD_494_U56 ; P3_ADD_494_U119
g24018 not P3_ADD_494_U58 ; P3_ADD_494_U120
g24019 not P3_ADD_494_U60 ; P3_ADD_494_U121
g24020 not P3_ADD_494_U93 ; P3_ADD_494_U122
g24021 nand P3_ADD_494_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_494_U123
g24022 nand P3_ADD_494_U100 P3_ADD_494_U18 ; P3_ADD_494_U124
g24023 nand P3_ADD_494_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_494_U125
g24024 nand P3_ADD_494_U99 P3_ADD_494_U17 ; P3_ADD_494_U126
g24025 nand P3_ADD_494_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_494_U127
g24026 nand P3_ADD_494_U98 P3_ADD_494_U15 ; P3_ADD_494_U128
g24027 nand P3_ADD_494_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_494_U129
g24028 nand P3_ADD_494_U97 P3_ADD_494_U13 ; P3_ADD_494_U130
g24029 nand P3_ADD_494_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_494_U131
g24030 nand P3_ADD_494_U96 P3_ADD_494_U11 ; P3_ADD_494_U132
g24031 nand P3_ADD_494_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_494_U133
g24032 nand P3_ADD_494_U95 P3_ADD_494_U9 ; P3_ADD_494_U134
g24033 nand P3_ADD_494_U6 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_494_U135
g24034 nand P3_ADD_494_U94 P3_ADD_494_U7 ; P3_ADD_494_U136
g24035 nand P3_ADD_494_U93 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_494_U137
g24036 nand P3_ADD_494_U122 P3_ADD_494_U92 ; P3_ADD_494_U138
g24037 nand P3_ADD_494_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_494_U139
g24038 nand P3_ADD_494_U121 P3_ADD_494_U61 ; P3_ADD_494_U140
g24039 nand P3_ADD_494_U4 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_494_U141
g24040 nand P3_ADD_494_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_494_U142
g24041 nand P3_ADD_494_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_494_U143
g24042 nand P3_ADD_494_U120 P3_ADD_494_U59 ; P3_ADD_494_U144
g24043 nand P3_ADD_494_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_494_U145
g24044 nand P3_ADD_494_U119 P3_ADD_494_U57 ; P3_ADD_494_U146
g24045 nand P3_ADD_494_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_494_U147
g24046 nand P3_ADD_494_U118 P3_ADD_494_U55 ; P3_ADD_494_U148
g24047 nand P3_ADD_494_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_494_U149
g24048 nand P3_ADD_494_U117 P3_ADD_494_U53 ; P3_ADD_494_U150
g24049 nand P3_ADD_494_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_494_U151
g24050 nand P3_ADD_494_U116 P3_ADD_494_U51 ; P3_ADD_494_U152
g24051 nand P3_ADD_494_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_494_U153
g24052 nand P3_ADD_494_U115 P3_ADD_494_U49 ; P3_ADD_494_U154
g24053 nand P3_ADD_494_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_494_U155
g24054 nand P3_ADD_494_U114 P3_ADD_494_U47 ; P3_ADD_494_U156
g24055 nand P3_ADD_494_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_494_U157
g24056 nand P3_ADD_494_U113 P3_ADD_494_U45 ; P3_ADD_494_U158
g24057 nand P3_ADD_494_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_494_U159
g24058 nand P3_ADD_494_U112 P3_ADD_494_U43 ; P3_ADD_494_U160
g24059 nand P3_ADD_494_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_494_U161
g24060 nand P3_ADD_494_U111 P3_ADD_494_U41 ; P3_ADD_494_U162
g24061 nand P3_ADD_494_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_494_U163
g24062 nand P3_ADD_494_U110 P3_ADD_494_U39 ; P3_ADD_494_U164
g24063 nand P3_ADD_494_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_494_U165
g24064 nand P3_ADD_494_U109 P3_ADD_494_U37 ; P3_ADD_494_U166
g24065 nand P3_ADD_494_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_494_U167
g24066 nand P3_ADD_494_U108 P3_ADD_494_U35 ; P3_ADD_494_U168
g24067 nand P3_ADD_494_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_494_U169
g24068 nand P3_ADD_494_U107 P3_ADD_494_U33 ; P3_ADD_494_U170
g24069 nand P3_ADD_494_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_494_U171
g24070 nand P3_ADD_494_U106 P3_ADD_494_U31 ; P3_ADD_494_U172
g24071 nand P3_ADD_494_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_494_U173
g24072 nand P3_ADD_494_U105 P3_ADD_494_U29 ; P3_ADD_494_U174
g24073 nand P3_ADD_494_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_494_U175
g24074 nand P3_ADD_494_U104 P3_ADD_494_U27 ; P3_ADD_494_U176
g24075 nand P3_ADD_494_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_494_U177
g24076 nand P3_ADD_494_U103 P3_ADD_494_U25 ; P3_ADD_494_U178
g24077 nand P3_ADD_494_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_494_U179
g24078 nand P3_ADD_494_U102 P3_ADD_494_U23 ; P3_ADD_494_U180
g24079 nand P3_ADD_494_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_494_U181
g24080 nand P3_ADD_494_U101 P3_ADD_494_U21 ; P3_ADD_494_U182
g24081 not P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_536_U4
g24082 not P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_536_U5
g24083 nand P3_INSTADDRPOINTER_REG_1__SCAN_IN P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_536_U6
g24084 not P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_536_U7
g24085 nand P3_ADD_536_U94 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_536_U8
g24086 not P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_536_U9
g24087 nand P3_ADD_536_U95 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_536_U10
g24088 not P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_536_U11
g24089 nand P3_ADD_536_U96 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_536_U12
g24090 not P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_536_U13
g24091 nand P3_ADD_536_U97 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_536_U14
g24092 not P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_536_U15
g24093 nand P3_ADD_536_U98 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_536_U16
g24094 not P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_536_U17
g24095 not P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_536_U18
g24096 nand P3_ADD_536_U99 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_536_U19
g24097 nand P3_ADD_536_U100 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_536_U20
g24098 not P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_536_U21
g24099 nand P3_ADD_536_U101 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_536_U22
g24100 not P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_536_U23
g24101 nand P3_ADD_536_U102 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_536_U24
g24102 not P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_536_U25
g24103 nand P3_ADD_536_U103 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_536_U26
g24104 not P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_536_U27
g24105 nand P3_ADD_536_U104 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_536_U28
g24106 not P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_536_U29
g24107 nand P3_ADD_536_U105 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_536_U30
g24108 not P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_536_U31
g24109 nand P3_ADD_536_U106 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_536_U32
g24110 not P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_536_U33
g24111 nand P3_ADD_536_U107 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_536_U34
g24112 not P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_536_U35
g24113 nand P3_ADD_536_U108 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_536_U36
g24114 not P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_536_U37
g24115 nand P3_ADD_536_U109 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_536_U38
g24116 not P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_536_U39
g24117 nand P3_ADD_536_U110 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_536_U40
g24118 not P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_536_U41
g24119 nand P3_ADD_536_U111 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_536_U42
g24120 not P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_536_U43
g24121 nand P3_ADD_536_U112 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_536_U44
g24122 not P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_536_U45
g24123 nand P3_ADD_536_U113 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_536_U46
g24124 not P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_536_U47
g24125 nand P3_ADD_536_U114 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_536_U48
g24126 not P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_536_U49
g24127 nand P3_ADD_536_U115 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_536_U50
g24128 not P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_536_U51
g24129 nand P3_ADD_536_U116 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_536_U52
g24130 not P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_536_U53
g24131 nand P3_ADD_536_U117 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_536_U54
g24132 not P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_536_U55
g24133 nand P3_ADD_536_U118 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_536_U56
g24134 not P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_536_U57
g24135 nand P3_ADD_536_U119 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_536_U58
g24136 not P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_536_U59
g24137 nand P3_ADD_536_U120 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_536_U60
g24138 not P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_536_U61
g24139 nand P3_ADD_536_U124 P3_ADD_536_U123 ; P3_ADD_536_U62
g24140 nand P3_ADD_536_U126 P3_ADD_536_U125 ; P3_ADD_536_U63
g24141 nand P3_ADD_536_U128 P3_ADD_536_U127 ; P3_ADD_536_U64
g24142 nand P3_ADD_536_U130 P3_ADD_536_U129 ; P3_ADD_536_U65
g24143 nand P3_ADD_536_U132 P3_ADD_536_U131 ; P3_ADD_536_U66
g24144 nand P3_ADD_536_U134 P3_ADD_536_U133 ; P3_ADD_536_U67
g24145 nand P3_ADD_536_U136 P3_ADD_536_U135 ; P3_ADD_536_U68
g24146 nand P3_ADD_536_U138 P3_ADD_536_U137 ; P3_ADD_536_U69
g24147 nand P3_ADD_536_U140 P3_ADD_536_U139 ; P3_ADD_536_U70
g24148 nand P3_ADD_536_U142 P3_ADD_536_U141 ; P3_ADD_536_U71
g24149 nand P3_ADD_536_U144 P3_ADD_536_U143 ; P3_ADD_536_U72
g24150 nand P3_ADD_536_U146 P3_ADD_536_U145 ; P3_ADD_536_U73
g24151 nand P3_ADD_536_U148 P3_ADD_536_U147 ; P3_ADD_536_U74
g24152 nand P3_ADD_536_U150 P3_ADD_536_U149 ; P3_ADD_536_U75
g24153 nand P3_ADD_536_U152 P3_ADD_536_U151 ; P3_ADD_536_U76
g24154 nand P3_ADD_536_U154 P3_ADD_536_U153 ; P3_ADD_536_U77
g24155 nand P3_ADD_536_U156 P3_ADD_536_U155 ; P3_ADD_536_U78
g24156 nand P3_ADD_536_U158 P3_ADD_536_U157 ; P3_ADD_536_U79
g24157 nand P3_ADD_536_U160 P3_ADD_536_U159 ; P3_ADD_536_U80
g24158 nand P3_ADD_536_U162 P3_ADD_536_U161 ; P3_ADD_536_U81
g24159 nand P3_ADD_536_U164 P3_ADD_536_U163 ; P3_ADD_536_U82
g24160 nand P3_ADD_536_U166 P3_ADD_536_U165 ; P3_ADD_536_U83
g24161 nand P3_ADD_536_U168 P3_ADD_536_U167 ; P3_ADD_536_U84
g24162 nand P3_ADD_536_U170 P3_ADD_536_U169 ; P3_ADD_536_U85
g24163 nand P3_ADD_536_U172 P3_ADD_536_U171 ; P3_ADD_536_U86
g24164 nand P3_ADD_536_U174 P3_ADD_536_U173 ; P3_ADD_536_U87
g24165 nand P3_ADD_536_U176 P3_ADD_536_U175 ; P3_ADD_536_U88
g24166 nand P3_ADD_536_U178 P3_ADD_536_U177 ; P3_ADD_536_U89
g24167 nand P3_ADD_536_U180 P3_ADD_536_U179 ; P3_ADD_536_U90
g24168 nand P3_ADD_536_U182 P3_ADD_536_U181 ; P3_ADD_536_U91
g24169 not P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_536_U92
g24170 nand P3_ADD_536_U121 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_536_U93
g24171 not P3_ADD_536_U6 ; P3_ADD_536_U94
g24172 not P3_ADD_536_U8 ; P3_ADD_536_U95
g24173 not P3_ADD_536_U10 ; P3_ADD_536_U96
g24174 not P3_ADD_536_U12 ; P3_ADD_536_U97
g24175 not P3_ADD_536_U14 ; P3_ADD_536_U98
g24176 not P3_ADD_536_U16 ; P3_ADD_536_U99
g24177 not P3_ADD_536_U19 ; P3_ADD_536_U100
g24178 not P3_ADD_536_U20 ; P3_ADD_536_U101
g24179 not P3_ADD_536_U22 ; P3_ADD_536_U102
g24180 not P3_ADD_536_U24 ; P3_ADD_536_U103
g24181 not P3_ADD_536_U26 ; P3_ADD_536_U104
g24182 not P3_ADD_536_U28 ; P3_ADD_536_U105
g24183 not P3_ADD_536_U30 ; P3_ADD_536_U106
g24184 not P3_ADD_536_U32 ; P3_ADD_536_U107
g24185 not P3_ADD_536_U34 ; P3_ADD_536_U108
g24186 not P3_ADD_536_U36 ; P3_ADD_536_U109
g24187 not P3_ADD_536_U38 ; P3_ADD_536_U110
g24188 not P3_ADD_536_U40 ; P3_ADD_536_U111
g24189 not P3_ADD_536_U42 ; P3_ADD_536_U112
g24190 not P3_ADD_536_U44 ; P3_ADD_536_U113
g24191 not P3_ADD_536_U46 ; P3_ADD_536_U114
g24192 not P3_ADD_536_U48 ; P3_ADD_536_U115
g24193 not P3_ADD_536_U50 ; P3_ADD_536_U116
g24194 not P3_ADD_536_U52 ; P3_ADD_536_U117
g24195 not P3_ADD_536_U54 ; P3_ADD_536_U118
g24196 not P3_ADD_536_U56 ; P3_ADD_536_U119
g24197 not P3_ADD_536_U58 ; P3_ADD_536_U120
g24198 not P3_ADD_536_U60 ; P3_ADD_536_U121
g24199 not P3_ADD_536_U93 ; P3_ADD_536_U122
g24200 nand P3_ADD_536_U19 P3_INSTADDRPOINTER_REG_9__SCAN_IN ; P3_ADD_536_U123
g24201 nand P3_ADD_536_U100 P3_ADD_536_U18 ; P3_ADD_536_U124
g24202 nand P3_ADD_536_U16 P3_INSTADDRPOINTER_REG_8__SCAN_IN ; P3_ADD_536_U125
g24203 nand P3_ADD_536_U99 P3_ADD_536_U17 ; P3_ADD_536_U126
g24204 nand P3_ADD_536_U14 P3_INSTADDRPOINTER_REG_7__SCAN_IN ; P3_ADD_536_U127
g24205 nand P3_ADD_536_U98 P3_ADD_536_U15 ; P3_ADD_536_U128
g24206 nand P3_ADD_536_U12 P3_INSTADDRPOINTER_REG_6__SCAN_IN ; P3_ADD_536_U129
g24207 nand P3_ADD_536_U97 P3_ADD_536_U13 ; P3_ADD_536_U130
g24208 nand P3_ADD_536_U10 P3_INSTADDRPOINTER_REG_5__SCAN_IN ; P3_ADD_536_U131
g24209 nand P3_ADD_536_U96 P3_ADD_536_U11 ; P3_ADD_536_U132
g24210 nand P3_ADD_536_U8 P3_INSTADDRPOINTER_REG_4__SCAN_IN ; P3_ADD_536_U133
g24211 nand P3_ADD_536_U95 P3_ADD_536_U9 ; P3_ADD_536_U134
g24212 nand P3_ADD_536_U6 P3_INSTADDRPOINTER_REG_3__SCAN_IN ; P3_ADD_536_U135
g24213 nand P3_ADD_536_U94 P3_ADD_536_U7 ; P3_ADD_536_U136
g24214 nand P3_ADD_536_U93 P3_INSTADDRPOINTER_REG_31__SCAN_IN ; P3_ADD_536_U137
g24215 nand P3_ADD_536_U122 P3_ADD_536_U92 ; P3_ADD_536_U138
g24216 nand P3_ADD_536_U60 P3_INSTADDRPOINTER_REG_30__SCAN_IN ; P3_ADD_536_U139
g24217 nand P3_ADD_536_U121 P3_ADD_536_U61 ; P3_ADD_536_U140
g24218 nand P3_ADD_536_U4 P3_INSTADDRPOINTER_REG_2__SCAN_IN ; P3_ADD_536_U141
g24219 nand P3_ADD_536_U5 P3_INSTADDRPOINTER_REG_1__SCAN_IN ; P3_ADD_536_U142
g24220 nand P3_ADD_536_U58 P3_INSTADDRPOINTER_REG_29__SCAN_IN ; P3_ADD_536_U143
g24221 nand P3_ADD_536_U120 P3_ADD_536_U59 ; P3_ADD_536_U144
g24222 nand P3_ADD_536_U56 P3_INSTADDRPOINTER_REG_28__SCAN_IN ; P3_ADD_536_U145
g24223 nand P3_ADD_536_U119 P3_ADD_536_U57 ; P3_ADD_536_U146
g24224 nand P3_ADD_536_U54 P3_INSTADDRPOINTER_REG_27__SCAN_IN ; P3_ADD_536_U147
g24225 nand P3_ADD_536_U118 P3_ADD_536_U55 ; P3_ADD_536_U148
g24226 nand P3_ADD_536_U52 P3_INSTADDRPOINTER_REG_26__SCAN_IN ; P3_ADD_536_U149
g24227 nand P3_ADD_536_U117 P3_ADD_536_U53 ; P3_ADD_536_U150
g24228 nand P3_ADD_536_U50 P3_INSTADDRPOINTER_REG_25__SCAN_IN ; P3_ADD_536_U151
g24229 nand P3_ADD_536_U116 P3_ADD_536_U51 ; P3_ADD_536_U152
g24230 nand P3_ADD_536_U48 P3_INSTADDRPOINTER_REG_24__SCAN_IN ; P3_ADD_536_U153
g24231 nand P3_ADD_536_U115 P3_ADD_536_U49 ; P3_ADD_536_U154
g24232 nand P3_ADD_536_U46 P3_INSTADDRPOINTER_REG_23__SCAN_IN ; P3_ADD_536_U155
g24233 nand P3_ADD_536_U114 P3_ADD_536_U47 ; P3_ADD_536_U156
g24234 nand P3_ADD_536_U44 P3_INSTADDRPOINTER_REG_22__SCAN_IN ; P3_ADD_536_U157
g24235 nand P3_ADD_536_U113 P3_ADD_536_U45 ; P3_ADD_536_U158
g24236 nand P3_ADD_536_U42 P3_INSTADDRPOINTER_REG_21__SCAN_IN ; P3_ADD_536_U159
g24237 nand P3_ADD_536_U112 P3_ADD_536_U43 ; P3_ADD_536_U160
g24238 nand P3_ADD_536_U40 P3_INSTADDRPOINTER_REG_20__SCAN_IN ; P3_ADD_536_U161
g24239 nand P3_ADD_536_U111 P3_ADD_536_U41 ; P3_ADD_536_U162
g24240 nand P3_ADD_536_U38 P3_INSTADDRPOINTER_REG_19__SCAN_IN ; P3_ADD_536_U163
g24241 nand P3_ADD_536_U110 P3_ADD_536_U39 ; P3_ADD_536_U164
g24242 nand P3_ADD_536_U36 P3_INSTADDRPOINTER_REG_18__SCAN_IN ; P3_ADD_536_U165
g24243 nand P3_ADD_536_U109 P3_ADD_536_U37 ; P3_ADD_536_U166
g24244 nand P3_ADD_536_U34 P3_INSTADDRPOINTER_REG_17__SCAN_IN ; P3_ADD_536_U167
g24245 nand P3_ADD_536_U108 P3_ADD_536_U35 ; P3_ADD_536_U168
g24246 nand P3_ADD_536_U32 P3_INSTADDRPOINTER_REG_16__SCAN_IN ; P3_ADD_536_U169
g24247 nand P3_ADD_536_U107 P3_ADD_536_U33 ; P3_ADD_536_U170
g24248 nand P3_ADD_536_U30 P3_INSTADDRPOINTER_REG_15__SCAN_IN ; P3_ADD_536_U171
g24249 nand P3_ADD_536_U106 P3_ADD_536_U31 ; P3_ADD_536_U172
g24250 nand P3_ADD_536_U28 P3_INSTADDRPOINTER_REG_14__SCAN_IN ; P3_ADD_536_U173
g24251 nand P3_ADD_536_U105 P3_ADD_536_U29 ; P3_ADD_536_U174
g24252 nand P3_ADD_536_U26 P3_INSTADDRPOINTER_REG_13__SCAN_IN ; P3_ADD_536_U175
g24253 nand P3_ADD_536_U104 P3_ADD_536_U27 ; P3_ADD_536_U176
g24254 nand P3_ADD_536_U24 P3_INSTADDRPOINTER_REG_12__SCAN_IN ; P3_ADD_536_U177
g24255 nand P3_ADD_536_U103 P3_ADD_536_U25 ; P3_ADD_536_U178
g24256 nand P3_ADD_536_U22 P3_INSTADDRPOINTER_REG_11__SCAN_IN ; P3_ADD_536_U179
g24257 nand P3_ADD_536_U102 P3_ADD_536_U23 ; P3_ADD_536_U180
g24258 nand P3_ADD_536_U20 P3_INSTADDRPOINTER_REG_10__SCAN_IN ; P3_ADD_536_U181
g24259 nand P3_ADD_536_U101 P3_ADD_536_U21 ; P3_ADD_536_U182
g24260 not P3_U2613 ; P3_ADD_402_1132_U4
g24261 not P3_U3069 ; P3_ADD_402_1132_U5
g24262 nand P3_U3069 P3_U2613 ; P3_ADD_402_1132_U6
g24263 not P3_U2614 ; P3_ADD_402_1132_U7
g24264 nand P3_U2614 P3_ADD_402_1132_U28 ; P3_ADD_402_1132_U8
g24265 not P3_U2615 ; P3_ADD_402_1132_U9
g24266 nand P3_U2615 P3_ADD_402_1132_U29 ; P3_ADD_402_1132_U10
g24267 not P3_U2616 ; P3_ADD_402_1132_U11
g24268 nand P3_U2616 P3_ADD_402_1132_U30 ; P3_ADD_402_1132_U12
g24269 not P3_U2617 ; P3_ADD_402_1132_U13
g24270 nand P3_U2617 P3_ADD_402_1132_U31 ; P3_ADD_402_1132_U14
g24271 not P3_U2618 ; P3_ADD_402_1132_U15
g24272 nand P3_U2618 P3_ADD_402_1132_U32 ; P3_ADD_402_1132_U16
g24273 not P3_U2619 ; P3_ADD_402_1132_U17
g24274 nand P3_ADD_402_1132_U36 P3_ADD_402_1132_U35 ; P3_ADD_402_1132_U18
g24275 nand P3_ADD_402_1132_U38 P3_ADD_402_1132_U37 ; P3_ADD_402_1132_U19
g24276 nand P3_ADD_402_1132_U40 P3_ADD_402_1132_U39 ; P3_ADD_402_1132_U20
g24277 nand P3_ADD_402_1132_U42 P3_ADD_402_1132_U41 ; P3_ADD_402_1132_U21
g24278 nand P3_ADD_402_1132_U44 P3_ADD_402_1132_U43 ; P3_ADD_402_1132_U22
g24279 nand P3_ADD_402_1132_U46 P3_ADD_402_1132_U45 ; P3_ADD_402_1132_U23
g24280 nand P3_ADD_402_1132_U48 P3_ADD_402_1132_U47 ; P3_ADD_402_1132_U24
g24281 nand P3_ADD_402_1132_U50 P3_ADD_402_1132_U49 ; P3_ADD_402_1132_U25
g24282 not P3_U2620 ; P3_ADD_402_1132_U26
g24283 nand P3_U2619 P3_ADD_402_1132_U33 ; P3_ADD_402_1132_U27
g24284 not P3_ADD_402_1132_U6 ; P3_ADD_402_1132_U28
g24285 not P3_ADD_402_1132_U8 ; P3_ADD_402_1132_U29
g24286 not P3_ADD_402_1132_U10 ; P3_ADD_402_1132_U30
g24287 not P3_ADD_402_1132_U12 ; P3_ADD_402_1132_U31
g24288 not P3_ADD_402_1132_U14 ; P3_ADD_402_1132_U32
g24289 not P3_ADD_402_1132_U16 ; P3_ADD_402_1132_U33
g24290 not P3_ADD_402_1132_U27 ; P3_ADD_402_1132_U34
g24291 nand P3_U2620 P3_ADD_402_1132_U27 ; P3_ADD_402_1132_U35
g24292 nand P3_ADD_402_1132_U34 P3_ADD_402_1132_U26 ; P3_ADD_402_1132_U36
g24293 nand P3_U2619 P3_ADD_402_1132_U16 ; P3_ADD_402_1132_U37
g24294 nand P3_ADD_402_1132_U33 P3_ADD_402_1132_U17 ; P3_ADD_402_1132_U38
g24295 nand P3_U2618 P3_ADD_402_1132_U14 ; P3_ADD_402_1132_U39
g24296 nand P3_ADD_402_1132_U32 P3_ADD_402_1132_U15 ; P3_ADD_402_1132_U40
g24297 nand P3_U2617 P3_ADD_402_1132_U12 ; P3_ADD_402_1132_U41
g24298 nand P3_ADD_402_1132_U31 P3_ADD_402_1132_U13 ; P3_ADD_402_1132_U42
g24299 nand P3_U2616 P3_ADD_402_1132_U10 ; P3_ADD_402_1132_U43
g24300 nand P3_ADD_402_1132_U30 P3_ADD_402_1132_U11 ; P3_ADD_402_1132_U44
g24301 nand P3_U2615 P3_ADD_402_1132_U8 ; P3_ADD_402_1132_U45
g24302 nand P3_ADD_402_1132_U29 P3_ADD_402_1132_U9 ; P3_ADD_402_1132_U46
g24303 nand P3_U2614 P3_ADD_402_1132_U6 ; P3_ADD_402_1132_U47
g24304 nand P3_ADD_402_1132_U28 P3_ADD_402_1132_U7 ; P3_ADD_402_1132_U48
g24305 nand P3_U3069 P3_ADD_402_1132_U4 ; P3_ADD_402_1132_U49
g24306 nand P3_U2613 P3_ADD_402_1132_U5 ; P3_ADD_402_1132_U50
g24307 nand P2_R2099_U107 P2_R2099_U148 ; P2_R2099_U5
g24308 not P2_U2747 ; P2_R2099_U6
g24309 not P2_U2751 ; P2_R2099_U7
g24310 not P2_U2750 ; P2_R2099_U8
g24311 not P2_U2746 ; P2_R2099_U9
g24312 not P2_U2749 ; P2_R2099_U10
g24313 not P2_U2745 ; P2_R2099_U11
g24314 not P2_U2748 ; P2_R2099_U12
g24315 not P2_U2744 ; P2_R2099_U13
g24316 not P2_U2743 ; P2_R2099_U14
g24317 nand P2_U2743 P2_R2099_U97 ; P2_R2099_U15
g24318 not P2_U2742 ; P2_R2099_U16
g24319 nand P2_U2742 P2_R2099_U120 ; P2_R2099_U17
g24320 not P2_U2741 ; P2_R2099_U18
g24321 nand P2_U2741 P2_R2099_U121 ; P2_R2099_U19
g24322 not P2_U2740 ; P2_R2099_U20
g24323 nand P2_U2740 P2_R2099_U122 ; P2_R2099_U21
g24324 not P2_U2739 ; P2_R2099_U22
g24325 not P2_U2738 ; P2_R2099_U23
g24326 nand P2_U2739 P2_R2099_U123 ; P2_R2099_U24
g24327 nand P2_R2099_U124 P2_U2738 ; P2_R2099_U25
g24328 not P2_U2737 ; P2_R2099_U26
g24329 nand P2_U2737 P2_R2099_U125 ; P2_R2099_U27
g24330 not P2_U2736 ; P2_R2099_U28
g24331 nand P2_U2736 P2_R2099_U126 ; P2_R2099_U29
g24332 not P2_U2735 ; P2_R2099_U30
g24333 nand P2_U2735 P2_R2099_U127 ; P2_R2099_U31
g24334 not P2_U2734 ; P2_R2099_U32
g24335 nand P2_U2734 P2_R2099_U128 ; P2_R2099_U33
g24336 not P2_U2733 ; P2_R2099_U34
g24337 nand P2_U2733 P2_R2099_U129 ; P2_R2099_U35
g24338 not P2_U2732 ; P2_R2099_U36
g24339 nand P2_U2732 P2_R2099_U130 ; P2_R2099_U37
g24340 not P2_U2731 ; P2_R2099_U38
g24341 nand P2_U2731 P2_R2099_U131 ; P2_R2099_U39
g24342 not P2_U2730 ; P2_R2099_U40
g24343 nand P2_U2730 P2_R2099_U132 ; P2_R2099_U41
g24344 not P2_U2729 ; P2_R2099_U42
g24345 nand P2_U2729 P2_R2099_U133 ; P2_R2099_U43
g24346 not P2_U2728 ; P2_R2099_U44
g24347 nand P2_U2728 P2_R2099_U134 ; P2_R2099_U45
g24348 not P2_U2727 ; P2_R2099_U46
g24349 nand P2_U2727 P2_R2099_U135 ; P2_R2099_U47
g24350 not P2_U2726 ; P2_R2099_U48
g24351 nand P2_U2726 P2_R2099_U136 ; P2_R2099_U49
g24352 not P2_U2725 ; P2_R2099_U50
g24353 nand P2_U2725 P2_R2099_U137 ; P2_R2099_U51
g24354 not P2_U2724 ; P2_R2099_U52
g24355 nand P2_U2724 P2_R2099_U138 ; P2_R2099_U53
g24356 not P2_U2723 ; P2_R2099_U54
g24357 nand P2_U2723 P2_R2099_U139 ; P2_R2099_U55
g24358 not P2_U2722 ; P2_R2099_U56
g24359 nand P2_U2722 P2_R2099_U140 ; P2_R2099_U57
g24360 not P2_U2721 ; P2_R2099_U58
g24361 nand P2_U2721 P2_R2099_U141 ; P2_R2099_U59
g24362 not P2_U2720 ; P2_R2099_U60
g24363 nand P2_U2720 P2_R2099_U142 ; P2_R2099_U61
g24364 not P2_U2719 ; P2_R2099_U62
g24365 nand P2_U2719 P2_R2099_U143 ; P2_R2099_U63
g24366 not P2_U2718 ; P2_R2099_U64
g24367 nand P2_U2718 P2_R2099_U144 ; P2_R2099_U65
g24368 not P2_U2717 ; P2_R2099_U66
g24369 nand P2_R2099_U150 P2_R2099_U149 ; P2_R2099_U67
g24370 nand P2_R2099_U152 P2_R2099_U151 ; P2_R2099_U68
g24371 nand P2_R2099_U154 P2_R2099_U153 ; P2_R2099_U69
g24372 nand P2_R2099_U156 P2_R2099_U155 ; P2_R2099_U70
g24373 nand P2_R2099_U158 P2_R2099_U157 ; P2_R2099_U71
g24374 nand P2_R2099_U169 P2_R2099_U168 ; P2_R2099_U72
g24375 nand P2_R2099_U171 P2_R2099_U170 ; P2_R2099_U73
g24376 nand P2_R2099_U180 P2_R2099_U179 ; P2_R2099_U74
g24377 nand P2_R2099_U182 P2_R2099_U181 ; P2_R2099_U75
g24378 nand P2_R2099_U184 P2_R2099_U183 ; P2_R2099_U76
g24379 nand P2_R2099_U186 P2_R2099_U185 ; P2_R2099_U77
g24380 nand P2_R2099_U188 P2_R2099_U187 ; P2_R2099_U78
g24381 nand P2_R2099_U190 P2_R2099_U189 ; P2_R2099_U79
g24382 nand P2_R2099_U192 P2_R2099_U191 ; P2_R2099_U80
g24383 nand P2_R2099_U194 P2_R2099_U193 ; P2_R2099_U81
g24384 nand P2_R2099_U196 P2_R2099_U195 ; P2_R2099_U82
g24385 nand P2_R2099_U198 P2_R2099_U197 ; P2_R2099_U83
g24386 nand P2_R2099_U205 P2_R2099_U204 ; P2_R2099_U84
g24387 nand P2_R2099_U207 P2_R2099_U206 ; P2_R2099_U85
g24388 nand P2_R2099_U209 P2_R2099_U208 ; P2_R2099_U86
g24389 nand P2_R2099_U211 P2_R2099_U210 ; P2_R2099_U87
g24390 nand P2_R2099_U213 P2_R2099_U212 ; P2_R2099_U88
g24391 nand P2_R2099_U215 P2_R2099_U214 ; P2_R2099_U89
g24392 nand P2_R2099_U217 P2_R2099_U216 ; P2_R2099_U90
g24393 nand P2_R2099_U219 P2_R2099_U218 ; P2_R2099_U91
g24394 nand P2_R2099_U221 P2_R2099_U220 ; P2_R2099_U92
g24395 nand P2_R2099_U223 P2_R2099_U222 ; P2_R2099_U93
g24396 nand P2_R2099_U225 P2_R2099_U224 ; P2_R2099_U94
g24397 nand P2_R2099_U167 P2_R2099_U166 ; P2_R2099_U95
g24398 nand P2_R2099_U178 P2_R2099_U177 ; P2_R2099_U96
g24399 nand P2_R2099_U118 P2_R2099_U117 ; P2_R2099_U97
g24400 and P2_R2099_U160 P2_R2099_U159 ; P2_R2099_U98
g24401 and P2_R2099_U162 P2_R2099_U161 ; P2_R2099_U99
g24402 nand P2_R2099_U114 P2_R2099_U113 ; P2_R2099_U100
g24403 not P2_U2716 ; P2_R2099_U101
g24404 nand P2_U2717 P2_R2099_U145 ; P2_R2099_U102
g24405 and P2_R2099_U173 P2_R2099_U172 ; P2_R2099_U103
g24406 nand P2_R2099_U106 P2_R2099_U110 ; P2_R2099_U104
g24407 nand P2_U2751 P2_U2747 ; P2_R2099_U105
g24408 nand P2_U2746 P2_U2747 P2_U2751 ; P2_R2099_U106
g24409 and P2_R2099_U203 P2_R2099_U202 ; P2_R2099_U107
g24410 not P2_R2099_U106 ; P2_R2099_U108
g24411 nand P2_R2099_U9 P2_R2099_U105 ; P2_R2099_U109
g24412 nand P2_U2750 P2_R2099_U109 ; P2_R2099_U110
g24413 not P2_R2099_U104 ; P2_R2099_U111
g24414 or P2_U2749 P2_U2745 ; P2_R2099_U112
g24415 nand P2_R2099_U112 P2_R2099_U104 ; P2_R2099_U113
g24416 nand P2_U2745 P2_U2749 ; P2_R2099_U114
g24417 not P2_R2099_U100 ; P2_R2099_U115
g24418 or P2_U2748 P2_U2744 ; P2_R2099_U116
g24419 nand P2_R2099_U116 P2_R2099_U100 ; P2_R2099_U117
g24420 nand P2_U2744 P2_U2748 ; P2_R2099_U118
g24421 not P2_R2099_U97 ; P2_R2099_U119
g24422 not P2_R2099_U15 ; P2_R2099_U120
g24423 not P2_R2099_U17 ; P2_R2099_U121
g24424 not P2_R2099_U19 ; P2_R2099_U122
g24425 not P2_R2099_U21 ; P2_R2099_U123
g24426 not P2_R2099_U24 ; P2_R2099_U124
g24427 not P2_R2099_U25 ; P2_R2099_U125
g24428 not P2_R2099_U27 ; P2_R2099_U126
g24429 not P2_R2099_U29 ; P2_R2099_U127
g24430 not P2_R2099_U31 ; P2_R2099_U128
g24431 not P2_R2099_U33 ; P2_R2099_U129
g24432 not P2_R2099_U35 ; P2_R2099_U130
g24433 not P2_R2099_U37 ; P2_R2099_U131
g24434 not P2_R2099_U39 ; P2_R2099_U132
g24435 not P2_R2099_U41 ; P2_R2099_U133
g24436 not P2_R2099_U43 ; P2_R2099_U134
g24437 not P2_R2099_U45 ; P2_R2099_U135
g24438 not P2_R2099_U47 ; P2_R2099_U136
g24439 not P2_R2099_U49 ; P2_R2099_U137
g24440 not P2_R2099_U51 ; P2_R2099_U138
g24441 not P2_R2099_U53 ; P2_R2099_U139
g24442 not P2_R2099_U55 ; P2_R2099_U140
g24443 not P2_R2099_U57 ; P2_R2099_U141
g24444 not P2_R2099_U59 ; P2_R2099_U142
g24445 not P2_R2099_U61 ; P2_R2099_U143
g24446 not P2_R2099_U63 ; P2_R2099_U144
g24447 not P2_R2099_U65 ; P2_R2099_U145
g24448 not P2_R2099_U102 ; P2_R2099_U146
g24449 not P2_R2099_U105 ; P2_R2099_U147
g24450 nand P2_R2099_U201 P2_R2099_U9 ; P2_R2099_U148
g24451 nand P2_U2738 P2_R2099_U24 ; P2_R2099_U149
g24452 nand P2_R2099_U124 P2_R2099_U23 ; P2_R2099_U150
g24453 nand P2_U2739 P2_R2099_U21 ; P2_R2099_U151
g24454 nand P2_R2099_U123 P2_R2099_U22 ; P2_R2099_U152
g24455 nand P2_U2740 P2_R2099_U19 ; P2_R2099_U153
g24456 nand P2_R2099_U122 P2_R2099_U20 ; P2_R2099_U154
g24457 nand P2_U2741 P2_R2099_U17 ; P2_R2099_U155
g24458 nand P2_R2099_U121 P2_R2099_U18 ; P2_R2099_U156
g24459 nand P2_U2742 P2_R2099_U15 ; P2_R2099_U157
g24460 nand P2_R2099_U120 P2_R2099_U16 ; P2_R2099_U158
g24461 nand P2_U2743 P2_R2099_U97 ; P2_R2099_U159
g24462 nand P2_R2099_U119 P2_R2099_U14 ; P2_R2099_U160
g24463 nand P2_U2744 P2_R2099_U12 ; P2_R2099_U161
g24464 nand P2_U2748 P2_R2099_U13 ; P2_R2099_U162
g24465 nand P2_U2744 P2_R2099_U12 ; P2_R2099_U163
g24466 nand P2_U2748 P2_R2099_U13 ; P2_R2099_U164
g24467 nand P2_R2099_U164 P2_R2099_U163 ; P2_R2099_U165
g24468 nand P2_R2099_U99 P2_R2099_U100 ; P2_R2099_U166
g24469 nand P2_R2099_U115 P2_R2099_U165 ; P2_R2099_U167
g24470 nand P2_U2716 P2_R2099_U102 ; P2_R2099_U168
g24471 nand P2_R2099_U146 P2_R2099_U101 ; P2_R2099_U169
g24472 nand P2_U2717 P2_R2099_U65 ; P2_R2099_U170
g24473 nand P2_R2099_U145 P2_R2099_U66 ; P2_R2099_U171
g24474 nand P2_U2745 P2_R2099_U10 ; P2_R2099_U172
g24475 nand P2_U2749 P2_R2099_U11 ; P2_R2099_U173
g24476 nand P2_U2745 P2_R2099_U10 ; P2_R2099_U174
g24477 nand P2_U2749 P2_R2099_U11 ; P2_R2099_U175
g24478 nand P2_R2099_U175 P2_R2099_U174 ; P2_R2099_U176
g24479 nand P2_R2099_U103 P2_R2099_U104 ; P2_R2099_U177
g24480 nand P2_R2099_U111 P2_R2099_U176 ; P2_R2099_U178
g24481 nand P2_U2718 P2_R2099_U63 ; P2_R2099_U179
g24482 nand P2_R2099_U144 P2_R2099_U64 ; P2_R2099_U180
g24483 nand P2_U2719 P2_R2099_U61 ; P2_R2099_U181
g24484 nand P2_R2099_U143 P2_R2099_U62 ; P2_R2099_U182
g24485 nand P2_U2720 P2_R2099_U59 ; P2_R2099_U183
g24486 nand P2_R2099_U142 P2_R2099_U60 ; P2_R2099_U184
g24487 nand P2_U2721 P2_R2099_U57 ; P2_R2099_U185
g24488 nand P2_R2099_U141 P2_R2099_U58 ; P2_R2099_U186
g24489 nand P2_U2722 P2_R2099_U55 ; P2_R2099_U187
g24490 nand P2_R2099_U140 P2_R2099_U56 ; P2_R2099_U188
g24491 nand P2_U2723 P2_R2099_U53 ; P2_R2099_U189
g24492 nand P2_R2099_U139 P2_R2099_U54 ; P2_R2099_U190
g24493 nand P2_U2724 P2_R2099_U51 ; P2_R2099_U191
g24494 nand P2_R2099_U138 P2_R2099_U52 ; P2_R2099_U192
g24495 nand P2_U2725 P2_R2099_U49 ; P2_R2099_U193
g24496 nand P2_R2099_U137 P2_R2099_U50 ; P2_R2099_U194
g24497 nand P2_U2726 P2_R2099_U47 ; P2_R2099_U195
g24498 nand P2_R2099_U136 P2_R2099_U48 ; P2_R2099_U196
g24499 nand P2_U2727 P2_R2099_U45 ; P2_R2099_U197
g24500 nand P2_R2099_U135 P2_R2099_U46 ; P2_R2099_U198
g24501 nand P2_U2750 P2_R2099_U105 ; P2_R2099_U199
g24502 nand P2_R2099_U147 P2_R2099_U8 ; P2_R2099_U200
g24503 nand P2_R2099_U200 P2_R2099_U199 ; P2_R2099_U201
g24504 nand P2_U2746 P2_R2099_U105 P2_R2099_U8 ; P2_R2099_U202
g24505 nand P2_R2099_U108 P2_U2750 ; P2_R2099_U203
g24506 nand P2_U2728 P2_R2099_U43 ; P2_R2099_U204
g24507 nand P2_R2099_U134 P2_R2099_U44 ; P2_R2099_U205
g24508 nand P2_U2729 P2_R2099_U41 ; P2_R2099_U206
g24509 nand P2_R2099_U133 P2_R2099_U42 ; P2_R2099_U207
g24510 nand P2_U2730 P2_R2099_U39 ; P2_R2099_U208
g24511 nand P2_R2099_U132 P2_R2099_U40 ; P2_R2099_U209
g24512 nand P2_U2731 P2_R2099_U37 ; P2_R2099_U210
g24513 nand P2_R2099_U131 P2_R2099_U38 ; P2_R2099_U211
g24514 nand P2_U2732 P2_R2099_U35 ; P2_R2099_U212
g24515 nand P2_R2099_U130 P2_R2099_U36 ; P2_R2099_U213
g24516 nand P2_U2733 P2_R2099_U33 ; P2_R2099_U214
g24517 nand P2_R2099_U129 P2_R2099_U34 ; P2_R2099_U215
g24518 nand P2_U2734 P2_R2099_U31 ; P2_R2099_U216
g24519 nand P2_R2099_U128 P2_R2099_U32 ; P2_R2099_U217
g24520 nand P2_U2735 P2_R2099_U29 ; P2_R2099_U218
g24521 nand P2_R2099_U127 P2_R2099_U30 ; P2_R2099_U219
g24522 nand P2_U2736 P2_R2099_U27 ; P2_R2099_U220
g24523 nand P2_R2099_U126 P2_R2099_U28 ; P2_R2099_U221
g24524 nand P2_U2737 P2_R2099_U25 ; P2_R2099_U222
g24525 nand P2_R2099_U125 P2_R2099_U26 ; P2_R2099_U223
g24526 nand P2_U2751 P2_R2099_U6 ; P2_R2099_U224
g24527 nand P2_U2747 P2_R2099_U7 ; P2_R2099_U225
g24528 and P2_ADD_391_1196_U301 P2_ADD_391_1196_U299 ; P2_ADD_391_1196_U5
g24529 and P2_ADD_391_1196_U296 P2_ADD_391_1196_U294 ; P2_ADD_391_1196_U6
g24530 and P2_ADD_391_1196_U292 P2_ADD_391_1196_U290 ; P2_ADD_391_1196_U7
g24531 and P2_ADD_391_1196_U287 P2_ADD_391_1196_U283 ; P2_ADD_391_1196_U8
g24532 and P2_ADD_391_1196_U205 P2_ADD_391_1196_U203 ; P2_ADD_391_1196_U9
g24533 and P2_ADD_391_1196_U201 P2_ADD_391_1196_U199 ; P2_ADD_391_1196_U10
g24534 and P2_ADD_391_1196_U196 P2_ADD_391_1196_U192 ; P2_ADD_391_1196_U11
g24535 nand P2_ADD_391_1196_U144 P2_ADD_391_1196_U306 ; P2_ADD_391_1196_U12
g24536 not P2_R2182_U72 ; P2_ADD_391_1196_U13
g24537 not P2_R2096_U71 ; P2_ADD_391_1196_U14
g24538 not P2_R2182_U73 ; P2_ADD_391_1196_U15
g24539 not P2_R2096_U72 ; P2_ADD_391_1196_U16
g24540 not P2_R2182_U74 ; P2_ADD_391_1196_U17
g24541 not P2_R2096_U73 ; P2_ADD_391_1196_U18
g24542 not P2_R2096_U68 ; P2_ADD_391_1196_U19
g24543 not P2_R2182_U69 ; P2_ADD_391_1196_U20
g24544 not P2_R2182_U68 ; P2_ADD_391_1196_U21
g24545 nand P2_R2182_U69 P2_R2096_U68 ; P2_ADD_391_1196_U22
g24546 not P2_R2096_U51 ; P2_ADD_391_1196_U23
g24547 not P2_R2182_U40 ; P2_ADD_391_1196_U24
g24548 not P2_R2096_U77 ; P2_ADD_391_1196_U25
g24549 not P2_R2182_U76 ; P2_ADD_391_1196_U26
g24550 not P2_R2096_U75 ; P2_ADD_391_1196_U27
g24551 not P2_R2182_U75 ; P2_ADD_391_1196_U28
g24552 not P2_R2096_U74 ; P2_ADD_391_1196_U29
g24553 nand P2_ADD_391_1196_U39 P2_ADD_391_1196_U180 ; P2_ADD_391_1196_U30
g24554 not P2_R2182_U71 ; P2_ADD_391_1196_U31
g24555 not P2_R2096_U70 ; P2_ADD_391_1196_U32
g24556 not P2_R2096_U69 ; P2_ADD_391_1196_U33
g24557 not P2_R2182_U70 ; P2_ADD_391_1196_U34
g24558 nand P2_ADD_391_1196_U190 P2_ADD_391_1196_U189 ; P2_ADD_391_1196_U35
g24559 nand P2_ADD_391_1196_U35 P2_ADD_391_1196_U193 ; P2_ADD_391_1196_U36
g24560 nand P2_ADD_391_1196_U184 P2_ADD_391_1196_U182 P2_ADD_391_1196_U183 ; P2_ADD_391_1196_U37
g24561 nand P2_ADD_391_1196_U176 P2_ADD_391_1196_U175 ; P2_ADD_391_1196_U38
g24562 nand P2_ADD_391_1196_U38 P2_ADD_391_1196_U178 ; P2_ADD_391_1196_U39
g24563 not P2_R2182_U91 ; P2_ADD_391_1196_U40
g24564 not P2_R2096_U92 ; P2_ADD_391_1196_U41
g24565 not P2_R2182_U92 ; P2_ADD_391_1196_U42
g24566 not P2_R2096_U93 ; P2_ADD_391_1196_U43
g24567 not P2_R2182_U93 ; P2_ADD_391_1196_U44
g24568 not P2_R2096_U94 ; P2_ADD_391_1196_U45
g24569 not P2_R2182_U95 ; P2_ADD_391_1196_U46
g24570 not P2_R2096_U96 ; P2_ADD_391_1196_U47
g24571 not P2_R2182_U96 ; P2_ADD_391_1196_U48
g24572 not P2_R2096_U97 ; P2_ADD_391_1196_U49
g24573 nand P2_ADD_391_1196_U36 P2_ADD_391_1196_U206 ; P2_ADD_391_1196_U50
g24574 not P2_R2182_U94 ; P2_ADD_391_1196_U51
g24575 not P2_R2096_U95 ; P2_ADD_391_1196_U52
g24576 nand P2_ADD_391_1196_U85 P2_ADD_391_1196_U220 ; P2_ADD_391_1196_U53
g24577 not P2_R2182_U90 ; P2_ADD_391_1196_U54
g24578 not P2_R2096_U91 ; P2_ADD_391_1196_U55
g24579 not P2_R2182_U89 ; P2_ADD_391_1196_U56
g24580 not P2_R2096_U90 ; P2_ADD_391_1196_U57
g24581 not P2_R2182_U88 ; P2_ADD_391_1196_U58
g24582 not P2_R2096_U89 ; P2_ADD_391_1196_U59
g24583 not P2_R2182_U87 ; P2_ADD_391_1196_U60
g24584 not P2_R2096_U88 ; P2_ADD_391_1196_U61
g24585 not P2_R2182_U86 ; P2_ADD_391_1196_U62
g24586 not P2_R2096_U87 ; P2_ADD_391_1196_U63
g24587 not P2_R2182_U85 ; P2_ADD_391_1196_U64
g24588 not P2_R2096_U86 ; P2_ADD_391_1196_U65
g24589 not P2_R2182_U84 ; P2_ADD_391_1196_U66
g24590 not P2_R2096_U85 ; P2_ADD_391_1196_U67
g24591 not P2_R2182_U83 ; P2_ADD_391_1196_U68
g24592 not P2_R2096_U84 ; P2_ADD_391_1196_U69
g24593 not P2_R2182_U82 ; P2_ADD_391_1196_U70
g24594 not P2_R2096_U83 ; P2_ADD_391_1196_U71
g24595 not P2_R2182_U81 ; P2_ADD_391_1196_U72
g24596 not P2_R2096_U82 ; P2_ADD_391_1196_U73
g24597 not P2_R2182_U80 ; P2_ADD_391_1196_U74
g24598 not P2_R2096_U81 ; P2_ADD_391_1196_U75
g24599 not P2_R2182_U79 ; P2_ADD_391_1196_U76
g24600 not P2_R2096_U80 ; P2_ADD_391_1196_U77
g24601 not P2_R2096_U79 ; P2_ADD_391_1196_U78
g24602 not P2_R2182_U78 ; P2_ADD_391_1196_U79
g24603 not P2_R2096_U78 ; P2_ADD_391_1196_U80
g24604 not P2_R2182_U77 ; P2_ADD_391_1196_U81
g24605 nand P2_ADD_391_1196_U278 P2_ADD_391_1196_U277 ; P2_ADD_391_1196_U82
g24606 nand P2_ADD_391_1196_U224 P2_ADD_391_1196_U222 P2_ADD_391_1196_U223 ; P2_ADD_391_1196_U83
g24607 nand P2_ADD_391_1196_U216 P2_ADD_391_1196_U215 ; P2_ADD_391_1196_U84
g24608 nand P2_ADD_391_1196_U84 P2_ADD_391_1196_U218 ; P2_ADD_391_1196_U85
g24609 nand P2_ADD_391_1196_U210 P2_ADD_391_1196_U208 P2_ADD_391_1196_U209 ; P2_ADD_391_1196_U86
g24610 nand P2_ADD_391_1196_U478 P2_ADD_391_1196_U477 ; P2_ADD_391_1196_U87
g24611 nand P2_ADD_391_1196_U315 P2_ADD_391_1196_U314 ; P2_ADD_391_1196_U88
g24612 nand P2_ADD_391_1196_U322 P2_ADD_391_1196_U321 ; P2_ADD_391_1196_U89
g24613 nand P2_ADD_391_1196_U331 P2_ADD_391_1196_U330 ; P2_ADD_391_1196_U90
g24614 nand P2_ADD_391_1196_U338 P2_ADD_391_1196_U337 ; P2_ADD_391_1196_U91
g24615 nand P2_ADD_391_1196_U350 P2_ADD_391_1196_U349 ; P2_ADD_391_1196_U92
g24616 nand P2_ADD_391_1196_U357 P2_ADD_391_1196_U356 ; P2_ADD_391_1196_U93
g24617 nand P2_ADD_391_1196_U364 P2_ADD_391_1196_U363 ; P2_ADD_391_1196_U94
g24618 nand P2_ADD_391_1196_U371 P2_ADD_391_1196_U370 ; P2_ADD_391_1196_U95
g24619 nand P2_ADD_391_1196_U378 P2_ADD_391_1196_U377 ; P2_ADD_391_1196_U96
g24620 nand P2_ADD_391_1196_U385 P2_ADD_391_1196_U384 ; P2_ADD_391_1196_U97
g24621 nand P2_ADD_391_1196_U392 P2_ADD_391_1196_U391 ; P2_ADD_391_1196_U98
g24622 nand P2_ADD_391_1196_U399 P2_ADD_391_1196_U398 ; P2_ADD_391_1196_U99
g24623 nand P2_ADD_391_1196_U406 P2_ADD_391_1196_U405 ; P2_ADD_391_1196_U100
g24624 nand P2_ADD_391_1196_U413 P2_ADD_391_1196_U412 ; P2_ADD_391_1196_U101
g24625 nand P2_ADD_391_1196_U420 P2_ADD_391_1196_U419 ; P2_ADD_391_1196_U102
g24626 nand P2_ADD_391_1196_U432 P2_ADD_391_1196_U431 ; P2_ADD_391_1196_U103
g24627 nand P2_ADD_391_1196_U439 P2_ADD_391_1196_U438 ; P2_ADD_391_1196_U104
g24628 nand P2_ADD_391_1196_U446 P2_ADD_391_1196_U445 ; P2_ADD_391_1196_U105
g24629 nand P2_ADD_391_1196_U453 P2_ADD_391_1196_U452 ; P2_ADD_391_1196_U106
g24630 nand P2_ADD_391_1196_U460 P2_ADD_391_1196_U459 ; P2_ADD_391_1196_U107
g24631 nand P2_ADD_391_1196_U469 P2_ADD_391_1196_U468 ; P2_ADD_391_1196_U108
g24632 nand P2_ADD_391_1196_U476 P2_ADD_391_1196_U475 ; P2_ADD_391_1196_U109
g24633 and P2_ADD_391_1196_U308 P2_ADD_391_1196_U307 ; P2_ADD_391_1196_U110
g24634 and P2_ADD_391_1196_U310 P2_ADD_391_1196_U309 ; P2_ADD_391_1196_U111
g24635 nand P2_ADD_391_1196_U37 P2_ADD_391_1196_U186 ; P2_ADD_391_1196_U112
g24636 and P2_ADD_391_1196_U317 P2_ADD_391_1196_U316 ; P2_ADD_391_1196_U113
g24637 and P2_ADD_391_1196_U324 P2_ADD_391_1196_U323 ; P2_ADD_391_1196_U114
g24638 and P2_ADD_391_1196_U326 P2_ADD_391_1196_U325 ; P2_ADD_391_1196_U115
g24639 nand P2_ADD_391_1196_U172 P2_ADD_391_1196_U171 ; P2_ADD_391_1196_U116
g24640 and P2_ADD_391_1196_U333 P2_ADD_391_1196_U332 ; P2_ADD_391_1196_U117
g24641 nand P2_ADD_391_1196_U168 P2_ADD_391_1196_U167 ; P2_ADD_391_1196_U118
g24642 not P2_R2182_U41 ; P2_ADD_391_1196_U119
g24643 not P2_R2096_U76 ; P2_ADD_391_1196_U120
g24644 and P2_ADD_391_1196_U340 P2_ADD_391_1196_U339 ; P2_ADD_391_1196_U121
g24645 and P2_ADD_391_1196_U345 P2_ADD_391_1196_U344 ; P2_ADD_391_1196_U122
g24646 nand P2_ADD_391_1196_U143 P2_ADD_391_1196_U164 ; P2_ADD_391_1196_U123
g24647 and P2_ADD_391_1196_U352 P2_ADD_391_1196_U351 ; P2_ADD_391_1196_U124
g24648 and P2_ADD_391_1196_U359 P2_ADD_391_1196_U358 ; P2_ADD_391_1196_U125
g24649 nand P2_ADD_391_1196_U274 P2_ADD_391_1196_U273 ; P2_ADD_391_1196_U126
g24650 and P2_ADD_391_1196_U366 P2_ADD_391_1196_U365 ; P2_ADD_391_1196_U127
g24651 nand P2_ADD_391_1196_U270 P2_ADD_391_1196_U269 ; P2_ADD_391_1196_U128
g24652 and P2_ADD_391_1196_U373 P2_ADD_391_1196_U372 ; P2_ADD_391_1196_U129
g24653 nand P2_ADD_391_1196_U266 P2_ADD_391_1196_U265 ; P2_ADD_391_1196_U130
g24654 and P2_ADD_391_1196_U380 P2_ADD_391_1196_U379 ; P2_ADD_391_1196_U131
g24655 nand P2_ADD_391_1196_U262 P2_ADD_391_1196_U261 ; P2_ADD_391_1196_U132
g24656 and P2_ADD_391_1196_U387 P2_ADD_391_1196_U386 ; P2_ADD_391_1196_U133
g24657 nand P2_ADD_391_1196_U258 P2_ADD_391_1196_U257 ; P2_ADD_391_1196_U134
g24658 and P2_ADD_391_1196_U394 P2_ADD_391_1196_U393 ; P2_ADD_391_1196_U135
g24659 nand P2_ADD_391_1196_U254 P2_ADD_391_1196_U253 ; P2_ADD_391_1196_U136
g24660 and P2_ADD_391_1196_U401 P2_ADD_391_1196_U400 ; P2_ADD_391_1196_U137
g24661 nand P2_ADD_391_1196_U250 P2_ADD_391_1196_U249 ; P2_ADD_391_1196_U138
g24662 and P2_ADD_391_1196_U408 P2_ADD_391_1196_U407 ; P2_ADD_391_1196_U139
g24663 nand P2_ADD_391_1196_U246 P2_ADD_391_1196_U245 ; P2_ADD_391_1196_U140
g24664 and P2_ADD_391_1196_U415 P2_ADD_391_1196_U414 ; P2_ADD_391_1196_U141
g24665 nand P2_ADD_391_1196_U242 P2_ADD_391_1196_U241 ; P2_ADD_391_1196_U142
g24666 nand P2_R2096_U51 P2_ADD_391_1196_U162 ; P2_ADD_391_1196_U143
g24667 and P2_ADD_391_1196_U425 P2_ADD_391_1196_U424 ; P2_ADD_391_1196_U144
g24668 and P2_ADD_391_1196_U427 P2_ADD_391_1196_U426 ; P2_ADD_391_1196_U145
g24669 nand P2_ADD_391_1196_U238 P2_ADD_391_1196_U237 ; P2_ADD_391_1196_U146
g24670 and P2_ADD_391_1196_U434 P2_ADD_391_1196_U433 ; P2_ADD_391_1196_U147
g24671 nand P2_ADD_391_1196_U234 P2_ADD_391_1196_U233 ; P2_ADD_391_1196_U148
g24672 and P2_ADD_391_1196_U441 P2_ADD_391_1196_U440 ; P2_ADD_391_1196_U149
g24673 nand P2_ADD_391_1196_U230 P2_ADD_391_1196_U229 ; P2_ADD_391_1196_U150
g24674 and P2_ADD_391_1196_U448 P2_ADD_391_1196_U447 ; P2_ADD_391_1196_U151
g24675 nand P2_ADD_391_1196_U83 P2_ADD_391_1196_U226 ; P2_ADD_391_1196_U152
g24676 and P2_ADD_391_1196_U455 P2_ADD_391_1196_U454 ; P2_ADD_391_1196_U153
g24677 and P2_ADD_391_1196_U462 P2_ADD_391_1196_U461 ; P2_ADD_391_1196_U154
g24678 and P2_ADD_391_1196_U464 P2_ADD_391_1196_U463 ; P2_ADD_391_1196_U155
g24679 nand P2_ADD_391_1196_U86 P2_ADD_391_1196_U212 ; P2_ADD_391_1196_U156
g24680 and P2_ADD_391_1196_U471 P2_ADD_391_1196_U470 ; P2_ADD_391_1196_U157
g24681 nand P2_R2096_U97 P2_R2182_U96 ; P2_ADD_391_1196_U158
g24682 nand P2_R2096_U93 P2_R2182_U92 ; P2_ADD_391_1196_U159
g24683 not P2_ADD_391_1196_U143 ; P2_ADD_391_1196_U160
g24684 nand P2_R2096_U72 P2_R2182_U73 ; P2_ADD_391_1196_U161
g24685 not P2_ADD_391_1196_U22 ; P2_ADD_391_1196_U162
g24686 nand P2_ADD_391_1196_U23 P2_ADD_391_1196_U22 ; P2_ADD_391_1196_U163
g24687 nand P2_R2182_U68 P2_ADD_391_1196_U163 ; P2_ADD_391_1196_U164
g24688 not P2_ADD_391_1196_U123 ; P2_ADD_391_1196_U165
g24689 or P2_R2182_U40 P2_R2096_U77 ; P2_ADD_391_1196_U166
g24690 nand P2_ADD_391_1196_U166 P2_ADD_391_1196_U123 ; P2_ADD_391_1196_U167
g24691 nand P2_R2096_U77 P2_R2182_U40 ; P2_ADD_391_1196_U168
g24692 not P2_ADD_391_1196_U118 ; P2_ADD_391_1196_U169
g24693 or P2_R2182_U76 P2_R2096_U75 ; P2_ADD_391_1196_U170
g24694 nand P2_ADD_391_1196_U170 P2_ADD_391_1196_U118 ; P2_ADD_391_1196_U171
g24695 nand P2_R2096_U75 P2_R2182_U76 ; P2_ADD_391_1196_U172
g24696 not P2_ADD_391_1196_U116 ; P2_ADD_391_1196_U173
g24697 or P2_R2182_U75 P2_R2096_U74 ; P2_ADD_391_1196_U174
g24698 nand P2_ADD_391_1196_U174 P2_ADD_391_1196_U116 ; P2_ADD_391_1196_U175
g24699 nand P2_R2096_U74 P2_R2182_U75 ; P2_ADD_391_1196_U176
g24700 not P2_ADD_391_1196_U38 ; P2_ADD_391_1196_U177
g24701 or P2_R2096_U73 P2_R2182_U74 ; P2_ADD_391_1196_U178
g24702 not P2_ADD_391_1196_U39 ; P2_ADD_391_1196_U179
g24703 nand P2_R2096_U73 P2_R2182_U74 ; P2_ADD_391_1196_U180
g24704 not P2_ADD_391_1196_U30 ; P2_ADD_391_1196_U181
g24705 nand P2_ADD_391_1196_U181 P2_ADD_391_1196_U161 ; P2_ADD_391_1196_U182
g24706 or P2_R2096_U71 P2_R2182_U72 ; P2_ADD_391_1196_U183
g24707 or P2_R2096_U72 P2_R2182_U73 ; P2_ADD_391_1196_U184
g24708 not P2_ADD_391_1196_U37 ; P2_ADD_391_1196_U185
g24709 nand P2_R2096_U71 P2_R2182_U72 ; P2_ADD_391_1196_U186
g24710 not P2_ADD_391_1196_U112 ; P2_ADD_391_1196_U187
g24711 or P2_R2182_U71 P2_R2096_U70 ; P2_ADD_391_1196_U188
g24712 nand P2_ADD_391_1196_U188 P2_ADD_391_1196_U112 ; P2_ADD_391_1196_U189
g24713 nand P2_R2096_U70 P2_R2182_U71 ; P2_ADD_391_1196_U190
g24714 not P2_ADD_391_1196_U35 ; P2_ADD_391_1196_U191
g24715 nand P2_ADD_391_1196_U110 P2_ADD_391_1196_U191 ; P2_ADD_391_1196_U192
g24716 or P2_R2096_U69 P2_R2182_U70 ; P2_ADD_391_1196_U193
g24717 not P2_ADD_391_1196_U36 ; P2_ADD_391_1196_U194
g24718 nand P2_R2182_U70 P2_R2096_U69 ; P2_ADD_391_1196_U195
g24719 nand P2_ADD_391_1196_U194 P2_ADD_391_1196_U195 ; P2_ADD_391_1196_U196
g24720 or P2_R2182_U73 P2_R2096_U72 ; P2_ADD_391_1196_U197
g24721 nand P2_ADD_391_1196_U197 P2_ADD_391_1196_U30 ; P2_ADD_391_1196_U198
g24722 nand P2_ADD_391_1196_U198 P2_ADD_391_1196_U161 P2_ADD_391_1196_U113 ; P2_ADD_391_1196_U199
g24723 nand P2_R2096_U71 P2_R2182_U72 ; P2_ADD_391_1196_U200
g24724 nand P2_ADD_391_1196_U185 P2_ADD_391_1196_U200 ; P2_ADD_391_1196_U201
g24725 or P2_R2096_U72 P2_R2182_U73 ; P2_ADD_391_1196_U202
g24726 nand P2_ADD_391_1196_U114 P2_ADD_391_1196_U177 ; P2_ADD_391_1196_U203
g24727 nand P2_R2096_U73 P2_R2182_U74 ; P2_ADD_391_1196_U204
g24728 nand P2_ADD_391_1196_U179 P2_ADD_391_1196_U204 ; P2_ADD_391_1196_U205
g24729 nand P2_R2182_U70 P2_R2096_U69 ; P2_ADD_391_1196_U206
g24730 not P2_ADD_391_1196_U50 ; P2_ADD_391_1196_U207
g24731 nand P2_ADD_391_1196_U207 P2_ADD_391_1196_U158 ; P2_ADD_391_1196_U208
g24732 or P2_R2096_U96 P2_R2182_U95 ; P2_ADD_391_1196_U209
g24733 or P2_R2096_U97 P2_R2182_U96 ; P2_ADD_391_1196_U210
g24734 not P2_ADD_391_1196_U86 ; P2_ADD_391_1196_U211
g24735 nand P2_R2096_U96 P2_R2182_U95 ; P2_ADD_391_1196_U212
g24736 not P2_ADD_391_1196_U156 ; P2_ADD_391_1196_U213
g24737 or P2_R2182_U94 P2_R2096_U95 ; P2_ADD_391_1196_U214
g24738 nand P2_ADD_391_1196_U214 P2_ADD_391_1196_U156 ; P2_ADD_391_1196_U215
g24739 nand P2_R2096_U95 P2_R2182_U94 ; P2_ADD_391_1196_U216
g24740 not P2_ADD_391_1196_U84 ; P2_ADD_391_1196_U217
g24741 or P2_R2096_U94 P2_R2182_U93 ; P2_ADD_391_1196_U218
g24742 not P2_ADD_391_1196_U85 ; P2_ADD_391_1196_U219
g24743 nand P2_R2096_U94 P2_R2182_U93 ; P2_ADD_391_1196_U220
g24744 not P2_ADD_391_1196_U53 ; P2_ADD_391_1196_U221
g24745 nand P2_ADD_391_1196_U221 P2_ADD_391_1196_U159 ; P2_ADD_391_1196_U222
g24746 or P2_R2096_U92 P2_R2182_U91 ; P2_ADD_391_1196_U223
g24747 or P2_R2096_U93 P2_R2182_U92 ; P2_ADD_391_1196_U224
g24748 not P2_ADD_391_1196_U83 ; P2_ADD_391_1196_U225
g24749 nand P2_R2096_U92 P2_R2182_U91 ; P2_ADD_391_1196_U226
g24750 not P2_ADD_391_1196_U152 ; P2_ADD_391_1196_U227
g24751 or P2_R2182_U90 P2_R2096_U91 ; P2_ADD_391_1196_U228
g24752 nand P2_ADD_391_1196_U228 P2_ADD_391_1196_U152 ; P2_ADD_391_1196_U229
g24753 nand P2_R2096_U91 P2_R2182_U90 ; P2_ADD_391_1196_U230
g24754 not P2_ADD_391_1196_U150 ; P2_ADD_391_1196_U231
g24755 or P2_R2182_U89 P2_R2096_U90 ; P2_ADD_391_1196_U232
g24756 nand P2_ADD_391_1196_U232 P2_ADD_391_1196_U150 ; P2_ADD_391_1196_U233
g24757 nand P2_R2096_U90 P2_R2182_U89 ; P2_ADD_391_1196_U234
g24758 not P2_ADD_391_1196_U148 ; P2_ADD_391_1196_U235
g24759 or P2_R2182_U88 P2_R2096_U89 ; P2_ADD_391_1196_U236
g24760 nand P2_ADD_391_1196_U236 P2_ADD_391_1196_U148 ; P2_ADD_391_1196_U237
g24761 nand P2_R2096_U89 P2_R2182_U88 ; P2_ADD_391_1196_U238
g24762 not P2_ADD_391_1196_U146 ; P2_ADD_391_1196_U239
g24763 or P2_R2182_U87 P2_R2096_U88 ; P2_ADD_391_1196_U240
g24764 nand P2_ADD_391_1196_U240 P2_ADD_391_1196_U146 ; P2_ADD_391_1196_U241
g24765 nand P2_R2096_U88 P2_R2182_U87 ; P2_ADD_391_1196_U242
g24766 not P2_ADD_391_1196_U142 ; P2_ADD_391_1196_U243
g24767 or P2_R2182_U86 P2_R2096_U87 ; P2_ADD_391_1196_U244
g24768 nand P2_ADD_391_1196_U244 P2_ADD_391_1196_U142 ; P2_ADD_391_1196_U245
g24769 nand P2_R2096_U87 P2_R2182_U86 ; P2_ADD_391_1196_U246
g24770 not P2_ADD_391_1196_U140 ; P2_ADD_391_1196_U247
g24771 or P2_R2182_U85 P2_R2096_U86 ; P2_ADD_391_1196_U248
g24772 nand P2_ADD_391_1196_U248 P2_ADD_391_1196_U140 ; P2_ADD_391_1196_U249
g24773 nand P2_R2096_U86 P2_R2182_U85 ; P2_ADD_391_1196_U250
g24774 not P2_ADD_391_1196_U138 ; P2_ADD_391_1196_U251
g24775 or P2_R2182_U84 P2_R2096_U85 ; P2_ADD_391_1196_U252
g24776 nand P2_ADD_391_1196_U252 P2_ADD_391_1196_U138 ; P2_ADD_391_1196_U253
g24777 nand P2_R2096_U85 P2_R2182_U84 ; P2_ADD_391_1196_U254
g24778 not P2_ADD_391_1196_U136 ; P2_ADD_391_1196_U255
g24779 or P2_R2182_U83 P2_R2096_U84 ; P2_ADD_391_1196_U256
g24780 nand P2_ADD_391_1196_U256 P2_ADD_391_1196_U136 ; P2_ADD_391_1196_U257
g24781 nand P2_R2096_U84 P2_R2182_U83 ; P2_ADD_391_1196_U258
g24782 not P2_ADD_391_1196_U134 ; P2_ADD_391_1196_U259
g24783 or P2_R2182_U82 P2_R2096_U83 ; P2_ADD_391_1196_U260
g24784 nand P2_ADD_391_1196_U260 P2_ADD_391_1196_U134 ; P2_ADD_391_1196_U261
g24785 nand P2_R2096_U83 P2_R2182_U82 ; P2_ADD_391_1196_U262
g24786 not P2_ADD_391_1196_U132 ; P2_ADD_391_1196_U263
g24787 or P2_R2182_U81 P2_R2096_U82 ; P2_ADD_391_1196_U264
g24788 nand P2_ADD_391_1196_U264 P2_ADD_391_1196_U132 ; P2_ADD_391_1196_U265
g24789 nand P2_R2096_U82 P2_R2182_U81 ; P2_ADD_391_1196_U266
g24790 not P2_ADD_391_1196_U130 ; P2_ADD_391_1196_U267
g24791 or P2_R2182_U80 P2_R2096_U81 ; P2_ADD_391_1196_U268
g24792 nand P2_ADD_391_1196_U268 P2_ADD_391_1196_U130 ; P2_ADD_391_1196_U269
g24793 nand P2_R2096_U81 P2_R2182_U80 ; P2_ADD_391_1196_U270
g24794 not P2_ADD_391_1196_U128 ; P2_ADD_391_1196_U271
g24795 or P2_R2182_U79 P2_R2096_U80 ; P2_ADD_391_1196_U272
g24796 nand P2_ADD_391_1196_U272 P2_ADD_391_1196_U128 ; P2_ADD_391_1196_U273
g24797 nand P2_R2096_U80 P2_R2182_U79 ; P2_ADD_391_1196_U274
g24798 not P2_ADD_391_1196_U126 ; P2_ADD_391_1196_U275
g24799 or P2_R2096_U79 P2_R2182_U78 ; P2_ADD_391_1196_U276
g24800 nand P2_ADD_391_1196_U276 P2_ADD_391_1196_U126 ; P2_ADD_391_1196_U277
g24801 nand P2_R2182_U78 P2_R2096_U79 ; P2_ADD_391_1196_U278
g24802 not P2_ADD_391_1196_U82 ; P2_ADD_391_1196_U279
g24803 or P2_R2096_U78 P2_R2182_U77 ; P2_ADD_391_1196_U280
g24804 nand P2_ADD_391_1196_U280 P2_ADD_391_1196_U82 ; P2_ADD_391_1196_U281
g24805 nand P2_R2182_U77 P2_R2096_U78 ; P2_ADD_391_1196_U282
g24806 nand P2_ADD_391_1196_U282 P2_ADD_391_1196_U281 P2_ADD_391_1196_U121 ; P2_ADD_391_1196_U283
g24807 nand P2_R2182_U77 P2_R2096_U78 ; P2_ADD_391_1196_U284
g24808 nand P2_ADD_391_1196_U279 P2_ADD_391_1196_U284 ; P2_ADD_391_1196_U285
g24809 or P2_R2182_U77 P2_R2096_U78 ; P2_ADD_391_1196_U286
g24810 nand P2_ADD_391_1196_U286 P2_ADD_391_1196_U285 P2_ADD_391_1196_U343 ; P2_ADD_391_1196_U287
g24811 or P2_R2182_U92 P2_R2096_U93 ; P2_ADD_391_1196_U288
g24812 nand P2_ADD_391_1196_U288 P2_ADD_391_1196_U53 ; P2_ADD_391_1196_U289
g24813 nand P2_ADD_391_1196_U289 P2_ADD_391_1196_U159 P2_ADD_391_1196_U153 ; P2_ADD_391_1196_U290
g24814 nand P2_R2096_U92 P2_R2182_U91 ; P2_ADD_391_1196_U291
g24815 nand P2_ADD_391_1196_U225 P2_ADD_391_1196_U291 ; P2_ADD_391_1196_U292
g24816 or P2_R2096_U93 P2_R2182_U92 ; P2_ADD_391_1196_U293
g24817 nand P2_ADD_391_1196_U154 P2_ADD_391_1196_U217 ; P2_ADD_391_1196_U294
g24818 nand P2_R2096_U94 P2_R2182_U93 ; P2_ADD_391_1196_U295
g24819 nand P2_ADD_391_1196_U219 P2_ADD_391_1196_U295 ; P2_ADD_391_1196_U296
g24820 or P2_R2182_U96 P2_R2096_U97 ; P2_ADD_391_1196_U297
g24821 nand P2_ADD_391_1196_U297 P2_ADD_391_1196_U50 ; P2_ADD_391_1196_U298
g24822 nand P2_ADD_391_1196_U298 P2_ADD_391_1196_U158 P2_ADD_391_1196_U157 ; P2_ADD_391_1196_U299
g24823 nand P2_R2096_U96 P2_R2182_U95 ; P2_ADD_391_1196_U300
g24824 nand P2_ADD_391_1196_U211 P2_ADD_391_1196_U300 ; P2_ADD_391_1196_U301
g24825 or P2_R2096_U97 P2_R2182_U96 ; P2_ADD_391_1196_U302
g24826 nand P2_ADD_391_1196_U202 P2_ADD_391_1196_U161 ; P2_ADD_391_1196_U303
g24827 nand P2_ADD_391_1196_U293 P2_ADD_391_1196_U159 ; P2_ADD_391_1196_U304
g24828 nand P2_ADD_391_1196_U302 P2_ADD_391_1196_U158 ; P2_ADD_391_1196_U305
g24829 nand P2_ADD_391_1196_U423 P2_ADD_391_1196_U23 ; P2_ADD_391_1196_U306
g24830 nand P2_R2096_U69 P2_ADD_391_1196_U34 ; P2_ADD_391_1196_U307
g24831 nand P2_R2182_U70 P2_ADD_391_1196_U33 ; P2_ADD_391_1196_U308
g24832 nand P2_R2096_U70 P2_ADD_391_1196_U31 ; P2_ADD_391_1196_U309
g24833 nand P2_R2182_U71 P2_ADD_391_1196_U32 ; P2_ADD_391_1196_U310
g24834 nand P2_R2096_U70 P2_ADD_391_1196_U31 ; P2_ADD_391_1196_U311
g24835 nand P2_R2182_U71 P2_ADD_391_1196_U32 ; P2_ADD_391_1196_U312
g24836 nand P2_ADD_391_1196_U312 P2_ADD_391_1196_U311 ; P2_ADD_391_1196_U313
g24837 nand P2_ADD_391_1196_U111 P2_ADD_391_1196_U112 ; P2_ADD_391_1196_U314
g24838 nand P2_ADD_391_1196_U187 P2_ADD_391_1196_U313 ; P2_ADD_391_1196_U315
g24839 nand P2_R2096_U71 P2_ADD_391_1196_U13 ; P2_ADD_391_1196_U316
g24840 nand P2_R2182_U72 P2_ADD_391_1196_U14 ; P2_ADD_391_1196_U317
g24841 nand P2_R2096_U72 P2_ADD_391_1196_U15 ; P2_ADD_391_1196_U318
g24842 nand P2_R2182_U73 P2_ADD_391_1196_U16 ; P2_ADD_391_1196_U319
g24843 nand P2_ADD_391_1196_U319 P2_ADD_391_1196_U318 ; P2_ADD_391_1196_U320
g24844 nand P2_ADD_391_1196_U303 P2_ADD_391_1196_U30 ; P2_ADD_391_1196_U321
g24845 nand P2_ADD_391_1196_U320 P2_ADD_391_1196_U181 ; P2_ADD_391_1196_U322
g24846 nand P2_R2096_U73 P2_ADD_391_1196_U17 ; P2_ADD_391_1196_U323
g24847 nand P2_R2182_U74 P2_ADD_391_1196_U18 ; P2_ADD_391_1196_U324
g24848 nand P2_R2096_U74 P2_ADD_391_1196_U28 ; P2_ADD_391_1196_U325
g24849 nand P2_R2182_U75 P2_ADD_391_1196_U29 ; P2_ADD_391_1196_U326
g24850 nand P2_R2096_U74 P2_ADD_391_1196_U28 ; P2_ADD_391_1196_U327
g24851 nand P2_R2182_U75 P2_ADD_391_1196_U29 ; P2_ADD_391_1196_U328
g24852 nand P2_ADD_391_1196_U328 P2_ADD_391_1196_U327 ; P2_ADD_391_1196_U329
g24853 nand P2_ADD_391_1196_U115 P2_ADD_391_1196_U116 ; P2_ADD_391_1196_U330
g24854 nand P2_ADD_391_1196_U173 P2_ADD_391_1196_U329 ; P2_ADD_391_1196_U331
g24855 nand P2_R2096_U75 P2_ADD_391_1196_U26 ; P2_ADD_391_1196_U332
g24856 nand P2_R2182_U76 P2_ADD_391_1196_U27 ; P2_ADD_391_1196_U333
g24857 nand P2_R2096_U75 P2_ADD_391_1196_U26 ; P2_ADD_391_1196_U334
g24858 nand P2_R2182_U76 P2_ADD_391_1196_U27 ; P2_ADD_391_1196_U335
g24859 nand P2_ADD_391_1196_U335 P2_ADD_391_1196_U334 ; P2_ADD_391_1196_U336
g24860 nand P2_ADD_391_1196_U117 P2_ADD_391_1196_U118 ; P2_ADD_391_1196_U337
g24861 nand P2_ADD_391_1196_U169 P2_ADD_391_1196_U336 ; P2_ADD_391_1196_U338
g24862 nand P2_R2182_U41 P2_ADD_391_1196_U120 ; P2_ADD_391_1196_U339
g24863 nand P2_R2096_U76 P2_ADD_391_1196_U119 ; P2_ADD_391_1196_U340
g24864 nand P2_R2182_U41 P2_ADD_391_1196_U120 ; P2_ADD_391_1196_U341
g24865 nand P2_R2096_U76 P2_ADD_391_1196_U119 ; P2_ADD_391_1196_U342
g24866 nand P2_ADD_391_1196_U342 P2_ADD_391_1196_U341 ; P2_ADD_391_1196_U343
g24867 nand P2_R2096_U77 P2_ADD_391_1196_U24 ; P2_ADD_391_1196_U344
g24868 nand P2_R2182_U40 P2_ADD_391_1196_U25 ; P2_ADD_391_1196_U345
g24869 nand P2_R2096_U77 P2_ADD_391_1196_U24 ; P2_ADD_391_1196_U346
g24870 nand P2_R2182_U40 P2_ADD_391_1196_U25 ; P2_ADD_391_1196_U347
g24871 nand P2_ADD_391_1196_U347 P2_ADD_391_1196_U346 ; P2_ADD_391_1196_U348
g24872 nand P2_ADD_391_1196_U122 P2_ADD_391_1196_U123 ; P2_ADD_391_1196_U349
g24873 nand P2_ADD_391_1196_U165 P2_ADD_391_1196_U348 ; P2_ADD_391_1196_U350
g24874 nand P2_R2182_U77 P2_ADD_391_1196_U80 ; P2_ADD_391_1196_U351
g24875 nand P2_R2096_U78 P2_ADD_391_1196_U81 ; P2_ADD_391_1196_U352
g24876 nand P2_R2182_U77 P2_ADD_391_1196_U80 ; P2_ADD_391_1196_U353
g24877 nand P2_R2096_U78 P2_ADD_391_1196_U81 ; P2_ADD_391_1196_U354
g24878 nand P2_ADD_391_1196_U354 P2_ADD_391_1196_U353 ; P2_ADD_391_1196_U355
g24879 nand P2_ADD_391_1196_U124 P2_ADD_391_1196_U82 ; P2_ADD_391_1196_U356
g24880 nand P2_ADD_391_1196_U355 P2_ADD_391_1196_U279 ; P2_ADD_391_1196_U357
g24881 nand P2_R2182_U78 P2_ADD_391_1196_U78 ; P2_ADD_391_1196_U358
g24882 nand P2_R2096_U79 P2_ADD_391_1196_U79 ; P2_ADD_391_1196_U359
g24883 nand P2_R2182_U78 P2_ADD_391_1196_U78 ; P2_ADD_391_1196_U360
g24884 nand P2_R2096_U79 P2_ADD_391_1196_U79 ; P2_ADD_391_1196_U361
g24885 nand P2_ADD_391_1196_U361 P2_ADD_391_1196_U360 ; P2_ADD_391_1196_U362
g24886 nand P2_ADD_391_1196_U125 P2_ADD_391_1196_U126 ; P2_ADD_391_1196_U363
g24887 nand P2_ADD_391_1196_U275 P2_ADD_391_1196_U362 ; P2_ADD_391_1196_U364
g24888 nand P2_R2096_U80 P2_ADD_391_1196_U76 ; P2_ADD_391_1196_U365
g24889 nand P2_R2182_U79 P2_ADD_391_1196_U77 ; P2_ADD_391_1196_U366
g24890 nand P2_R2096_U80 P2_ADD_391_1196_U76 ; P2_ADD_391_1196_U367
g24891 nand P2_R2182_U79 P2_ADD_391_1196_U77 ; P2_ADD_391_1196_U368
g24892 nand P2_ADD_391_1196_U368 P2_ADD_391_1196_U367 ; P2_ADD_391_1196_U369
g24893 nand P2_ADD_391_1196_U127 P2_ADD_391_1196_U128 ; P2_ADD_391_1196_U370
g24894 nand P2_ADD_391_1196_U271 P2_ADD_391_1196_U369 ; P2_ADD_391_1196_U371
g24895 nand P2_R2096_U81 P2_ADD_391_1196_U74 ; P2_ADD_391_1196_U372
g24896 nand P2_R2182_U80 P2_ADD_391_1196_U75 ; P2_ADD_391_1196_U373
g24897 nand P2_R2096_U81 P2_ADD_391_1196_U74 ; P2_ADD_391_1196_U374
g24898 nand P2_R2182_U80 P2_ADD_391_1196_U75 ; P2_ADD_391_1196_U375
g24899 nand P2_ADD_391_1196_U375 P2_ADD_391_1196_U374 ; P2_ADD_391_1196_U376
g24900 nand P2_ADD_391_1196_U129 P2_ADD_391_1196_U130 ; P2_ADD_391_1196_U377
g24901 nand P2_ADD_391_1196_U267 P2_ADD_391_1196_U376 ; P2_ADD_391_1196_U378
g24902 nand P2_R2096_U82 P2_ADD_391_1196_U72 ; P2_ADD_391_1196_U379
g24903 nand P2_R2182_U81 P2_ADD_391_1196_U73 ; P2_ADD_391_1196_U380
g24904 nand P2_R2096_U82 P2_ADD_391_1196_U72 ; P2_ADD_391_1196_U381
g24905 nand P2_R2182_U81 P2_ADD_391_1196_U73 ; P2_ADD_391_1196_U382
g24906 nand P2_ADD_391_1196_U382 P2_ADD_391_1196_U381 ; P2_ADD_391_1196_U383
g24907 nand P2_ADD_391_1196_U131 P2_ADD_391_1196_U132 ; P2_ADD_391_1196_U384
g24908 nand P2_ADD_391_1196_U263 P2_ADD_391_1196_U383 ; P2_ADD_391_1196_U385
g24909 nand P2_R2096_U83 P2_ADD_391_1196_U70 ; P2_ADD_391_1196_U386
g24910 nand P2_R2182_U82 P2_ADD_391_1196_U71 ; P2_ADD_391_1196_U387
g24911 nand P2_R2096_U83 P2_ADD_391_1196_U70 ; P2_ADD_391_1196_U388
g24912 nand P2_R2182_U82 P2_ADD_391_1196_U71 ; P2_ADD_391_1196_U389
g24913 nand P2_ADD_391_1196_U389 P2_ADD_391_1196_U388 ; P2_ADD_391_1196_U390
g24914 nand P2_ADD_391_1196_U133 P2_ADD_391_1196_U134 ; P2_ADD_391_1196_U391
g24915 nand P2_ADD_391_1196_U259 P2_ADD_391_1196_U390 ; P2_ADD_391_1196_U392
g24916 nand P2_R2096_U84 P2_ADD_391_1196_U68 ; P2_ADD_391_1196_U393
g24917 nand P2_R2182_U83 P2_ADD_391_1196_U69 ; P2_ADD_391_1196_U394
g24918 nand P2_R2096_U84 P2_ADD_391_1196_U68 ; P2_ADD_391_1196_U395
g24919 nand P2_R2182_U83 P2_ADD_391_1196_U69 ; P2_ADD_391_1196_U396
g24920 nand P2_ADD_391_1196_U396 P2_ADD_391_1196_U395 ; P2_ADD_391_1196_U397
g24921 nand P2_ADD_391_1196_U135 P2_ADD_391_1196_U136 ; P2_ADD_391_1196_U398
g24922 nand P2_ADD_391_1196_U255 P2_ADD_391_1196_U397 ; P2_ADD_391_1196_U399
g24923 nand P2_R2096_U85 P2_ADD_391_1196_U66 ; P2_ADD_391_1196_U400
g24924 nand P2_R2182_U84 P2_ADD_391_1196_U67 ; P2_ADD_391_1196_U401
g24925 nand P2_R2096_U85 P2_ADD_391_1196_U66 ; P2_ADD_391_1196_U402
g24926 nand P2_R2182_U84 P2_ADD_391_1196_U67 ; P2_ADD_391_1196_U403
g24927 nand P2_ADD_391_1196_U403 P2_ADD_391_1196_U402 ; P2_ADD_391_1196_U404
g24928 nand P2_ADD_391_1196_U137 P2_ADD_391_1196_U138 ; P2_ADD_391_1196_U405
g24929 nand P2_ADD_391_1196_U251 P2_ADD_391_1196_U404 ; P2_ADD_391_1196_U406
g24930 nand P2_R2096_U86 P2_ADD_391_1196_U64 ; P2_ADD_391_1196_U407
g24931 nand P2_R2182_U85 P2_ADD_391_1196_U65 ; P2_ADD_391_1196_U408
g24932 nand P2_R2096_U86 P2_ADD_391_1196_U64 ; P2_ADD_391_1196_U409
g24933 nand P2_R2182_U85 P2_ADD_391_1196_U65 ; P2_ADD_391_1196_U410
g24934 nand P2_ADD_391_1196_U410 P2_ADD_391_1196_U409 ; P2_ADD_391_1196_U411
g24935 nand P2_ADD_391_1196_U139 P2_ADD_391_1196_U140 ; P2_ADD_391_1196_U412
g24936 nand P2_ADD_391_1196_U247 P2_ADD_391_1196_U411 ; P2_ADD_391_1196_U413
g24937 nand P2_R2096_U87 P2_ADD_391_1196_U62 ; P2_ADD_391_1196_U414
g24938 nand P2_R2182_U86 P2_ADD_391_1196_U63 ; P2_ADD_391_1196_U415
g24939 nand P2_R2096_U87 P2_ADD_391_1196_U62 ; P2_ADD_391_1196_U416
g24940 nand P2_R2182_U86 P2_ADD_391_1196_U63 ; P2_ADD_391_1196_U417
g24941 nand P2_ADD_391_1196_U417 P2_ADD_391_1196_U416 ; P2_ADD_391_1196_U418
g24942 nand P2_ADD_391_1196_U141 P2_ADD_391_1196_U142 ; P2_ADD_391_1196_U419
g24943 nand P2_ADD_391_1196_U243 P2_ADD_391_1196_U418 ; P2_ADD_391_1196_U420
g24944 nand P2_R2182_U68 P2_ADD_391_1196_U22 ; P2_ADD_391_1196_U421
g24945 nand P2_ADD_391_1196_U162 P2_ADD_391_1196_U21 ; P2_ADD_391_1196_U422
g24946 nand P2_ADD_391_1196_U422 P2_ADD_391_1196_U421 ; P2_ADD_391_1196_U423
g24947 nand P2_R2096_U51 P2_ADD_391_1196_U22 P2_ADD_391_1196_U21 ; P2_ADD_391_1196_U424
g24948 nand P2_ADD_391_1196_U160 P2_R2182_U68 ; P2_ADD_391_1196_U425
g24949 nand P2_R2096_U88 P2_ADD_391_1196_U60 ; P2_ADD_391_1196_U426
g24950 nand P2_R2182_U87 P2_ADD_391_1196_U61 ; P2_ADD_391_1196_U427
g24951 nand P2_R2096_U88 P2_ADD_391_1196_U60 ; P2_ADD_391_1196_U428
g24952 nand P2_R2182_U87 P2_ADD_391_1196_U61 ; P2_ADD_391_1196_U429
g24953 nand P2_ADD_391_1196_U429 P2_ADD_391_1196_U428 ; P2_ADD_391_1196_U430
g24954 nand P2_ADD_391_1196_U145 P2_ADD_391_1196_U146 ; P2_ADD_391_1196_U431
g24955 nand P2_ADD_391_1196_U239 P2_ADD_391_1196_U430 ; P2_ADD_391_1196_U432
g24956 nand P2_R2096_U89 P2_ADD_391_1196_U58 ; P2_ADD_391_1196_U433
g24957 nand P2_R2182_U88 P2_ADD_391_1196_U59 ; P2_ADD_391_1196_U434
g24958 nand P2_R2096_U89 P2_ADD_391_1196_U58 ; P2_ADD_391_1196_U435
g24959 nand P2_R2182_U88 P2_ADD_391_1196_U59 ; P2_ADD_391_1196_U436
g24960 nand P2_ADD_391_1196_U436 P2_ADD_391_1196_U435 ; P2_ADD_391_1196_U437
g24961 nand P2_ADD_391_1196_U147 P2_ADD_391_1196_U148 ; P2_ADD_391_1196_U438
g24962 nand P2_ADD_391_1196_U235 P2_ADD_391_1196_U437 ; P2_ADD_391_1196_U439
g24963 nand P2_R2096_U90 P2_ADD_391_1196_U56 ; P2_ADD_391_1196_U440
g24964 nand P2_R2182_U89 P2_ADD_391_1196_U57 ; P2_ADD_391_1196_U441
g24965 nand P2_R2096_U90 P2_ADD_391_1196_U56 ; P2_ADD_391_1196_U442
g24966 nand P2_R2182_U89 P2_ADD_391_1196_U57 ; P2_ADD_391_1196_U443
g24967 nand P2_ADD_391_1196_U443 P2_ADD_391_1196_U442 ; P2_ADD_391_1196_U444
g24968 nand P2_ADD_391_1196_U149 P2_ADD_391_1196_U150 ; P2_ADD_391_1196_U445
g24969 nand P2_ADD_391_1196_U231 P2_ADD_391_1196_U444 ; P2_ADD_391_1196_U446
g24970 nand P2_R2096_U91 P2_ADD_391_1196_U54 ; P2_ADD_391_1196_U447
g24971 nand P2_R2182_U90 P2_ADD_391_1196_U55 ; P2_ADD_391_1196_U448
g24972 nand P2_R2096_U91 P2_ADD_391_1196_U54 ; P2_ADD_391_1196_U449
g24973 nand P2_R2182_U90 P2_ADD_391_1196_U55 ; P2_ADD_391_1196_U450
g24974 nand P2_ADD_391_1196_U450 P2_ADD_391_1196_U449 ; P2_ADD_391_1196_U451
g24975 nand P2_ADD_391_1196_U151 P2_ADD_391_1196_U152 ; P2_ADD_391_1196_U452
g24976 nand P2_ADD_391_1196_U227 P2_ADD_391_1196_U451 ; P2_ADD_391_1196_U453
g24977 nand P2_R2096_U92 P2_ADD_391_1196_U40 ; P2_ADD_391_1196_U454
g24978 nand P2_R2182_U91 P2_ADD_391_1196_U41 ; P2_ADD_391_1196_U455
g24979 nand P2_R2096_U93 P2_ADD_391_1196_U42 ; P2_ADD_391_1196_U456
g24980 nand P2_R2182_U92 P2_ADD_391_1196_U43 ; P2_ADD_391_1196_U457
g24981 nand P2_ADD_391_1196_U457 P2_ADD_391_1196_U456 ; P2_ADD_391_1196_U458
g24982 nand P2_ADD_391_1196_U304 P2_ADD_391_1196_U53 ; P2_ADD_391_1196_U459
g24983 nand P2_ADD_391_1196_U458 P2_ADD_391_1196_U221 ; P2_ADD_391_1196_U460
g24984 nand P2_R2096_U94 P2_ADD_391_1196_U44 ; P2_ADD_391_1196_U461
g24985 nand P2_R2182_U93 P2_ADD_391_1196_U45 ; P2_ADD_391_1196_U462
g24986 nand P2_R2096_U95 P2_ADD_391_1196_U51 ; P2_ADD_391_1196_U463
g24987 nand P2_R2182_U94 P2_ADD_391_1196_U52 ; P2_ADD_391_1196_U464
g24988 nand P2_R2096_U95 P2_ADD_391_1196_U51 ; P2_ADD_391_1196_U465
g24989 nand P2_R2182_U94 P2_ADD_391_1196_U52 ; P2_ADD_391_1196_U466
g24990 nand P2_ADD_391_1196_U466 P2_ADD_391_1196_U465 ; P2_ADD_391_1196_U467
g24991 nand P2_ADD_391_1196_U155 P2_ADD_391_1196_U156 ; P2_ADD_391_1196_U468
g24992 nand P2_ADD_391_1196_U213 P2_ADD_391_1196_U467 ; P2_ADD_391_1196_U469
g24993 nand P2_R2096_U96 P2_ADD_391_1196_U46 ; P2_ADD_391_1196_U470
g24994 nand P2_R2182_U95 P2_ADD_391_1196_U47 ; P2_ADD_391_1196_U471
g24995 nand P2_R2096_U97 P2_ADD_391_1196_U48 ; P2_ADD_391_1196_U472
g24996 nand P2_R2182_U96 P2_ADD_391_1196_U49 ; P2_ADD_391_1196_U473
g24997 nand P2_ADD_391_1196_U473 P2_ADD_391_1196_U472 ; P2_ADD_391_1196_U474
g24998 nand P2_ADD_391_1196_U305 P2_ADD_391_1196_U50 ; P2_ADD_391_1196_U475
g24999 nand P2_ADD_391_1196_U474 P2_ADD_391_1196_U207 ; P2_ADD_391_1196_U476
g25000 nand P2_R2182_U69 P2_ADD_391_1196_U19 ; P2_ADD_391_1196_U477
g25001 nand P2_R2096_U68 P2_ADD_391_1196_U20 ; P2_ADD_391_1196_U478
g25002 not P2_U2606 ; P2_ADD_402_1132_U4
g25003 not P2_U2591 ; P2_ADD_402_1132_U5
g25004 nand P2_U2591 P2_U2606 ; P2_ADD_402_1132_U6
g25005 not P2_U2592 ; P2_ADD_402_1132_U7
g25006 nand P2_U2592 P2_ADD_402_1132_U28 ; P2_ADD_402_1132_U8
g25007 not P2_U2593 ; P2_ADD_402_1132_U9
g25008 nand P2_U2593 P2_ADD_402_1132_U29 ; P2_ADD_402_1132_U10
g25009 not P2_U2594 ; P2_ADD_402_1132_U11
g25010 nand P2_U2594 P2_ADD_402_1132_U30 ; P2_ADD_402_1132_U12
g25011 not P2_U2595 ; P2_ADD_402_1132_U13
g25012 nand P2_U2595 P2_ADD_402_1132_U31 ; P2_ADD_402_1132_U14
g25013 not P2_U2596 ; P2_ADD_402_1132_U15
g25014 nand P2_U2596 P2_ADD_402_1132_U32 ; P2_ADD_402_1132_U16
g25015 not P2_U2597 ; P2_ADD_402_1132_U17
g25016 nand P2_ADD_402_1132_U36 P2_ADD_402_1132_U35 ; P2_ADD_402_1132_U18
g25017 nand P2_ADD_402_1132_U38 P2_ADD_402_1132_U37 ; P2_ADD_402_1132_U19
g25018 nand P2_ADD_402_1132_U40 P2_ADD_402_1132_U39 ; P2_ADD_402_1132_U20
g25019 nand P2_ADD_402_1132_U42 P2_ADD_402_1132_U41 ; P2_ADD_402_1132_U21
g25020 nand P2_ADD_402_1132_U44 P2_ADD_402_1132_U43 ; P2_ADD_402_1132_U22
g25021 nand P2_ADD_402_1132_U46 P2_ADD_402_1132_U45 ; P2_ADD_402_1132_U23
g25022 nand P2_ADD_402_1132_U48 P2_ADD_402_1132_U47 ; P2_ADD_402_1132_U24
g25023 nand P2_ADD_402_1132_U50 P2_ADD_402_1132_U49 ; P2_ADD_402_1132_U25
g25024 not P2_U2598 ; P2_ADD_402_1132_U26
g25025 nand P2_U2597 P2_ADD_402_1132_U33 ; P2_ADD_402_1132_U27
g25026 not P2_ADD_402_1132_U6 ; P2_ADD_402_1132_U28
g25027 not P2_ADD_402_1132_U8 ; P2_ADD_402_1132_U29
g25028 not P2_ADD_402_1132_U10 ; P2_ADD_402_1132_U30
g25029 not P2_ADD_402_1132_U12 ; P2_ADD_402_1132_U31
g25030 not P2_ADD_402_1132_U14 ; P2_ADD_402_1132_U32
g25031 not P2_ADD_402_1132_U16 ; P2_ADD_402_1132_U33
g25032 not P2_ADD_402_1132_U27 ; P2_ADD_402_1132_U34
g25033 nand P2_U2598 P2_ADD_402_1132_U27 ; P2_ADD_402_1132_U35
g25034 nand P2_ADD_402_1132_U34 P2_ADD_402_1132_U26 ; P2_ADD_402_1132_U36
g25035 nand P2_U2597 P2_ADD_402_1132_U16 ; P2_ADD_402_1132_U37
g25036 nand P2_ADD_402_1132_U33 P2_ADD_402_1132_U17 ; P2_ADD_402_1132_U38
g25037 nand P2_U2592 P2_ADD_402_1132_U6 ; P2_ADD_402_1132_U39
g25038 nand P2_ADD_402_1132_U28 P2_ADD_402_1132_U7 ; P2_ADD_402_1132_U40
g25039 nand P2_U2594 P2_ADD_402_1132_U10 ; P2_ADD_402_1132_U41
g25040 nand P2_ADD_402_1132_U30 P2_ADD_402_1132_U11 ; P2_ADD_402_1132_U42
g25041 nand P2_U2595 P2_ADD_402_1132_U12 ; P2_ADD_402_1132_U43
g25042 nand P2_ADD_402_1132_U31 P2_ADD_402_1132_U13 ; P2_ADD_402_1132_U44
g25043 nand P2_U2591 P2_ADD_402_1132_U4 ; P2_ADD_402_1132_U45
g25044 nand P2_U2606 P2_ADD_402_1132_U5 ; P2_ADD_402_1132_U46
g25045 nand P2_U2596 P2_ADD_402_1132_U14 ; P2_ADD_402_1132_U47
g25046 nand P2_ADD_402_1132_U32 P2_ADD_402_1132_U15 ; P2_ADD_402_1132_U48
g25047 nand P2_U2593 P2_ADD_402_1132_U8 ; P2_ADD_402_1132_U49
g25048 nand P2_ADD_402_1132_U29 P2_ADD_402_1132_U9 ; P2_ADD_402_1132_U50
g25049 not P2_U3618 ; P2_SUB_563_U6
g25050 not P2_U3619 ; P2_SUB_563_U7
g25051 and P2_U2671 P2_R2182_U20 ; P2_R2182_U4
g25052 and P2_U2670 P2_R2182_U4 ; P2_R2182_U5
g25053 and P2_U2669 P2_R2182_U5 ; P2_R2182_U6
g25054 and P2_U2690 P2_R2182_U8 ; P2_R2182_U7
g25055 and P2_U2691 P2_R2182_U11 ; P2_R2182_U8
g25056 and P2_U2675 P2_R2182_U21 ; P2_R2182_U9
g25057 and P2_U2674 P2_R2182_U9 ; P2_R2182_U10
g25058 and P2_U2692 P2_R2182_U13 ; P2_R2182_U11
g25059 and P2_U2694 P2_R2182_U18 ; P2_R2182_U12
g25060 and P2_U2693 P2_R2182_U12 ; P2_R2182_U13
g25061 and P2_U2668 P2_R2182_U6 ; P2_R2182_U14
g25062 and P2_U2667 P2_R2182_U14 ; P2_R2182_U15
g25063 and P2_U2666 P2_R2182_U15 ; P2_R2182_U16
g25064 and P2_U2696 P2_R2182_U16 ; P2_R2182_U17
g25065 and P2_U2695 P2_R2182_U17 ; P2_R2182_U18
g25066 and P2_U2673 P2_R2182_U10 ; P2_R2182_U19
g25067 and P2_U2672 P2_R2182_U19 ; P2_R2182_U20
g25068 and P2_U2676 P2_R2182_U102 ; P2_R2182_U21
g25069 not P2_U2675 ; P2_R2182_U22
g25070 not P2_U2671 ; P2_R2182_U23
g25071 not P2_U2676 ; P2_R2182_U24
g25072 not P2_U2666 ; P2_R2182_U25
g25073 not P2_U2667 ; P2_R2182_U26
g25074 not P2_U2696 ; P2_R2182_U27
g25075 not P2_U2695 ; P2_R2182_U28
g25076 not P2_U2694 ; P2_R2182_U29
g25077 not P2_U2693 ; P2_R2182_U30
g25078 not P2_U2692 ; P2_R2182_U31
g25079 not P2_U2691 ; P2_R2182_U32
g25080 not P2_U2670 ; P2_R2182_U33
g25081 not P2_U2672 ; P2_R2182_U34
g25082 not P2_U2674 ; P2_R2182_U35
g25083 not P2_U2673 ; P2_R2182_U36
g25084 not P2_U2690 ; P2_R2182_U37
g25085 not P2_U2668 ; P2_R2182_U38
g25086 not P2_U2669 ; P2_R2182_U39
g25087 and P2_R2182_U192 P2_R2182_U190 ; P2_R2182_U40
g25088 and P2_R2182_U186 P2_R2182_U182 ; P2_R2182_U41
g25089 not P2_U2700 ; P2_R2182_U42
g25090 not P2_U2679 ; P2_R2182_U43
g25091 not P2_U2702 ; P2_R2182_U44
g25092 not P2_U2681 ; P2_R2182_U45
g25093 nand P2_U2681 P2_U2702 ; P2_R2182_U46
g25094 not P2_U2680 ; P2_R2182_U47
g25095 not P2_U2699 ; P2_R2182_U48
g25096 not P2_U2678 ; P2_R2182_U49
g25097 not P2_U2698 ; P2_R2182_U50
g25098 not P2_U2677 ; P2_R2182_U51
g25099 not P2_U2689 ; P2_R2182_U52
g25100 not P2_U2665 ; P2_R2182_U53
g25101 not P2_U2688 ; P2_R2182_U54
g25102 not P2_U2664 ; P2_R2182_U55
g25103 not P2_U2687 ; P2_R2182_U56
g25104 not P2_U2663 ; P2_R2182_U57
g25105 not P2_U2686 ; P2_R2182_U58
g25106 not P2_U2662 ; P2_R2182_U59
g25107 not P2_U2685 ; P2_R2182_U60
g25108 not P2_U2661 ; P2_R2182_U61
g25109 not P2_U2684 ; P2_R2182_U62
g25110 not P2_U2660 ; P2_R2182_U63
g25111 not P2_U2683 ; P2_R2182_U64
g25112 not P2_U2659 ; P2_R2182_U65
g25113 nand P2_R2182_U177 P2_R2182_U176 ; P2_R2182_U66
g25114 not P2_U2701 ; P2_R2182_U67
g25115 nand P2_R2182_U283 P2_R2182_U282 ; P2_R2182_U68
g25116 nand P2_R2182_U305 P2_R2182_U304 ; P2_R2182_U69
g25117 nand P2_R2182_U194 P2_R2182_U193 ; P2_R2182_U70
g25118 nand P2_R2182_U196 P2_R2182_U195 ; P2_R2182_U71
g25119 nand P2_R2182_U198 P2_R2182_U197 ; P2_R2182_U72
g25120 nand P2_R2182_U200 P2_R2182_U199 ; P2_R2182_U73
g25121 nand P2_R2182_U202 P2_R2182_U201 ; P2_R2182_U74
g25122 nand P2_R2182_U209 P2_R2182_U208 ; P2_R2182_U75
g25123 nand P2_R2182_U216 P2_R2182_U215 ; P2_R2182_U76
g25124 nand P2_R2182_U230 P2_R2182_U229 ; P2_R2182_U77
g25125 nand P2_R2182_U237 P2_R2182_U236 ; P2_R2182_U78
g25126 nand P2_R2182_U244 P2_R2182_U243 ; P2_R2182_U79
g25127 nand P2_R2182_U251 P2_R2182_U250 ; P2_R2182_U80
g25128 nand P2_R2182_U258 P2_R2182_U257 ; P2_R2182_U81
g25129 nand P2_R2182_U265 P2_R2182_U264 ; P2_R2182_U82
g25130 nand P2_R2182_U272 P2_R2182_U271 ; P2_R2182_U83
g25131 nand P2_R2182_U274 P2_R2182_U273 ; P2_R2182_U84
g25132 nand P2_R2182_U276 P2_R2182_U275 ; P2_R2182_U85
g25133 nand P2_R2182_U278 P2_R2182_U277 ; P2_R2182_U86
g25134 nand P2_R2182_U285 P2_R2182_U284 ; P2_R2182_U87
g25135 nand P2_R2182_U287 P2_R2182_U286 ; P2_R2182_U88
g25136 nand P2_R2182_U289 P2_R2182_U288 ; P2_R2182_U89
g25137 nand P2_R2182_U291 P2_R2182_U290 ; P2_R2182_U90
g25138 nand P2_R2182_U293 P2_R2182_U292 ; P2_R2182_U91
g25139 nand P2_R2182_U295 P2_R2182_U294 ; P2_R2182_U92
g25140 nand P2_R2182_U297 P2_R2182_U296 ; P2_R2182_U93
g25141 nand P2_R2182_U299 P2_R2182_U298 ; P2_R2182_U94
g25142 nand P2_R2182_U301 P2_R2182_U300 ; P2_R2182_U95
g25143 nand P2_R2182_U303 P2_R2182_U302 ; P2_R2182_U96
g25144 and P2_R2182_U218 P2_R2182_U217 P2_R2182_U181 ; P2_R2182_U97
g25145 and P2_R2182_U185 P2_R2182_U221 ; P2_R2182_U98
g25146 and P2_R2182_U223 P2_R2182_U222 P2_R2182_U189 ; P2_R2182_U99
g25147 and P2_R2182_U191 P2_R2182_U125 ; P2_R2182_U100
g25148 nand P2_R2182_U280 P2_R2182_U279 ; P2_R2182_U101
g25149 nand P2_R2182_U135 P2_R2182_U134 ; P2_R2182_U102
g25150 and P2_R2182_U204 P2_R2182_U203 ; P2_R2182_U103
g25151 nand P2_R2182_U131 P2_R2182_U130 ; P2_R2182_U104
g25152 and P2_R2182_U211 P2_R2182_U210 ; P2_R2182_U105
g25153 nand P2_R2182_U126 P2_R2182_U127 ; P2_R2182_U106
g25154 not P2_U2658 ; P2_R2182_U107
g25155 not P2_U2682 ; P2_R2182_U108
g25156 and P2_R2182_U225 P2_R2182_U224 ; P2_R2182_U109
g25157 and P2_R2182_U232 P2_R2182_U231 ; P2_R2182_U110
g25158 nand P2_R2182_U173 P2_R2182_U172 ; P2_R2182_U111
g25159 and P2_R2182_U239 P2_R2182_U238 ; P2_R2182_U112
g25160 nand P2_R2182_U169 P2_R2182_U168 ; P2_R2182_U113
g25161 and P2_R2182_U246 P2_R2182_U245 ; P2_R2182_U114
g25162 nand P2_R2182_U165 P2_R2182_U164 ; P2_R2182_U115
g25163 and P2_R2182_U253 P2_R2182_U252 ; P2_R2182_U116
g25164 nand P2_R2182_U161 P2_R2182_U160 ; P2_R2182_U117
g25165 and P2_R2182_U260 P2_R2182_U259 ; P2_R2182_U118
g25166 nand P2_R2182_U157 P2_R2182_U156 ; P2_R2182_U119
g25167 and P2_R2182_U267 P2_R2182_U266 ; P2_R2182_U120
g25168 not P2_R2182_U46 ; P2_R2182_U121
g25169 nand P2_U2680 P2_R2182_U121 ; P2_R2182_U122
g25170 nand P2_R2182_U122 P2_R2182_U67 ; P2_R2182_U123
g25171 or P2_U2679 P2_U2700 ; P2_R2182_U124
g25172 nand P2_R2182_U46 P2_R2182_U47 ; P2_R2182_U125
g25173 nand P2_R2182_U125 P2_R2182_U123 P2_R2182_U124 ; P2_R2182_U126
g25174 nand P2_U2679 P2_U2700 ; P2_R2182_U127
g25175 not P2_R2182_U106 ; P2_R2182_U128
g25176 or P2_U2699 P2_U2678 ; P2_R2182_U129
g25177 nand P2_R2182_U129 P2_R2182_U106 ; P2_R2182_U130
g25178 nand P2_U2678 P2_U2699 ; P2_R2182_U131
g25179 not P2_R2182_U104 ; P2_R2182_U132
g25180 or P2_U2698 P2_U2677 ; P2_R2182_U133
g25181 nand P2_R2182_U133 P2_R2182_U104 ; P2_R2182_U134
g25182 nand P2_U2677 P2_U2698 ; P2_R2182_U135
g25183 not P2_R2182_U102 ; P2_R2182_U136
g25184 not P2_R2182_U21 ; P2_R2182_U137
g25185 not P2_R2182_U9 ; P2_R2182_U138
g25186 not P2_R2182_U10 ; P2_R2182_U139
g25187 not P2_R2182_U19 ; P2_R2182_U140
g25188 not P2_R2182_U20 ; P2_R2182_U141
g25189 not P2_R2182_U4 ; P2_R2182_U142
g25190 not P2_R2182_U5 ; P2_R2182_U143
g25191 not P2_R2182_U6 ; P2_R2182_U144
g25192 not P2_R2182_U14 ; P2_R2182_U145
g25193 not P2_R2182_U15 ; P2_R2182_U146
g25194 not P2_R2182_U16 ; P2_R2182_U147
g25195 not P2_R2182_U17 ; P2_R2182_U148
g25196 not P2_R2182_U18 ; P2_R2182_U149
g25197 not P2_R2182_U12 ; P2_R2182_U150
g25198 not P2_R2182_U13 ; P2_R2182_U151
g25199 not P2_R2182_U11 ; P2_R2182_U152
g25200 not P2_R2182_U8 ; P2_R2182_U153
g25201 not P2_R2182_U7 ; P2_R2182_U154
g25202 or P2_U2689 P2_U2665 ; P2_R2182_U155
g25203 nand P2_R2182_U155 P2_R2182_U7 ; P2_R2182_U156
g25204 nand P2_U2665 P2_U2689 ; P2_R2182_U157
g25205 not P2_R2182_U119 ; P2_R2182_U158
g25206 or P2_U2688 P2_U2664 ; P2_R2182_U159
g25207 nand P2_R2182_U159 P2_R2182_U119 ; P2_R2182_U160
g25208 nand P2_U2664 P2_U2688 ; P2_R2182_U161
g25209 not P2_R2182_U117 ; P2_R2182_U162
g25210 or P2_U2687 P2_U2663 ; P2_R2182_U163
g25211 nand P2_R2182_U163 P2_R2182_U117 ; P2_R2182_U164
g25212 nand P2_U2663 P2_U2687 ; P2_R2182_U165
g25213 not P2_R2182_U115 ; P2_R2182_U166
g25214 or P2_U2686 P2_U2662 ; P2_R2182_U167
g25215 nand P2_R2182_U167 P2_R2182_U115 ; P2_R2182_U168
g25216 nand P2_U2662 P2_U2686 ; P2_R2182_U169
g25217 not P2_R2182_U113 ; P2_R2182_U170
g25218 or P2_U2685 P2_U2661 ; P2_R2182_U171
g25219 nand P2_R2182_U171 P2_R2182_U113 ; P2_R2182_U172
g25220 nand P2_U2661 P2_U2685 ; P2_R2182_U173
g25221 not P2_R2182_U111 ; P2_R2182_U174
g25222 or P2_U2684 P2_U2660 ; P2_R2182_U175
g25223 nand P2_R2182_U175 P2_R2182_U111 ; P2_R2182_U176
g25224 nand P2_U2660 P2_U2684 ; P2_R2182_U177
g25225 not P2_R2182_U66 ; P2_R2182_U178
g25226 or P2_U2683 P2_U2659 ; P2_R2182_U179
g25227 nand P2_R2182_U179 P2_R2182_U66 ; P2_R2182_U180
g25228 nand P2_U2659 P2_U2683 ; P2_R2182_U181
g25229 nand P2_R2182_U97 P2_R2182_U180 ; P2_R2182_U182
g25230 nand P2_U2659 P2_U2683 ; P2_R2182_U183
g25231 nand P2_R2182_U178 P2_R2182_U183 ; P2_R2182_U184
g25232 or P2_U2659 P2_U2683 ; P2_R2182_U185
g25233 nand P2_R2182_U98 P2_R2182_U184 ; P2_R2182_U186
g25234 nand P2_R2182_U47 P2_R2182_U46 ; P2_R2182_U187
g25235 nand P2_U2701 P2_R2182_U187 ; P2_R2182_U188
g25236 nand P2_U2680 P2_R2182_U121 ; P2_R2182_U189
g25237 nand P2_R2182_U99 P2_R2182_U188 ; P2_R2182_U190
g25238 nand P2_U2679 P2_U2700 ; P2_R2182_U191
g25239 nand P2_R2182_U124 P2_R2182_U123 P2_R2182_U100 ; P2_R2182_U192
g25240 nand P2_R2182_U34 P2_R2182_U19 ; P2_R2182_U193
g25241 nand P2_R2182_U140 P2_U2672 ; P2_R2182_U194
g25242 nand P2_R2182_U36 P2_R2182_U10 ; P2_R2182_U195
g25243 nand P2_R2182_U139 P2_U2673 ; P2_R2182_U196
g25244 nand P2_R2182_U35 P2_R2182_U9 ; P2_R2182_U197
g25245 nand P2_R2182_U138 P2_U2674 ; P2_R2182_U198
g25246 nand P2_R2182_U22 P2_R2182_U21 ; P2_R2182_U199
g25247 nand P2_R2182_U137 P2_U2675 ; P2_R2182_U200
g25248 nand P2_R2182_U24 P2_R2182_U102 ; P2_R2182_U201
g25249 nand P2_R2182_U136 P2_U2676 ; P2_R2182_U202
g25250 nand P2_U2677 P2_R2182_U50 ; P2_R2182_U203
g25251 nand P2_U2698 P2_R2182_U51 ; P2_R2182_U204
g25252 nand P2_U2677 P2_R2182_U50 ; P2_R2182_U205
g25253 nand P2_U2698 P2_R2182_U51 ; P2_R2182_U206
g25254 nand P2_R2182_U206 P2_R2182_U205 ; P2_R2182_U207
g25255 nand P2_R2182_U103 P2_R2182_U104 ; P2_R2182_U208
g25256 nand P2_R2182_U132 P2_R2182_U207 ; P2_R2182_U209
g25257 nand P2_U2678 P2_R2182_U48 ; P2_R2182_U210
g25258 nand P2_U2699 P2_R2182_U49 ; P2_R2182_U211
g25259 nand P2_U2678 P2_R2182_U48 ; P2_R2182_U212
g25260 nand P2_U2699 P2_R2182_U49 ; P2_R2182_U213
g25261 nand P2_R2182_U213 P2_R2182_U212 ; P2_R2182_U214
g25262 nand P2_R2182_U105 P2_R2182_U106 ; P2_R2182_U215
g25263 nand P2_R2182_U128 P2_R2182_U214 ; P2_R2182_U216
g25264 nand P2_U2658 P2_R2182_U108 ; P2_R2182_U217
g25265 nand P2_U2682 P2_R2182_U107 ; P2_R2182_U218
g25266 nand P2_U2658 P2_R2182_U108 ; P2_R2182_U219
g25267 nand P2_U2682 P2_R2182_U107 ; P2_R2182_U220
g25268 nand P2_R2182_U220 P2_R2182_U219 ; P2_R2182_U221
g25269 nand P2_U2679 P2_R2182_U42 ; P2_R2182_U222
g25270 nand P2_U2700 P2_R2182_U43 ; P2_R2182_U223
g25271 nand P2_U2659 P2_R2182_U64 ; P2_R2182_U224
g25272 nand P2_U2683 P2_R2182_U65 ; P2_R2182_U225
g25273 nand P2_U2659 P2_R2182_U64 ; P2_R2182_U226
g25274 nand P2_U2683 P2_R2182_U65 ; P2_R2182_U227
g25275 nand P2_R2182_U227 P2_R2182_U226 ; P2_R2182_U228
g25276 nand P2_R2182_U109 P2_R2182_U66 ; P2_R2182_U229
g25277 nand P2_R2182_U228 P2_R2182_U178 ; P2_R2182_U230
g25278 nand P2_U2660 P2_R2182_U62 ; P2_R2182_U231
g25279 nand P2_U2684 P2_R2182_U63 ; P2_R2182_U232
g25280 nand P2_U2660 P2_R2182_U62 ; P2_R2182_U233
g25281 nand P2_U2684 P2_R2182_U63 ; P2_R2182_U234
g25282 nand P2_R2182_U234 P2_R2182_U233 ; P2_R2182_U235
g25283 nand P2_R2182_U110 P2_R2182_U111 ; P2_R2182_U236
g25284 nand P2_R2182_U174 P2_R2182_U235 ; P2_R2182_U237
g25285 nand P2_U2661 P2_R2182_U60 ; P2_R2182_U238
g25286 nand P2_U2685 P2_R2182_U61 ; P2_R2182_U239
g25287 nand P2_U2661 P2_R2182_U60 ; P2_R2182_U240
g25288 nand P2_U2685 P2_R2182_U61 ; P2_R2182_U241
g25289 nand P2_R2182_U241 P2_R2182_U240 ; P2_R2182_U242
g25290 nand P2_R2182_U112 P2_R2182_U113 ; P2_R2182_U243
g25291 nand P2_R2182_U170 P2_R2182_U242 ; P2_R2182_U244
g25292 nand P2_U2662 P2_R2182_U58 ; P2_R2182_U245
g25293 nand P2_U2686 P2_R2182_U59 ; P2_R2182_U246
g25294 nand P2_U2662 P2_R2182_U58 ; P2_R2182_U247
g25295 nand P2_U2686 P2_R2182_U59 ; P2_R2182_U248
g25296 nand P2_R2182_U248 P2_R2182_U247 ; P2_R2182_U249
g25297 nand P2_R2182_U114 P2_R2182_U115 ; P2_R2182_U250
g25298 nand P2_R2182_U166 P2_R2182_U249 ; P2_R2182_U251
g25299 nand P2_U2663 P2_R2182_U56 ; P2_R2182_U252
g25300 nand P2_U2687 P2_R2182_U57 ; P2_R2182_U253
g25301 nand P2_U2663 P2_R2182_U56 ; P2_R2182_U254
g25302 nand P2_U2687 P2_R2182_U57 ; P2_R2182_U255
g25303 nand P2_R2182_U255 P2_R2182_U254 ; P2_R2182_U256
g25304 nand P2_R2182_U116 P2_R2182_U117 ; P2_R2182_U257
g25305 nand P2_R2182_U162 P2_R2182_U256 ; P2_R2182_U258
g25306 nand P2_U2664 P2_R2182_U54 ; P2_R2182_U259
g25307 nand P2_U2688 P2_R2182_U55 ; P2_R2182_U260
g25308 nand P2_U2664 P2_R2182_U54 ; P2_R2182_U261
g25309 nand P2_U2688 P2_R2182_U55 ; P2_R2182_U262
g25310 nand P2_R2182_U262 P2_R2182_U261 ; P2_R2182_U263
g25311 nand P2_R2182_U118 P2_R2182_U119 ; P2_R2182_U264
g25312 nand P2_R2182_U158 P2_R2182_U263 ; P2_R2182_U265
g25313 nand P2_U2665 P2_R2182_U52 ; P2_R2182_U266
g25314 nand P2_U2689 P2_R2182_U53 ; P2_R2182_U267
g25315 nand P2_U2665 P2_R2182_U52 ; P2_R2182_U268
g25316 nand P2_U2689 P2_R2182_U53 ; P2_R2182_U269
g25317 nand P2_R2182_U269 P2_R2182_U268 ; P2_R2182_U270
g25318 nand P2_R2182_U120 P2_R2182_U7 ; P2_R2182_U271
g25319 nand P2_R2182_U154 P2_R2182_U270 ; P2_R2182_U272
g25320 nand P2_R2182_U37 P2_R2182_U8 ; P2_R2182_U273
g25321 nand P2_R2182_U153 P2_U2690 ; P2_R2182_U274
g25322 nand P2_R2182_U32 P2_R2182_U11 ; P2_R2182_U275
g25323 nand P2_R2182_U152 P2_U2691 ; P2_R2182_U276
g25324 nand P2_R2182_U31 P2_R2182_U13 ; P2_R2182_U277
g25325 nand P2_R2182_U151 P2_U2692 ; P2_R2182_U278
g25326 nand P2_R2182_U121 P2_R2182_U47 ; P2_R2182_U279
g25327 nand P2_U2680 P2_R2182_U46 ; P2_R2182_U280
g25328 not P2_R2182_U101 ; P2_R2182_U281
g25329 nand P2_R2182_U281 P2_U2701 ; P2_R2182_U282
g25330 nand P2_R2182_U101 P2_R2182_U67 ; P2_R2182_U283
g25331 nand P2_R2182_U30 P2_R2182_U12 ; P2_R2182_U284
g25332 nand P2_R2182_U150 P2_U2693 ; P2_R2182_U285
g25333 nand P2_R2182_U29 P2_R2182_U18 ; P2_R2182_U286
g25334 nand P2_R2182_U149 P2_U2694 ; P2_R2182_U287
g25335 nand P2_R2182_U28 P2_R2182_U17 ; P2_R2182_U288
g25336 nand P2_R2182_U148 P2_U2695 ; P2_R2182_U289
g25337 nand P2_R2182_U27 P2_R2182_U16 ; P2_R2182_U290
g25338 nand P2_R2182_U147 P2_U2696 ; P2_R2182_U291
g25339 nand P2_R2182_U25 P2_R2182_U15 ; P2_R2182_U292
g25340 nand P2_R2182_U146 P2_U2666 ; P2_R2182_U293
g25341 nand P2_R2182_U26 P2_R2182_U14 ; P2_R2182_U294
g25342 nand P2_R2182_U145 P2_U2667 ; P2_R2182_U295
g25343 nand P2_R2182_U38 P2_R2182_U6 ; P2_R2182_U296
g25344 nand P2_R2182_U144 P2_U2668 ; P2_R2182_U297
g25345 nand P2_R2182_U39 P2_R2182_U5 ; P2_R2182_U298
g25346 nand P2_R2182_U143 P2_U2669 ; P2_R2182_U299
g25347 nand P2_R2182_U33 P2_R2182_U4 ; P2_R2182_U300
g25348 nand P2_R2182_U142 P2_U2670 ; P2_R2182_U301
g25349 nand P2_R2182_U23 P2_R2182_U20 ; P2_R2182_U302
g25350 nand P2_R2182_U141 P2_U2671 ; P2_R2182_U303
g25351 nand P2_U2681 P2_R2182_U44 ; P2_R2182_U304
g25352 nand P2_U2702 P2_R2182_U45 ; P2_R2182_U305
g25353 nand P2_R2167_U42 P2_R2167_U41 P2_R2167_U38 ; P2_R2167_U6
g25354 not P2_U2706 ; P2_R2167_U7
g25355 not P2_U2713 ; P2_R2167_U8
g25356 not P2_U2712 ; P2_R2167_U9
g25357 not P2_U2705 ; P2_R2167_U10
g25358 not P2_U2704 ; P2_R2167_U11
g25359 not P2_U2711 ; P2_R2167_U12
g25360 not P2_U2710 ; P2_R2167_U13
g25361 not P2_U2703 ; P2_R2167_U14
g25362 not P2_U2361 ; P2_R2167_U15
g25363 not P2_U2709 ; P2_R2167_U16
g25364 not P2_STATE2_REG_0__SCAN_IN ; P2_R2167_U17
g25365 not P2_U2708 ; P2_R2167_U18
g25366 nand P2_U2714 P2_U2715 ; P2_R2167_U19
g25367 nand P2_U2707 P2_R2167_U19 ; P2_R2167_U20
g25368 or P2_U2714 P2_U2715 ; P2_R2167_U21
g25369 nand P2_U2706 P2_R2167_U8 ; P2_R2167_U22
g25370 nand P2_R2167_U21 P2_R2167_U20 P2_R2167_U22 ; P2_R2167_U23
g25371 nand P2_U2713 P2_R2167_U7 ; P2_R2167_U24
g25372 nand P2_U2712 P2_R2167_U10 ; P2_R2167_U25
g25373 nand P2_R2167_U24 P2_R2167_U25 P2_R2167_U23 ; P2_R2167_U26
g25374 nand P2_U2705 P2_R2167_U9 ; P2_R2167_U27
g25375 nand P2_U2704 P2_R2167_U12 ; P2_R2167_U28
g25376 nand P2_R2167_U27 P2_R2167_U28 P2_R2167_U26 ; P2_R2167_U29
g25377 nand P2_U2711 P2_R2167_U11 ; P2_R2167_U30
g25378 nand P2_U2710 P2_R2167_U14 ; P2_R2167_U31
g25379 nand P2_R2167_U30 P2_R2167_U29 P2_R2167_U31 ; P2_R2167_U32
g25380 nand P2_U2703 P2_R2167_U13 ; P2_R2167_U33
g25381 nand P2_U2361 P2_R2167_U16 ; P2_R2167_U34
g25382 nand P2_R2167_U33 P2_R2167_U32 P2_R2167_U34 ; P2_R2167_U35
g25383 nand P2_U2709 P2_R2167_U15 ; P2_R2167_U36
g25384 nand P2_R2167_U36 P2_R2167_U35 ; P2_R2167_U37
g25385 nand P2_R2167_U40 P2_R2167_U39 P2_R2167_U37 ; P2_R2167_U38
g25386 nand P2_U2361 P2_R2167_U18 ; P2_R2167_U39
g25387 nand P2_U2708 P2_R2167_U15 ; P2_R2167_U40
g25388 nand P2_U2361 P2_R2167_U18 P2_STATE2_REG_0__SCAN_IN ; P2_R2167_U41
g25389 nand P2_R2167_U17 P2_R2167_U15 P2_U2708 ; P2_R2167_U42
g25390 not P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_R2027_U5
g25391 not P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2027_U6
g25392 nand P2_INSTADDRPOINTER_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2027_U7
g25393 not P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2027_U8
g25394 nand P2_R2027_U98 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2027_U9
g25395 not P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2027_U10
g25396 nand P2_R2027_U99 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2027_U11
g25397 not P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2027_U12
g25398 nand P2_R2027_U100 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2027_U13
g25399 not P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2027_U14
g25400 nand P2_R2027_U101 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2027_U15
g25401 not P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2027_U16
g25402 nand P2_R2027_U102 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2027_U17
g25403 not P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2027_U18
g25404 nand P2_R2027_U103 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2027_U19
g25405 not P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2027_U20
g25406 not P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2027_U21
g25407 nand P2_R2027_U104 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2027_U22
g25408 nand P2_R2027_U105 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2027_U23
g25409 not P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2027_U24
g25410 nand P2_R2027_U106 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2027_U25
g25411 not P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2027_U26
g25412 nand P2_R2027_U107 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2027_U27
g25413 not P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2027_U28
g25414 nand P2_R2027_U108 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2027_U29
g25415 not P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2027_U30
g25416 nand P2_R2027_U109 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2027_U31
g25417 not P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2027_U32
g25418 nand P2_R2027_U110 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2027_U33
g25419 not P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2027_U34
g25420 nand P2_R2027_U111 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2027_U35
g25421 not P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2027_U36
g25422 nand P2_R2027_U112 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2027_U37
g25423 not P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2027_U38
g25424 nand P2_R2027_U113 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2027_U39
g25425 not P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2027_U40
g25426 nand P2_R2027_U114 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2027_U41
g25427 not P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2027_U42
g25428 nand P2_R2027_U115 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2027_U43
g25429 not P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2027_U44
g25430 nand P2_R2027_U116 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2027_U45
g25431 not P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2027_U46
g25432 nand P2_R2027_U117 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2027_U47
g25433 not P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2027_U48
g25434 nand P2_R2027_U118 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2027_U49
g25435 not P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2027_U50
g25436 nand P2_R2027_U119 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2027_U51
g25437 not P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2027_U52
g25438 nand P2_R2027_U120 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2027_U53
g25439 not P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2027_U54
g25440 nand P2_R2027_U121 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2027_U55
g25441 not P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2027_U56
g25442 nand P2_R2027_U122 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2027_U57
g25443 not P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2027_U58
g25444 nand P2_R2027_U123 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2027_U59
g25445 not P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2027_U60
g25446 nand P2_R2027_U124 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2027_U61
g25447 not P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2027_U62
g25448 nand P2_R2027_U125 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2027_U63
g25449 not P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2027_U64
g25450 nand P2_R2027_U129 P2_R2027_U128 ; P2_R2027_U65
g25451 nand P2_R2027_U131 P2_R2027_U130 ; P2_R2027_U66
g25452 nand P2_R2027_U133 P2_R2027_U132 ; P2_R2027_U67
g25453 nand P2_R2027_U135 P2_R2027_U134 ; P2_R2027_U68
g25454 nand P2_R2027_U137 P2_R2027_U136 ; P2_R2027_U69
g25455 nand P2_R2027_U139 P2_R2027_U138 ; P2_R2027_U70
g25456 nand P2_R2027_U141 P2_R2027_U140 ; P2_R2027_U71
g25457 nand P2_R2027_U143 P2_R2027_U142 ; P2_R2027_U72
g25458 nand P2_R2027_U145 P2_R2027_U144 ; P2_R2027_U73
g25459 nand P2_R2027_U147 P2_R2027_U146 ; P2_R2027_U74
g25460 nand P2_R2027_U149 P2_R2027_U148 ; P2_R2027_U75
g25461 nand P2_R2027_U151 P2_R2027_U150 ; P2_R2027_U76
g25462 nand P2_R2027_U153 P2_R2027_U152 ; P2_R2027_U77
g25463 nand P2_R2027_U155 P2_R2027_U154 ; P2_R2027_U78
g25464 nand P2_R2027_U157 P2_R2027_U156 ; P2_R2027_U79
g25465 nand P2_R2027_U159 P2_R2027_U158 ; P2_R2027_U80
g25466 nand P2_R2027_U161 P2_R2027_U160 ; P2_R2027_U81
g25467 nand P2_R2027_U163 P2_R2027_U162 ; P2_R2027_U82
g25468 nand P2_R2027_U165 P2_R2027_U164 ; P2_R2027_U83
g25469 nand P2_R2027_U167 P2_R2027_U166 ; P2_R2027_U84
g25470 nand P2_R2027_U169 P2_R2027_U168 ; P2_R2027_U85
g25471 nand P2_R2027_U171 P2_R2027_U170 ; P2_R2027_U86
g25472 nand P2_R2027_U173 P2_R2027_U172 ; P2_R2027_U87
g25473 nand P2_R2027_U175 P2_R2027_U174 ; P2_R2027_U88
g25474 nand P2_R2027_U177 P2_R2027_U176 ; P2_R2027_U89
g25475 nand P2_R2027_U179 P2_R2027_U178 ; P2_R2027_U90
g25476 nand P2_R2027_U181 P2_R2027_U180 ; P2_R2027_U91
g25477 nand P2_R2027_U183 P2_R2027_U182 ; P2_R2027_U92
g25478 nand P2_R2027_U185 P2_R2027_U184 ; P2_R2027_U93
g25479 nand P2_R2027_U187 P2_R2027_U186 ; P2_R2027_U94
g25480 nand P2_R2027_U189 P2_R2027_U188 ; P2_R2027_U95
g25481 not P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_R2027_U96
g25482 nand P2_R2027_U126 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2027_U97
g25483 not P2_R2027_U7 ; P2_R2027_U98
g25484 not P2_R2027_U9 ; P2_R2027_U99
g25485 not P2_R2027_U11 ; P2_R2027_U100
g25486 not P2_R2027_U13 ; P2_R2027_U101
g25487 not P2_R2027_U15 ; P2_R2027_U102
g25488 not P2_R2027_U17 ; P2_R2027_U103
g25489 not P2_R2027_U19 ; P2_R2027_U104
g25490 not P2_R2027_U22 ; P2_R2027_U105
g25491 not P2_R2027_U23 ; P2_R2027_U106
g25492 not P2_R2027_U25 ; P2_R2027_U107
g25493 not P2_R2027_U27 ; P2_R2027_U108
g25494 not P2_R2027_U29 ; P2_R2027_U109
g25495 not P2_R2027_U31 ; P2_R2027_U110
g25496 not P2_R2027_U33 ; P2_R2027_U111
g25497 not P2_R2027_U35 ; P2_R2027_U112
g25498 not P2_R2027_U37 ; P2_R2027_U113
g25499 not P2_R2027_U39 ; P2_R2027_U114
g25500 not P2_R2027_U41 ; P2_R2027_U115
g25501 not P2_R2027_U43 ; P2_R2027_U116
g25502 not P2_R2027_U45 ; P2_R2027_U117
g25503 not P2_R2027_U47 ; P2_R2027_U118
g25504 not P2_R2027_U49 ; P2_R2027_U119
g25505 not P2_R2027_U51 ; P2_R2027_U120
g25506 not P2_R2027_U53 ; P2_R2027_U121
g25507 not P2_R2027_U55 ; P2_R2027_U122
g25508 not P2_R2027_U57 ; P2_R2027_U123
g25509 not P2_R2027_U59 ; P2_R2027_U124
g25510 not P2_R2027_U61 ; P2_R2027_U125
g25511 not P2_R2027_U63 ; P2_R2027_U126
g25512 not P2_R2027_U97 ; P2_R2027_U127
g25513 nand P2_R2027_U22 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2027_U128
g25514 nand P2_R2027_U105 P2_R2027_U21 ; P2_R2027_U129
g25515 nand P2_R2027_U19 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2027_U130
g25516 nand P2_R2027_U104 P2_R2027_U20 ; P2_R2027_U131
g25517 nand P2_R2027_U17 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2027_U132
g25518 nand P2_R2027_U103 P2_R2027_U18 ; P2_R2027_U133
g25519 nand P2_R2027_U15 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2027_U134
g25520 nand P2_R2027_U102 P2_R2027_U16 ; P2_R2027_U135
g25521 nand P2_R2027_U13 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2027_U136
g25522 nand P2_R2027_U101 P2_R2027_U14 ; P2_R2027_U137
g25523 nand P2_R2027_U11 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2027_U138
g25524 nand P2_R2027_U100 P2_R2027_U12 ; P2_R2027_U139
g25525 nand P2_R2027_U9 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2027_U140
g25526 nand P2_R2027_U99 P2_R2027_U10 ; P2_R2027_U141
g25527 nand P2_R2027_U97 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_R2027_U142
g25528 nand P2_R2027_U127 P2_R2027_U96 ; P2_R2027_U143
g25529 nand P2_R2027_U63 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2027_U144
g25530 nand P2_R2027_U126 P2_R2027_U64 ; P2_R2027_U145
g25531 nand P2_R2027_U7 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2027_U146
g25532 nand P2_R2027_U98 P2_R2027_U8 ; P2_R2027_U147
g25533 nand P2_R2027_U61 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2027_U148
g25534 nand P2_R2027_U125 P2_R2027_U62 ; P2_R2027_U149
g25535 nand P2_R2027_U59 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2027_U150
g25536 nand P2_R2027_U124 P2_R2027_U60 ; P2_R2027_U151
g25537 nand P2_R2027_U57 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2027_U152
g25538 nand P2_R2027_U123 P2_R2027_U58 ; P2_R2027_U153
g25539 nand P2_R2027_U55 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2027_U154
g25540 nand P2_R2027_U122 P2_R2027_U56 ; P2_R2027_U155
g25541 nand P2_R2027_U53 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2027_U156
g25542 nand P2_R2027_U121 P2_R2027_U54 ; P2_R2027_U157
g25543 nand P2_R2027_U51 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2027_U158
g25544 nand P2_R2027_U120 P2_R2027_U52 ; P2_R2027_U159
g25545 nand P2_R2027_U49 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2027_U160
g25546 nand P2_R2027_U119 P2_R2027_U50 ; P2_R2027_U161
g25547 nand P2_R2027_U47 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2027_U162
g25548 nand P2_R2027_U118 P2_R2027_U48 ; P2_R2027_U163
g25549 nand P2_R2027_U45 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2027_U164
g25550 nand P2_R2027_U117 P2_R2027_U46 ; P2_R2027_U165
g25551 nand P2_R2027_U43 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2027_U166
g25552 nand P2_R2027_U116 P2_R2027_U44 ; P2_R2027_U167
g25553 nand P2_R2027_U5 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2027_U168
g25554 nand P2_R2027_U6 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_R2027_U169
g25555 nand P2_R2027_U41 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2027_U170
g25556 nand P2_R2027_U115 P2_R2027_U42 ; P2_R2027_U171
g25557 nand P2_R2027_U39 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2027_U172
g25558 nand P2_R2027_U114 P2_R2027_U40 ; P2_R2027_U173
g25559 nand P2_R2027_U37 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2027_U174
g25560 nand P2_R2027_U113 P2_R2027_U38 ; P2_R2027_U175
g25561 nand P2_R2027_U35 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2027_U176
g25562 nand P2_R2027_U112 P2_R2027_U36 ; P2_R2027_U177
g25563 nand P2_R2027_U33 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2027_U178
g25564 nand P2_R2027_U111 P2_R2027_U34 ; P2_R2027_U179
g25565 nand P2_R2027_U31 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2027_U180
g25566 nand P2_R2027_U110 P2_R2027_U32 ; P2_R2027_U181
g25567 nand P2_R2027_U29 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2027_U182
g25568 nand P2_R2027_U109 P2_R2027_U30 ; P2_R2027_U183
g25569 nand P2_R2027_U27 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2027_U184
g25570 nand P2_R2027_U108 P2_R2027_U28 ; P2_R2027_U185
g25571 nand P2_R2027_U25 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2027_U186
g25572 nand P2_R2027_U107 P2_R2027_U26 ; P2_R2027_U187
g25573 nand P2_R2027_U23 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2027_U188
g25574 nand P2_R2027_U106 P2_R2027_U24 ; P2_R2027_U189
g25575 or P2_LT_563_1260_U7 P2_U3617 ; P2_LT_563_1260_U6
g25576 nor P2_SUB_563_U6 P2_SUB_563_U7 ; P2_LT_563_1260_U7
g25577 not P2_PHYADDRPOINTER_REG_1__SCAN_IN ; P2_R2337_U4
g25578 not P2_PHYADDRPOINTER_REG_3__SCAN_IN ; P2_R2337_U5
g25579 not P2_PHYADDRPOINTER_REG_2__SCAN_IN ; P2_R2337_U6
g25580 nand P2_PHYADDRPOINTER_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_2__SCAN_IN P2_PHYADDRPOINTER_REG_3__SCAN_IN ; P2_R2337_U7
g25581 not P2_PHYADDRPOINTER_REG_4__SCAN_IN ; P2_R2337_U8
g25582 nand P2_R2337_U95 P2_PHYADDRPOINTER_REG_4__SCAN_IN ; P2_R2337_U9
g25583 not P2_PHYADDRPOINTER_REG_5__SCAN_IN ; P2_R2337_U10
g25584 nand P2_R2337_U96 P2_PHYADDRPOINTER_REG_5__SCAN_IN ; P2_R2337_U11
g25585 not P2_PHYADDRPOINTER_REG_6__SCAN_IN ; P2_R2337_U12
g25586 nand P2_R2337_U97 P2_PHYADDRPOINTER_REG_6__SCAN_IN ; P2_R2337_U13
g25587 not P2_PHYADDRPOINTER_REG_7__SCAN_IN ; P2_R2337_U14
g25588 nand P2_R2337_U98 P2_PHYADDRPOINTER_REG_7__SCAN_IN ; P2_R2337_U15
g25589 not P2_PHYADDRPOINTER_REG_8__SCAN_IN ; P2_R2337_U16
g25590 not P2_PHYADDRPOINTER_REG_9__SCAN_IN ; P2_R2337_U17
g25591 nand P2_R2337_U99 P2_PHYADDRPOINTER_REG_8__SCAN_IN ; P2_R2337_U18
g25592 nand P2_R2337_U100 P2_PHYADDRPOINTER_REG_9__SCAN_IN ; P2_R2337_U19
g25593 not P2_PHYADDRPOINTER_REG_10__SCAN_IN ; P2_R2337_U20
g25594 nand P2_R2337_U101 P2_PHYADDRPOINTER_REG_10__SCAN_IN ; P2_R2337_U21
g25595 not P2_PHYADDRPOINTER_REG_11__SCAN_IN ; P2_R2337_U22
g25596 nand P2_R2337_U102 P2_PHYADDRPOINTER_REG_11__SCAN_IN ; P2_R2337_U23
g25597 not P2_PHYADDRPOINTER_REG_12__SCAN_IN ; P2_R2337_U24
g25598 nand P2_R2337_U103 P2_PHYADDRPOINTER_REG_12__SCAN_IN ; P2_R2337_U25
g25599 not P2_PHYADDRPOINTER_REG_13__SCAN_IN ; P2_R2337_U26
g25600 nand P2_R2337_U104 P2_PHYADDRPOINTER_REG_13__SCAN_IN ; P2_R2337_U27
g25601 not P2_PHYADDRPOINTER_REG_14__SCAN_IN ; P2_R2337_U28
g25602 nand P2_R2337_U105 P2_PHYADDRPOINTER_REG_14__SCAN_IN ; P2_R2337_U29
g25603 not P2_PHYADDRPOINTER_REG_15__SCAN_IN ; P2_R2337_U30
g25604 nand P2_R2337_U106 P2_PHYADDRPOINTER_REG_15__SCAN_IN ; P2_R2337_U31
g25605 not P2_PHYADDRPOINTER_REG_16__SCAN_IN ; P2_R2337_U32
g25606 nand P2_R2337_U107 P2_PHYADDRPOINTER_REG_16__SCAN_IN ; P2_R2337_U33
g25607 not P2_PHYADDRPOINTER_REG_17__SCAN_IN ; P2_R2337_U34
g25608 nand P2_R2337_U108 P2_PHYADDRPOINTER_REG_17__SCAN_IN ; P2_R2337_U35
g25609 not P2_PHYADDRPOINTER_REG_18__SCAN_IN ; P2_R2337_U36
g25610 nand P2_R2337_U109 P2_PHYADDRPOINTER_REG_18__SCAN_IN ; P2_R2337_U37
g25611 not P2_PHYADDRPOINTER_REG_19__SCAN_IN ; P2_R2337_U38
g25612 nand P2_R2337_U110 P2_PHYADDRPOINTER_REG_19__SCAN_IN ; P2_R2337_U39
g25613 not P2_PHYADDRPOINTER_REG_20__SCAN_IN ; P2_R2337_U40
g25614 nand P2_R2337_U111 P2_PHYADDRPOINTER_REG_20__SCAN_IN ; P2_R2337_U41
g25615 not P2_PHYADDRPOINTER_REG_21__SCAN_IN ; P2_R2337_U42
g25616 nand P2_R2337_U112 P2_PHYADDRPOINTER_REG_21__SCAN_IN ; P2_R2337_U43
g25617 not P2_PHYADDRPOINTER_REG_22__SCAN_IN ; P2_R2337_U44
g25618 nand P2_R2337_U113 P2_PHYADDRPOINTER_REG_22__SCAN_IN ; P2_R2337_U45
g25619 not P2_PHYADDRPOINTER_REG_23__SCAN_IN ; P2_R2337_U46
g25620 nand P2_R2337_U114 P2_PHYADDRPOINTER_REG_23__SCAN_IN ; P2_R2337_U47
g25621 not P2_PHYADDRPOINTER_REG_24__SCAN_IN ; P2_R2337_U48
g25622 nand P2_R2337_U115 P2_PHYADDRPOINTER_REG_24__SCAN_IN ; P2_R2337_U49
g25623 not P2_PHYADDRPOINTER_REG_25__SCAN_IN ; P2_R2337_U50
g25624 nand P2_R2337_U116 P2_PHYADDRPOINTER_REG_25__SCAN_IN ; P2_R2337_U51
g25625 not P2_PHYADDRPOINTER_REG_26__SCAN_IN ; P2_R2337_U52
g25626 nand P2_R2337_U117 P2_PHYADDRPOINTER_REG_26__SCAN_IN ; P2_R2337_U53
g25627 not P2_PHYADDRPOINTER_REG_27__SCAN_IN ; P2_R2337_U54
g25628 nand P2_R2337_U118 P2_PHYADDRPOINTER_REG_27__SCAN_IN ; P2_R2337_U55
g25629 not P2_PHYADDRPOINTER_REG_28__SCAN_IN ; P2_R2337_U56
g25630 nand P2_R2337_U119 P2_PHYADDRPOINTER_REG_28__SCAN_IN ; P2_R2337_U57
g25631 not P2_PHYADDRPOINTER_REG_29__SCAN_IN ; P2_R2337_U58
g25632 nand P2_R2337_U120 P2_PHYADDRPOINTER_REG_29__SCAN_IN ; P2_R2337_U59
g25633 not P2_PHYADDRPOINTER_REG_30__SCAN_IN ; P2_R2337_U60
g25634 nand P2_R2337_U124 P2_R2337_U123 ; P2_R2337_U61
g25635 nand P2_R2337_U126 P2_R2337_U125 ; P2_R2337_U62
g25636 nand P2_R2337_U128 P2_R2337_U127 ; P2_R2337_U63
g25637 nand P2_R2337_U130 P2_R2337_U129 ; P2_R2337_U64
g25638 nand P2_R2337_U132 P2_R2337_U131 ; P2_R2337_U65
g25639 nand P2_R2337_U134 P2_R2337_U133 ; P2_R2337_U66
g25640 nand P2_R2337_U136 P2_R2337_U135 ; P2_R2337_U67
g25641 nand P2_R2337_U138 P2_R2337_U137 ; P2_R2337_U68
g25642 nand P2_R2337_U140 P2_R2337_U139 ; P2_R2337_U69
g25643 nand P2_R2337_U142 P2_R2337_U141 ; P2_R2337_U70
g25644 nand P2_R2337_U144 P2_R2337_U143 ; P2_R2337_U71
g25645 nand P2_R2337_U146 P2_R2337_U145 ; P2_R2337_U72
g25646 nand P2_R2337_U148 P2_R2337_U147 ; P2_R2337_U73
g25647 nand P2_R2337_U150 P2_R2337_U149 ; P2_R2337_U74
g25648 nand P2_R2337_U152 P2_R2337_U151 ; P2_R2337_U75
g25649 nand P2_R2337_U154 P2_R2337_U153 ; P2_R2337_U76
g25650 nand P2_R2337_U156 P2_R2337_U155 ; P2_R2337_U77
g25651 nand P2_R2337_U158 P2_R2337_U157 ; P2_R2337_U78
g25652 nand P2_R2337_U160 P2_R2337_U159 ; P2_R2337_U79
g25653 nand P2_R2337_U162 P2_R2337_U161 ; P2_R2337_U80
g25654 nand P2_R2337_U164 P2_R2337_U163 ; P2_R2337_U81
g25655 nand P2_R2337_U166 P2_R2337_U165 ; P2_R2337_U82
g25656 nand P2_R2337_U168 P2_R2337_U167 ; P2_R2337_U83
g25657 nand P2_R2337_U170 P2_R2337_U169 ; P2_R2337_U84
g25658 nand P2_R2337_U172 P2_R2337_U171 ; P2_R2337_U85
g25659 nand P2_R2337_U174 P2_R2337_U173 ; P2_R2337_U86
g25660 nand P2_R2337_U176 P2_R2337_U175 ; P2_R2337_U87
g25661 nand P2_R2337_U178 P2_R2337_U177 ; P2_R2337_U88
g25662 nand P2_R2337_U180 P2_R2337_U179 ; P2_R2337_U89
g25663 nand P2_R2337_U182 P2_R2337_U181 ; P2_R2337_U90
g25664 nand P2_PHYADDRPOINTER_REG_1__SCAN_IN P2_PHYADDRPOINTER_REG_2__SCAN_IN ; P2_R2337_U91
g25665 not P2_PHYADDRPOINTER_REG_31__SCAN_IN ; P2_R2337_U92
g25666 nand P2_R2337_U121 P2_PHYADDRPOINTER_REG_30__SCAN_IN ; P2_R2337_U93
g25667 not P2_R2337_U91 ; P2_R2337_U94
g25668 not P2_R2337_U7 ; P2_R2337_U95
g25669 not P2_R2337_U9 ; P2_R2337_U96
g25670 not P2_R2337_U11 ; P2_R2337_U97
g25671 not P2_R2337_U13 ; P2_R2337_U98
g25672 not P2_R2337_U15 ; P2_R2337_U99
g25673 not P2_R2337_U18 ; P2_R2337_U100
g25674 not P2_R2337_U19 ; P2_R2337_U101
g25675 not P2_R2337_U21 ; P2_R2337_U102
g25676 not P2_R2337_U23 ; P2_R2337_U103
g25677 not P2_R2337_U25 ; P2_R2337_U104
g25678 not P2_R2337_U27 ; P2_R2337_U105
g25679 not P2_R2337_U29 ; P2_R2337_U106
g25680 not P2_R2337_U31 ; P2_R2337_U107
g25681 not P2_R2337_U33 ; P2_R2337_U108
g25682 not P2_R2337_U35 ; P2_R2337_U109
g25683 not P2_R2337_U37 ; P2_R2337_U110
g25684 not P2_R2337_U39 ; P2_R2337_U111
g25685 not P2_R2337_U41 ; P2_R2337_U112
g25686 not P2_R2337_U43 ; P2_R2337_U113
g25687 not P2_R2337_U45 ; P2_R2337_U114
g25688 not P2_R2337_U47 ; P2_R2337_U115
g25689 not P2_R2337_U49 ; P2_R2337_U116
g25690 not P2_R2337_U51 ; P2_R2337_U117
g25691 not P2_R2337_U53 ; P2_R2337_U118
g25692 not P2_R2337_U55 ; P2_R2337_U119
g25693 not P2_R2337_U57 ; P2_R2337_U120
g25694 not P2_R2337_U59 ; P2_R2337_U121
g25695 not P2_R2337_U93 ; P2_R2337_U122
g25696 nand P2_R2337_U18 P2_PHYADDRPOINTER_REG_9__SCAN_IN ; P2_R2337_U123
g25697 nand P2_R2337_U100 P2_R2337_U17 ; P2_R2337_U124
g25698 nand P2_R2337_U15 P2_PHYADDRPOINTER_REG_8__SCAN_IN ; P2_R2337_U125
g25699 nand P2_R2337_U99 P2_R2337_U16 ; P2_R2337_U126
g25700 nand P2_R2337_U13 P2_PHYADDRPOINTER_REG_7__SCAN_IN ; P2_R2337_U127
g25701 nand P2_R2337_U98 P2_R2337_U14 ; P2_R2337_U128
g25702 nand P2_R2337_U11 P2_PHYADDRPOINTER_REG_6__SCAN_IN ; P2_R2337_U129
g25703 nand P2_R2337_U97 P2_R2337_U12 ; P2_R2337_U130
g25704 nand P2_R2337_U9 P2_PHYADDRPOINTER_REG_5__SCAN_IN ; P2_R2337_U131
g25705 nand P2_R2337_U96 P2_R2337_U10 ; P2_R2337_U132
g25706 nand P2_R2337_U7 P2_PHYADDRPOINTER_REG_4__SCAN_IN ; P2_R2337_U133
g25707 nand P2_R2337_U95 P2_R2337_U8 ; P2_R2337_U134
g25708 nand P2_R2337_U91 P2_PHYADDRPOINTER_REG_3__SCAN_IN ; P2_R2337_U135
g25709 nand P2_R2337_U94 P2_R2337_U5 ; P2_R2337_U136
g25710 nand P2_R2337_U93 P2_PHYADDRPOINTER_REG_31__SCAN_IN ; P2_R2337_U137
g25711 nand P2_R2337_U122 P2_R2337_U92 ; P2_R2337_U138
g25712 nand P2_R2337_U59 P2_PHYADDRPOINTER_REG_30__SCAN_IN ; P2_R2337_U139
g25713 nand P2_R2337_U121 P2_R2337_U60 ; P2_R2337_U140
g25714 nand P2_R2337_U4 P2_PHYADDRPOINTER_REG_2__SCAN_IN ; P2_R2337_U141
g25715 nand P2_R2337_U6 P2_PHYADDRPOINTER_REG_1__SCAN_IN ; P2_R2337_U142
g25716 nand P2_R2337_U57 P2_PHYADDRPOINTER_REG_29__SCAN_IN ; P2_R2337_U143
g25717 nand P2_R2337_U120 P2_R2337_U58 ; P2_R2337_U144
g25718 nand P2_R2337_U55 P2_PHYADDRPOINTER_REG_28__SCAN_IN ; P2_R2337_U145
g25719 nand P2_R2337_U119 P2_R2337_U56 ; P2_R2337_U146
g25720 nand P2_R2337_U53 P2_PHYADDRPOINTER_REG_27__SCAN_IN ; P2_R2337_U147
g25721 nand P2_R2337_U118 P2_R2337_U54 ; P2_R2337_U148
g25722 nand P2_R2337_U51 P2_PHYADDRPOINTER_REG_26__SCAN_IN ; P2_R2337_U149
g25723 nand P2_R2337_U117 P2_R2337_U52 ; P2_R2337_U150
g25724 nand P2_R2337_U49 P2_PHYADDRPOINTER_REG_25__SCAN_IN ; P2_R2337_U151
g25725 nand P2_R2337_U116 P2_R2337_U50 ; P2_R2337_U152
g25726 nand P2_R2337_U47 P2_PHYADDRPOINTER_REG_24__SCAN_IN ; P2_R2337_U153
g25727 nand P2_R2337_U115 P2_R2337_U48 ; P2_R2337_U154
g25728 nand P2_R2337_U45 P2_PHYADDRPOINTER_REG_23__SCAN_IN ; P2_R2337_U155
g25729 nand P2_R2337_U114 P2_R2337_U46 ; P2_R2337_U156
g25730 nand P2_R2337_U43 P2_PHYADDRPOINTER_REG_22__SCAN_IN ; P2_R2337_U157
g25731 nand P2_R2337_U113 P2_R2337_U44 ; P2_R2337_U158
g25732 nand P2_R2337_U41 P2_PHYADDRPOINTER_REG_21__SCAN_IN ; P2_R2337_U159
g25733 nand P2_R2337_U112 P2_R2337_U42 ; P2_R2337_U160
g25734 nand P2_R2337_U39 P2_PHYADDRPOINTER_REG_20__SCAN_IN ; P2_R2337_U161
g25735 nand P2_R2337_U111 P2_R2337_U40 ; P2_R2337_U162
g25736 nand P2_R2337_U37 P2_PHYADDRPOINTER_REG_19__SCAN_IN ; P2_R2337_U163
g25737 nand P2_R2337_U110 P2_R2337_U38 ; P2_R2337_U164
g25738 nand P2_R2337_U35 P2_PHYADDRPOINTER_REG_18__SCAN_IN ; P2_R2337_U165
g25739 nand P2_R2337_U109 P2_R2337_U36 ; P2_R2337_U166
g25740 nand P2_R2337_U33 P2_PHYADDRPOINTER_REG_17__SCAN_IN ; P2_R2337_U167
g25741 nand P2_R2337_U108 P2_R2337_U34 ; P2_R2337_U168
g25742 nand P2_R2337_U31 P2_PHYADDRPOINTER_REG_16__SCAN_IN ; P2_R2337_U169
g25743 nand P2_R2337_U107 P2_R2337_U32 ; P2_R2337_U170
g25744 nand P2_R2337_U29 P2_PHYADDRPOINTER_REG_15__SCAN_IN ; P2_R2337_U171
g25745 nand P2_R2337_U106 P2_R2337_U30 ; P2_R2337_U172
g25746 nand P2_R2337_U27 P2_PHYADDRPOINTER_REG_14__SCAN_IN ; P2_R2337_U173
g25747 nand P2_R2337_U105 P2_R2337_U28 ; P2_R2337_U174
g25748 nand P2_R2337_U25 P2_PHYADDRPOINTER_REG_13__SCAN_IN ; P2_R2337_U175
g25749 nand P2_R2337_U104 P2_R2337_U26 ; P2_R2337_U176
g25750 nand P2_R2337_U23 P2_PHYADDRPOINTER_REG_12__SCAN_IN ; P2_R2337_U177
g25751 nand P2_R2337_U103 P2_R2337_U24 ; P2_R2337_U178
g25752 nand P2_R2337_U21 P2_PHYADDRPOINTER_REG_11__SCAN_IN ; P2_R2337_U179
g25753 nand P2_R2337_U102 P2_R2337_U22 ; P2_R2337_U180
g25754 nand P2_R2337_U19 P2_PHYADDRPOINTER_REG_10__SCAN_IN ; P2_R2337_U181
g25755 nand P2_R2337_U101 P2_R2337_U20 ; P2_R2337_U182
g25756 not P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_R2147_U4
g25757 not P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_R2147_U5
g25758 not P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_R2147_U6
g25759 nand P2_R2147_U16 P2_R2147_U15 ; P2_R2147_U7
g25760 nand P2_R2147_U18 P2_R2147_U17 ; P2_R2147_U8
g25761 nand P2_R2147_U20 P2_R2147_U19 ; P2_R2147_U9
g25762 not P2_U2752 ; P2_R2147_U10
g25763 nand P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_R2147_U11
g25764 nand P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_R2147_U12
g25765 not P2_R2147_U11 ; P2_R2147_U13
g25766 not P2_R2147_U12 ; P2_R2147_U14
g25767 nand P2_U2752 P2_R2147_U11 ; P2_R2147_U15
g25768 nand P2_R2147_U13 P2_R2147_U10 ; P2_R2147_U16
g25769 nand P2_R2147_U12 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_R2147_U17
g25770 nand P2_R2147_U14 P2_R2147_U5 ; P2_R2147_U18
g25771 nand P2_R2147_U4 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_R2147_U19
g25772 nand P2_R2147_U6 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_R2147_U20
g25773 and P2_R2219_U52 P2_R2219_U48 ; P2_R2219_U6
g25774 and P2_R2219_U68 P2_R2219_U66 ; P2_R2219_U7
g25775 nand P2_R2219_U45 P2_R2219_U69 ; P2_R2219_U8
g25776 not P2_U4428 ; P2_R2219_U9
g25777 not P2_U2753 ; P2_R2219_U10
g25778 not P2_U2761 ; P2_R2219_U11
g25779 not P2_U2763 ; P2_R2219_U12
g25780 not P2_U2762 ; P2_R2219_U13
g25781 not P2_U2756 ; P2_R2219_U14
g25782 not P2_U2765 ; P2_R2219_U15
g25783 not P2_U2764 ; P2_R2219_U16
g25784 not P2_U2755 ; P2_R2219_U17
g25785 not P2_U2754 ; P2_R2219_U18
g25786 nand P2_R2219_U72 P2_R2219_U76 ; P2_R2219_U19
g25787 not P2_U2760 ; P2_R2219_U20
g25788 not P2_U2759 ; P2_R2219_U21
g25789 not P2_U2758 ; P2_R2219_U22
g25790 not P2_U2757 ; P2_R2219_U23
g25791 nand P2_R2219_U86 P2_R2219_U85 ; P2_R2219_U24
g25792 nand P2_R2219_U91 P2_R2219_U90 ; P2_R2219_U25
g25793 nand P2_R2219_U96 P2_R2219_U95 ; P2_R2219_U26
g25794 nand P2_R2219_U101 P2_R2219_U100 ; P2_R2219_U27
g25795 nand P2_R2219_U106 P2_R2219_U105 ; P2_R2219_U28
g25796 nand P2_R2219_U111 P2_R2219_U110 ; P2_R2219_U29
g25797 nand P2_R2219_U116 P2_R2219_U115 ; P2_R2219_U30
g25798 and P2_R2219_U6 P2_R2219_U55 ; P2_R2219_U31
g25799 nand P2_R2219_U83 P2_R2219_U82 ; P2_R2219_U32
g25800 nand P2_R2219_U88 P2_R2219_U87 ; P2_R2219_U33
g25801 nand P2_R2219_U93 P2_R2219_U92 ; P2_R2219_U34
g25802 nand P2_R2219_U98 P2_R2219_U97 ; P2_R2219_U35
g25803 nand P2_R2219_U103 P2_R2219_U102 ; P2_R2219_U36
g25804 nand P2_R2219_U108 P2_R2219_U107 ; P2_R2219_U37
g25805 nand P2_R2219_U113 P2_R2219_U112 ; P2_R2219_U38
g25806 nand P2_R2219_U64 P2_R2219_U63 ; P2_R2219_U39
g25807 nand P2_R2219_U60 P2_R2219_U59 ; P2_R2219_U40
g25808 nand P2_R2219_U75 P2_R2219_U56 P2_R2219_U74 ; P2_R2219_U41
g25809 nand P2_R2219_U19 P2_R2219_U71 ; P2_R2219_U42
g25810 nand P2_R2219_U50 P2_R2219_U49 ; P2_R2219_U43
g25811 nand P2_R2219_U78 P2_R2219_U70 ; P2_R2219_U44
g25812 nand P2_U2765 P2_R2219_U23 ; P2_R2219_U45
g25813 not P2_R2219_U45 ; P2_R2219_U46
g25814 nand P2_U2764 P2_R2219_U14 ; P2_R2219_U47
g25815 nand P2_U2763 P2_R2219_U17 ; P2_R2219_U48
g25816 nand P2_R2219_U48 P2_R2219_U81 ; P2_R2219_U49
g25817 nand P2_U2755 P2_R2219_U12 ; P2_R2219_U50
g25818 not P2_R2219_U43 ; P2_R2219_U51
g25819 nand P2_U2762 P2_R2219_U18 ; P2_R2219_U52
g25820 nand P2_U2754 P2_R2219_U13 ; P2_R2219_U53
g25821 not P2_R2219_U42 ; P2_R2219_U54
g25822 nand P2_U2761 P2_R2219_U10 ; P2_R2219_U55
g25823 nand P2_U2753 P2_R2219_U11 ; P2_R2219_U56
g25824 not P2_R2219_U41 ; P2_R2219_U57
g25825 nand P2_U2760 P2_R2219_U9 ; P2_R2219_U58
g25826 nand P2_R2219_U58 P2_R2219_U41 ; P2_R2219_U59
g25827 nand P2_U4428 P2_R2219_U20 ; P2_R2219_U60
g25828 not P2_R2219_U40 ; P2_R2219_U61
g25829 nand P2_U2759 P2_R2219_U9 ; P2_R2219_U62
g25830 nand P2_R2219_U62 P2_R2219_U40 ; P2_R2219_U63
g25831 nand P2_U4428 P2_R2219_U21 ; P2_R2219_U64
g25832 not P2_R2219_U39 ; P2_R2219_U65
g25833 nand P2_U4428 P2_R2219_U22 ; P2_R2219_U66
g25834 nand P2_U2758 P2_R2219_U9 ; P2_R2219_U67
g25835 nand P2_R2219_U67 P2_R2219_U39 ; P2_R2219_U68
g25836 nand P2_U2757 P2_R2219_U15 ; P2_R2219_U69
g25837 nand P2_U2756 P2_R2219_U16 ; P2_R2219_U70
g25838 nand P2_R2219_U6 P2_R2219_U44 ; P2_R2219_U71
g25839 nand P2_R2219_U53 P2_R2219_U50 ; P2_R2219_U72
g25840 not P2_R2219_U19 ; P2_R2219_U73
g25841 nand P2_R2219_U31 P2_R2219_U44 ; P2_R2219_U74
g25842 nand P2_R2219_U73 P2_R2219_U55 ; P2_R2219_U75
g25843 nand P2_U2762 P2_R2219_U18 ; P2_R2219_U76
g25844 nand P2_U2764 P2_R2219_U14 ; P2_R2219_U77
g25845 nand P2_R2219_U47 P2_R2219_U45 ; P2_R2219_U78
g25846 not P2_R2219_U44 ; P2_R2219_U79
g25847 nand P2_R2219_U77 P2_R2219_U45 ; P2_R2219_U80
g25848 nand P2_R2219_U80 P2_R2219_U70 ; P2_R2219_U81
g25849 nand P2_U2758 P2_R2219_U9 ; P2_R2219_U82
g25850 nand P2_U4428 P2_R2219_U22 ; P2_R2219_U83
g25851 not P2_R2219_U32 ; P2_R2219_U84
g25852 nand P2_R2219_U65 P2_R2219_U84 ; P2_R2219_U85
g25853 nand P2_R2219_U32 P2_R2219_U39 ; P2_R2219_U86
g25854 nand P2_U2759 P2_R2219_U9 ; P2_R2219_U87
g25855 nand P2_U4428 P2_R2219_U21 ; P2_R2219_U88
g25856 not P2_R2219_U33 ; P2_R2219_U89
g25857 nand P2_R2219_U61 P2_R2219_U89 ; P2_R2219_U90
g25858 nand P2_R2219_U33 P2_R2219_U40 ; P2_R2219_U91
g25859 nand P2_U2760 P2_R2219_U9 ; P2_R2219_U92
g25860 nand P2_U4428 P2_R2219_U20 ; P2_R2219_U93
g25861 not P2_R2219_U34 ; P2_R2219_U94
g25862 nand P2_R2219_U57 P2_R2219_U94 ; P2_R2219_U95
g25863 nand P2_R2219_U34 P2_R2219_U41 ; P2_R2219_U96
g25864 nand P2_U2761 P2_R2219_U10 ; P2_R2219_U97
g25865 nand P2_U2753 P2_R2219_U11 ; P2_R2219_U98
g25866 not P2_R2219_U35 ; P2_R2219_U99
g25867 nand P2_R2219_U54 P2_R2219_U99 ; P2_R2219_U100
g25868 nand P2_R2219_U35 P2_R2219_U42 ; P2_R2219_U101
g25869 nand P2_U2762 P2_R2219_U18 ; P2_R2219_U102
g25870 nand P2_U2754 P2_R2219_U13 ; P2_R2219_U103
g25871 not P2_R2219_U36 ; P2_R2219_U104
g25872 nand P2_R2219_U51 P2_R2219_U104 ; P2_R2219_U105
g25873 nand P2_R2219_U36 P2_R2219_U43 ; P2_R2219_U106
g25874 nand P2_U2763 P2_R2219_U17 ; P2_R2219_U107
g25875 nand P2_U2755 P2_R2219_U12 ; P2_R2219_U108
g25876 not P2_R2219_U37 ; P2_R2219_U109
g25877 nand P2_R2219_U79 P2_R2219_U109 ; P2_R2219_U110
g25878 nand P2_R2219_U37 P2_R2219_U44 ; P2_R2219_U111
g25879 nand P2_U2764 P2_R2219_U14 ; P2_R2219_U112
g25880 nand P2_U2756 P2_R2219_U16 ; P2_R2219_U113
g25881 not P2_R2219_U38 ; P2_R2219_U114
g25882 nand P2_R2219_U46 P2_R2219_U114 ; P2_R2219_U115
g25883 nand P2_R2219_U38 P2_R2219_U45 ; P2_R2219_U116
g25884 nor P2_U3686 P2_U3685 P2_U3684 P2_U3687 ; P2_R2243_U6
g25885 nor P2_U3684 P2_R2243_U9 ; P2_R2243_U7
g25886 nand P2_R2243_U7 P2_R2243_U11 ; P2_R2243_U8
g25887 nor P2_U3689 P2_U3687 P2_U3684 P2_U3686 P2_U3685 ; P2_R2243_U9
g25888 not P2_U3688 ; P2_R2243_U10
g25889 nand P2_R2243_U6 P2_R2243_U10 ; P2_R2243_U11
g25890 not P2_U3614 ; P2_SUB_589_U6
g25891 not P2_U3615 ; P2_SUB_589_U7
g25892 not P2_U2813 ; P2_SUB_589_U8
g25893 not P2_U3613 ; P2_SUB_589_U9
g25894 and P2_U2640 P2_R2096_U23 ; P2_R2096_U4
g25895 and P2_U2633 P2_R2096_U18 ; P2_R2096_U5
g25896 and P2_U2631 P2_R2096_U25 ; P2_R2096_U6
g25897 and P2_U2629 P2_R2096_U16 ; P2_R2096_U7
g25898 and P2_U2628 P2_R2096_U7 ; P2_R2096_U8
g25899 and P2_U2627 P2_R2096_U8 ; P2_R2096_U9
g25900 and P2_U2626 P2_R2096_U9 ; P2_R2096_U10
g25901 and P2_U2625 P2_R2096_U10 ; P2_R2096_U11
g25902 and P2_U2624 P2_R2096_U11 ; P2_R2096_U12
g25903 and P2_U2622 P2_R2096_U15 ; P2_R2096_U13
g25904 and P2_U2621 P2_R2096_U13 ; P2_R2096_U14
g25905 and P2_U2623 P2_R2096_U12 ; P2_R2096_U15
g25906 and P2_U2630 P2_R2096_U6 ; P2_R2096_U16
g25907 and P2_U2635 P2_R2096_U21 ; P2_R2096_U17
g25908 and P2_U2634 P2_R2096_U17 ; P2_R2096_U18
g25909 and P2_U2638 P2_R2096_U24 ; P2_R2096_U19
g25910 and P2_U2637 P2_R2096_U19 ; P2_R2096_U20
g25911 and P2_U2636 P2_R2096_U20 ; P2_R2096_U21
g25912 and P2_U2620 P2_R2096_U14 ; P2_R2096_U22
g25913 and P2_U2641 P2_R2096_U99 ; P2_R2096_U23
g25914 and P2_U2639 P2_R2096_U4 ; P2_R2096_U24
g25915 and P2_U2632 P2_R2096_U5 ; P2_R2096_U25
g25916 not P2_U2631 ; P2_R2096_U26
g25917 not P2_U2638 ; P2_R2096_U27
g25918 not P2_U2640 ; P2_R2096_U28
g25919 not P2_U2618 ; P2_R2096_U29
g25920 not P2_U2619 ; P2_R2096_U30
g25921 not P2_U2635 ; P2_R2096_U31
g25922 not P2_U2636 ; P2_R2096_U32
g25923 not P2_U2637 ; P2_R2096_U33
g25924 not P2_U2633 ; P2_R2096_U34
g25925 not P2_U2634 ; P2_R2096_U35
g25926 not P2_U2629 ; P2_R2096_U36
g25927 not P2_U2641 ; P2_R2096_U37
g25928 not P2_U2622 ; P2_R2096_U38
g25929 not P2_U2627 ; P2_R2096_U39
g25930 not P2_U2620 ; P2_R2096_U40
g25931 not P2_U2621 ; P2_R2096_U41
g25932 not P2_U2623 ; P2_R2096_U42
g25933 not P2_U2624 ; P2_R2096_U43
g25934 not P2_U2625 ; P2_R2096_U44
g25935 not P2_U2626 ; P2_R2096_U45
g25936 not P2_U2628 ; P2_R2096_U46
g25937 not P2_U2630 ; P2_R2096_U47
g25938 not P2_U2632 ; P2_R2096_U48
g25939 not P2_U2639 ; P2_R2096_U49
g25940 and P2_R2096_U168 P2_R2096_U167 ; P2_R2096_U50
g25941 nand P2_R2096_U114 P2_R2096_U170 ; P2_R2096_U51
g25942 not P2_U2657 ; P2_R2096_U52
g25943 not P2_U2649 ; P2_R2096_U53
g25944 not P2_U2648 ; P2_R2096_U54
g25945 not P2_U2656 ; P2_R2096_U55
g25946 not P2_U2655 ; P2_R2096_U56
g25947 not P2_U2647 ; P2_R2096_U57
g25948 not P2_U2654 ; P2_R2096_U58
g25949 not P2_U2646 ; P2_R2096_U59
g25950 not P2_U2653 ; P2_R2096_U60
g25951 not P2_U2645 ; P2_R2096_U61
g25952 not P2_U2652 ; P2_R2096_U62
g25953 not P2_U2644 ; P2_R2096_U63
g25954 not P2_U2651 ; P2_R2096_U64
g25955 not P2_U2643 ; P2_R2096_U65
g25956 not P2_U2650 ; P2_R2096_U66
g25957 not P2_U2642 ; P2_R2096_U67
g25958 nand P2_R2096_U265 P2_R2096_U264 ; P2_R2096_U68
g25959 nand P2_R2096_U172 P2_R2096_U171 ; P2_R2096_U69
g25960 nand P2_R2096_U174 P2_R2096_U173 ; P2_R2096_U70
g25961 nand P2_R2096_U181 P2_R2096_U180 ; P2_R2096_U71
g25962 nand P2_R2096_U188 P2_R2096_U187 ; P2_R2096_U72
g25963 nand P2_R2096_U195 P2_R2096_U194 ; P2_R2096_U73
g25964 nand P2_R2096_U202 P2_R2096_U201 ; P2_R2096_U74
g25965 nand P2_R2096_U209 P2_R2096_U208 ; P2_R2096_U75
g25966 nand P2_R2096_U211 P2_R2096_U210 ; P2_R2096_U76
g25967 nand P2_R2096_U218 P2_R2096_U217 ; P2_R2096_U77
g25968 nand P2_R2096_U220 P2_R2096_U219 ; P2_R2096_U78
g25969 nand P2_R2096_U222 P2_R2096_U221 ; P2_R2096_U79
g25970 nand P2_R2096_U224 P2_R2096_U223 ; P2_R2096_U80
g25971 nand P2_R2096_U226 P2_R2096_U225 ; P2_R2096_U81
g25972 nand P2_R2096_U228 P2_R2096_U227 ; P2_R2096_U82
g25973 nand P2_R2096_U230 P2_R2096_U229 ; P2_R2096_U83
g25974 nand P2_R2096_U232 P2_R2096_U231 ; P2_R2096_U84
g25975 nand P2_R2096_U234 P2_R2096_U233 ; P2_R2096_U85
g25976 nand P2_R2096_U236 P2_R2096_U235 ; P2_R2096_U86
g25977 nand P2_R2096_U238 P2_R2096_U237 ; P2_R2096_U87
g25978 nand P2_R2096_U245 P2_R2096_U244 ; P2_R2096_U88
g25979 nand P2_R2096_U247 P2_R2096_U246 ; P2_R2096_U89
g25980 nand P2_R2096_U249 P2_R2096_U248 ; P2_R2096_U90
g25981 nand P2_R2096_U251 P2_R2096_U250 ; P2_R2096_U91
g25982 nand P2_R2096_U253 P2_R2096_U252 ; P2_R2096_U92
g25983 nand P2_R2096_U255 P2_R2096_U254 ; P2_R2096_U93
g25984 nand P2_R2096_U257 P2_R2096_U256 ; P2_R2096_U94
g25985 nand P2_R2096_U259 P2_R2096_U258 ; P2_R2096_U95
g25986 nand P2_R2096_U261 P2_R2096_U260 ; P2_R2096_U96
g25987 nand P2_R2096_U263 P2_R2096_U262 ; P2_R2096_U97
g25988 and P2_U2619 P2_U2618 ; P2_R2096_U98
g25989 nand P2_R2096_U142 P2_R2096_U141 ; P2_R2096_U99
g25990 and P2_R2096_U176 P2_R2096_U175 ; P2_R2096_U100
g25991 nand P2_R2096_U138 P2_R2096_U137 ; P2_R2096_U101
g25992 and P2_R2096_U183 P2_R2096_U182 ; P2_R2096_U102
g25993 nand P2_R2096_U134 P2_R2096_U133 ; P2_R2096_U103
g25994 and P2_R2096_U190 P2_R2096_U189 ; P2_R2096_U104
g25995 nand P2_R2096_U130 P2_R2096_U129 ; P2_R2096_U105
g25996 and P2_R2096_U197 P2_R2096_U196 ; P2_R2096_U106
g25997 nand P2_R2096_U126 P2_R2096_U125 ; P2_R2096_U107
g25998 and P2_R2096_U204 P2_R2096_U203 ; P2_R2096_U108
g25999 nand P2_R2096_U122 P2_R2096_U121 ; P2_R2096_U109
g26000 and P2_R2096_U213 P2_R2096_U212 ; P2_R2096_U110
g26001 nand P2_R2096_U113 P2_R2096_U118 ; P2_R2096_U111
g26002 nand P2_U2649 P2_U2657 ; P2_R2096_U112
g26003 nand P2_U2649 P2_U2657 P2_U2656 ; P2_R2096_U113
g26004 and P2_R2096_U243 P2_R2096_U242 ; P2_R2096_U114
g26005 not P2_R2096_U113 ; P2_R2096_U115
g26006 nand P2_U2649 P2_U2657 ; P2_R2096_U116
g26007 nand P2_R2096_U55 P2_R2096_U116 ; P2_R2096_U117
g26008 nand P2_U2648 P2_R2096_U117 ; P2_R2096_U118
g26009 not P2_R2096_U111 ; P2_R2096_U119
g26010 or P2_U2655 P2_U2647 ; P2_R2096_U120
g26011 nand P2_R2096_U120 P2_R2096_U111 ; P2_R2096_U121
g26012 nand P2_U2647 P2_U2655 ; P2_R2096_U122
g26013 not P2_R2096_U109 ; P2_R2096_U123
g26014 or P2_U2654 P2_U2646 ; P2_R2096_U124
g26015 nand P2_R2096_U124 P2_R2096_U109 ; P2_R2096_U125
g26016 nand P2_U2646 P2_U2654 ; P2_R2096_U126
g26017 not P2_R2096_U107 ; P2_R2096_U127
g26018 or P2_U2653 P2_U2645 ; P2_R2096_U128
g26019 nand P2_R2096_U128 P2_R2096_U107 ; P2_R2096_U129
g26020 nand P2_U2645 P2_U2653 ; P2_R2096_U130
g26021 not P2_R2096_U105 ; P2_R2096_U131
g26022 or P2_U2652 P2_U2644 ; P2_R2096_U132
g26023 nand P2_R2096_U132 P2_R2096_U105 ; P2_R2096_U133
g26024 nand P2_U2644 P2_U2652 ; P2_R2096_U134
g26025 not P2_R2096_U103 ; P2_R2096_U135
g26026 or P2_U2651 P2_U2643 ; P2_R2096_U136
g26027 nand P2_R2096_U136 P2_R2096_U103 ; P2_R2096_U137
g26028 nand P2_U2643 P2_U2651 ; P2_R2096_U138
g26029 not P2_R2096_U101 ; P2_R2096_U139
g26030 or P2_U2650 P2_U2642 ; P2_R2096_U140
g26031 nand P2_R2096_U140 P2_R2096_U101 ; P2_R2096_U141
g26032 nand P2_U2642 P2_U2650 ; P2_R2096_U142
g26033 not P2_R2096_U99 ; P2_R2096_U143
g26034 not P2_R2096_U23 ; P2_R2096_U144
g26035 not P2_R2096_U4 ; P2_R2096_U145
g26036 not P2_R2096_U24 ; P2_R2096_U146
g26037 not P2_R2096_U19 ; P2_R2096_U147
g26038 not P2_R2096_U20 ; P2_R2096_U148
g26039 not P2_R2096_U21 ; P2_R2096_U149
g26040 not P2_R2096_U17 ; P2_R2096_U150
g26041 not P2_R2096_U18 ; P2_R2096_U151
g26042 not P2_R2096_U5 ; P2_R2096_U152
g26043 not P2_R2096_U25 ; P2_R2096_U153
g26044 not P2_R2096_U6 ; P2_R2096_U154
g26045 not P2_R2096_U16 ; P2_R2096_U155
g26046 not P2_R2096_U7 ; P2_R2096_U156
g26047 not P2_R2096_U8 ; P2_R2096_U157
g26048 not P2_R2096_U9 ; P2_R2096_U158
g26049 not P2_R2096_U10 ; P2_R2096_U159
g26050 not P2_R2096_U11 ; P2_R2096_U160
g26051 not P2_R2096_U12 ; P2_R2096_U161
g26052 not P2_R2096_U15 ; P2_R2096_U162
g26053 not P2_R2096_U13 ; P2_R2096_U163
g26054 not P2_R2096_U14 ; P2_R2096_U164
g26055 not P2_R2096_U22 ; P2_R2096_U165
g26056 nand P2_U2619 P2_R2096_U22 ; P2_R2096_U166
g26057 nand P2_R2096_U29 P2_R2096_U166 ; P2_R2096_U167
g26058 nand P2_R2096_U98 P2_R2096_U22 ; P2_R2096_U168
g26059 not P2_R2096_U112 ; P2_R2096_U169
g26060 nand P2_R2096_U241 P2_R2096_U55 ; P2_R2096_U170
g26061 nand P2_R2096_U28 P2_R2096_U23 ; P2_R2096_U171
g26062 nand P2_R2096_U144 P2_U2640 ; P2_R2096_U172
g26063 nand P2_R2096_U37 P2_R2096_U99 ; P2_R2096_U173
g26064 nand P2_R2096_U143 P2_U2641 ; P2_R2096_U174
g26065 nand P2_U2642 P2_R2096_U66 ; P2_R2096_U175
g26066 nand P2_U2650 P2_R2096_U67 ; P2_R2096_U176
g26067 nand P2_U2642 P2_R2096_U66 ; P2_R2096_U177
g26068 nand P2_U2650 P2_R2096_U67 ; P2_R2096_U178
g26069 nand P2_R2096_U178 P2_R2096_U177 ; P2_R2096_U179
g26070 nand P2_R2096_U100 P2_R2096_U101 ; P2_R2096_U180
g26071 nand P2_R2096_U139 P2_R2096_U179 ; P2_R2096_U181
g26072 nand P2_U2643 P2_R2096_U64 ; P2_R2096_U182
g26073 nand P2_U2651 P2_R2096_U65 ; P2_R2096_U183
g26074 nand P2_U2643 P2_R2096_U64 ; P2_R2096_U184
g26075 nand P2_U2651 P2_R2096_U65 ; P2_R2096_U185
g26076 nand P2_R2096_U185 P2_R2096_U184 ; P2_R2096_U186
g26077 nand P2_R2096_U102 P2_R2096_U103 ; P2_R2096_U187
g26078 nand P2_R2096_U135 P2_R2096_U186 ; P2_R2096_U188
g26079 nand P2_U2644 P2_R2096_U62 ; P2_R2096_U189
g26080 nand P2_U2652 P2_R2096_U63 ; P2_R2096_U190
g26081 nand P2_U2644 P2_R2096_U62 ; P2_R2096_U191
g26082 nand P2_U2652 P2_R2096_U63 ; P2_R2096_U192
g26083 nand P2_R2096_U192 P2_R2096_U191 ; P2_R2096_U193
g26084 nand P2_R2096_U104 P2_R2096_U105 ; P2_R2096_U194
g26085 nand P2_R2096_U131 P2_R2096_U193 ; P2_R2096_U195
g26086 nand P2_U2645 P2_R2096_U60 ; P2_R2096_U196
g26087 nand P2_U2653 P2_R2096_U61 ; P2_R2096_U197
g26088 nand P2_U2645 P2_R2096_U60 ; P2_R2096_U198
g26089 nand P2_U2653 P2_R2096_U61 ; P2_R2096_U199
g26090 nand P2_R2096_U199 P2_R2096_U198 ; P2_R2096_U200
g26091 nand P2_R2096_U106 P2_R2096_U107 ; P2_R2096_U201
g26092 nand P2_R2096_U127 P2_R2096_U200 ; P2_R2096_U202
g26093 nand P2_U2646 P2_R2096_U58 ; P2_R2096_U203
g26094 nand P2_U2654 P2_R2096_U59 ; P2_R2096_U204
g26095 nand P2_U2646 P2_R2096_U58 ; P2_R2096_U205
g26096 nand P2_U2654 P2_R2096_U59 ; P2_R2096_U206
g26097 nand P2_R2096_U206 P2_R2096_U205 ; P2_R2096_U207
g26098 nand P2_R2096_U108 P2_R2096_U109 ; P2_R2096_U208
g26099 nand P2_R2096_U123 P2_R2096_U207 ; P2_R2096_U209
g26100 nand P2_R2096_U30 P2_R2096_U22 ; P2_R2096_U210
g26101 nand P2_U2619 P2_R2096_U165 ; P2_R2096_U211
g26102 nand P2_U2647 P2_R2096_U56 ; P2_R2096_U212
g26103 nand P2_U2655 P2_R2096_U57 ; P2_R2096_U213
g26104 nand P2_U2647 P2_R2096_U56 ; P2_R2096_U214
g26105 nand P2_U2655 P2_R2096_U57 ; P2_R2096_U215
g26106 nand P2_R2096_U215 P2_R2096_U214 ; P2_R2096_U216
g26107 nand P2_R2096_U110 P2_R2096_U111 ; P2_R2096_U217
g26108 nand P2_R2096_U119 P2_R2096_U216 ; P2_R2096_U218
g26109 nand P2_R2096_U40 P2_R2096_U14 ; P2_R2096_U219
g26110 nand P2_R2096_U164 P2_U2620 ; P2_R2096_U220
g26111 nand P2_R2096_U41 P2_R2096_U13 ; P2_R2096_U221
g26112 nand P2_R2096_U163 P2_U2621 ; P2_R2096_U222
g26113 nand P2_R2096_U38 P2_R2096_U15 ; P2_R2096_U223
g26114 nand P2_R2096_U162 P2_U2622 ; P2_R2096_U224
g26115 nand P2_R2096_U42 P2_R2096_U12 ; P2_R2096_U225
g26116 nand P2_R2096_U161 P2_U2623 ; P2_R2096_U226
g26117 nand P2_R2096_U43 P2_R2096_U11 ; P2_R2096_U227
g26118 nand P2_R2096_U160 P2_U2624 ; P2_R2096_U228
g26119 nand P2_R2096_U44 P2_R2096_U10 ; P2_R2096_U229
g26120 nand P2_R2096_U159 P2_U2625 ; P2_R2096_U230
g26121 nand P2_R2096_U45 P2_R2096_U9 ; P2_R2096_U231
g26122 nand P2_R2096_U158 P2_U2626 ; P2_R2096_U232
g26123 nand P2_R2096_U39 P2_R2096_U8 ; P2_R2096_U233
g26124 nand P2_R2096_U157 P2_U2627 ; P2_R2096_U234
g26125 nand P2_R2096_U46 P2_R2096_U7 ; P2_R2096_U235
g26126 nand P2_R2096_U156 P2_U2628 ; P2_R2096_U236
g26127 nand P2_R2096_U36 P2_R2096_U16 ; P2_R2096_U237
g26128 nand P2_R2096_U155 P2_U2629 ; P2_R2096_U238
g26129 nand P2_U2648 P2_R2096_U112 ; P2_R2096_U239
g26130 nand P2_R2096_U169 P2_R2096_U54 ; P2_R2096_U240
g26131 nand P2_R2096_U240 P2_R2096_U239 ; P2_R2096_U241
g26132 nand P2_U2656 P2_R2096_U116 P2_R2096_U54 ; P2_R2096_U242
g26133 nand P2_R2096_U115 P2_U2648 ; P2_R2096_U243
g26134 nand P2_R2096_U47 P2_R2096_U6 ; P2_R2096_U244
g26135 nand P2_R2096_U154 P2_U2630 ; P2_R2096_U245
g26136 nand P2_R2096_U26 P2_R2096_U25 ; P2_R2096_U246
g26137 nand P2_R2096_U153 P2_U2631 ; P2_R2096_U247
g26138 nand P2_R2096_U48 P2_R2096_U5 ; P2_R2096_U248
g26139 nand P2_R2096_U152 P2_U2632 ; P2_R2096_U249
g26140 nand P2_R2096_U34 P2_R2096_U18 ; P2_R2096_U250
g26141 nand P2_R2096_U151 P2_U2633 ; P2_R2096_U251
g26142 nand P2_R2096_U35 P2_R2096_U17 ; P2_R2096_U252
g26143 nand P2_R2096_U150 P2_U2634 ; P2_R2096_U253
g26144 nand P2_R2096_U31 P2_R2096_U21 ; P2_R2096_U254
g26145 nand P2_R2096_U149 P2_U2635 ; P2_R2096_U255
g26146 nand P2_R2096_U32 P2_R2096_U20 ; P2_R2096_U256
g26147 nand P2_R2096_U148 P2_U2636 ; P2_R2096_U257
g26148 nand P2_R2096_U33 P2_R2096_U19 ; P2_R2096_U258
g26149 nand P2_R2096_U147 P2_U2637 ; P2_R2096_U259
g26150 nand P2_R2096_U27 P2_R2096_U24 ; P2_R2096_U260
g26151 nand P2_R2096_U146 P2_U2638 ; P2_R2096_U261
g26152 nand P2_R2096_U49 P2_R2096_U4 ; P2_R2096_U262
g26153 nand P2_R2096_U145 P2_U2639 ; P2_R2096_U263
g26154 nand P2_U2649 P2_R2096_U52 ; P2_R2096_U264
g26155 nand P2_U2657 P2_R2096_U53 ; P2_R2096_U265
g26156 nor P2_R2219_U25 P2_GTE_370_U8 ; P2_GTE_370_U6
g26157 and P2_R2219_U29 P2_GTE_370_U9 ; P2_GTE_370_U7
g26158 nor P2_R2219_U26 P2_R2219_U27 P2_R2219_U28 P2_GTE_370_U7 ; P2_GTE_370_U8
g26159 or P2_R2219_U8 P2_R2219_U30 ; P2_GTE_370_U9
g26160 and P2_LT_563_U27 P2_LT_563_U26 ; P2_LT_563_U6
g26161 not P2_U3620 ; P2_LT_563_U7
g26162 not P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_LT_563_U8
g26163 not P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_LT_563_U9
g26164 not P2_U3619 ; P2_LT_563_U10
g26165 not P2_U3618 ; P2_LT_563_U11
g26166 not P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_LT_563_U12
g26167 not P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_LT_563_U13
g26168 not P2_U3617 ; P2_LT_563_U14
g26169 not P2_U3621 ; P2_LT_563_U15
g26170 nand P2_U3620 P2_LT_563_U8 ; P2_LT_563_U16
g26171 nand P2_LT_563_U15 P2_LT_563_U16 P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_LT_563_U17
g26172 nand P2_LT_563_U7 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_LT_563_U18
g26173 nand P2_LT_563_U10 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_LT_563_U19
g26174 nand P2_LT_563_U18 P2_LT_563_U19 P2_LT_563_U17 ; P2_LT_563_U20
g26175 nand P2_U3619 P2_LT_563_U9 ; P2_LT_563_U21
g26176 nand P2_U3618 P2_LT_563_U12 ; P2_LT_563_U22
g26177 nand P2_LT_563_U21 P2_LT_563_U22 P2_LT_563_U20 ; P2_LT_563_U23
g26178 nand P2_LT_563_U11 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_LT_563_U24
g26179 nand P2_LT_563_U14 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_LT_563_U25
g26180 nand P2_LT_563_U24 P2_LT_563_U25 P2_LT_563_U23 ; P2_LT_563_U26
g26181 nand P2_U3617 P2_LT_563_U13 ; P2_LT_563_U27
g26182 nand P2_R2256_U31 P2_R2256_U46 ; P2_R2256_U4
g26183 and P2_R2256_U23 P2_R2256_U43 ; P2_R2256_U5
g26184 not P2_U3629 ; P2_R2256_U6
g26185 not P2_U3628 ; P2_R2256_U7
g26186 not P2_U3627 ; P2_R2256_U8
g26187 not P2_U3626 ; P2_R2256_U9
g26188 nand P2_U3626 P2_R2256_U25 ; P2_R2256_U10
g26189 not P2_U3625 ; P2_R2256_U11
g26190 nand P2_U3625 P2_R2256_U41 ; P2_R2256_U12
g26191 not P2_U3624 ; P2_R2256_U13
g26192 nand P2_U3624 P2_R2256_U42 ; P2_R2256_U14
g26193 not P2_U3622 ; P2_R2256_U15
g26194 not P2_U3623 ; P2_R2256_U16
g26195 nand P2_R2256_U48 P2_R2256_U47 ; P2_R2256_U17
g26196 nand P2_R2256_U50 P2_R2256_U49 ; P2_R2256_U18
g26197 nand P2_R2256_U52 P2_R2256_U51 ; P2_R2256_U19
g26198 nand P2_R2256_U54 P2_R2256_U53 ; P2_R2256_U20
g26199 nand P2_R2256_U70 P2_R2256_U69 ; P2_R2256_U21
g26200 nand P2_R2256_U63 P2_R2256_U62 ; P2_R2256_U22
g26201 and P2_U3622 P2_U3623 ; P2_R2256_U23
g26202 nand P2_U3623 P2_R2256_U43 ; P2_R2256_U24
g26203 nand P2_R2256_U39 P2_R2256_U38 ; P2_R2256_U25
g26204 and P2_R2256_U56 P2_R2256_U55 ; P2_R2256_U26
g26205 and P2_R2256_U58 P2_R2256_U57 ; P2_R2256_U27
g26206 nand P2_R2256_U30 P2_R2256_U35 ; P2_R2256_U28
g26207 nand P2_U7873 P2_U3629 ; P2_R2256_U29
g26208 nand P2_U7873 P2_U3629 P2_U3628 ; P2_R2256_U30
g26209 and P2_R2256_U68 P2_R2256_U67 ; P2_R2256_U31
g26210 not P2_R2256_U30 ; P2_R2256_U32
g26211 nand P2_U7873 P2_U3629 ; P2_R2256_U33
g26212 nand P2_R2256_U7 P2_R2256_U33 ; P2_R2256_U34
g26213 nand P2_U2616 P2_R2256_U34 ; P2_R2256_U35
g26214 not P2_R2256_U28 ; P2_R2256_U36
g26215 or P2_U3627 P2_U7873 ; P2_R2256_U37
g26216 nand P2_R2256_U37 P2_R2256_U28 ; P2_R2256_U38
g26217 nand P2_U7873 P2_U3627 ; P2_R2256_U39
g26218 not P2_R2256_U25 ; P2_R2256_U40
g26219 not P2_R2256_U10 ; P2_R2256_U41
g26220 not P2_R2256_U12 ; P2_R2256_U42
g26221 not P2_R2256_U14 ; P2_R2256_U43
g26222 not P2_R2256_U24 ; P2_R2256_U44
g26223 not P2_R2256_U29 ; P2_R2256_U45
g26224 nand P2_R2256_U66 P2_R2256_U7 ; P2_R2256_U46
g26225 nand P2_U3622 P2_R2256_U24 ; P2_R2256_U47
g26226 nand P2_R2256_U44 P2_R2256_U15 ; P2_R2256_U48
g26227 nand P2_U3623 P2_R2256_U14 ; P2_R2256_U49
g26228 nand P2_R2256_U43 P2_R2256_U16 ; P2_R2256_U50
g26229 nand P2_U3624 P2_R2256_U12 ; P2_R2256_U51
g26230 nand P2_R2256_U42 P2_R2256_U13 ; P2_R2256_U52
g26231 nand P2_U3625 P2_R2256_U10 ; P2_R2256_U53
g26232 nand P2_R2256_U41 P2_R2256_U11 ; P2_R2256_U54
g26233 nand P2_U3626 P2_R2256_U25 ; P2_R2256_U55
g26234 nand P2_R2256_U40 P2_R2256_U9 ; P2_R2256_U56
g26235 nand P2_U7873 P2_R2256_U8 ; P2_R2256_U57
g26236 nand P2_U3627 P2_U2616 ; P2_R2256_U58
g26237 nand P2_U7873 P2_R2256_U8 ; P2_R2256_U59
g26238 nand P2_U3627 P2_U2616 ; P2_R2256_U60
g26239 nand P2_R2256_U60 P2_R2256_U59 ; P2_R2256_U61
g26240 nand P2_R2256_U27 P2_R2256_U28 ; P2_R2256_U62
g26241 nand P2_R2256_U36 P2_R2256_U61 ; P2_R2256_U63
g26242 nand P2_U2616 P2_R2256_U29 ; P2_R2256_U64
g26243 nand P2_R2256_U45 P2_U7873 ; P2_R2256_U65
g26244 nand P2_R2256_U65 P2_R2256_U64 ; P2_R2256_U66
g26245 nand P2_U3628 P2_R2256_U33 P2_U7873 ; P2_R2256_U67
g26246 nand P2_R2256_U32 P2_U2616 ; P2_R2256_U68
g26247 nand P2_U7873 P2_R2256_U6 ; P2_R2256_U69
g26248 nand P2_U3629 P2_U2616 ; P2_R2256_U70
g26249 nand P2_R2238_U45 P2_R2238_U44 ; P2_R2238_U6
g26250 nand P2_R2238_U9 P2_R2238_U46 ; P2_R2238_U7
g26251 not P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_R2238_U8
g26252 nand P2_R2238_U18 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_R2238_U9
g26253 not P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_R2238_U10
g26254 not P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_R2238_U11
g26255 not P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_R2238_U12
g26256 not P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_R2238_U13
g26257 not P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_R2238_U14
g26258 not P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_R2238_U15
g26259 nand P2_R2238_U41 P2_R2238_U40 ; P2_R2238_U16
g26260 not P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_R2238_U17
g26261 not P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_R2238_U18
g26262 nand P2_R2238_U51 P2_R2238_U50 ; P2_R2238_U19
g26263 nand P2_R2238_U56 P2_R2238_U55 ; P2_R2238_U20
g26264 nand P2_R2238_U61 P2_R2238_U60 ; P2_R2238_U21
g26265 nand P2_R2238_U66 P2_R2238_U65 ; P2_R2238_U22
g26266 nand P2_R2238_U48 P2_R2238_U47 ; P2_R2238_U23
g26267 nand P2_R2238_U53 P2_R2238_U52 ; P2_R2238_U24
g26268 nand P2_R2238_U58 P2_R2238_U57 ; P2_R2238_U25
g26269 nand P2_R2238_U63 P2_R2238_U62 ; P2_R2238_U26
g26270 nand P2_R2238_U37 P2_R2238_U36 ; P2_R2238_U27
g26271 nand P2_R2238_U33 P2_R2238_U32 ; P2_R2238_U28
g26272 not P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_R2238_U29
g26273 not P2_R2238_U9 ; P2_R2238_U30
g26274 nand P2_R2238_U30 P2_R2238_U10 ; P2_R2238_U31
g26275 nand P2_R2238_U31 P2_R2238_U29 ; P2_R2238_U32
g26276 nand P2_R2238_U9 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_R2238_U33
g26277 not P2_R2238_U28 ; P2_R2238_U34
g26278 nand P2_R2238_U12 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_R2238_U35
g26279 nand P2_R2238_U35 P2_R2238_U28 ; P2_R2238_U36
g26280 nand P2_R2238_U11 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_R2238_U37
g26281 not P2_R2238_U27 ; P2_R2238_U38
g26282 nand P2_R2238_U14 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_R2238_U39
g26283 nand P2_R2238_U39 P2_R2238_U27 ; P2_R2238_U40
g26284 nand P2_R2238_U13 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_R2238_U41
g26285 not P2_R2238_U16 ; P2_R2238_U42
g26286 nand P2_R2238_U17 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_R2238_U43
g26287 nand P2_R2238_U42 P2_R2238_U43 ; P2_R2238_U44
g26288 nand P2_R2238_U15 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_R2238_U45
g26289 nand P2_R2238_U8 P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_R2238_U46
g26290 nand P2_R2238_U15 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_R2238_U47
g26291 nand P2_R2238_U17 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_R2238_U48
g26292 not P2_R2238_U23 ; P2_R2238_U49
g26293 nand P2_R2238_U49 P2_R2238_U42 ; P2_R2238_U50
g26294 nand P2_R2238_U23 P2_R2238_U16 ; P2_R2238_U51
g26295 nand P2_R2238_U14 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_R2238_U52
g26296 nand P2_R2238_U13 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_R2238_U53
g26297 not P2_R2238_U24 ; P2_R2238_U54
g26298 nand P2_R2238_U38 P2_R2238_U54 ; P2_R2238_U55
g26299 nand P2_R2238_U24 P2_R2238_U27 ; P2_R2238_U56
g26300 nand P2_R2238_U12 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_R2238_U57
g26301 nand P2_R2238_U11 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_R2238_U58
g26302 not P2_R2238_U25 ; P2_R2238_U59
g26303 nand P2_R2238_U34 P2_R2238_U59 ; P2_R2238_U60
g26304 nand P2_R2238_U25 P2_R2238_U28 ; P2_R2238_U61
g26305 nand P2_R2238_U10 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_R2238_U62
g26306 nand P2_R2238_U29 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_R2238_U63
g26307 not P2_R2238_U26 ; P2_R2238_U64
g26308 nand P2_R2238_U64 P2_R2238_U30 ; P2_R2238_U65
g26309 nand P2_R2238_U26 P2_R2238_U9 ; P2_R2238_U66
g26310 and P2_R1957_U126 P2_R1957_U27 ; P2_R1957_U6
g26311 and P2_R1957_U124 P2_R1957_U28 ; P2_R1957_U7
g26312 and P2_R1957_U122 P2_R1957_U29 ; P2_R1957_U8
g26313 and P2_R1957_U120 P2_R1957_U30 ; P2_R1957_U9
g26314 and P2_R1957_U118 P2_R1957_U31 ; P2_R1957_U10
g26315 and P2_R1957_U116 P2_R1957_U32 ; P2_R1957_U11
g26316 and P2_R1957_U114 P2_R1957_U33 ; P2_R1957_U12
g26317 and P2_R1957_U112 P2_R1957_U34 ; P2_R1957_U13
g26318 and P2_R1957_U110 P2_R1957_U35 ; P2_R1957_U14
g26319 and P2_R1957_U108 P2_R1957_U36 ; P2_R1957_U15
g26320 and P2_R1957_U106 P2_R1957_U37 ; P2_R1957_U16
g26321 and P2_R1957_U105 P2_R1957_U21 ; P2_R1957_U17
g26322 and P2_R1957_U92 P2_R1957_U22 ; P2_R1957_U18
g26323 and P2_R1957_U90 P2_R1957_U23 ; P2_R1957_U19
g26324 and P2_R1957_U88 P2_R1957_U24 ; P2_R1957_U20
g26325 or P2_U3682 P2_U3683 P2_U3671 ; P2_R1957_U21
g26326 nand P2_R1957_U51 P2_R1957_U83 ; P2_R1957_U22
g26327 nand P2_R1957_U84 P2_R1957_U56 P2_R1957_U26 ; P2_R1957_U23
g26328 nand P2_R1957_U85 P2_R1957_U54 P2_R1957_U25 ; P2_R1957_U24
g26329 not P2_U3654 ; P2_R1957_U25
g26330 not P2_U3656 ; P2_R1957_U26
g26331 nand P2_R1957_U52 P2_R1957_U86 P2_R1957_U48 ; P2_R1957_U27
g26332 nand P2_R1957_U93 P2_R1957_U81 P2_R1957_U47 ; P2_R1957_U28
g26333 nand P2_R1957_U94 P2_R1957_U79 P2_R1957_U46 ; P2_R1957_U29
g26334 nand P2_R1957_U95 P2_R1957_U77 P2_R1957_U45 ; P2_R1957_U30
g26335 nand P2_R1957_U96 P2_R1957_U75 P2_R1957_U44 ; P2_R1957_U31
g26336 nand P2_R1957_U97 P2_R1957_U73 P2_R1957_U43 ; P2_R1957_U32
g26337 nand P2_R1957_U98 P2_R1957_U69 P2_R1957_U42 ; P2_R1957_U33
g26338 nand P2_R1957_U99 P2_R1957_U67 P2_R1957_U41 ; P2_R1957_U34
g26339 nand P2_R1957_U100 P2_R1957_U65 P2_R1957_U40 ; P2_R1957_U35
g26340 nand P2_R1957_U101 P2_R1957_U63 P2_R1957_U39 ; P2_R1957_U36
g26341 nand P2_R1957_U102 P2_R1957_U38 ; P2_R1957_U37
g26342 not P2_U3661 ; P2_R1957_U38
g26343 not P2_U3662 ; P2_R1957_U39
g26344 not P2_U3664 ; P2_R1957_U40
g26345 not P2_U3666 ; P2_R1957_U41
g26346 not P2_U3668 ; P2_R1957_U42
g26347 not P2_U3670 ; P2_R1957_U43
g26348 not P2_U3673 ; P2_R1957_U44
g26349 not P2_U3675 ; P2_R1957_U45
g26350 not P2_U3677 ; P2_R1957_U46
g26351 not P2_U3679 ; P2_R1957_U47
g26352 not P2_U3681 ; P2_R1957_U48
g26353 nand P2_R1957_U149 P2_R1957_U148 ; P2_R1957_U49
g26354 nand P2_R1957_U137 P2_R1957_U136 ; P2_R1957_U50
g26355 nor P2_U3660 P2_U3658 ; P2_R1957_U51
g26356 not P2_U3653 ; P2_R1957_U52
g26357 and P2_R1957_U129 P2_R1957_U128 ; P2_R1957_U53
g26358 not P2_U3655 ; P2_R1957_U54
g26359 and P2_R1957_U131 P2_R1957_U130 ; P2_R1957_U55
g26360 not P2_U3657 ; P2_R1957_U56
g26361 and P2_R1957_U133 P2_R1957_U132 ; P2_R1957_U57
g26362 not P2_U3660 ; P2_R1957_U58
g26363 and P2_R1957_U135 P2_R1957_U134 ; P2_R1957_U59
g26364 not P2_U3647 ; P2_R1957_U60
g26365 not P2_U3659 ; P2_R1957_U61
g26366 and P2_R1957_U139 P2_R1957_U138 ; P2_R1957_U62
g26367 not P2_U3663 ; P2_R1957_U63
g26368 and P2_R1957_U141 P2_R1957_U140 ; P2_R1957_U64
g26369 not P2_U3665 ; P2_R1957_U65
g26370 and P2_R1957_U143 P2_R1957_U142 ; P2_R1957_U66
g26371 not P2_U3667 ; P2_R1957_U67
g26372 and P2_R1957_U145 P2_R1957_U144 ; P2_R1957_U68
g26373 not P2_U3669 ; P2_R1957_U69
g26374 and P2_R1957_U147 P2_R1957_U146 ; P2_R1957_U70
g26375 not P2_U3682 ; P2_R1957_U71
g26376 not P2_U3683 ; P2_R1957_U72
g26377 not P2_U3672 ; P2_R1957_U73
g26378 and P2_R1957_U151 P2_R1957_U150 ; P2_R1957_U74
g26379 not P2_U3674 ; P2_R1957_U75
g26380 and P2_R1957_U153 P2_R1957_U152 ; P2_R1957_U76
g26381 not P2_U3676 ; P2_R1957_U77
g26382 and P2_R1957_U155 P2_R1957_U154 ; P2_R1957_U78
g26383 not P2_U3678 ; P2_R1957_U79
g26384 and P2_R1957_U157 P2_R1957_U156 ; P2_R1957_U80
g26385 not P2_U3680 ; P2_R1957_U81
g26386 and P2_R1957_U159 P2_R1957_U158 ; P2_R1957_U82
g26387 not P2_R1957_U21 ; P2_R1957_U83
g26388 not P2_R1957_U22 ; P2_R1957_U84
g26389 not P2_R1957_U23 ; P2_R1957_U85
g26390 not P2_R1957_U24 ; P2_R1957_U86
g26391 nand P2_R1957_U85 P2_R1957_U54 ; P2_R1957_U87
g26392 nand P2_U3654 P2_R1957_U87 ; P2_R1957_U88
g26393 nand P2_R1957_U84 P2_R1957_U56 ; P2_R1957_U89
g26394 nand P2_U3656 P2_R1957_U89 ; P2_R1957_U90
g26395 nand P2_R1957_U83 P2_R1957_U58 ; P2_R1957_U91
g26396 nand P2_U3658 P2_R1957_U91 ; P2_R1957_U92
g26397 not P2_R1957_U27 ; P2_R1957_U93
g26398 not P2_R1957_U28 ; P2_R1957_U94
g26399 not P2_R1957_U29 ; P2_R1957_U95
g26400 not P2_R1957_U30 ; P2_R1957_U96
g26401 not P2_R1957_U31 ; P2_R1957_U97
g26402 not P2_R1957_U32 ; P2_R1957_U98
g26403 not P2_R1957_U33 ; P2_R1957_U99
g26404 not P2_R1957_U34 ; P2_R1957_U100
g26405 not P2_R1957_U35 ; P2_R1957_U101
g26406 not P2_R1957_U36 ; P2_R1957_U102
g26407 not P2_R1957_U37 ; P2_R1957_U103
g26408 or P2_U3682 P2_U3683 ; P2_R1957_U104
g26409 nand P2_U3671 P2_R1957_U104 ; P2_R1957_U105
g26410 nand P2_U3661 P2_R1957_U36 ; P2_R1957_U106
g26411 nand P2_R1957_U101 P2_R1957_U63 ; P2_R1957_U107
g26412 nand P2_U3662 P2_R1957_U107 ; P2_R1957_U108
g26413 nand P2_R1957_U100 P2_R1957_U65 ; P2_R1957_U109
g26414 nand P2_U3664 P2_R1957_U109 ; P2_R1957_U110
g26415 nand P2_R1957_U99 P2_R1957_U67 ; P2_R1957_U111
g26416 nand P2_U3666 P2_R1957_U111 ; P2_R1957_U112
g26417 nand P2_R1957_U98 P2_R1957_U69 ; P2_R1957_U113
g26418 nand P2_U3668 P2_R1957_U113 ; P2_R1957_U114
g26419 nand P2_R1957_U97 P2_R1957_U73 ; P2_R1957_U115
g26420 nand P2_U3670 P2_R1957_U115 ; P2_R1957_U116
g26421 nand P2_R1957_U96 P2_R1957_U75 ; P2_R1957_U117
g26422 nand P2_U3673 P2_R1957_U117 ; P2_R1957_U118
g26423 nand P2_R1957_U95 P2_R1957_U77 ; P2_R1957_U119
g26424 nand P2_U3675 P2_R1957_U119 ; P2_R1957_U120
g26425 nand P2_R1957_U94 P2_R1957_U79 ; P2_R1957_U121
g26426 nand P2_U3677 P2_R1957_U121 ; P2_R1957_U122
g26427 nand P2_R1957_U93 P2_R1957_U81 ; P2_R1957_U123
g26428 nand P2_U3679 P2_R1957_U123 ; P2_R1957_U124
g26429 nand P2_R1957_U86 P2_R1957_U52 ; P2_R1957_U125
g26430 nand P2_U3681 P2_R1957_U125 ; P2_R1957_U126
g26431 nand P2_R1957_U103 P2_R1957_U61 ; P2_R1957_U127
g26432 nand P2_U3653 P2_R1957_U24 ; P2_R1957_U128
g26433 nand P2_R1957_U86 P2_R1957_U52 ; P2_R1957_U129
g26434 nand P2_U3655 P2_R1957_U23 ; P2_R1957_U130
g26435 nand P2_R1957_U85 P2_R1957_U54 ; P2_R1957_U131
g26436 nand P2_U3657 P2_R1957_U22 ; P2_R1957_U132
g26437 nand P2_R1957_U84 P2_R1957_U56 ; P2_R1957_U133
g26438 nand P2_U3660 P2_R1957_U21 ; P2_R1957_U134
g26439 nand P2_R1957_U83 P2_R1957_U58 ; P2_R1957_U135
g26440 nand P2_R1957_U127 P2_R1957_U60 ; P2_R1957_U136
g26441 nand P2_R1957_U103 P2_R1957_U61 P2_U3647 ; P2_R1957_U137
g26442 nand P2_U3659 P2_R1957_U37 ; P2_R1957_U138
g26443 nand P2_R1957_U103 P2_R1957_U61 ; P2_R1957_U139
g26444 nand P2_U3663 P2_R1957_U35 ; P2_R1957_U140
g26445 nand P2_R1957_U101 P2_R1957_U63 ; P2_R1957_U141
g26446 nand P2_U3665 P2_R1957_U34 ; P2_R1957_U142
g26447 nand P2_R1957_U100 P2_R1957_U65 ; P2_R1957_U143
g26448 nand P2_U3667 P2_R1957_U33 ; P2_R1957_U144
g26449 nand P2_R1957_U99 P2_R1957_U67 ; P2_R1957_U145
g26450 nand P2_U3669 P2_R1957_U32 ; P2_R1957_U146
g26451 nand P2_R1957_U98 P2_R1957_U69 ; P2_R1957_U147
g26452 nand P2_U3682 P2_R1957_U72 ; P2_R1957_U148
g26453 nand P2_U3683 P2_R1957_U71 ; P2_R1957_U149
g26454 nand P2_U3672 P2_R1957_U31 ; P2_R1957_U150
g26455 nand P2_R1957_U97 P2_R1957_U73 ; P2_R1957_U151
g26456 nand P2_U3674 P2_R1957_U30 ; P2_R1957_U152
g26457 nand P2_R1957_U96 P2_R1957_U75 ; P2_R1957_U153
g26458 nand P2_U3676 P2_R1957_U29 ; P2_R1957_U154
g26459 nand P2_R1957_U95 P2_R1957_U77 ; P2_R1957_U155
g26460 nand P2_U3678 P2_R1957_U28 ; P2_R1957_U156
g26461 nand P2_R1957_U94 P2_R1957_U79 ; P2_R1957_U157
g26462 nand P2_U3680 P2_R1957_U27 ; P2_R1957_U158
g26463 nand P2_R1957_U93 P2_R1957_U81 ; P2_R1957_U159
g26464 and P2_R2278_U399 P2_R2278_U398 ; P2_R2278_U4
g26465 and P2_R2278_U161 P2_R2278_U309 P2_R2278_U206 ; P2_R2278_U5
g26466 nand P2_R2278_U490 P2_R2278_U489 P2_R2278_U345 ; P2_R2278_U6
g26467 not P2_U3631 ; P2_R2278_U7
g26468 not P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2278_U8
g26469 not P2_U3633 ; P2_R2278_U9
g26470 not P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2278_U10
g26471 not P2_U3635 ; P2_R2278_U11
g26472 not P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2278_U12
g26473 not P2_U3638 ; P2_R2278_U13
g26474 not P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_R2278_U14
g26475 nand P2_U3638 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_R2278_U15
g26476 not P2_U3637 ; P2_R2278_U16
g26477 not P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2278_U17
g26478 not P2_U3636 ; P2_R2278_U18
g26479 not P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2278_U19
g26480 nand P2_U3636 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2278_U20
g26481 not P2_U3634 ; P2_R2278_U21
g26482 not P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2278_U22
g26483 nand P2_U3634 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2278_U23
g26484 not P2_U3632 ; P2_R2278_U24
g26485 not P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2278_U25
g26486 nand P2_U3632 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2278_U26
g26487 not P2_U3630 ; P2_R2278_U27
g26488 not P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2278_U28
g26489 not P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2278_U29
g26490 not P2_U2812 ; P2_R2278_U30
g26491 not P2_U2793 ; P2_R2278_U31
g26492 not P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2278_U32
g26493 not P2_U2792 ; P2_R2278_U33
g26494 not P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2278_U34
g26495 not P2_U2797 ; P2_R2278_U35
g26496 not P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2278_U36
g26497 not P2_U2799 ; P2_R2278_U37
g26498 not P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2278_U38
g26499 not P2_U2801 ; P2_R2278_U39
g26500 not P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2278_U40
g26501 not P2_U2804 ; P2_R2278_U41
g26502 not P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2278_U42
g26503 not P2_U2806 ; P2_R2278_U43
g26504 not P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2278_U44
g26505 not P2_U2808 ; P2_R2278_U45
g26506 not P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2278_U46
g26507 not P2_U2810 ; P2_R2278_U47
g26508 not P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2278_U48
g26509 nand P2_U3630 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2278_U49
g26510 not P2_U2811 ; P2_R2278_U50
g26511 not P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2278_U51
g26512 nand P2_U2811 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2278_U52
g26513 not P2_U2809 ; P2_R2278_U53
g26514 not P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2278_U54
g26515 nand P2_U2809 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2278_U55
g26516 not P2_U2807 ; P2_R2278_U56
g26517 not P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2278_U57
g26518 nand P2_U2807 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2278_U58
g26519 not P2_U2805 ; P2_R2278_U59
g26520 not P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2278_U60
g26521 nand P2_U2805 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2278_U61
g26522 not P2_U2802 ; P2_R2278_U62
g26523 not P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2278_U63
g26524 not P2_U2803 ; P2_R2278_U64
g26525 not P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2278_U65
g26526 not P2_U2800 ; P2_R2278_U66
g26527 not P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2278_U67
g26528 nand P2_U2800 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2278_U68
g26529 not P2_U2798 ; P2_R2278_U69
g26530 not P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2278_U70
g26531 nand P2_U2798 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2278_U71
g26532 not P2_U2796 ; P2_R2278_U72
g26533 not P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2278_U73
g26534 not P2_U2794 ; P2_R2278_U74
g26535 not P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2278_U75
g26536 not P2_U2795 ; P2_R2278_U76
g26537 not P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2278_U77
g26538 nand P2_U2795 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2278_U78
g26539 not P2_U2791 ; P2_R2278_U79
g26540 not P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2278_U80
g26541 nand P2_R2278_U340 P2_R2278_U297 ; P2_R2278_U81
g26542 nand P2_U3637 P2_R2278_U208 ; P2_R2278_U82
g26543 nand P2_R2278_U562 P2_R2278_U561 ; P2_R2278_U83
g26544 nand P2_R2278_U352 P2_R2278_U351 ; P2_R2278_U84
g26545 nand P2_R2278_U359 P2_R2278_U358 ; P2_R2278_U85
g26546 nand P2_R2278_U366 P2_R2278_U365 ; P2_R2278_U86
g26547 nand P2_R2278_U373 P2_R2278_U372 ; P2_R2278_U87
g26548 nand P2_R2278_U380 P2_R2278_U379 ; P2_R2278_U88
g26549 nand P2_R2278_U387 P2_R2278_U386 ; P2_R2278_U89
g26550 nand P2_R2278_U394 P2_R2278_U393 ; P2_R2278_U90
g26551 nand P2_R2278_U408 P2_R2278_U407 ; P2_R2278_U91
g26552 nand P2_R2278_U415 P2_R2278_U414 ; P2_R2278_U92
g26553 nand P2_R2278_U422 P2_R2278_U421 ; P2_R2278_U93
g26554 nand P2_R2278_U429 P2_R2278_U428 ; P2_R2278_U94
g26555 nand P2_R2278_U436 P2_R2278_U435 ; P2_R2278_U95
g26556 nand P2_R2278_U443 P2_R2278_U442 ; P2_R2278_U96
g26557 nand P2_R2278_U450 P2_R2278_U449 ; P2_R2278_U97
g26558 nand P2_R2278_U457 P2_R2278_U456 ; P2_R2278_U98
g26559 nand P2_R2278_U464 P2_R2278_U463 ; P2_R2278_U99
g26560 nand P2_R2278_U471 P2_R2278_U470 ; P2_R2278_U100
g26561 nand P2_R2278_U478 P2_R2278_U477 ; P2_R2278_U101
g26562 nand P2_R2278_U485 P2_R2278_U484 ; P2_R2278_U102
g26563 nand P2_R2278_U497 P2_R2278_U496 ; P2_R2278_U103
g26564 nand P2_R2278_U504 P2_R2278_U503 ; P2_R2278_U104
g26565 nand P2_R2278_U511 P2_R2278_U510 ; P2_R2278_U105
g26566 nand P2_R2278_U518 P2_R2278_U517 ; P2_R2278_U106
g26567 nand P2_R2278_U525 P2_R2278_U524 ; P2_R2278_U107
g26568 nand P2_R2278_U532 P2_R2278_U531 ; P2_R2278_U108
g26569 nand P2_R2278_U539 P2_R2278_U538 ; P2_R2278_U109
g26570 nand P2_R2278_U546 P2_R2278_U545 ; P2_R2278_U110
g26571 nand P2_R2278_U553 P2_R2278_U552 ; P2_R2278_U111
g26572 nand P2_R2278_U560 P2_R2278_U559 ; P2_R2278_U112
g26573 and P2_R2278_U210 P2_R2278_U314 ; P2_R2278_U113
g26574 and P2_R2278_U313 P2_R2278_U215 ; P2_R2278_U114
g26575 and P2_R2278_U217 P2_R2278_U221 ; P2_R2278_U115
g26576 and P2_R2278_U316 P2_R2278_U222 ; P2_R2278_U116
g26577 and P2_R2278_U224 P2_R2278_U228 ; P2_R2278_U117
g26578 and P2_R2278_U318 P2_R2278_U229 ; P2_R2278_U118
g26579 and P2_R2278_U231 P2_R2278_U235 ; P2_R2278_U119
g26580 and P2_R2278_U320 P2_R2278_U236 ; P2_R2278_U120
g26581 and P2_R2278_U238 P2_R2278_U242 ; P2_R2278_U121
g26582 and P2_R2278_U322 P2_R2278_U243 ; P2_R2278_U122
g26583 and P2_R2278_U245 P2_R2278_U249 ; P2_R2278_U123
g26584 and P2_R2278_U324 P2_R2278_U250 ; P2_R2278_U124
g26585 and P2_R2278_U252 P2_R2278_U256 ; P2_R2278_U125
g26586 and P2_R2278_U326 P2_R2278_U257 ; P2_R2278_U126
g26587 and P2_R2278_U259 P2_R2278_U263 ; P2_R2278_U127
g26588 and P2_R2278_U328 P2_R2278_U264 ; P2_R2278_U128
g26589 and P2_R2278_U273 P2_R2278_U270 ; P2_R2278_U129
g26590 and P2_R2278_U331 P2_R2278_U273 ; P2_R2278_U130
g26591 and P2_R2278_U334 P2_R2278_U274 ; P2_R2278_U131
g26592 and P2_R2278_U276 P2_R2278_U280 ; P2_R2278_U132
g26593 and P2_R2278_U336 P2_R2278_U281 ; P2_R2278_U133
g26594 and P2_R2278_U283 P2_R2278_U287 ; P2_R2278_U134
g26595 and P2_R2278_U338 P2_R2278_U288 ; P2_R2278_U135
g26596 and P2_R2278_U299 P2_R2278_U296 P2_R2278_U292 ; P2_R2278_U136
g26597 and P2_R2278_U304 P2_R2278_U300 ; P2_R2278_U137
g26598 and P2_R2278_U307 P2_R2278_U302 ; P2_R2278_U138
g26599 and P2_R2278_U397 P2_R2278_U138 ; P2_R2278_U139
g26600 and P2_R2278_U343 P2_R2278_U300 ; P2_R2278_U140
g26601 and P2_R2278_U4 P2_R2278_U142 ; P2_R2278_U141
g26602 and P2_R2278_U304 P2_R2278_U306 ; P2_R2278_U142
g26603 and P2_R2278_U292 P2_R2278_U296 ; P2_R2278_U143
g26604 and P2_R2278_U266 P2_R2278_U270 ; P2_R2278_U144
g26605 and P2_R2278_U347 P2_R2278_U346 ; P2_R2278_U145
g26606 nand P2_R2278_U49 P2_R2278_U232 ; P2_R2278_U146
g26607 and P2_R2278_U354 P2_R2278_U353 ; P2_R2278_U147
g26608 nand P2_R2278_U118 P2_R2278_U317 ; P2_R2278_U148
g26609 and P2_R2278_U361 P2_R2278_U360 ; P2_R2278_U149
g26610 nand P2_R2278_U26 P2_R2278_U225 ; P2_R2278_U150
g26611 and P2_R2278_U368 P2_R2278_U367 ; P2_R2278_U151
g26612 nand P2_R2278_U116 P2_R2278_U315 ; P2_R2278_U152
g26613 and P2_R2278_U375 P2_R2278_U374 ; P2_R2278_U153
g26614 nand P2_R2278_U23 P2_R2278_U218 ; P2_R2278_U154
g26615 and P2_R2278_U382 P2_R2278_U381 ; P2_R2278_U155
g26616 nand P2_R2278_U114 P2_R2278_U312 ; P2_R2278_U156
g26617 and P2_R2278_U389 P2_R2278_U388 ; P2_R2278_U157
g26618 nand P2_R2278_U20 P2_R2278_U211 ; P2_R2278_U158
g26619 not P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_R2278_U159
g26620 not P2_U2790 ; P2_R2278_U160
g26621 and P2_R2278_U401 P2_R2278_U400 ; P2_R2278_U161
g26622 and P2_R2278_U403 P2_R2278_U402 ; P2_R2278_U162
g26623 nand P2_R2278_U304 P2_R2278_U303 ; P2_R2278_U163
g26624 and P2_R2278_U410 P2_R2278_U409 ; P2_R2278_U164
g26625 nand P2_R2278_U310 P2_R2278_U82 P2_R2278_U311 ; P2_R2278_U165
g26626 and P2_R2278_U417 P2_R2278_U416 ; P2_R2278_U166
g26627 nand P2_R2278_U140 P2_R2278_U342 ; P2_R2278_U167
g26628 and P2_R2278_U424 P2_R2278_U423 ; P2_R2278_U168
g26629 nand P2_R2278_U341 P2_R2278_U339 ; P2_R2278_U169
g26630 and P2_R2278_U431 P2_R2278_U430 ; P2_R2278_U170
g26631 nand P2_R2278_U78 P2_R2278_U293 ; P2_R2278_U171
g26632 and P2_R2278_U438 P2_R2278_U437 ; P2_R2278_U172
g26633 nand P2_R2278_U290 P2_R2278_U205 P2_R2278_U308 ; P2_R2278_U173
g26634 nand P2_R2278_U135 P2_R2278_U337 ; P2_R2278_U174
g26635 and P2_R2278_U452 P2_R2278_U451 ; P2_R2278_U175
g26636 nand P2_R2278_U71 P2_R2278_U284 ; P2_R2278_U176
g26637 and P2_R2278_U459 P2_R2278_U458 ; P2_R2278_U177
g26638 nand P2_R2278_U133 P2_R2278_U335 ; P2_R2278_U178
g26639 and P2_R2278_U466 P2_R2278_U465 ; P2_R2278_U179
g26640 nand P2_R2278_U68 P2_R2278_U277 ; P2_R2278_U180
g26641 and P2_R2278_U473 P2_R2278_U472 ; P2_R2278_U181
g26642 nand P2_R2278_U131 P2_R2278_U333 ; P2_R2278_U182
g26643 and P2_R2278_U480 P2_R2278_U479 ; P2_R2278_U183
g26644 nand P2_R2278_U330 P2_R2278_U329 ; P2_R2278_U184
g26645 and P2_R2278_U492 P2_R2278_U491 ; P2_R2278_U185
g26646 nand P2_R2278_U268 P2_R2278_U267 ; P2_R2278_U186
g26647 and P2_R2278_U499 P2_R2278_U498 ; P2_R2278_U187
g26648 nand P2_R2278_U128 P2_R2278_U327 ; P2_R2278_U188
g26649 and P2_R2278_U506 P2_R2278_U505 ; P2_R2278_U189
g26650 nand P2_R2278_U61 P2_R2278_U260 ; P2_R2278_U190
g26651 and P2_R2278_U513 P2_R2278_U512 ; P2_R2278_U191
g26652 nand P2_R2278_U126 P2_R2278_U325 ; P2_R2278_U192
g26653 and P2_R2278_U520 P2_R2278_U519 ; P2_R2278_U193
g26654 nand P2_R2278_U58 P2_R2278_U253 ; P2_R2278_U194
g26655 and P2_R2278_U527 P2_R2278_U526 ; P2_R2278_U195
g26656 nand P2_R2278_U124 P2_R2278_U323 ; P2_R2278_U196
g26657 and P2_R2278_U534 P2_R2278_U533 ; P2_R2278_U197
g26658 nand P2_R2278_U55 P2_R2278_U246 ; P2_R2278_U198
g26659 and P2_R2278_U541 P2_R2278_U540 ; P2_R2278_U199
g26660 nand P2_R2278_U122 P2_R2278_U321 ; P2_R2278_U200
g26661 and P2_R2278_U548 P2_R2278_U547 ; P2_R2278_U201
g26662 nand P2_R2278_U52 P2_R2278_U239 ; P2_R2278_U202
g26663 and P2_R2278_U555 P2_R2278_U554 ; P2_R2278_U203
g26664 nand P2_R2278_U120 P2_R2278_U319 ; P2_R2278_U204
g26665 nand P2_U2796 P2_R2278_U174 ; P2_R2278_U205
g26666 nand P2_R2278_U139 P2_R2278_U344 ; P2_R2278_U206
g26667 not P2_R2278_U82 ; P2_R2278_U207
g26668 not P2_R2278_U15 ; P2_R2278_U208
g26669 not P2_R2278_U165 ; P2_R2278_U209
g26670 or P2_U3636 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2278_U210
g26671 nand P2_R2278_U210 P2_R2278_U165 ; P2_R2278_U211
g26672 not P2_R2278_U20 ; P2_R2278_U212
g26673 not P2_R2278_U158 ; P2_R2278_U213
g26674 or P2_U3635 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2278_U214
g26675 nand P2_U3635 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2278_U215
g26676 not P2_R2278_U156 ; P2_R2278_U216
g26677 or P2_U3634 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2278_U217
g26678 nand P2_R2278_U217 P2_R2278_U156 ; P2_R2278_U218
g26679 not P2_R2278_U23 ; P2_R2278_U219
g26680 not P2_R2278_U154 ; P2_R2278_U220
g26681 or P2_U3633 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2278_U221
g26682 nand P2_U3633 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2278_U222
g26683 not P2_R2278_U152 ; P2_R2278_U223
g26684 or P2_U3632 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2278_U224
g26685 nand P2_R2278_U224 P2_R2278_U152 ; P2_R2278_U225
g26686 not P2_R2278_U26 ; P2_R2278_U226
g26687 not P2_R2278_U150 ; P2_R2278_U227
g26688 or P2_U3631 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2278_U228
g26689 nand P2_U3631 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2278_U229
g26690 not P2_R2278_U148 ; P2_R2278_U230
g26691 or P2_U3630 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2278_U231
g26692 nand P2_R2278_U231 P2_R2278_U148 ; P2_R2278_U232
g26693 not P2_R2278_U49 ; P2_R2278_U233
g26694 not P2_R2278_U146 ; P2_R2278_U234
g26695 or P2_U2812 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2278_U235
g26696 nand P2_U2812 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2278_U236
g26697 not P2_R2278_U204 ; P2_R2278_U237
g26698 or P2_U2811 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2278_U238
g26699 nand P2_R2278_U238 P2_R2278_U204 ; P2_R2278_U239
g26700 not P2_R2278_U52 ; P2_R2278_U240
g26701 not P2_R2278_U202 ; P2_R2278_U241
g26702 or P2_U2810 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2278_U242
g26703 nand P2_U2810 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2278_U243
g26704 not P2_R2278_U200 ; P2_R2278_U244
g26705 or P2_U2809 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2278_U245
g26706 nand P2_R2278_U245 P2_R2278_U200 ; P2_R2278_U246
g26707 not P2_R2278_U55 ; P2_R2278_U247
g26708 not P2_R2278_U198 ; P2_R2278_U248
g26709 or P2_U2808 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2278_U249
g26710 nand P2_U2808 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2278_U250
g26711 not P2_R2278_U196 ; P2_R2278_U251
g26712 or P2_U2807 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2278_U252
g26713 nand P2_R2278_U252 P2_R2278_U196 ; P2_R2278_U253
g26714 not P2_R2278_U58 ; P2_R2278_U254
g26715 not P2_R2278_U194 ; P2_R2278_U255
g26716 or P2_U2806 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2278_U256
g26717 nand P2_U2806 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2278_U257
g26718 not P2_R2278_U192 ; P2_R2278_U258
g26719 or P2_U2805 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2278_U259
g26720 nand P2_R2278_U259 P2_R2278_U192 ; P2_R2278_U260
g26721 not P2_R2278_U61 ; P2_R2278_U261
g26722 not P2_R2278_U190 ; P2_R2278_U262
g26723 or P2_U2804 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2278_U263
g26724 nand P2_U2804 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2278_U264
g26725 not P2_R2278_U188 ; P2_R2278_U265
g26726 or P2_U2803 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2278_U266
g26727 nand P2_R2278_U266 P2_R2278_U188 ; P2_R2278_U267
g26728 nand P2_U2803 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2278_U268
g26729 not P2_R2278_U186 ; P2_R2278_U269
g26730 or P2_U2802 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2278_U270
g26731 nand P2_U2802 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2278_U271
g26732 not P2_R2278_U184 ; P2_R2278_U272
g26733 or P2_U2801 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2278_U273
g26734 nand P2_U2801 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2278_U274
g26735 not P2_R2278_U182 ; P2_R2278_U275
g26736 or P2_U2800 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2278_U276
g26737 nand P2_R2278_U276 P2_R2278_U182 ; P2_R2278_U277
g26738 not P2_R2278_U68 ; P2_R2278_U278
g26739 not P2_R2278_U180 ; P2_R2278_U279
g26740 or P2_U2799 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2278_U280
g26741 nand P2_U2799 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2278_U281
g26742 not P2_R2278_U178 ; P2_R2278_U282
g26743 or P2_U2798 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2278_U283
g26744 nand P2_R2278_U283 P2_R2278_U178 ; P2_R2278_U284
g26745 not P2_R2278_U71 ; P2_R2278_U285
g26746 not P2_R2278_U176 ; P2_R2278_U286
g26747 or P2_U2797 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2278_U287
g26748 nand P2_U2797 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2278_U288
g26749 not P2_R2278_U174 ; P2_R2278_U289
g26750 nand P2_R2278_U174 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2278_U290
g26751 not P2_R2278_U173 ; P2_R2278_U291
g26752 or P2_U2795 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2278_U292
g26753 nand P2_R2278_U292 P2_R2278_U173 ; P2_R2278_U293
g26754 not P2_R2278_U78 ; P2_R2278_U294
g26755 not P2_R2278_U171 ; P2_R2278_U295
g26756 or P2_U2794 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2278_U296
g26757 nand P2_U2794 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2278_U297
g26758 not P2_R2278_U169 ; P2_R2278_U298
g26759 or P2_U2793 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2278_U299
g26760 nand P2_U2793 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2278_U300
g26761 not P2_R2278_U167 ; P2_R2278_U301
g26762 or P2_U2792 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2278_U302
g26763 nand P2_R2278_U302 P2_R2278_U167 ; P2_R2278_U303
g26764 nand P2_U2792 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2278_U304
g26765 not P2_R2278_U163 ; P2_R2278_U305
g26766 nand P2_U2791 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2278_U306
g26767 or P2_U2791 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2278_U307
g26768 nand P2_U2796 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2278_U308
g26769 nand P2_R2278_U303 P2_R2278_U141 ; P2_R2278_U309
g26770 nand P2_R2278_U208 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2278_U310
g26771 nand P2_U3637 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2278_U311
g26772 nand P2_R2278_U113 P2_R2278_U165 ; P2_R2278_U312
g26773 nand P2_R2278_U212 P2_R2278_U214 ; P2_R2278_U313
g26774 or P2_U3635 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2278_U314
g26775 nand P2_R2278_U115 P2_R2278_U156 ; P2_R2278_U315
g26776 nand P2_R2278_U219 P2_R2278_U221 ; P2_R2278_U316
g26777 nand P2_R2278_U117 P2_R2278_U152 ; P2_R2278_U317
g26778 nand P2_R2278_U226 P2_R2278_U228 ; P2_R2278_U318
g26779 nand P2_R2278_U119 P2_R2278_U148 ; P2_R2278_U319
g26780 nand P2_R2278_U233 P2_R2278_U235 ; P2_R2278_U320
g26781 nand P2_R2278_U121 P2_R2278_U204 ; P2_R2278_U321
g26782 nand P2_R2278_U240 P2_R2278_U242 ; P2_R2278_U322
g26783 nand P2_R2278_U123 P2_R2278_U200 ; P2_R2278_U323
g26784 nand P2_R2278_U247 P2_R2278_U249 ; P2_R2278_U324
g26785 nand P2_R2278_U125 P2_R2278_U196 ; P2_R2278_U325
g26786 nand P2_R2278_U254 P2_R2278_U256 ; P2_R2278_U326
g26787 nand P2_R2278_U127 P2_R2278_U192 ; P2_R2278_U327
g26788 nand P2_R2278_U261 P2_R2278_U263 ; P2_R2278_U328
g26789 nand P2_R2278_U144 P2_R2278_U188 ; P2_R2278_U329
g26790 nand P2_R2278_U331 P2_R2278_U332 ; P2_R2278_U330
g26791 or P2_U2802 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2278_U331
g26792 nand P2_R2278_U268 P2_R2278_U271 ; P2_R2278_U332
g26793 nand P2_R2278_U266 P2_R2278_U188 P2_R2278_U129 ; P2_R2278_U333
g26794 nand P2_R2278_U130 P2_R2278_U332 ; P2_R2278_U334
g26795 nand P2_R2278_U132 P2_R2278_U182 ; P2_R2278_U335
g26796 nand P2_R2278_U278 P2_R2278_U280 ; P2_R2278_U336
g26797 nand P2_R2278_U134 P2_R2278_U178 ; P2_R2278_U337
g26798 nand P2_R2278_U285 P2_R2278_U287 ; P2_R2278_U338
g26799 nand P2_R2278_U143 P2_R2278_U173 ; P2_R2278_U339
g26800 nand P2_R2278_U294 P2_R2278_U296 ; P2_R2278_U340
g26801 not P2_R2278_U81 ; P2_R2278_U341
g26802 nand P2_R2278_U173 P2_R2278_U136 ; P2_R2278_U342
g26803 nand P2_R2278_U81 P2_R2278_U299 ; P2_R2278_U343
g26804 nand P2_R2278_U343 P2_R2278_U342 P2_R2278_U137 ; P2_R2278_U344
g26805 nand P2_R2278_U207 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2278_U345
g26806 nand P2_R2278_U30 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2278_U346
g26807 nand P2_U2812 P2_R2278_U29 ; P2_R2278_U347
g26808 nand P2_R2278_U30 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_R2278_U348
g26809 nand P2_U2812 P2_R2278_U29 ; P2_R2278_U349
g26810 nand P2_R2278_U349 P2_R2278_U348 ; P2_R2278_U350
g26811 nand P2_R2278_U145 P2_R2278_U146 ; P2_R2278_U351
g26812 nand P2_R2278_U234 P2_R2278_U350 ; P2_R2278_U352
g26813 nand P2_R2278_U27 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2278_U353
g26814 nand P2_U3630 P2_R2278_U28 ; P2_R2278_U354
g26815 nand P2_R2278_U27 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_R2278_U355
g26816 nand P2_U3630 P2_R2278_U28 ; P2_R2278_U356
g26817 nand P2_R2278_U356 P2_R2278_U355 ; P2_R2278_U357
g26818 nand P2_R2278_U147 P2_R2278_U148 ; P2_R2278_U358
g26819 nand P2_R2278_U230 P2_R2278_U357 ; P2_R2278_U359
g26820 nand P2_R2278_U7 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2278_U360
g26821 nand P2_U3631 P2_R2278_U8 ; P2_R2278_U361
g26822 nand P2_R2278_U7 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_R2278_U362
g26823 nand P2_U3631 P2_R2278_U8 ; P2_R2278_U363
g26824 nand P2_R2278_U363 P2_R2278_U362 ; P2_R2278_U364
g26825 nand P2_R2278_U149 P2_R2278_U150 ; P2_R2278_U365
g26826 nand P2_R2278_U227 P2_R2278_U364 ; P2_R2278_U366
g26827 nand P2_R2278_U24 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2278_U367
g26828 nand P2_U3632 P2_R2278_U25 ; P2_R2278_U368
g26829 nand P2_R2278_U24 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_R2278_U369
g26830 nand P2_U3632 P2_R2278_U25 ; P2_R2278_U370
g26831 nand P2_R2278_U370 P2_R2278_U369 ; P2_R2278_U371
g26832 nand P2_R2278_U151 P2_R2278_U152 ; P2_R2278_U372
g26833 nand P2_R2278_U223 P2_R2278_U371 ; P2_R2278_U373
g26834 nand P2_R2278_U9 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2278_U374
g26835 nand P2_U3633 P2_R2278_U10 ; P2_R2278_U375
g26836 nand P2_R2278_U9 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_R2278_U376
g26837 nand P2_U3633 P2_R2278_U10 ; P2_R2278_U377
g26838 nand P2_R2278_U377 P2_R2278_U376 ; P2_R2278_U378
g26839 nand P2_R2278_U153 P2_R2278_U154 ; P2_R2278_U379
g26840 nand P2_R2278_U220 P2_R2278_U378 ; P2_R2278_U380
g26841 nand P2_R2278_U21 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2278_U381
g26842 nand P2_U3634 P2_R2278_U22 ; P2_R2278_U382
g26843 nand P2_R2278_U21 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_R2278_U383
g26844 nand P2_U3634 P2_R2278_U22 ; P2_R2278_U384
g26845 nand P2_R2278_U384 P2_R2278_U383 ; P2_R2278_U385
g26846 nand P2_R2278_U155 P2_R2278_U156 ; P2_R2278_U386
g26847 nand P2_R2278_U216 P2_R2278_U385 ; P2_R2278_U387
g26848 nand P2_R2278_U11 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2278_U388
g26849 nand P2_U3635 P2_R2278_U12 ; P2_R2278_U389
g26850 nand P2_R2278_U11 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_R2278_U390
g26851 nand P2_U3635 P2_R2278_U12 ; P2_R2278_U391
g26852 nand P2_R2278_U391 P2_R2278_U390 ; P2_R2278_U392
g26853 nand P2_R2278_U157 P2_R2278_U158 ; P2_R2278_U393
g26854 nand P2_R2278_U213 P2_R2278_U392 ; P2_R2278_U394
g26855 nand P2_R2278_U160 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_R2278_U395
g26856 nand P2_U2790 P2_R2278_U159 ; P2_R2278_U396
g26857 nand P2_R2278_U396 P2_R2278_U395 ; P2_R2278_U397
g26858 nand P2_R2278_U160 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_R2278_U398
g26859 nand P2_U2790 P2_R2278_U159 ; P2_R2278_U399
g26860 nand P2_R2278_U4 P2_R2278_U79 P2_R2278_U80 ; P2_R2278_U400
g26861 nand P2_U2791 P2_R2278_U397 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2278_U401
g26862 nand P2_R2278_U79 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2278_U402
g26863 nand P2_U2791 P2_R2278_U80 ; P2_R2278_U403
g26864 nand P2_R2278_U79 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_R2278_U404
g26865 nand P2_U2791 P2_R2278_U80 ; P2_R2278_U405
g26866 nand P2_R2278_U405 P2_R2278_U404 ; P2_R2278_U406
g26867 nand P2_R2278_U162 P2_R2278_U163 ; P2_R2278_U407
g26868 nand P2_R2278_U305 P2_R2278_U406 ; P2_R2278_U408
g26869 nand P2_R2278_U18 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2278_U409
g26870 nand P2_U3636 P2_R2278_U19 ; P2_R2278_U410
g26871 nand P2_R2278_U18 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_R2278_U411
g26872 nand P2_U3636 P2_R2278_U19 ; P2_R2278_U412
g26873 nand P2_R2278_U412 P2_R2278_U411 ; P2_R2278_U413
g26874 nand P2_R2278_U164 P2_R2278_U165 ; P2_R2278_U414
g26875 nand P2_R2278_U209 P2_R2278_U413 ; P2_R2278_U415
g26876 nand P2_R2278_U33 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2278_U416
g26877 nand P2_U2792 P2_R2278_U34 ; P2_R2278_U417
g26878 nand P2_R2278_U33 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_R2278_U418
g26879 nand P2_U2792 P2_R2278_U34 ; P2_R2278_U419
g26880 nand P2_R2278_U419 P2_R2278_U418 ; P2_R2278_U420
g26881 nand P2_R2278_U166 P2_R2278_U167 ; P2_R2278_U421
g26882 nand P2_R2278_U301 P2_R2278_U420 ; P2_R2278_U422
g26883 nand P2_R2278_U31 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2278_U423
g26884 nand P2_U2793 P2_R2278_U32 ; P2_R2278_U424
g26885 nand P2_R2278_U31 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_R2278_U425
g26886 nand P2_U2793 P2_R2278_U32 ; P2_R2278_U426
g26887 nand P2_R2278_U426 P2_R2278_U425 ; P2_R2278_U427
g26888 nand P2_R2278_U168 P2_R2278_U169 ; P2_R2278_U428
g26889 nand P2_R2278_U298 P2_R2278_U427 ; P2_R2278_U429
g26890 nand P2_R2278_U74 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2278_U430
g26891 nand P2_U2794 P2_R2278_U75 ; P2_R2278_U431
g26892 nand P2_R2278_U74 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_R2278_U432
g26893 nand P2_U2794 P2_R2278_U75 ; P2_R2278_U433
g26894 nand P2_R2278_U433 P2_R2278_U432 ; P2_R2278_U434
g26895 nand P2_R2278_U170 P2_R2278_U171 ; P2_R2278_U435
g26896 nand P2_R2278_U295 P2_R2278_U434 ; P2_R2278_U436
g26897 nand P2_R2278_U76 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2278_U437
g26898 nand P2_U2795 P2_R2278_U77 ; P2_R2278_U438
g26899 nand P2_R2278_U76 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_R2278_U439
g26900 nand P2_U2795 P2_R2278_U77 ; P2_R2278_U440
g26901 nand P2_R2278_U440 P2_R2278_U439 ; P2_R2278_U441
g26902 nand P2_R2278_U172 P2_R2278_U173 ; P2_R2278_U442
g26903 nand P2_R2278_U291 P2_R2278_U441 ; P2_R2278_U443
g26904 nand P2_R2278_U174 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2278_U444
g26905 nand P2_R2278_U289 P2_R2278_U73 ; P2_R2278_U445
g26906 nand P2_R2278_U174 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_R2278_U446
g26907 nand P2_R2278_U289 P2_R2278_U73 ; P2_R2278_U447
g26908 nand P2_R2278_U447 P2_R2278_U446 ; P2_R2278_U448
g26909 nand P2_R2278_U445 P2_R2278_U444 P2_R2278_U72 ; P2_R2278_U449
g26910 nand P2_R2278_U448 P2_U2796 ; P2_R2278_U450
g26911 nand P2_R2278_U35 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2278_U451
g26912 nand P2_U2797 P2_R2278_U36 ; P2_R2278_U452
g26913 nand P2_R2278_U35 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_R2278_U453
g26914 nand P2_U2797 P2_R2278_U36 ; P2_R2278_U454
g26915 nand P2_R2278_U454 P2_R2278_U453 ; P2_R2278_U455
g26916 nand P2_R2278_U175 P2_R2278_U176 ; P2_R2278_U456
g26917 nand P2_R2278_U286 P2_R2278_U455 ; P2_R2278_U457
g26918 nand P2_R2278_U69 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2278_U458
g26919 nand P2_U2798 P2_R2278_U70 ; P2_R2278_U459
g26920 nand P2_R2278_U69 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_R2278_U460
g26921 nand P2_U2798 P2_R2278_U70 ; P2_R2278_U461
g26922 nand P2_R2278_U461 P2_R2278_U460 ; P2_R2278_U462
g26923 nand P2_R2278_U177 P2_R2278_U178 ; P2_R2278_U463
g26924 nand P2_R2278_U282 P2_R2278_U462 ; P2_R2278_U464
g26925 nand P2_R2278_U37 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2278_U465
g26926 nand P2_U2799 P2_R2278_U38 ; P2_R2278_U466
g26927 nand P2_R2278_U37 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_R2278_U467
g26928 nand P2_U2799 P2_R2278_U38 ; P2_R2278_U468
g26929 nand P2_R2278_U468 P2_R2278_U467 ; P2_R2278_U469
g26930 nand P2_R2278_U179 P2_R2278_U180 ; P2_R2278_U470
g26931 nand P2_R2278_U279 P2_R2278_U469 ; P2_R2278_U471
g26932 nand P2_R2278_U66 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2278_U472
g26933 nand P2_U2800 P2_R2278_U67 ; P2_R2278_U473
g26934 nand P2_R2278_U66 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_R2278_U474
g26935 nand P2_U2800 P2_R2278_U67 ; P2_R2278_U475
g26936 nand P2_R2278_U475 P2_R2278_U474 ; P2_R2278_U476
g26937 nand P2_R2278_U181 P2_R2278_U182 ; P2_R2278_U477
g26938 nand P2_R2278_U275 P2_R2278_U476 ; P2_R2278_U478
g26939 nand P2_R2278_U39 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2278_U479
g26940 nand P2_U2801 P2_R2278_U40 ; P2_R2278_U480
g26941 nand P2_R2278_U39 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_R2278_U481
g26942 nand P2_U2801 P2_R2278_U40 ; P2_R2278_U482
g26943 nand P2_R2278_U482 P2_R2278_U481 ; P2_R2278_U483
g26944 nand P2_R2278_U183 P2_R2278_U184 ; P2_R2278_U484
g26945 nand P2_R2278_U272 P2_R2278_U483 ; P2_R2278_U485
g26946 nand P2_R2278_U15 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_R2278_U486
g26947 nand P2_R2278_U208 P2_R2278_U17 ; P2_R2278_U487
g26948 nand P2_R2278_U487 P2_R2278_U486 ; P2_R2278_U488
g26949 nand P2_R2278_U15 P2_R2278_U17 P2_U3637 ; P2_R2278_U489
g26950 nand P2_R2278_U488 P2_R2278_U16 ; P2_R2278_U490
g26951 nand P2_R2278_U62 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2278_U491
g26952 nand P2_U2802 P2_R2278_U63 ; P2_R2278_U492
g26953 nand P2_R2278_U62 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_R2278_U493
g26954 nand P2_U2802 P2_R2278_U63 ; P2_R2278_U494
g26955 nand P2_R2278_U494 P2_R2278_U493 ; P2_R2278_U495
g26956 nand P2_R2278_U185 P2_R2278_U186 ; P2_R2278_U496
g26957 nand P2_R2278_U269 P2_R2278_U495 ; P2_R2278_U497
g26958 nand P2_R2278_U64 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2278_U498
g26959 nand P2_U2803 P2_R2278_U65 ; P2_R2278_U499
g26960 nand P2_R2278_U64 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_R2278_U500
g26961 nand P2_U2803 P2_R2278_U65 ; P2_R2278_U501
g26962 nand P2_R2278_U501 P2_R2278_U500 ; P2_R2278_U502
g26963 nand P2_R2278_U187 P2_R2278_U188 ; P2_R2278_U503
g26964 nand P2_R2278_U265 P2_R2278_U502 ; P2_R2278_U504
g26965 nand P2_R2278_U41 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2278_U505
g26966 nand P2_U2804 P2_R2278_U42 ; P2_R2278_U506
g26967 nand P2_R2278_U41 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_R2278_U507
g26968 nand P2_U2804 P2_R2278_U42 ; P2_R2278_U508
g26969 nand P2_R2278_U508 P2_R2278_U507 ; P2_R2278_U509
g26970 nand P2_R2278_U189 P2_R2278_U190 ; P2_R2278_U510
g26971 nand P2_R2278_U262 P2_R2278_U509 ; P2_R2278_U511
g26972 nand P2_R2278_U59 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2278_U512
g26973 nand P2_U2805 P2_R2278_U60 ; P2_R2278_U513
g26974 nand P2_R2278_U59 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_R2278_U514
g26975 nand P2_U2805 P2_R2278_U60 ; P2_R2278_U515
g26976 nand P2_R2278_U515 P2_R2278_U514 ; P2_R2278_U516
g26977 nand P2_R2278_U191 P2_R2278_U192 ; P2_R2278_U517
g26978 nand P2_R2278_U258 P2_R2278_U516 ; P2_R2278_U518
g26979 nand P2_R2278_U43 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2278_U519
g26980 nand P2_U2806 P2_R2278_U44 ; P2_R2278_U520
g26981 nand P2_R2278_U43 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_R2278_U521
g26982 nand P2_U2806 P2_R2278_U44 ; P2_R2278_U522
g26983 nand P2_R2278_U522 P2_R2278_U521 ; P2_R2278_U523
g26984 nand P2_R2278_U193 P2_R2278_U194 ; P2_R2278_U524
g26985 nand P2_R2278_U255 P2_R2278_U523 ; P2_R2278_U525
g26986 nand P2_R2278_U56 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2278_U526
g26987 nand P2_U2807 P2_R2278_U57 ; P2_R2278_U527
g26988 nand P2_R2278_U56 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_R2278_U528
g26989 nand P2_U2807 P2_R2278_U57 ; P2_R2278_U529
g26990 nand P2_R2278_U529 P2_R2278_U528 ; P2_R2278_U530
g26991 nand P2_R2278_U195 P2_R2278_U196 ; P2_R2278_U531
g26992 nand P2_R2278_U251 P2_R2278_U530 ; P2_R2278_U532
g26993 nand P2_R2278_U45 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2278_U533
g26994 nand P2_U2808 P2_R2278_U46 ; P2_R2278_U534
g26995 nand P2_R2278_U45 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_R2278_U535
g26996 nand P2_U2808 P2_R2278_U46 ; P2_R2278_U536
g26997 nand P2_R2278_U536 P2_R2278_U535 ; P2_R2278_U537
g26998 nand P2_R2278_U197 P2_R2278_U198 ; P2_R2278_U538
g26999 nand P2_R2278_U248 P2_R2278_U537 ; P2_R2278_U539
g27000 nand P2_R2278_U53 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2278_U540
g27001 nand P2_U2809 P2_R2278_U54 ; P2_R2278_U541
g27002 nand P2_R2278_U53 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_R2278_U542
g27003 nand P2_U2809 P2_R2278_U54 ; P2_R2278_U543
g27004 nand P2_R2278_U543 P2_R2278_U542 ; P2_R2278_U544
g27005 nand P2_R2278_U199 P2_R2278_U200 ; P2_R2278_U545
g27006 nand P2_R2278_U244 P2_R2278_U544 ; P2_R2278_U546
g27007 nand P2_R2278_U47 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2278_U547
g27008 nand P2_U2810 P2_R2278_U48 ; P2_R2278_U548
g27009 nand P2_R2278_U47 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_R2278_U549
g27010 nand P2_U2810 P2_R2278_U48 ; P2_R2278_U550
g27011 nand P2_R2278_U550 P2_R2278_U549 ; P2_R2278_U551
g27012 nand P2_R2278_U201 P2_R2278_U202 ; P2_R2278_U552
g27013 nand P2_R2278_U241 P2_R2278_U551 ; P2_R2278_U553
g27014 nand P2_R2278_U50 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2278_U554
g27015 nand P2_U2811 P2_R2278_U51 ; P2_R2278_U555
g27016 nand P2_R2278_U50 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_R2278_U556
g27017 nand P2_U2811 P2_R2278_U51 ; P2_R2278_U557
g27018 nand P2_R2278_U557 P2_R2278_U556 ; P2_R2278_U558
g27019 nand P2_R2278_U203 P2_R2278_U204 ; P2_R2278_U559
g27020 nand P2_R2278_U237 P2_R2278_U558 ; P2_R2278_U560
g27021 nand P2_R2278_U13 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_R2278_U561
g27022 nand P2_U3638 P2_R2278_U14 ; P2_R2278_U562
g27023 nand P2_SUB_450_U43 P2_SUB_450_U42 ; P2_SUB_450_U6
g27024 nand P2_SUB_450_U16 P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P2_SUB_450_U7
g27025 not P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_SUB_450_U8
g27026 not P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_SUB_450_U9
g27027 not P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_SUB_450_U10
g27028 not P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_SUB_450_U11
g27029 not P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_SUB_450_U12
g27030 not P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_SUB_450_U13
g27031 nand P2_SUB_450_U39 P2_SUB_450_U38 ; P2_SUB_450_U14
g27032 not P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_SUB_450_U15
g27033 not P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P2_SUB_450_U16
g27034 nand P2_SUB_450_U48 P2_SUB_450_U47 ; P2_SUB_450_U17
g27035 nand P2_SUB_450_U53 P2_SUB_450_U52 ; P2_SUB_450_U18
g27036 nand P2_SUB_450_U58 P2_SUB_450_U57 ; P2_SUB_450_U19
g27037 nand P2_SUB_450_U63 P2_SUB_450_U62 ; P2_SUB_450_U20
g27038 nand P2_SUB_450_U45 P2_SUB_450_U44 ; P2_SUB_450_U21
g27039 nand P2_SUB_450_U50 P2_SUB_450_U49 ; P2_SUB_450_U22
g27040 nand P2_SUB_450_U55 P2_SUB_450_U54 ; P2_SUB_450_U23
g27041 nand P2_SUB_450_U60 P2_SUB_450_U59 ; P2_SUB_450_U24
g27042 nand P2_SUB_450_U35 P2_SUB_450_U34 ; P2_SUB_450_U25
g27043 nand P2_SUB_450_U31 P2_SUB_450_U30 ; P2_SUB_450_U26
g27044 not P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_SUB_450_U27
g27045 not P2_SUB_450_U7 ; P2_SUB_450_U28
g27046 nand P2_SUB_450_U28 P2_SUB_450_U8 ; P2_SUB_450_U29
g27047 nand P2_SUB_450_U29 P2_SUB_450_U27 ; P2_SUB_450_U30
g27048 nand P2_SUB_450_U7 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_SUB_450_U31
g27049 not P2_SUB_450_U26 ; P2_SUB_450_U32
g27050 nand P2_SUB_450_U10 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_SUB_450_U33
g27051 nand P2_SUB_450_U33 P2_SUB_450_U26 ; P2_SUB_450_U34
g27052 nand P2_SUB_450_U9 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_SUB_450_U35
g27053 not P2_SUB_450_U25 ; P2_SUB_450_U36
g27054 nand P2_SUB_450_U12 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_SUB_450_U37
g27055 nand P2_SUB_450_U37 P2_SUB_450_U25 ; P2_SUB_450_U38
g27056 nand P2_SUB_450_U11 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_SUB_450_U39
g27057 not P2_SUB_450_U14 ; P2_SUB_450_U40
g27058 nand P2_SUB_450_U15 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_SUB_450_U41
g27059 nand P2_SUB_450_U40 P2_SUB_450_U41 ; P2_SUB_450_U42
g27060 nand P2_SUB_450_U13 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_SUB_450_U43
g27061 nand P2_SUB_450_U13 P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P2_SUB_450_U44
g27062 nand P2_SUB_450_U15 P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P2_SUB_450_U45
g27063 not P2_SUB_450_U21 ; P2_SUB_450_U46
g27064 nand P2_SUB_450_U46 P2_SUB_450_U40 ; P2_SUB_450_U47
g27065 nand P2_SUB_450_U21 P2_SUB_450_U14 ; P2_SUB_450_U48
g27066 nand P2_SUB_450_U12 P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P2_SUB_450_U49
g27067 nand P2_SUB_450_U11 P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P2_SUB_450_U50
g27068 not P2_SUB_450_U22 ; P2_SUB_450_U51
g27069 nand P2_SUB_450_U36 P2_SUB_450_U51 ; P2_SUB_450_U52
g27070 nand P2_SUB_450_U22 P2_SUB_450_U25 ; P2_SUB_450_U53
g27071 nand P2_SUB_450_U10 P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P2_SUB_450_U54
g27072 nand P2_SUB_450_U9 P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P2_SUB_450_U55
g27073 not P2_SUB_450_U23 ; P2_SUB_450_U56
g27074 nand P2_SUB_450_U32 P2_SUB_450_U56 ; P2_SUB_450_U57
g27075 nand P2_SUB_450_U23 P2_SUB_450_U26 ; P2_SUB_450_U58
g27076 nand P2_SUB_450_U8 P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P2_SUB_450_U59
g27077 nand P2_SUB_450_U27 P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P2_SUB_450_U60
g27078 not P2_SUB_450_U24 ; P2_SUB_450_U61
g27079 nand P2_SUB_450_U61 P2_SUB_450_U28 ; P2_SUB_450_U62
g27080 nand P2_SUB_450_U24 P2_SUB_450_U7 ; P2_SUB_450_U63
g27081 nor P2_U3648 P2_R2088_U7 ; P2_R2088_U6
g27082 nor P2_U3648 P2_U3649 P2_U3650 P2_U3652 P2_U3651 ; P2_R2088_U7
g27083 not P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_ADD_394_U4
g27084 nand P2_ADD_394_U94 P2_ADD_394_U125 ; P2_ADD_394_U5
g27085 not P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_394_U6
g27086 not P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_394_U7
g27087 nand P2_ADD_394_U94 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_394_U8
g27088 not P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_394_U9
g27089 nand P2_ADD_394_U98 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_394_U10
g27090 not P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_394_U11
g27091 not P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_394_U12
g27092 nand P2_ADD_394_U99 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_394_U13
g27093 nand P2_ADD_394_U100 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_394_U14
g27094 not P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_394_U15
g27095 nand P2_ADD_394_U101 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_394_U16
g27096 not P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_394_U17
g27097 nand P2_ADD_394_U102 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_394_U18
g27098 not P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_ADD_394_U19
g27099 nand P2_ADD_394_U103 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_ADD_394_U20
g27100 not P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_ADD_394_U21
g27101 nand P2_ADD_394_U104 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_ADD_394_U22
g27102 not P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_ADD_394_U23
g27103 nand P2_ADD_394_U105 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_ADD_394_U24
g27104 not P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_ADD_394_U25
g27105 nand P2_ADD_394_U106 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_ADD_394_U26
g27106 not P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_ADD_394_U27
g27107 nand P2_ADD_394_U107 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_ADD_394_U28
g27108 not P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_ADD_394_U29
g27109 nand P2_ADD_394_U108 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_ADD_394_U30
g27110 not P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_ADD_394_U31
g27111 nand P2_ADD_394_U109 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_ADD_394_U32
g27112 not P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_ADD_394_U33
g27113 nand P2_ADD_394_U110 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_ADD_394_U34
g27114 not P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_ADD_394_U35
g27115 nand P2_ADD_394_U111 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_ADD_394_U36
g27116 not P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_ADD_394_U37
g27117 nand P2_ADD_394_U112 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_ADD_394_U38
g27118 not P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_ADD_394_U39
g27119 nand P2_ADD_394_U113 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_ADD_394_U40
g27120 not P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_ADD_394_U41
g27121 nand P2_ADD_394_U114 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_ADD_394_U42
g27122 not P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_ADD_394_U43
g27123 nand P2_ADD_394_U115 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_ADD_394_U44
g27124 not P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_ADD_394_U45
g27125 nand P2_ADD_394_U116 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_ADD_394_U46
g27126 not P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_ADD_394_U47
g27127 nand P2_ADD_394_U117 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_ADD_394_U48
g27128 not P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_ADD_394_U49
g27129 nand P2_ADD_394_U118 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_ADD_394_U50
g27130 not P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_ADD_394_U51
g27131 nand P2_ADD_394_U119 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_ADD_394_U52
g27132 not P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_ADD_394_U53
g27133 nand P2_ADD_394_U120 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_ADD_394_U54
g27134 not P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_ADD_394_U55
g27135 nand P2_ADD_394_U121 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_ADD_394_U56
g27136 not P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_ADD_394_U57
g27137 nand P2_ADD_394_U122 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_ADD_394_U58
g27138 not P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_ADD_394_U59
g27139 not P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_394_U60
g27140 nand P2_ADD_394_U123 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_ADD_394_U61
g27141 not P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_394_U62
g27142 nand P2_ADD_394_U128 P2_ADD_394_U127 ; P2_ADD_394_U63
g27143 nand P2_ADD_394_U130 P2_ADD_394_U129 ; P2_ADD_394_U64
g27144 nand P2_ADD_394_U132 P2_ADD_394_U131 ; P2_ADD_394_U65
g27145 nand P2_ADD_394_U134 P2_ADD_394_U133 ; P2_ADD_394_U66
g27146 nand P2_ADD_394_U136 P2_ADD_394_U135 ; P2_ADD_394_U67
g27147 nand P2_ADD_394_U138 P2_ADD_394_U137 ; P2_ADD_394_U68
g27148 nand P2_ADD_394_U140 P2_ADD_394_U139 ; P2_ADD_394_U69
g27149 nand P2_ADD_394_U142 P2_ADD_394_U141 ; P2_ADD_394_U70
g27150 nand P2_ADD_394_U144 P2_ADD_394_U143 ; P2_ADD_394_U71
g27151 nand P2_ADD_394_U146 P2_ADD_394_U145 ; P2_ADD_394_U72
g27152 nand P2_ADD_394_U148 P2_ADD_394_U147 ; P2_ADD_394_U73
g27153 nand P2_ADD_394_U150 P2_ADD_394_U149 ; P2_ADD_394_U74
g27154 nand P2_ADD_394_U152 P2_ADD_394_U151 ; P2_ADD_394_U75
g27155 nand P2_ADD_394_U154 P2_ADD_394_U153 ; P2_ADD_394_U76
g27156 nand P2_ADD_394_U156 P2_ADD_394_U155 ; P2_ADD_394_U77
g27157 nand P2_ADD_394_U158 P2_ADD_394_U157 ; P2_ADD_394_U78
g27158 nand P2_ADD_394_U160 P2_ADD_394_U159 ; P2_ADD_394_U79
g27159 nand P2_ADD_394_U162 P2_ADD_394_U161 ; P2_ADD_394_U80
g27160 nand P2_ADD_394_U164 P2_ADD_394_U163 ; P2_ADD_394_U81
g27161 nand P2_ADD_394_U166 P2_ADD_394_U165 ; P2_ADD_394_U82
g27162 nand P2_ADD_394_U168 P2_ADD_394_U167 ; P2_ADD_394_U83
g27163 nand P2_ADD_394_U170 P2_ADD_394_U169 ; P2_ADD_394_U84
g27164 nand P2_ADD_394_U174 P2_ADD_394_U173 ; P2_ADD_394_U85
g27165 nand P2_ADD_394_U176 P2_ADD_394_U175 ; P2_ADD_394_U86
g27166 nand P2_ADD_394_U178 P2_ADD_394_U177 ; P2_ADD_394_U87
g27167 nand P2_ADD_394_U180 P2_ADD_394_U179 ; P2_ADD_394_U88
g27168 nand P2_ADD_394_U182 P2_ADD_394_U181 ; P2_ADD_394_U89
g27169 nand P2_ADD_394_U184 P2_ADD_394_U183 ; P2_ADD_394_U90
g27170 nand P2_ADD_394_U186 P2_ADD_394_U185 ; P2_ADD_394_U91
g27171 not P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_ADD_394_U92
g27172 nand P2_ADD_394_U124 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_394_U93
g27173 nand P2_ADD_394_U62 P2_ADD_394_U96 ; P2_ADD_394_U94
g27174 and P2_ADD_394_U172 P2_ADD_394_U171 ; P2_ADD_394_U95
g27175 nand P2_INSTADDRPOINTER_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_394_U96
g27176 not P2_ADD_394_U94 ; P2_ADD_394_U97
g27177 not P2_ADD_394_U8 ; P2_ADD_394_U98
g27178 not P2_ADD_394_U10 ; P2_ADD_394_U99
g27179 not P2_ADD_394_U13 ; P2_ADD_394_U100
g27180 not P2_ADD_394_U14 ; P2_ADD_394_U101
g27181 not P2_ADD_394_U16 ; P2_ADD_394_U102
g27182 not P2_ADD_394_U18 ; P2_ADD_394_U103
g27183 not P2_ADD_394_U20 ; P2_ADD_394_U104
g27184 not P2_ADD_394_U22 ; P2_ADD_394_U105
g27185 not P2_ADD_394_U24 ; P2_ADD_394_U106
g27186 not P2_ADD_394_U26 ; P2_ADD_394_U107
g27187 not P2_ADD_394_U28 ; P2_ADD_394_U108
g27188 not P2_ADD_394_U30 ; P2_ADD_394_U109
g27189 not P2_ADD_394_U32 ; P2_ADD_394_U110
g27190 not P2_ADD_394_U34 ; P2_ADD_394_U111
g27191 not P2_ADD_394_U36 ; P2_ADD_394_U112
g27192 not P2_ADD_394_U38 ; P2_ADD_394_U113
g27193 not P2_ADD_394_U40 ; P2_ADD_394_U114
g27194 not P2_ADD_394_U42 ; P2_ADD_394_U115
g27195 not P2_ADD_394_U44 ; P2_ADD_394_U116
g27196 not P2_ADD_394_U46 ; P2_ADD_394_U117
g27197 not P2_ADD_394_U48 ; P2_ADD_394_U118
g27198 not P2_ADD_394_U50 ; P2_ADD_394_U119
g27199 not P2_ADD_394_U52 ; P2_ADD_394_U120
g27200 not P2_ADD_394_U54 ; P2_ADD_394_U121
g27201 not P2_ADD_394_U56 ; P2_ADD_394_U122
g27202 not P2_ADD_394_U58 ; P2_ADD_394_U123
g27203 not P2_ADD_394_U61 ; P2_ADD_394_U124
g27204 nand P2_INSTADDRPOINTER_REG_0__SCAN_IN P2_INSTADDRPOINTER_REG_1__SCAN_IN P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_394_U125
g27205 not P2_ADD_394_U93 ; P2_ADD_394_U126
g27206 nand P2_ADD_394_U13 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_394_U127
g27207 nand P2_ADD_394_U100 P2_ADD_394_U12 ; P2_ADD_394_U128
g27208 nand P2_ADD_394_U61 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_394_U129
g27209 nand P2_ADD_394_U124 P2_ADD_394_U60 ; P2_ADD_394_U130
g27210 nand P2_ADD_394_U58 P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_ADD_394_U131
g27211 nand P2_ADD_394_U123 P2_ADD_394_U59 ; P2_ADD_394_U132
g27212 nand P2_ADD_394_U48 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_ADD_394_U133
g27213 nand P2_ADD_394_U118 P2_ADD_394_U49 ; P2_ADD_394_U134
g27214 nand P2_ADD_394_U34 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_ADD_394_U135
g27215 nand P2_ADD_394_U111 P2_ADD_394_U35 ; P2_ADD_394_U136
g27216 nand P2_ADD_394_U40 P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_ADD_394_U137
g27217 nand P2_ADD_394_U114 P2_ADD_394_U41 ; P2_ADD_394_U138
g27218 nand P2_ADD_394_U26 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_ADD_394_U139
g27219 nand P2_ADD_394_U107 P2_ADD_394_U27 ; P2_ADD_394_U140
g27220 nand P2_ADD_394_U18 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_ADD_394_U141
g27221 nand P2_ADD_394_U103 P2_ADD_394_U19 ; P2_ADD_394_U142
g27222 nand P2_ADD_394_U44 P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_ADD_394_U143
g27223 nand P2_ADD_394_U116 P2_ADD_394_U45 ; P2_ADD_394_U144
g27224 nand P2_ADD_394_U36 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_ADD_394_U145
g27225 nand P2_ADD_394_U112 P2_ADD_394_U37 ; P2_ADD_394_U146
g27226 nand P2_ADD_394_U22 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_ADD_394_U147
g27227 nand P2_ADD_394_U105 P2_ADD_394_U23 ; P2_ADD_394_U148
g27228 nand P2_ADD_394_U52 P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_ADD_394_U149
g27229 nand P2_ADD_394_U120 P2_ADD_394_U53 ; P2_ADD_394_U150
g27230 nand P2_ADD_394_U30 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_ADD_394_U151
g27231 nand P2_ADD_394_U109 P2_ADD_394_U31 ; P2_ADD_394_U152
g27232 nand P2_ADD_394_U8 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_394_U153
g27233 nand P2_ADD_394_U98 P2_ADD_394_U9 ; P2_ADD_394_U154
g27234 nand P2_ADD_394_U54 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_ADD_394_U155
g27235 nand P2_ADD_394_U121 P2_ADD_394_U55 ; P2_ADD_394_U156
g27236 nand P2_ADD_394_U28 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_ADD_394_U157
g27237 nand P2_ADD_394_U108 P2_ADD_394_U29 ; P2_ADD_394_U158
g27238 nand P2_ADD_394_U10 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_394_U159
g27239 nand P2_ADD_394_U99 P2_ADD_394_U11 ; P2_ADD_394_U160
g27240 nand P2_ADD_394_U16 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_394_U161
g27241 nand P2_ADD_394_U102 P2_ADD_394_U17 ; P2_ADD_394_U162
g27242 nand P2_ADD_394_U46 P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_ADD_394_U163
g27243 nand P2_ADD_394_U117 P2_ADD_394_U47 ; P2_ADD_394_U164
g27244 nand P2_ADD_394_U38 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_ADD_394_U165
g27245 nand P2_ADD_394_U113 P2_ADD_394_U39 ; P2_ADD_394_U166
g27246 nand P2_ADD_394_U20 P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_ADD_394_U167
g27247 nand P2_ADD_394_U104 P2_ADD_394_U21 ; P2_ADD_394_U168
g27248 nand P2_ADD_394_U93 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_ADD_394_U169
g27249 nand P2_ADD_394_U126 P2_ADD_394_U92 ; P2_ADD_394_U170
g27250 nand P2_ADD_394_U94 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_394_U171
g27251 nand P2_ADD_394_U97 P2_ADD_394_U7 ; P2_ADD_394_U172
g27252 nand P2_ADD_394_U4 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_394_U173
g27253 nand P2_ADD_394_U6 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_ADD_394_U174
g27254 nand P2_ADD_394_U56 P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_ADD_394_U175
g27255 nand P2_ADD_394_U122 P2_ADD_394_U57 ; P2_ADD_394_U176
g27256 nand P2_ADD_394_U42 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_ADD_394_U177
g27257 nand P2_ADD_394_U115 P2_ADD_394_U43 ; P2_ADD_394_U178
g27258 nand P2_ADD_394_U24 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_ADD_394_U179
g27259 nand P2_ADD_394_U106 P2_ADD_394_U25 ; P2_ADD_394_U180
g27260 nand P2_ADD_394_U14 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_394_U181
g27261 nand P2_ADD_394_U101 P2_ADD_394_U15 ; P2_ADD_394_U182
g27262 nand P2_ADD_394_U50 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_ADD_394_U183
g27263 nand P2_ADD_394_U119 P2_ADD_394_U51 ; P2_ADD_394_U184
g27264 nand P2_ADD_394_U32 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_ADD_394_U185
g27265 nand P2_ADD_394_U110 P2_ADD_394_U33 ; P2_ADD_394_U186
g27266 and P2_R2267_U133 P2_R2267_U31 ; P2_R2267_U6
g27267 and P2_R2267_U131 P2_R2267_U32 ; P2_R2267_U7
g27268 and P2_R2267_U129 P2_R2267_U33 ; P2_R2267_U8
g27269 and P2_R2267_U127 P2_R2267_U34 ; P2_R2267_U9
g27270 and P2_R2267_U125 P2_R2267_U35 ; P2_R2267_U10
g27271 and P2_R2267_U123 P2_R2267_U36 ; P2_R2267_U11
g27272 and P2_R2267_U121 P2_R2267_U37 ; P2_R2267_U12
g27273 and P2_R2267_U119 P2_R2267_U38 ; P2_R2267_U13
g27274 and P2_R2267_U117 P2_R2267_U39 ; P2_R2267_U14
g27275 and P2_R2267_U115 P2_R2267_U40 ; P2_R2267_U15
g27276 and P2_R2267_U113 P2_R2267_U62 ; P2_R2267_U16
g27277 and P2_R2267_U101 P2_R2267_U24 ; P2_R2267_U17
g27278 and P2_R2267_U99 P2_R2267_U25 ; P2_R2267_U18
g27279 and P2_R2267_U97 P2_R2267_U26 ; P2_R2267_U19
g27280 and P2_R2267_U95 P2_R2267_U30 ; P2_R2267_U20
g27281 nand P2_R2267_U77 P2_R2267_U134 ; P2_R2267_U21
g27282 not P2_U3646 ; P2_R2267_U22
g27283 nand P2_R2267_U76 P2_R2267_U77 ; P2_R2267_U23
g27284 nand P2_R2267_U89 P2_R2267_U64 P2_R2267_U29 ; P2_R2267_U24
g27285 nand P2_R2267_U90 P2_R2267_U59 P2_R2267_U28 ; P2_R2267_U25
g27286 nand P2_R2267_U91 P2_R2267_U57 P2_R2267_U27 ; P2_R2267_U26
g27287 not P2_U3639 ; P2_R2267_U27
g27288 not P2_U3641 ; P2_R2267_U28
g27289 not P2_U3643 ; P2_R2267_U29
g27290 nand P2_R2267_U44 P2_R2267_U92 ; P2_R2267_U30
g27291 nand P2_R2267_U45 P2_R2267_U93 ; P2_R2267_U31
g27292 nand P2_R2267_U46 P2_R2267_U102 ; P2_R2267_U32
g27293 nand P2_R2267_U47 P2_R2267_U103 ; P2_R2267_U33
g27294 nand P2_R2267_U48 P2_R2267_U104 ; P2_R2267_U34
g27295 nand P2_R2267_U49 P2_R2267_U105 ; P2_R2267_U35
g27296 nand P2_R2267_U50 P2_R2267_U106 ; P2_R2267_U36
g27297 nand P2_R2267_U51 P2_R2267_U107 ; P2_R2267_U37
g27298 nand P2_R2267_U52 P2_R2267_U108 ; P2_R2267_U38
g27299 nand P2_R2267_U53 P2_R2267_U109 ; P2_R2267_U39
g27300 nand P2_R2267_U54 P2_R2267_U110 ; P2_R2267_U40
g27301 not P2_U2767 ; P2_R2267_U41
g27302 not P2_U2617 ; P2_R2267_U42
g27303 nand P2_R2267_U156 P2_R2267_U155 ; P2_R2267_U43
g27304 nor P2_U2789 P2_U2788 ; P2_R2267_U44
g27305 nor P2_U2787 P2_U2786 ; P2_R2267_U45
g27306 nor P2_U2785 P2_U2784 ; P2_R2267_U46
g27307 nor P2_U2783 P2_U2782 ; P2_R2267_U47
g27308 nor P2_U2781 P2_U2780 ; P2_R2267_U48
g27309 nor P2_U2779 P2_U2778 ; P2_R2267_U49
g27310 nor P2_U2777 P2_U2776 ; P2_R2267_U50
g27311 nor P2_U2775 P2_U2774 ; P2_R2267_U51
g27312 nor P2_U2773 P2_U2772 ; P2_R2267_U52
g27313 nor P2_U2771 P2_U2770 ; P2_R2267_U53
g27314 nor P2_U2769 P2_U2768 ; P2_R2267_U54
g27315 not P2_U2789 ; P2_R2267_U55
g27316 and P2_R2267_U136 P2_R2267_U135 ; P2_R2267_U56
g27317 not P2_U3640 ; P2_R2267_U57
g27318 and P2_R2267_U138 P2_R2267_U137 ; P2_R2267_U58
g27319 not P2_U3642 ; P2_R2267_U59
g27320 and P2_R2267_U140 P2_R2267_U139 ; P2_R2267_U60
g27321 not P2_U2766 ; P2_R2267_U61
g27322 nand P2_R2267_U111 P2_R2267_U41 ; P2_R2267_U62
g27323 and P2_R2267_U142 P2_R2267_U141 ; P2_R2267_U63
g27324 not P2_U3644 ; P2_R2267_U64
g27325 and P2_R2267_U144 P2_R2267_U143 ; P2_R2267_U65
g27326 not P2_U2769 ; P2_R2267_U66
g27327 and P2_R2267_U146 P2_R2267_U145 ; P2_R2267_U67
g27328 not P2_U2771 ; P2_R2267_U68
g27329 and P2_R2267_U148 P2_R2267_U147 ; P2_R2267_U69
g27330 not P2_U2773 ; P2_R2267_U70
g27331 and P2_R2267_U150 P2_R2267_U149 ; P2_R2267_U71
g27332 not P2_U2775 ; P2_R2267_U72
g27333 and P2_R2267_U152 P2_R2267_U151 ; P2_R2267_U73
g27334 not P2_U2777 ; P2_R2267_U74
g27335 and P2_R2267_U154 P2_R2267_U153 ; P2_R2267_U75
g27336 not P2_U3645 ; P2_R2267_U76
g27337 nand P2_U3646 P2_R2267_U42 ; P2_R2267_U77
g27338 not P2_U2779 ; P2_R2267_U78
g27339 and P2_R2267_U158 P2_R2267_U157 ; P2_R2267_U79
g27340 not P2_U2781 ; P2_R2267_U80
g27341 and P2_R2267_U160 P2_R2267_U159 ; P2_R2267_U81
g27342 not P2_U2783 ; P2_R2267_U82
g27343 and P2_R2267_U162 P2_R2267_U161 ; P2_R2267_U83
g27344 not P2_U2785 ; P2_R2267_U84
g27345 and P2_R2267_U164 P2_R2267_U163 ; P2_R2267_U85
g27346 not P2_U2787 ; P2_R2267_U86
g27347 and P2_R2267_U166 P2_R2267_U165 ; P2_R2267_U87
g27348 not P2_R2267_U77 ; P2_R2267_U88
g27349 not P2_R2267_U23 ; P2_R2267_U89
g27350 not P2_R2267_U24 ; P2_R2267_U90
g27351 not P2_R2267_U25 ; P2_R2267_U91
g27352 not P2_R2267_U26 ; P2_R2267_U92
g27353 not P2_R2267_U30 ; P2_R2267_U93
g27354 nand P2_R2267_U92 P2_R2267_U55 ; P2_R2267_U94
g27355 nand P2_U2788 P2_R2267_U94 ; P2_R2267_U95
g27356 nand P2_R2267_U91 P2_R2267_U57 ; P2_R2267_U96
g27357 nand P2_U3639 P2_R2267_U96 ; P2_R2267_U97
g27358 nand P2_R2267_U90 P2_R2267_U59 ; P2_R2267_U98
g27359 nand P2_U3641 P2_R2267_U98 ; P2_R2267_U99
g27360 nand P2_R2267_U89 P2_R2267_U64 ; P2_R2267_U100
g27361 nand P2_U3643 P2_R2267_U100 ; P2_R2267_U101
g27362 not P2_R2267_U31 ; P2_R2267_U102
g27363 not P2_R2267_U32 ; P2_R2267_U103
g27364 not P2_R2267_U33 ; P2_R2267_U104
g27365 not P2_R2267_U34 ; P2_R2267_U105
g27366 not P2_R2267_U35 ; P2_R2267_U106
g27367 not P2_R2267_U36 ; P2_R2267_U107
g27368 not P2_R2267_U37 ; P2_R2267_U108
g27369 not P2_R2267_U38 ; P2_R2267_U109
g27370 not P2_R2267_U39 ; P2_R2267_U110
g27371 not P2_R2267_U40 ; P2_R2267_U111
g27372 not P2_R2267_U62 ; P2_R2267_U112
g27373 nand P2_U2767 P2_R2267_U40 ; P2_R2267_U113
g27374 nand P2_R2267_U110 P2_R2267_U66 ; P2_R2267_U114
g27375 nand P2_U2768 P2_R2267_U114 ; P2_R2267_U115
g27376 nand P2_R2267_U109 P2_R2267_U68 ; P2_R2267_U116
g27377 nand P2_U2770 P2_R2267_U116 ; P2_R2267_U117
g27378 nand P2_R2267_U108 P2_R2267_U70 ; P2_R2267_U118
g27379 nand P2_U2772 P2_R2267_U118 ; P2_R2267_U119
g27380 nand P2_R2267_U107 P2_R2267_U72 ; P2_R2267_U120
g27381 nand P2_U2774 P2_R2267_U120 ; P2_R2267_U121
g27382 nand P2_R2267_U106 P2_R2267_U74 ; P2_R2267_U122
g27383 nand P2_U2776 P2_R2267_U122 ; P2_R2267_U123
g27384 nand P2_R2267_U105 P2_R2267_U78 ; P2_R2267_U124
g27385 nand P2_U2778 P2_R2267_U124 ; P2_R2267_U125
g27386 nand P2_R2267_U104 P2_R2267_U80 ; P2_R2267_U126
g27387 nand P2_U2780 P2_R2267_U126 ; P2_R2267_U127
g27388 nand P2_R2267_U103 P2_R2267_U82 ; P2_R2267_U128
g27389 nand P2_U2782 P2_R2267_U128 ; P2_R2267_U129
g27390 nand P2_R2267_U102 P2_R2267_U84 ; P2_R2267_U130
g27391 nand P2_U2784 P2_R2267_U130 ; P2_R2267_U131
g27392 nand P2_R2267_U93 P2_R2267_U86 ; P2_R2267_U132
g27393 nand P2_U2786 P2_R2267_U132 ; P2_R2267_U133
g27394 nand P2_U2617 P2_R2267_U22 ; P2_R2267_U134
g27395 nand P2_U2789 P2_R2267_U26 ; P2_R2267_U135
g27396 nand P2_R2267_U92 P2_R2267_U55 ; P2_R2267_U136
g27397 nand P2_U3640 P2_R2267_U25 ; P2_R2267_U137
g27398 nand P2_R2267_U91 P2_R2267_U57 ; P2_R2267_U138
g27399 nand P2_U3642 P2_R2267_U24 ; P2_R2267_U139
g27400 nand P2_R2267_U90 P2_R2267_U59 ; P2_R2267_U140
g27401 nand P2_U2766 P2_R2267_U62 ; P2_R2267_U141
g27402 nand P2_R2267_U112 P2_R2267_U61 ; P2_R2267_U142
g27403 nand P2_U3644 P2_R2267_U23 ; P2_R2267_U143
g27404 nand P2_R2267_U89 P2_R2267_U64 ; P2_R2267_U144
g27405 nand P2_U2769 P2_R2267_U39 ; P2_R2267_U145
g27406 nand P2_R2267_U110 P2_R2267_U66 ; P2_R2267_U146
g27407 nand P2_U2771 P2_R2267_U38 ; P2_R2267_U147
g27408 nand P2_R2267_U109 P2_R2267_U68 ; P2_R2267_U148
g27409 nand P2_U2773 P2_R2267_U37 ; P2_R2267_U149
g27410 nand P2_R2267_U108 P2_R2267_U70 ; P2_R2267_U150
g27411 nand P2_U2775 P2_R2267_U36 ; P2_R2267_U151
g27412 nand P2_R2267_U107 P2_R2267_U72 ; P2_R2267_U152
g27413 nand P2_U2777 P2_R2267_U35 ; P2_R2267_U153
g27414 nand P2_R2267_U106 P2_R2267_U74 ; P2_R2267_U154
g27415 nand P2_U3645 P2_R2267_U77 ; P2_R2267_U155
g27416 nand P2_R2267_U88 P2_R2267_U76 ; P2_R2267_U156
g27417 nand P2_U2779 P2_R2267_U34 ; P2_R2267_U157
g27418 nand P2_R2267_U105 P2_R2267_U78 ; P2_R2267_U158
g27419 nand P2_U2781 P2_R2267_U33 ; P2_R2267_U159
g27420 nand P2_R2267_U104 P2_R2267_U80 ; P2_R2267_U160
g27421 nand P2_U2783 P2_R2267_U32 ; P2_R2267_U161
g27422 nand P2_R2267_U103 P2_R2267_U82 ; P2_R2267_U162
g27423 nand P2_U2785 P2_R2267_U31 ; P2_R2267_U163
g27424 nand P2_R2267_U102 P2_R2267_U84 ; P2_R2267_U164
g27425 nand P2_U2787 P2_R2267_U30 ; P2_R2267_U165
g27426 nand P2_R2267_U93 P2_R2267_U86 ; P2_R2267_U166
g27427 and P2_ADD_371_1212_U10 P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_ADD_371_1212_U4
g27428 and P2_INSTADDRPOINTER_REG_9__SCAN_IN P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_ADD_371_1212_U5
g27429 and P2_ADD_371_1212_U89 P2_ADD_371_1212_U11 ; P2_ADD_371_1212_U6
g27430 and P2_ADD_371_1212_U10 P2_ADD_371_1212_U87 ; P2_ADD_371_1212_U7
g27431 and P2_ADD_371_1212_U9 P2_ADD_371_1212_U91 ; P2_ADD_371_1212_U8
g27432 and P2_ADD_371_1212_U6 P2_ADD_371_1212_U90 ; P2_ADD_371_1212_U9
g27433 and P2_INSTADDRPOINTER_REG_9__SCAN_IN P2_INSTADDRPOINTER_REG_10__SCAN_IN P2_INSTADDRPOINTER_REG_11__SCAN_IN P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_ADD_371_1212_U10
g27434 and P2_ADD_371_1212_U7 P2_ADD_371_1212_U88 ; P2_ADD_371_1212_U11
g27435 and P2_ADD_371_1212_U8 P2_ADD_371_1212_U92 ; P2_ADD_371_1212_U12
g27436 and P2_ADD_371_1212_U196 P2_ADD_371_1212_U168 ; P2_ADD_371_1212_U13
g27437 and P2_ADD_371_1212_U188 P2_ADD_371_1212_U132 ; P2_ADD_371_1212_U14
g27438 and P2_ADD_371_1212_U185 P2_ADD_371_1212_U170 ; P2_ADD_371_1212_U15
g27439 and P2_ADD_371_1212_U191 P2_ADD_371_1212_U120 ; P2_ADD_371_1212_U16
g27440 and P2_ADD_371_1212_U200 P2_ADD_371_1212_U114 ; P2_ADD_371_1212_U17
g27441 and P2_ADD_371_1212_U194 P2_ADD_371_1212_U174 ; P2_ADD_371_1212_U18
g27442 and P2_ADD_371_1212_U183 P2_ADD_371_1212_U131 ; P2_ADD_371_1212_U19
g27443 and P2_ADD_371_1212_U187 P2_ADD_371_1212_U176 ; P2_ADD_371_1212_U20
g27444 and P2_ADD_371_1212_U192 P2_ADD_371_1212_U113 ; P2_ADD_371_1212_U21
g27445 and P2_ADD_371_1212_U190 P2_ADD_371_1212_U123 ; P2_ADD_371_1212_U22
g27446 and P2_ADD_371_1212_U198 P2_ADD_371_1212_U180 ; P2_ADD_371_1212_U23
g27447 and P2_ADD_371_1212_U182 P2_ADD_371_1212_U112 ; P2_ADD_371_1212_U24
g27448 nand P2_ADD_371_1212_U269 P2_ADD_371_1212_U268 P2_ADD_371_1212_U204 ; P2_ADD_371_1212_U25
g27449 not P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_ADD_371_1212_U26
g27450 not P2_R2256_U21 ; P2_ADD_371_1212_U27
g27451 not P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_371_1212_U28
g27452 nand P2_R2256_U21 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_ADD_371_1212_U29
g27453 not P2_R2256_U4 ; P2_ADD_371_1212_U30
g27454 not P2_R2256_U22 ; P2_ADD_371_1212_U31
g27455 not P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_371_1212_U32
g27456 not P2_R2256_U26 ; P2_ADD_371_1212_U33
g27457 not P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_371_1212_U34
g27458 not P2_R2256_U20 ; P2_ADD_371_1212_U35
g27459 not P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_371_1212_U36
g27460 not P2_R2256_U19 ; P2_ADD_371_1212_U37
g27461 not P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_371_1212_U38
g27462 not P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_371_1212_U39
g27463 not P2_R2256_U18 ; P2_ADD_371_1212_U40
g27464 not P2_R2256_U5 ; P2_ADD_371_1212_U41
g27465 not P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_371_1212_U42
g27466 not P2_R2256_U17 ; P2_ADD_371_1212_U43
g27467 not P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_371_1212_U44
g27468 not P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_ADD_371_1212_U45
g27469 not P2_INSTADDRPOINTER_REG_10__SCAN_IN ; P2_ADD_371_1212_U46
g27470 not P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_ADD_371_1212_U47
g27471 not P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_ADD_371_1212_U48
g27472 not P2_INSTADDRPOINTER_REG_13__SCAN_IN ; P2_ADD_371_1212_U49
g27473 not P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_ADD_371_1212_U50
g27474 not P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_ADD_371_1212_U51
g27475 not P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_ADD_371_1212_U52
g27476 not P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_ADD_371_1212_U53
g27477 not P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_ADD_371_1212_U54
g27478 not P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_ADD_371_1212_U55
g27479 not P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_ADD_371_1212_U56
g27480 not P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_ADD_371_1212_U57
g27481 not P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_ADD_371_1212_U58
g27482 not P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_ADD_371_1212_U59
g27483 not P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_ADD_371_1212_U60
g27484 not P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_ADD_371_1212_U61
g27485 not P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_ADD_371_1212_U62
g27486 not P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_ADD_371_1212_U63
g27487 not P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_ADD_371_1212_U64
g27488 not P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_ADD_371_1212_U65
g27489 not P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_371_1212_U66
g27490 nand P2_R2256_U4 P2_ADD_371_1212_U137 ; P2_ADD_371_1212_U67
g27491 nand P2_ADD_371_1212_U206 P2_ADD_371_1212_U205 ; P2_ADD_371_1212_U68
g27492 nand P2_ADD_371_1212_U215 P2_ADD_371_1212_U214 ; P2_ADD_371_1212_U69
g27493 nand P2_ADD_371_1212_U217 P2_ADD_371_1212_U216 ; P2_ADD_371_1212_U70
g27494 nand P2_ADD_371_1212_U219 P2_ADD_371_1212_U218 ; P2_ADD_371_1212_U71
g27495 nand P2_ADD_371_1212_U230 P2_ADD_371_1212_U229 ; P2_ADD_371_1212_U72
g27496 nand P2_ADD_371_1212_U232 P2_ADD_371_1212_U231 ; P2_ADD_371_1212_U73
g27497 nand P2_ADD_371_1212_U241 P2_ADD_371_1212_U240 ; P2_ADD_371_1212_U74
g27498 nand P2_ADD_371_1212_U271 P2_ADD_371_1212_U270 ; P2_ADD_371_1212_U75
g27499 nand P2_ADD_371_1212_U273 P2_ADD_371_1212_U272 ; P2_ADD_371_1212_U76
g27500 nand P2_ADD_371_1212_U282 P2_ADD_371_1212_U281 ; P2_ADD_371_1212_U77
g27501 nand P2_ADD_371_1212_U213 P2_ADD_371_1212_U212 ; P2_ADD_371_1212_U78
g27502 nand P2_ADD_371_1212_U226 P2_ADD_371_1212_U225 ; P2_ADD_371_1212_U79
g27503 nand P2_ADD_371_1212_U239 P2_ADD_371_1212_U238 ; P2_ADD_371_1212_U80
g27504 nand P2_ADD_371_1212_U248 P2_ADD_371_1212_U247 ; P2_ADD_371_1212_U81
g27505 nand P2_ADD_371_1212_U255 P2_ADD_371_1212_U254 ; P2_ADD_371_1212_U82
g27506 nand P2_ADD_371_1212_U257 P2_ADD_371_1212_U256 ; P2_ADD_371_1212_U83
g27507 nand P2_ADD_371_1212_U264 P2_ADD_371_1212_U263 ; P2_ADD_371_1212_U84
g27508 nand P2_ADD_371_1212_U280 P2_ADD_371_1212_U279 ; P2_ADD_371_1212_U85
g27509 and P2_ADD_371_1212_U203 P2_ADD_371_1212_U166 ; P2_ADD_371_1212_U86
g27510 and P2_INSTADDRPOINTER_REG_13__SCAN_IN P2_INSTADDRPOINTER_REG_14__SCAN_IN P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_ADD_371_1212_U87
g27511 and P2_INSTADDRPOINTER_REG_16__SCAN_IN P2_INSTADDRPOINTER_REG_17__SCAN_IN P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_ADD_371_1212_U88
g27512 and P2_INSTADDRPOINTER_REG_19__SCAN_IN P2_INSTADDRPOINTER_REG_20__SCAN_IN ; P2_ADD_371_1212_U89
g27513 and P2_INSTADDRPOINTER_REG_21__SCAN_IN P2_INSTADDRPOINTER_REG_22__SCAN_IN P2_INSTADDRPOINTER_REG_23__SCAN_IN ; P2_ADD_371_1212_U90
g27514 and P2_INSTADDRPOINTER_REG_24__SCAN_IN P2_INSTADDRPOINTER_REG_25__SCAN_IN P2_INSTADDRPOINTER_REG_26__SCAN_IN ; P2_ADD_371_1212_U91
g27515 and P2_INSTADDRPOINTER_REG_27__SCAN_IN P2_INSTADDRPOINTER_REG_28__SCAN_IN P2_INSTADDRPOINTER_REG_29__SCAN_IN ; P2_ADD_371_1212_U92
g27516 and P2_ADD_371_1212_U8 P2_ADD_371_1212_U94 ; P2_ADD_371_1212_U93
g27517 and P2_INSTADDRPOINTER_REG_27__SCAN_IN P2_INSTADDRPOINTER_REG_28__SCAN_IN ; P2_ADD_371_1212_U94
g27518 and P2_ADD_371_1212_U7 P2_INSTADDRPOINTER_REG_16__SCAN_IN ; P2_ADD_371_1212_U95
g27519 and P2_ADD_371_1212_U11 P2_INSTADDRPOINTER_REG_19__SCAN_IN ; P2_ADD_371_1212_U96
g27520 and P2_ADD_371_1212_U6 P2_ADD_371_1212_U98 ; P2_ADD_371_1212_U97
g27521 and P2_INSTADDRPOINTER_REG_21__SCAN_IN P2_INSTADDRPOINTER_REG_22__SCAN_IN ; P2_ADD_371_1212_U98
g27522 and P2_ADD_371_1212_U6 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_ADD_371_1212_U99
g27523 and P2_ADD_371_1212_U7 P2_ADD_371_1212_U101 ; P2_ADD_371_1212_U100
g27524 and P2_INSTADDRPOINTER_REG_16__SCAN_IN P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_ADD_371_1212_U101
g27525 and P2_ADD_371_1212_U5 P2_INSTADDRPOINTER_REG_11__SCAN_IN ; P2_ADD_371_1212_U102
g27526 and P2_ADD_371_1212_U9 P2_ADD_371_1212_U104 ; P2_ADD_371_1212_U103
g27527 and P2_INSTADDRPOINTER_REG_24__SCAN_IN P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_ADD_371_1212_U104
g27528 and P2_ADD_371_1212_U4 P2_INSTADDRPOINTER_REG_14__SCAN_IN ; P2_ADD_371_1212_U105
g27529 and P2_ADD_371_1212_U12 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_371_1212_U106
g27530 and P2_ADD_371_1212_U12 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_371_1212_U107
g27531 and P2_ADD_371_1212_U8 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_ADD_371_1212_U108
g27532 and P2_ADD_371_1212_U9 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_ADD_371_1212_U109
g27533 and P2_ADD_371_1212_U208 P2_ADD_371_1212_U207 ; P2_ADD_371_1212_U110
g27534 nand P2_ADD_371_1212_U155 P2_ADD_371_1212_U154 ; P2_ADD_371_1212_U111
g27535 nand P2_ADD_371_1212_U12 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U112
g27536 nand P2_ADD_371_1212_U9 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U113
g27537 nand P2_ADD_371_1212_U95 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U114
g27538 and P2_ADD_371_1212_U221 P2_ADD_371_1212_U220 ; P2_ADD_371_1212_U115
g27539 nand P2_ADD_371_1212_U67 P2_ADD_371_1212_U139 ; P2_ADD_371_1212_U116
g27540 nand P2_ADD_371_1212_U86 P2_ADD_371_1212_U202 ; P2_ADD_371_1212_U117
g27541 and P2_ADD_371_1212_U228 P2_ADD_371_1212_U227 ; P2_ADD_371_1212_U118
g27542 nand P2_ADD_371_1212_U117 P2_ADD_371_1212_U100 ; P2_ADD_371_1212_U119
g27543 nand P2_ADD_371_1212_U105 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U120
g27544 and P2_ADD_371_1212_U234 P2_ADD_371_1212_U233 ; P2_ADD_371_1212_U121
g27545 nand P2_ADD_371_1212_U147 P2_ADD_371_1212_U146 ; P2_ADD_371_1212_U122
g27546 nand P2_ADD_371_1212_U8 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U123
g27547 and P2_ADD_371_1212_U243 P2_ADD_371_1212_U242 ; P2_ADD_371_1212_U124
g27548 nand P2_ADD_371_1212_U151 P2_ADD_371_1212_U150 ; P2_ADD_371_1212_U125
g27549 and P2_ADD_371_1212_U250 P2_ADD_371_1212_U249 ; P2_ADD_371_1212_U126
g27550 nand P2_ADD_371_1212_U163 P2_ADD_371_1212_U162 ; P2_ADD_371_1212_U127
g27551 not P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_ADD_371_1212_U128
g27552 and P2_ADD_371_1212_U259 P2_ADD_371_1212_U258 ; P2_ADD_371_1212_U129
g27553 nand P2_ADD_371_1212_U143 P2_ADD_371_1212_U142 ; P2_ADD_371_1212_U130
g27554 nand P2_ADD_371_1212_U6 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U131
g27555 nand P2_ADD_371_1212_U102 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U132
g27556 and P2_ADD_371_1212_U275 P2_ADD_371_1212_U274 ; P2_ADD_371_1212_U133
g27557 nand P2_ADD_371_1212_U159 P2_ADD_371_1212_U158 ; P2_ADD_371_1212_U134
g27558 nand P2_ADD_371_1212_U109 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U135
g27559 not P2_ADD_371_1212_U67 ; P2_ADD_371_1212_U136
g27560 not P2_ADD_371_1212_U29 ; P2_ADD_371_1212_U137
g27561 nand P2_ADD_371_1212_U30 P2_ADD_371_1212_U29 ; P2_ADD_371_1212_U138
g27562 nand P2_ADD_371_1212_U138 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_371_1212_U139
g27563 not P2_ADD_371_1212_U116 ; P2_ADD_371_1212_U140
g27564 or P2_R2256_U22 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_371_1212_U141
g27565 nand P2_ADD_371_1212_U141 P2_ADD_371_1212_U116 ; P2_ADD_371_1212_U142
g27566 nand P2_R2256_U22 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_371_1212_U143
g27567 not P2_ADD_371_1212_U130 ; P2_ADD_371_1212_U144
g27568 or P2_R2256_U26 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_371_1212_U145
g27569 nand P2_ADD_371_1212_U145 P2_ADD_371_1212_U130 ; P2_ADD_371_1212_U146
g27570 nand P2_R2256_U26 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_371_1212_U147
g27571 not P2_ADD_371_1212_U122 ; P2_ADD_371_1212_U148
g27572 or P2_R2256_U20 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_371_1212_U149
g27573 nand P2_ADD_371_1212_U149 P2_ADD_371_1212_U122 ; P2_ADD_371_1212_U150
g27574 nand P2_R2256_U20 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_371_1212_U151
g27575 not P2_ADD_371_1212_U125 ; P2_ADD_371_1212_U152
g27576 or P2_R2256_U19 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_371_1212_U153
g27577 nand P2_ADD_371_1212_U153 P2_ADD_371_1212_U125 ; P2_ADD_371_1212_U154
g27578 nand P2_R2256_U19 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_371_1212_U155
g27579 not P2_ADD_371_1212_U111 ; P2_ADD_371_1212_U156
g27580 or P2_R2256_U18 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_371_1212_U157
g27581 nand P2_ADD_371_1212_U157 P2_ADD_371_1212_U111 ; P2_ADD_371_1212_U158
g27582 nand P2_R2256_U18 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_371_1212_U159
g27583 not P2_ADD_371_1212_U134 ; P2_ADD_371_1212_U160
g27584 or P2_R2256_U17 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_371_1212_U161
g27585 nand P2_ADD_371_1212_U161 P2_ADD_371_1212_U134 ; P2_ADD_371_1212_U162
g27586 nand P2_R2256_U17 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_371_1212_U163
g27587 not P2_ADD_371_1212_U127 ; P2_ADD_371_1212_U164
g27588 or P2_R2256_U5 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_371_1212_U165
g27589 nand P2_R2256_U5 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_371_1212_U166
g27590 not P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U167
g27591 nand P2_ADD_371_1212_U5 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U168
g27592 not P2_ADD_371_1212_U132 ; P2_ADD_371_1212_U169
g27593 nand P2_ADD_371_1212_U4 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U170
g27594 not P2_ADD_371_1212_U120 ; P2_ADD_371_1212_U171
g27595 not P2_ADD_371_1212_U114 ; P2_ADD_371_1212_U172
g27596 not P2_ADD_371_1212_U119 ; P2_ADD_371_1212_U173
g27597 nand P2_ADD_371_1212_U96 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U174
g27598 not P2_ADD_371_1212_U131 ; P2_ADD_371_1212_U175
g27599 nand P2_ADD_371_1212_U117 P2_ADD_371_1212_U97 ; P2_ADD_371_1212_U176
g27600 not P2_ADD_371_1212_U113 ; P2_ADD_371_1212_U177
g27601 not P2_ADD_371_1212_U135 ; P2_ADD_371_1212_U178
g27602 not P2_ADD_371_1212_U123 ; P2_ADD_371_1212_U179
g27603 nand P2_ADD_371_1212_U117 P2_ADD_371_1212_U93 ; P2_ADD_371_1212_U180
g27604 not P2_ADD_371_1212_U112 ; P2_ADD_371_1212_U181
g27605 nand P2_ADD_371_1212_U65 P2_ADD_371_1212_U180 ; P2_ADD_371_1212_U182
g27606 nand P2_ADD_371_1212_U56 P2_ADD_371_1212_U174 ; P2_ADD_371_1212_U183
g27607 nand P2_ADD_371_1212_U10 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U184
g27608 nand P2_ADD_371_1212_U49 P2_ADD_371_1212_U184 ; P2_ADD_371_1212_U185
g27609 nand P2_ADD_371_1212_U99 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U186
g27610 nand P2_ADD_371_1212_U58 P2_ADD_371_1212_U186 ; P2_ADD_371_1212_U187
g27611 nand P2_ADD_371_1212_U47 P2_ADD_371_1212_U168 ; P2_ADD_371_1212_U188
g27612 nand P2_ADD_371_1212_U117 P2_ADD_371_1212_U103 ; P2_ADD_371_1212_U189
g27613 nand P2_ADD_371_1212_U61 P2_ADD_371_1212_U189 ; P2_ADD_371_1212_U190
g27614 nand P2_ADD_371_1212_U50 P2_ADD_371_1212_U170 ; P2_ADD_371_1212_U191
g27615 nand P2_ADD_371_1212_U59 P2_ADD_371_1212_U176 ; P2_ADD_371_1212_U192
g27616 nand P2_ADD_371_1212_U11 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U193
g27617 nand P2_ADD_371_1212_U55 P2_ADD_371_1212_U193 ; P2_ADD_371_1212_U194
g27618 nand P2_ADD_371_1212_U117 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_ADD_371_1212_U195
g27619 nand P2_ADD_371_1212_U46 P2_ADD_371_1212_U195 ; P2_ADD_371_1212_U196
g27620 nand P2_ADD_371_1212_U108 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U197
g27621 nand P2_ADD_371_1212_U64 P2_ADD_371_1212_U197 ; P2_ADD_371_1212_U198
g27622 nand P2_ADD_371_1212_U7 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U199
g27623 nand P2_ADD_371_1212_U52 P2_ADD_371_1212_U199 ; P2_ADD_371_1212_U200
g27624 nand P2_ADD_371_1212_U107 P2_ADD_371_1212_U117 ; P2_ADD_371_1212_U201
g27625 nand P2_ADD_371_1212_U165 P2_ADD_371_1212_U134 P2_ADD_371_1212_U161 ; P2_ADD_371_1212_U202
g27626 nand P2_ADD_371_1212_U165 P2_R2256_U17 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_371_1212_U203
g27627 nand P2_ADD_371_1212_U136 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_371_1212_U204
g27628 nand P2_ADD_371_1212_U27 P2_INSTADDRPOINTER_REG_0__SCAN_IN ; P2_ADD_371_1212_U205
g27629 nand P2_R2256_U21 P2_ADD_371_1212_U26 ; P2_ADD_371_1212_U206
g27630 nand P2_ADD_371_1212_U40 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_371_1212_U207
g27631 nand P2_R2256_U18 P2_ADD_371_1212_U39 ; P2_ADD_371_1212_U208
g27632 nand P2_ADD_371_1212_U40 P2_INSTADDRPOINTER_REG_6__SCAN_IN ; P2_ADD_371_1212_U209
g27633 nand P2_R2256_U18 P2_ADD_371_1212_U39 ; P2_ADD_371_1212_U210
g27634 nand P2_ADD_371_1212_U210 P2_ADD_371_1212_U209 ; P2_ADD_371_1212_U211
g27635 nand P2_ADD_371_1212_U110 P2_ADD_371_1212_U111 ; P2_ADD_371_1212_U212
g27636 nand P2_ADD_371_1212_U156 P2_ADD_371_1212_U211 ; P2_ADD_371_1212_U213
g27637 nand P2_ADD_371_1212_U112 P2_INSTADDRPOINTER_REG_30__SCAN_IN ; P2_ADD_371_1212_U214
g27638 nand P2_ADD_371_1212_U181 P2_ADD_371_1212_U66 ; P2_ADD_371_1212_U215
g27639 nand P2_ADD_371_1212_U113 P2_INSTADDRPOINTER_REG_24__SCAN_IN ; P2_ADD_371_1212_U216
g27640 nand P2_ADD_371_1212_U177 P2_ADD_371_1212_U60 ; P2_ADD_371_1212_U217
g27641 nand P2_ADD_371_1212_U114 P2_INSTADDRPOINTER_REG_17__SCAN_IN ; P2_ADD_371_1212_U218
g27642 nand P2_ADD_371_1212_U172 P2_ADD_371_1212_U54 ; P2_ADD_371_1212_U219
g27643 nand P2_ADD_371_1212_U31 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_371_1212_U220
g27644 nand P2_R2256_U22 P2_ADD_371_1212_U32 ; P2_ADD_371_1212_U221
g27645 nand P2_ADD_371_1212_U31 P2_INSTADDRPOINTER_REG_2__SCAN_IN ; P2_ADD_371_1212_U222
g27646 nand P2_R2256_U22 P2_ADD_371_1212_U32 ; P2_ADD_371_1212_U223
g27647 nand P2_ADD_371_1212_U223 P2_ADD_371_1212_U222 ; P2_ADD_371_1212_U224
g27648 nand P2_ADD_371_1212_U115 P2_ADD_371_1212_U116 ; P2_ADD_371_1212_U225
g27649 nand P2_ADD_371_1212_U140 P2_ADD_371_1212_U224 ; P2_ADD_371_1212_U226
g27650 nand P2_ADD_371_1212_U117 P2_INSTADDRPOINTER_REG_9__SCAN_IN ; P2_ADD_371_1212_U227
g27651 nand P2_ADD_371_1212_U167 P2_ADD_371_1212_U45 ; P2_ADD_371_1212_U228
g27652 nand P2_ADD_371_1212_U119 P2_INSTADDRPOINTER_REG_18__SCAN_IN ; P2_ADD_371_1212_U229
g27653 nand P2_ADD_371_1212_U173 P2_ADD_371_1212_U53 ; P2_ADD_371_1212_U230
g27654 nand P2_ADD_371_1212_U120 P2_INSTADDRPOINTER_REG_15__SCAN_IN ; P2_ADD_371_1212_U231
g27655 nand P2_ADD_371_1212_U171 P2_ADD_371_1212_U51 ; P2_ADD_371_1212_U232
g27656 nand P2_ADD_371_1212_U35 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_371_1212_U233
g27657 nand P2_R2256_U20 P2_ADD_371_1212_U36 ; P2_ADD_371_1212_U234
g27658 nand P2_ADD_371_1212_U35 P2_INSTADDRPOINTER_REG_4__SCAN_IN ; P2_ADD_371_1212_U235
g27659 nand P2_R2256_U20 P2_ADD_371_1212_U36 ; P2_ADD_371_1212_U236
g27660 nand P2_ADD_371_1212_U236 P2_ADD_371_1212_U235 ; P2_ADD_371_1212_U237
g27661 nand P2_ADD_371_1212_U121 P2_ADD_371_1212_U122 ; P2_ADD_371_1212_U238
g27662 nand P2_ADD_371_1212_U148 P2_ADD_371_1212_U237 ; P2_ADD_371_1212_U239
g27663 nand P2_ADD_371_1212_U123 P2_INSTADDRPOINTER_REG_27__SCAN_IN ; P2_ADD_371_1212_U240
g27664 nand P2_ADD_371_1212_U179 P2_ADD_371_1212_U63 ; P2_ADD_371_1212_U241
g27665 nand P2_ADD_371_1212_U37 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_371_1212_U242
g27666 nand P2_R2256_U19 P2_ADD_371_1212_U38 ; P2_ADD_371_1212_U243
g27667 nand P2_ADD_371_1212_U37 P2_INSTADDRPOINTER_REG_5__SCAN_IN ; P2_ADD_371_1212_U244
g27668 nand P2_R2256_U19 P2_ADD_371_1212_U38 ; P2_ADD_371_1212_U245
g27669 nand P2_ADD_371_1212_U245 P2_ADD_371_1212_U244 ; P2_ADD_371_1212_U246
g27670 nand P2_ADD_371_1212_U124 P2_ADD_371_1212_U125 ; P2_ADD_371_1212_U247
g27671 nand P2_ADD_371_1212_U152 P2_ADD_371_1212_U246 ; P2_ADD_371_1212_U248
g27672 nand P2_ADD_371_1212_U41 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_371_1212_U249
g27673 nand P2_R2256_U5 P2_ADD_371_1212_U42 ; P2_ADD_371_1212_U250
g27674 nand P2_ADD_371_1212_U41 P2_INSTADDRPOINTER_REG_8__SCAN_IN ; P2_ADD_371_1212_U251
g27675 nand P2_R2256_U5 P2_ADD_371_1212_U42 ; P2_ADD_371_1212_U252
g27676 nand P2_ADD_371_1212_U252 P2_ADD_371_1212_U251 ; P2_ADD_371_1212_U253
g27677 nand P2_ADD_371_1212_U126 P2_ADD_371_1212_U127 ; P2_ADD_371_1212_U254
g27678 nand P2_ADD_371_1212_U164 P2_ADD_371_1212_U253 ; P2_ADD_371_1212_U255
g27679 nand P2_ADD_371_1212_U201 P2_INSTADDRPOINTER_REG_31__SCAN_IN ; P2_ADD_371_1212_U256
g27680 nand P2_ADD_371_1212_U106 P2_ADD_371_1212_U117 P2_ADD_371_1212_U128 ; P2_ADD_371_1212_U257
g27681 nand P2_ADD_371_1212_U33 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_371_1212_U258
g27682 nand P2_R2256_U26 P2_ADD_371_1212_U34 ; P2_ADD_371_1212_U259
g27683 nand P2_ADD_371_1212_U33 P2_INSTADDRPOINTER_REG_3__SCAN_IN ; P2_ADD_371_1212_U260
g27684 nand P2_R2256_U26 P2_ADD_371_1212_U34 ; P2_ADD_371_1212_U261
g27685 nand P2_ADD_371_1212_U261 P2_ADD_371_1212_U260 ; P2_ADD_371_1212_U262
g27686 nand P2_ADD_371_1212_U129 P2_ADD_371_1212_U130 ; P2_ADD_371_1212_U263
g27687 nand P2_ADD_371_1212_U144 P2_ADD_371_1212_U262 ; P2_ADD_371_1212_U264
g27688 nand P2_ADD_371_1212_U29 P2_INSTADDRPOINTER_REG_1__SCAN_IN ; P2_ADD_371_1212_U265
g27689 nand P2_ADD_371_1212_U137 P2_ADD_371_1212_U28 ; P2_ADD_371_1212_U266
g27690 nand P2_ADD_371_1212_U266 P2_ADD_371_1212_U265 ; P2_ADD_371_1212_U267
g27691 nand P2_ADD_371_1212_U29 P2_ADD_371_1212_U28 P2_R2256_U4 ; P2_ADD_371_1212_U268
g27692 nand P2_ADD_371_1212_U267 P2_ADD_371_1212_U30 ; P2_ADD_371_1212_U269
g27693 nand P2_ADD_371_1212_U131 P2_INSTADDRPOINTER_REG_21__SCAN_IN ; P2_ADD_371_1212_U270
g27694 nand P2_ADD_371_1212_U175 P2_ADD_371_1212_U57 ; P2_ADD_371_1212_U271
g27695 nand P2_ADD_371_1212_U132 P2_INSTADDRPOINTER_REG_12__SCAN_IN ; P2_ADD_371_1212_U272
g27696 nand P2_ADD_371_1212_U169 P2_ADD_371_1212_U48 ; P2_ADD_371_1212_U273
g27697 nand P2_ADD_371_1212_U43 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_371_1212_U274
g27698 nand P2_R2256_U17 P2_ADD_371_1212_U44 ; P2_ADD_371_1212_U275
g27699 nand P2_ADD_371_1212_U43 P2_INSTADDRPOINTER_REG_7__SCAN_IN ; P2_ADD_371_1212_U276
g27700 nand P2_R2256_U17 P2_ADD_371_1212_U44 ; P2_ADD_371_1212_U277
g27701 nand P2_ADD_371_1212_U277 P2_ADD_371_1212_U276 ; P2_ADD_371_1212_U278
g27702 nand P2_ADD_371_1212_U133 P2_ADD_371_1212_U134 ; P2_ADD_371_1212_U279
g27703 nand P2_ADD_371_1212_U160 P2_ADD_371_1212_U278 ; P2_ADD_371_1212_U280
g27704 nand P2_ADD_371_1212_U135 P2_INSTADDRPOINTER_REG_25__SCAN_IN ; P2_ADD_371_1212_U281
g27705 nand P2_ADD_371_1212_U178 P2_ADD_371_1212_U62 ; P2_ADD_371_1212_U282
g27706 not P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_R2027_U5
g27707 not P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2027_U6
g27708 not P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2027_U7
g27709 not P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2027_U8
g27710 not P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2027_U9
g27711 nand P1_INSTADDRPOINTER_REG_0__SCAN_IN P1_INSTADDRPOINTER_REG_1__SCAN_IN P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2027_U10
g27712 not P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2027_U11
g27713 not P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2027_U12
g27714 nand P1_R2027_U82 P1_R2027_U111 ; P1_R2027_U13
g27715 not P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2027_U14
g27716 not P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2027_U15
g27717 nand P1_R2027_U83 P1_R2027_U112 ; P1_R2027_U16
g27718 nand P1_R2027_U84 P1_R2027_U118 ; P1_R2027_U17
g27719 not P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2027_U18
g27720 not P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2027_U19
g27721 not P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_R2027_U20
g27722 not P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2027_U21
g27723 nand P1_R2027_U85 P1_R2027_U120 ; P1_R2027_U22
g27724 not P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2027_U23
g27725 not P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2027_U24
g27726 nand P1_R2027_U86 P1_R2027_U113 ; P1_R2027_U25
g27727 not P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2027_U26
g27728 nand P1_R2027_U87 P1_R2027_U119 ; P1_R2027_U27
g27729 not P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2027_U28
g27730 not P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2027_U29
g27731 not P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2027_U30
g27732 nand P1_R2027_U88 P1_R2027_U124 ; P1_R2027_U31
g27733 not P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2027_U32
g27734 not P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2027_U33
g27735 nand P1_R2027_U89 P1_R2027_U117 ; P1_R2027_U34
g27736 not P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2027_U35
g27737 nand P1_R2027_U90 P1_R2027_U114 ; P1_R2027_U36
g27738 not P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2027_U37
g27739 not P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2027_U38
g27740 not P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2027_U39
g27741 nand P1_R2027_U91 P1_R2027_U121 ; P1_R2027_U40
g27742 not P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2027_U41
g27743 not P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2027_U42
g27744 nand P1_R2027_U92 P1_R2027_U115 ; P1_R2027_U43
g27745 not P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2027_U44
g27746 not P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2027_U45
g27747 nand P1_R2027_U93 P1_R2027_U116 ; P1_R2027_U46
g27748 not P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2027_U47
g27749 nand P1_R2027_U94 P1_R2027_U122 ; P1_R2027_U48
g27750 nand P1_R2027_U123 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2027_U49
g27751 not P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2027_U50
g27752 nand P1_R2027_U142 P1_R2027_U141 ; P1_R2027_U51
g27753 nand P1_R2027_U144 P1_R2027_U143 ; P1_R2027_U52
g27754 nand P1_R2027_U146 P1_R2027_U145 ; P1_R2027_U53
g27755 nand P1_R2027_U148 P1_R2027_U147 ; P1_R2027_U54
g27756 nand P1_R2027_U150 P1_R2027_U149 ; P1_R2027_U55
g27757 nand P1_R2027_U152 P1_R2027_U151 ; P1_R2027_U56
g27758 nand P1_R2027_U154 P1_R2027_U153 ; P1_R2027_U57
g27759 nand P1_R2027_U156 P1_R2027_U155 ; P1_R2027_U58
g27760 nand P1_R2027_U158 P1_R2027_U157 ; P1_R2027_U59
g27761 nand P1_R2027_U160 P1_R2027_U159 ; P1_R2027_U60
g27762 nand P1_R2027_U162 P1_R2027_U161 ; P1_R2027_U61
g27763 nand P1_R2027_U164 P1_R2027_U163 ; P1_R2027_U62
g27764 nand P1_R2027_U166 P1_R2027_U165 ; P1_R2027_U63
g27765 nand P1_R2027_U168 P1_R2027_U167 ; P1_R2027_U64
g27766 nand P1_R2027_U170 P1_R2027_U169 ; P1_R2027_U65
g27767 nand P1_R2027_U172 P1_R2027_U171 ; P1_R2027_U66
g27768 nand P1_R2027_U174 P1_R2027_U173 ; P1_R2027_U67
g27769 nand P1_R2027_U176 P1_R2027_U175 ; P1_R2027_U68
g27770 nand P1_R2027_U178 P1_R2027_U177 ; P1_R2027_U69
g27771 nand P1_R2027_U180 P1_R2027_U179 ; P1_R2027_U70
g27772 nand P1_R2027_U182 P1_R2027_U181 ; P1_R2027_U71
g27773 nand P1_R2027_U184 P1_R2027_U183 ; P1_R2027_U72
g27774 nand P1_R2027_U186 P1_R2027_U185 ; P1_R2027_U73
g27775 nand P1_R2027_U188 P1_R2027_U187 ; P1_R2027_U74
g27776 nand P1_R2027_U190 P1_R2027_U189 ; P1_R2027_U75
g27777 nand P1_R2027_U192 P1_R2027_U191 ; P1_R2027_U76
g27778 nand P1_R2027_U194 P1_R2027_U193 ; P1_R2027_U77
g27779 nand P1_R2027_U196 P1_R2027_U195 ; P1_R2027_U78
g27780 nand P1_R2027_U198 P1_R2027_U197 ; P1_R2027_U79
g27781 nand P1_R2027_U200 P1_R2027_U199 ; P1_R2027_U80
g27782 nand P1_R2027_U202 P1_R2027_U201 ; P1_R2027_U81
g27783 and P1_INSTADDRPOINTER_REG_3__SCAN_IN P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2027_U82
g27784 and P1_INSTADDRPOINTER_REG_5__SCAN_IN P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2027_U83
g27785 and P1_INSTADDRPOINTER_REG_7__SCAN_IN P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2027_U84
g27786 and P1_INSTADDRPOINTER_REG_9__SCAN_IN P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2027_U85
g27787 and P1_INSTADDRPOINTER_REG_11__SCAN_IN P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_R2027_U86
g27788 and P1_INSTADDRPOINTER_REG_13__SCAN_IN P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2027_U87
g27789 and P1_INSTADDRPOINTER_REG_15__SCAN_IN P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2027_U88
g27790 and P1_INSTADDRPOINTER_REG_17__SCAN_IN P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2027_U89
g27791 and P1_INSTADDRPOINTER_REG_19__SCAN_IN P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2027_U90
g27792 and P1_INSTADDRPOINTER_REG_21__SCAN_IN P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2027_U91
g27793 and P1_INSTADDRPOINTER_REG_23__SCAN_IN P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2027_U92
g27794 and P1_INSTADDRPOINTER_REG_25__SCAN_IN P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2027_U93
g27795 and P1_INSTADDRPOINTER_REG_27__SCAN_IN P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2027_U94
g27796 nand P1_R2027_U118 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2027_U95
g27797 nand P1_R2027_U112 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2027_U96
g27798 nand P1_R2027_U111 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2027_U97
g27799 not P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_R2027_U98
g27800 nand P1_R2027_U128 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2027_U99
g27801 nand P1_INSTADDRPOINTER_REG_0__SCAN_IN P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2027_U100
g27802 nand P1_R2027_U122 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2027_U101
g27803 nand P1_R2027_U116 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2027_U102
g27804 nand P1_R2027_U115 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2027_U103
g27805 nand P1_R2027_U121 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2027_U104
g27806 nand P1_R2027_U114 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2027_U105
g27807 nand P1_R2027_U117 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2027_U106
g27808 nand P1_R2027_U124 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2027_U107
g27809 nand P1_R2027_U119 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2027_U108
g27810 nand P1_R2027_U113 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2027_U109
g27811 nand P1_R2027_U120 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2027_U110
g27812 not P1_R2027_U10 ; P1_R2027_U111
g27813 not P1_R2027_U13 ; P1_R2027_U112
g27814 not P1_R2027_U22 ; P1_R2027_U113
g27815 not P1_R2027_U34 ; P1_R2027_U114
g27816 not P1_R2027_U40 ; P1_R2027_U115
g27817 not P1_R2027_U43 ; P1_R2027_U116
g27818 not P1_R2027_U31 ; P1_R2027_U117
g27819 not P1_R2027_U16 ; P1_R2027_U118
g27820 not P1_R2027_U25 ; P1_R2027_U119
g27821 not P1_R2027_U17 ; P1_R2027_U120
g27822 not P1_R2027_U36 ; P1_R2027_U121
g27823 not P1_R2027_U46 ; P1_R2027_U122
g27824 not P1_R2027_U48 ; P1_R2027_U123
g27825 not P1_R2027_U27 ; P1_R2027_U124
g27826 not P1_R2027_U95 ; P1_R2027_U125
g27827 not P1_R2027_U96 ; P1_R2027_U126
g27828 not P1_R2027_U97 ; P1_R2027_U127
g27829 not P1_R2027_U49 ; P1_R2027_U128
g27830 not P1_R2027_U99 ; P1_R2027_U129
g27831 not P1_R2027_U100 ; P1_R2027_U130
g27832 not P1_R2027_U101 ; P1_R2027_U131
g27833 not P1_R2027_U102 ; P1_R2027_U132
g27834 not P1_R2027_U103 ; P1_R2027_U133
g27835 not P1_R2027_U104 ; P1_R2027_U134
g27836 not P1_R2027_U105 ; P1_R2027_U135
g27837 not P1_R2027_U106 ; P1_R2027_U136
g27838 not P1_R2027_U107 ; P1_R2027_U137
g27839 not P1_R2027_U108 ; P1_R2027_U138
g27840 not P1_R2027_U109 ; P1_R2027_U139
g27841 not P1_R2027_U110 ; P1_R2027_U140
g27842 nand P1_R2027_U120 P1_R2027_U18 ; P1_R2027_U141
g27843 nand P1_R2027_U17 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2027_U142
g27844 nand P1_R2027_U95 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2027_U143
g27845 nand P1_R2027_U125 P1_R2027_U14 ; P1_R2027_U144
g27846 nand P1_R2027_U118 P1_R2027_U15 ; P1_R2027_U145
g27847 nand P1_R2027_U16 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2027_U146
g27848 nand P1_R2027_U96 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2027_U147
g27849 nand P1_R2027_U126 P1_R2027_U11 ; P1_R2027_U148
g27850 nand P1_R2027_U112 P1_R2027_U12 ; P1_R2027_U149
g27851 nand P1_R2027_U13 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2027_U150
g27852 nand P1_R2027_U97 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2027_U151
g27853 nand P1_R2027_U127 P1_R2027_U8 ; P1_R2027_U152
g27854 nand P1_R2027_U111 P1_R2027_U9 ; P1_R2027_U153
g27855 nand P1_R2027_U10 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2027_U154
g27856 nand P1_R2027_U99 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_R2027_U155
g27857 nand P1_R2027_U129 P1_R2027_U98 ; P1_R2027_U156
g27858 nand P1_R2027_U49 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2027_U157
g27859 nand P1_R2027_U128 P1_R2027_U50 ; P1_R2027_U158
g27860 nand P1_R2027_U100 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2027_U159
g27861 nand P1_R2027_U130 P1_R2027_U6 ; P1_R2027_U160
g27862 nand P1_R2027_U123 P1_R2027_U47 ; P1_R2027_U161
g27863 nand P1_R2027_U48 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2027_U162
g27864 nand P1_R2027_U101 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2027_U163
g27865 nand P1_R2027_U131 P1_R2027_U45 ; P1_R2027_U164
g27866 nand P1_R2027_U122 P1_R2027_U44 ; P1_R2027_U165
g27867 nand P1_R2027_U46 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2027_U166
g27868 nand P1_R2027_U102 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2027_U167
g27869 nand P1_R2027_U132 P1_R2027_U41 ; P1_R2027_U168
g27870 nand P1_R2027_U116 P1_R2027_U42 ; P1_R2027_U169
g27871 nand P1_R2027_U43 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2027_U170
g27872 nand P1_R2027_U103 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2027_U171
g27873 nand P1_R2027_U133 P1_R2027_U38 ; P1_R2027_U172
g27874 nand P1_R2027_U115 P1_R2027_U39 ; P1_R2027_U173
g27875 nand P1_R2027_U40 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2027_U174
g27876 nand P1_R2027_U104 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2027_U175
g27877 nand P1_R2027_U134 P1_R2027_U37 ; P1_R2027_U176
g27878 nand P1_R2027_U121 P1_R2027_U35 ; P1_R2027_U177
g27879 nand P1_R2027_U36 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2027_U178
g27880 nand P1_R2027_U105 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2027_U179
g27881 nand P1_R2027_U135 P1_R2027_U32 ; P1_R2027_U180
g27882 nand P1_R2027_U7 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_R2027_U181
g27883 nand P1_R2027_U5 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2027_U182
g27884 nand P1_R2027_U114 P1_R2027_U33 ; P1_R2027_U183
g27885 nand P1_R2027_U34 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2027_U184
g27886 nand P1_R2027_U106 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2027_U185
g27887 nand P1_R2027_U136 P1_R2027_U29 ; P1_R2027_U186
g27888 nand P1_R2027_U117 P1_R2027_U30 ; P1_R2027_U187
g27889 nand P1_R2027_U31 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2027_U188
g27890 nand P1_R2027_U107 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2027_U189
g27891 nand P1_R2027_U137 P1_R2027_U28 ; P1_R2027_U190
g27892 nand P1_R2027_U124 P1_R2027_U26 ; P1_R2027_U191
g27893 nand P1_R2027_U27 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2027_U192
g27894 nand P1_R2027_U108 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2027_U193
g27895 nand P1_R2027_U138 P1_R2027_U23 ; P1_R2027_U194
g27896 nand P1_R2027_U119 P1_R2027_U24 ; P1_R2027_U195
g27897 nand P1_R2027_U25 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2027_U196
g27898 nand P1_R2027_U109 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_R2027_U197
g27899 nand P1_R2027_U139 P1_R2027_U20 ; P1_R2027_U198
g27900 nand P1_R2027_U113 P1_R2027_U21 ; P1_R2027_U199
g27901 nand P1_R2027_U22 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2027_U200
g27902 nand P1_R2027_U110 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2027_U201
g27903 nand P1_R2027_U140 P1_R2027_U19 ; P1_R2027_U202
g27904 and P1_R2182_U47 P1_U2740 ; P1_R2182_U5
g27905 and P1_R2182_U60 P1_R2182_U16 ; P1_R2182_U6
g27906 not P1_U2744 ; P1_R2182_U7
g27907 not P1_U3246 ; P1_R2182_U8
g27908 nand P1_U3246 P1_U2744 ; P1_R2182_U9
g27909 not P1_U2742 ; P1_R2182_U10
g27910 not P1_U2741 ; P1_R2182_U11
g27911 not P1_U2740 ; P1_R2182_U12
g27912 nand P1_R2182_U35 P1_R2182_U41 ; P1_R2182_U13
g27913 not P1_U2737 ; P1_R2182_U14
g27914 not P1_U2738 ; P1_R2182_U15
g27915 nand P1_U2723 P1_U2739 ; P1_R2182_U16
g27916 not P1_U2736 ; P1_R2182_U17
g27917 not P1_U2735 ; P1_R2182_U18
g27918 nand P1_R2182_U36 P1_R2182_U49 ; P1_R2182_U19
g27919 not P1_U2734 ; P1_R2182_U20
g27920 nand P1_R2182_U37 P1_R2182_U46 ; P1_R2182_U21
g27921 nand P1_R2182_U48 P1_U2734 ; P1_R2182_U22
g27922 not P1_U2733 ; P1_R2182_U23
g27923 nand P1_R2182_U64 P1_R2182_U63 ; P1_R2182_U24
g27924 nand P1_R2182_U66 P1_R2182_U65 ; P1_R2182_U25
g27925 nand P1_R2182_U68 P1_R2182_U67 ; P1_R2182_U26
g27926 nand P1_R2182_U72 P1_R2182_U71 ; P1_R2182_U27
g27927 nand P1_R2182_U74 P1_R2182_U73 ; P1_R2182_U28
g27928 nand P1_R2182_U76 P1_R2182_U75 ; P1_R2182_U29
g27929 nand P1_R2182_U78 P1_R2182_U77 ; P1_R2182_U30
g27930 nand P1_R2182_U80 P1_R2182_U79 ; P1_R2182_U31
g27931 nand P1_R2182_U82 P1_R2182_U81 ; P1_R2182_U32
g27932 nand P1_R2182_U84 P1_R2182_U83 ; P1_R2182_U33
g27933 nand P1_R2182_U86 P1_R2182_U85 ; P1_R2182_U34
g27934 and P1_U2742 P1_U2741 ; P1_R2182_U35
g27935 and P1_U2738 P1_U2737 ; P1_R2182_U36
g27936 and P1_U2735 P1_U2736 ; P1_R2182_U37
g27937 nand P1_U2742 P1_R2182_U41 ; P1_R2182_U38
g27938 not P1_U2732 ; P1_R2182_U39
g27939 nand P1_U2733 P1_R2182_U56 ; P1_R2182_U40
g27940 nand P1_R2182_U52 P1_R2182_U53 ; P1_R2182_U41
g27941 and P1_R2182_U70 P1_R2182_U69 ; P1_R2182_U42
g27942 nand P1_R2182_U46 P1_U2736 ; P1_R2182_U43
g27943 nand P1_R2182_U49 P1_U2738 ; P1_R2182_U44
g27944 nand P1_R2182_U51 P1_R2182_U62 ; P1_R2182_U45
g27945 not P1_R2182_U19 ; P1_R2182_U46
g27946 not P1_R2182_U13 ; P1_R2182_U47
g27947 not P1_R2182_U21 ; P1_R2182_U48
g27948 not P1_R2182_U16 ; P1_R2182_U49
g27949 not P1_R2182_U9 ; P1_R2182_U50
g27950 or P1_U2743 P1_U2731 ; P1_R2182_U51
g27951 nand P1_U2731 P1_U2743 ; P1_R2182_U52
g27952 nand P1_R2182_U50 P1_R2182_U51 ; P1_R2182_U53
g27953 not P1_R2182_U41 ; P1_R2182_U54
g27954 not P1_R2182_U38 ; P1_R2182_U55
g27955 not P1_R2182_U22 ; P1_R2182_U56
g27956 not P1_R2182_U40 ; P1_R2182_U57
g27957 not P1_R2182_U43 ; P1_R2182_U58
g27958 not P1_R2182_U44 ; P1_R2182_U59
g27959 or P1_U2739 P1_U2723 ; P1_R2182_U60
g27960 not P1_R2182_U45 ; P1_R2182_U61
g27961 nand P1_U2731 P1_U2743 ; P1_R2182_U62
g27962 nand P1_R2182_U47 P1_R2182_U12 ; P1_R2182_U63
g27963 nand P1_U2740 P1_R2182_U13 ; P1_R2182_U64
g27964 nand P1_U2741 P1_R2182_U38 ; P1_R2182_U65
g27965 nand P1_R2182_U55 P1_R2182_U11 ; P1_R2182_U66
g27966 nand P1_U2732 P1_R2182_U40 ; P1_R2182_U67
g27967 nand P1_R2182_U57 P1_R2182_U39 ; P1_R2182_U68
g27968 nand P1_U2742 P1_R2182_U41 ; P1_R2182_U69
g27969 nand P1_R2182_U54 P1_R2182_U10 ; P1_R2182_U70
g27970 nand P1_U2733 P1_R2182_U22 ; P1_R2182_U71
g27971 nand P1_R2182_U56 P1_R2182_U23 ; P1_R2182_U72
g27972 nand P1_R2182_U48 P1_R2182_U20 ; P1_R2182_U73
g27973 nand P1_U2734 P1_R2182_U21 ; P1_R2182_U74
g27974 nand P1_U2735 P1_R2182_U43 ; P1_R2182_U75
g27975 nand P1_R2182_U58 P1_R2182_U18 ; P1_R2182_U76
g27976 nand P1_R2182_U46 P1_R2182_U17 ; P1_R2182_U77
g27977 nand P1_U2736 P1_R2182_U19 ; P1_R2182_U78
g27978 nand P1_U2737 P1_R2182_U44 ; P1_R2182_U79
g27979 nand P1_R2182_U59 P1_R2182_U14 ; P1_R2182_U80
g27980 nand P1_R2182_U49 P1_R2182_U15 ; P1_R2182_U81
g27981 nand P1_U2738 P1_R2182_U16 ; P1_R2182_U82
g27982 nand P1_R2182_U50 P1_R2182_U45 ; P1_R2182_U83
g27983 nand P1_R2182_U61 P1_R2182_U9 ; P1_R2182_U84
g27984 nand P1_U3246 P1_R2182_U7 ; P1_R2182_U85
g27985 nand P1_U2744 P1_R2182_U8 ; P1_R2182_U86
g27986 and P1_R2144_U104 P1_R2144_U103 ; P1_R2144_U5
g27987 and P1_R2144_U36 P1_R2144_U35 P1_R2144_U27 P1_R2144_U29 ; P1_R2144_U6
g27988 and P1_R2144_U104 P1_R2144_U81 ; P1_R2144_U7
g27989 and P1_R2144_U138 P1_R2144_U136 ; P1_R2144_U8
g27990 and P1_R2144_U128 P1_R2144_U127 ; P1_R2144_U9
g27991 and P1_R2144_U213 P1_R2144_U212 P1_R2144_U82 ; P1_R2144_U10
g27992 nand P1_R2144_U144 P1_R2144_U146 ; P1_R2144_U11
g27993 not P1_U2355 ; P1_R2144_U12
g27994 not P1_U2750 ; P1_R2144_U13
g27995 not P1_U2751 ; P1_R2144_U14
g27996 not P1_U2752 ; P1_R2144_U15
g27997 not P1_U2749 ; P1_R2144_U16
g27998 not P1_U2745 ; P1_R2144_U17
g27999 not P1_U2748 ; P1_R2144_U18
g28000 nand P1_U2748 P1_R2144_U178 ; P1_R2144_U19
g28001 not P1_U2747 ; P1_R2144_U20
g28002 nand P1_U2747 P1_R2144_U170 ; P1_R2144_U21
g28003 not P1_U2746 ; P1_R2144_U22
g28004 nand P1_U2746 P1_R2144_U173 ; P1_R2144_U23
g28005 nand P1_R2144_U79 P1_R2144_U63 ; P1_R2144_U24
g28006 nand P1_R2144_U6 P1_R2144_U79 ; P1_R2144_U25
g28007 nand P1_R2144_U65 P1_R2144_U141 ; P1_R2144_U26
g28008 nand P1_R2144_U206 P1_R2144_U205 ; P1_R2144_U27
g28009 nand P1_R2144_U186 P1_R2144_U185 ; P1_R2144_U28
g28010 nand P1_R2144_U203 P1_R2144_U202 ; P1_R2144_U29
g28011 nand P1_R2144_U209 P1_R2144_U208 ; P1_R2144_U30
g28012 nand P1_R2144_U224 P1_R2144_U223 ; P1_R2144_U31
g28013 nand P1_R2144_U221 P1_R2144_U220 ; P1_R2144_U32
g28014 nand P1_R2144_U227 P1_R2144_U226 ; P1_R2144_U33
g28015 nand P1_R2144_U230 P1_R2144_U229 ; P1_R2144_U34
g28016 nand P1_R2144_U233 P1_R2144_U232 ; P1_R2144_U35
g28017 nand P1_R2144_U236 P1_R2144_U235 ; P1_R2144_U36
g28018 nand P1_R2144_U248 P1_R2144_U247 ; P1_R2144_U37
g28019 nand P1_R2144_U250 P1_R2144_U249 ; P1_R2144_U38
g28020 nand P1_R2144_U252 P1_R2144_U251 ; P1_R2144_U39
g28021 nand P1_R2144_U254 P1_R2144_U253 ; P1_R2144_U40
g28022 nand P1_R2144_U256 P1_R2144_U255 ; P1_R2144_U41
g28023 nand P1_R2144_U258 P1_R2144_U257 ; P1_R2144_U42
g28024 nand P1_R2144_U260 P1_R2144_U259 ; P1_R2144_U43
g28025 and P1_R2144_U21 P1_R2144_U105 ; P1_R2144_U44
g28026 nand P1_R2144_U217 P1_R2144_U216 ; P1_R2144_U45
g28027 and P1_R2144_U19 P1_R2144_U106 ; P1_R2144_U46
g28028 nand P1_R2144_U219 P1_R2144_U218 ; P1_R2144_U47
g28029 and P1_R2144_U162 P1_R2144_U109 ; P1_R2144_U48
g28030 nand P1_R2144_U239 P1_R2144_U238 ; P1_R2144_U49
g28031 nand P1_R2144_U246 P1_R2144_U245 ; P1_R2144_U50
g28032 and P1_R2144_U110 P1_R2144_U109 ; P1_R2144_U51
g28033 and P1_R2144_U106 P1_R2144_U105 ; P1_R2144_U52
g28034 and P1_R2144_U7 P1_R2144_U52 ; P1_R2144_U53
g28035 and P1_R2144_U103 P1_R2144_U151 P1_R2144_U153 P1_R2144_U152 ; P1_R2144_U54
g28036 and P1_R2144_U109 P1_R2144_U106 ; P1_R2144_U55
g28037 and P1_R2144_U159 P1_R2144_U19 ; P1_R2144_U56
g28038 and P1_R2144_U156 P1_R2144_U21 ; P1_R2144_U57
g28039 and P1_R2144_U19 P1_R2144_U21 P1_R2144_U159 ; P1_R2144_U58
g28040 and P1_R2144_U5 P1_R2144_U105 ; P1_R2144_U59
g28041 and P1_R2144_U126 P1_R2144_U21 ; P1_R2144_U60
g28042 and P1_R2144_U23 P1_R2144_U81 ; P1_R2144_U61
g28043 and P1_R2144_U111 P1_R2144_U110 ; P1_R2144_U62
g28044 and P1_R2144_U6 P1_R2144_U64 ; P1_R2144_U63
g28045 and P1_R2144_U34 P1_R2144_U33 P1_R2144_U31 P1_R2144_U32 ; P1_R2144_U64
g28046 and P1_R2144_U34 P1_R2144_U33 ; P1_R2144_U65
g28047 and P1_R2144_U36 P1_R2144_U27 P1_R2144_U29 ; P1_R2144_U66
g28048 and P1_R2144_U29 P1_R2144_U27 ; P1_R2144_U67
g28049 not P1_U2762 ; P1_R2144_U68
g28050 not P1_U2761 ; P1_R2144_U69
g28051 not P1_U2763 ; P1_R2144_U70
g28052 not P1_U2764 ; P1_R2144_U71
g28053 not P1_U2766 ; P1_R2144_U72
g28054 not P1_U2767 ; P1_R2144_U73
g28055 not P1_U2768 ; P1_R2144_U74
g28056 not P1_U2765 ; P1_R2144_U75
g28057 not P1_U2760 ; P1_R2144_U76
g28058 not P1_U2759 ; P1_R2144_U77
g28059 nand P1_R2144_U29 P1_R2144_U79 ; P1_R2144_U78
g28060 nand P1_R2144_U99 P1_R2144_U54 ; P1_R2144_U79
g28061 and P1_R2144_U211 P1_R2144_U210 ; P1_R2144_U80
g28062 nand P1_R2144_U165 P1_R2144_U164 P1_R2144_U22 ; P1_R2144_U81
g28063 and P1_R2144_U215 P1_R2144_U214 ; P1_R2144_U82
g28064 nand P1_R2144_U56 P1_R2144_U158 ; P1_R2144_U83
g28065 nand P1_R2144_U111 P1_R2144_U118 ; P1_R2144_U84
g28066 not P1_U2754 ; P1_R2144_U85
g28067 not P1_U2753 ; P1_R2144_U86
g28068 not P1_U2755 ; P1_R2144_U87
g28069 not P1_U2756 ; P1_R2144_U88
g28070 not P1_U2757 ; P1_R2144_U89
g28071 not P1_U2758 ; P1_R2144_U90
g28072 nand P1_R2144_U100 P1_R2144_U132 ; P1_R2144_U91
g28073 and P1_R2144_U241 P1_R2144_U240 ; P1_R2144_U92
g28074 nand P1_R2144_U129 P1_R2144_U113 ; P1_R2144_U93
g28075 nand P1_R2144_U143 P1_R2144_U32 ; P1_R2144_U94
g28076 nand P1_R2144_U141 P1_R2144_U34 ; P1_R2144_U95
g28077 nand P1_R2144_U79 P1_R2144_U66 ; P1_R2144_U96
g28078 nand P1_R2144_U67 P1_R2144_U79 ; P1_R2144_U97
g28079 nand P1_R2144_U113 P1_R2144_U112 ; P1_R2144_U98
g28080 nand P1_R2144_U53 P1_R2144_U84 ; P1_R2144_U99
g28081 nand P1_U2751 P1_R2144_U28 ; P1_R2144_U100
g28082 not P1_R2144_U24 ; P1_R2144_U101
g28083 not P1_R2144_U81 ; P1_R2144_U102
g28084 nand P1_U2745 P1_R2144_U181 ; P1_R2144_U103
g28085 nand P1_R2144_U167 P1_R2144_U166 P1_R2144_U17 ; P1_R2144_U104
g28086 nand P1_R2144_U175 P1_R2144_U174 P1_R2144_U20 ; P1_R2144_U105
g28087 nand P1_R2144_U201 P1_R2144_U200 P1_R2144_U18 ; P1_R2144_U106
g28088 not P1_R2144_U21 ; P1_R2144_U107
g28089 not P1_R2144_U23 ; P1_R2144_U108
g28090 nand P1_R2144_U194 P1_R2144_U193 P1_R2144_U13 ; P1_R2144_U109
g28091 nand P1_R2144_U196 P1_R2144_U195 P1_R2144_U16 ; P1_R2144_U110
g28092 nand P1_U2749 P1_R2144_U199 ; P1_R2144_U111
g28093 nand P1_R2144_U189 P1_R2144_U188 P1_R2144_U15 ; P1_R2144_U112
g28094 nand P1_U2752 P1_R2144_U192 ; P1_R2144_U113
g28095 nand P1_R2144_U187 P1_R2144_U14 ; P1_R2144_U114
g28096 nand P1_U2355 P1_R2144_U112 ; P1_R2144_U115
g28097 nand P1_U2750 P1_R2144_U184 ; P1_R2144_U116
g28098 nand P1_R2144_U155 P1_R2144_U157 ; P1_R2144_U117
g28099 nand P1_R2144_U51 P1_R2144_U117 ; P1_R2144_U118
g28100 not P1_R2144_U84 ; P1_R2144_U119
g28101 not P1_R2144_U19 ; P1_R2144_U120
g28102 not P1_R2144_U79 ; P1_R2144_U121
g28103 not P1_R2144_U78 ; P1_R2144_U122
g28104 not P1_R2144_U83 ; P1_R2144_U123
g28105 nand P1_R2144_U83 P1_R2144_U105 ; P1_R2144_U124
g28106 nand P1_R2144_U21 P1_R2144_U124 ; P1_R2144_U125
g28107 nand P1_R2144_U23 P1_R2144_U81 ; P1_R2144_U126
g28108 nand P1_R2144_U60 P1_R2144_U124 ; P1_R2144_U127
g28109 nand P1_R2144_U61 P1_R2144_U125 ; P1_R2144_U128
g28110 nand P1_U2355 P1_R2144_U112 ; P1_R2144_U129
g28111 not P1_R2144_U93 ; P1_R2144_U130
g28112 nand P1_R2144_U187 P1_R2144_U14 ; P1_R2144_U131
g28113 nand P1_R2144_U131 P1_R2144_U93 ; P1_R2144_U132
g28114 not P1_R2144_U91 ; P1_R2144_U133
g28115 nand P1_R2144_U91 P1_R2144_U109 ; P1_R2144_U134
g28116 nand P1_R2144_U134 P1_R2144_U116 ; P1_R2144_U135
g28117 nand P1_R2144_U62 P1_R2144_U135 ; P1_R2144_U136
g28118 nand P1_R2144_U161 P1_R2144_U110 ; P1_R2144_U137
g28119 nand P1_R2144_U134 P1_R2144_U116 P1_R2144_U137 ; P1_R2144_U138
g28120 not P1_R2144_U97 ; P1_R2144_U139
g28121 not P1_R2144_U96 ; P1_R2144_U140
g28122 not P1_R2144_U25 ; P1_R2144_U141
g28123 not P1_R2144_U95 ; P1_R2144_U142
g28124 not P1_R2144_U26 ; P1_R2144_U143
g28125 nand P1_U2355 P1_R2144_U24 ; P1_R2144_U144
g28126 not P1_R2144_U144 ; P1_R2144_U145
g28127 nand P1_R2144_U101 P1_R2144_U12 ; P1_R2144_U146
g28128 not P1_R2144_U94 ; P1_R2144_U147
g28129 not P1_R2144_U98 ; P1_R2144_U148
g28130 nand P1_R2144_U21 P1_R2144_U105 ; P1_R2144_U149
g28131 nand P1_R2144_U19 P1_R2144_U106 ; P1_R2144_U150
g28132 nand P1_R2144_U120 P1_R2144_U105 P1_R2144_U7 ; P1_R2144_U151
g28133 nand P1_R2144_U107 P1_R2144_U7 ; P1_R2144_U152
g28134 nand P1_R2144_U108 P1_R2144_U7 ; P1_R2144_U153
g28135 nand P1_R2144_U113 P1_R2144_U115 P1_R2144_U100 ; P1_R2144_U154
g28136 nand P1_R2144_U154 P1_R2144_U114 ; P1_R2144_U155
g28137 nand P1_R2144_U104 P1_R2144_U103 ; P1_R2144_U156
g28138 nand P1_U2750 P1_R2144_U184 ; P1_R2144_U157
g28139 nand P1_R2144_U117 P1_R2144_U110 P1_R2144_U55 ; P1_R2144_U158
g28140 nand P1_U2749 P1_R2144_U106 P1_R2144_U199 ; P1_R2144_U159
g28141 nand P1_R2144_U58 P1_R2144_U158 ; P1_R2144_U160
g28142 nand P1_U2749 P1_R2144_U199 ; P1_R2144_U161
g28143 nand P1_U2750 P1_R2144_U184 ; P1_R2144_U162
g28144 nand P1_R2144_U116 P1_R2144_U109 ; P1_R2144_U163
g28145 nand P1_U2355 P1_R2144_U68 ; P1_R2144_U164
g28146 nand P1_U2762 P1_R2144_U12 ; P1_R2144_U165
g28147 nand P1_U2355 P1_R2144_U69 ; P1_R2144_U166
g28148 nand P1_U2761 P1_R2144_U12 ; P1_R2144_U167
g28149 nand P1_U2355 P1_R2144_U70 ; P1_R2144_U168
g28150 nand P1_U2763 P1_R2144_U12 ; P1_R2144_U169
g28151 nand P1_R2144_U169 P1_R2144_U168 ; P1_R2144_U170
g28152 nand P1_U2355 P1_R2144_U68 ; P1_R2144_U171
g28153 nand P1_U2762 P1_R2144_U12 ; P1_R2144_U172
g28154 nand P1_R2144_U172 P1_R2144_U171 ; P1_R2144_U173
g28155 nand P1_U2355 P1_R2144_U70 ; P1_R2144_U174
g28156 nand P1_U2763 P1_R2144_U12 ; P1_R2144_U175
g28157 nand P1_U2355 P1_R2144_U71 ; P1_R2144_U176
g28158 nand P1_U2764 P1_R2144_U12 ; P1_R2144_U177
g28159 nand P1_R2144_U177 P1_R2144_U176 ; P1_R2144_U178
g28160 nand P1_U2355 P1_R2144_U69 ; P1_R2144_U179
g28161 nand P1_U2761 P1_R2144_U12 ; P1_R2144_U180
g28162 nand P1_R2144_U180 P1_R2144_U179 ; P1_R2144_U181
g28163 nand P1_U2355 P1_R2144_U72 ; P1_R2144_U182
g28164 nand P1_U2766 P1_R2144_U12 ; P1_R2144_U183
g28165 nand P1_R2144_U183 P1_R2144_U182 ; P1_R2144_U184
g28166 nand P1_U2355 P1_R2144_U73 ; P1_R2144_U185
g28167 nand P1_U2767 P1_R2144_U12 ; P1_R2144_U186
g28168 not P1_R2144_U28 ; P1_R2144_U187
g28169 nand P1_U2355 P1_R2144_U74 ; P1_R2144_U188
g28170 nand P1_U2768 P1_R2144_U12 ; P1_R2144_U189
g28171 nand P1_U2355 P1_R2144_U74 ; P1_R2144_U190
g28172 nand P1_U2768 P1_R2144_U12 ; P1_R2144_U191
g28173 nand P1_R2144_U191 P1_R2144_U190 ; P1_R2144_U192
g28174 nand P1_U2355 P1_R2144_U72 ; P1_R2144_U193
g28175 nand P1_U2766 P1_R2144_U12 ; P1_R2144_U194
g28176 nand P1_U2355 P1_R2144_U75 ; P1_R2144_U195
g28177 nand P1_U2765 P1_R2144_U12 ; P1_R2144_U196
g28178 nand P1_U2355 P1_R2144_U75 ; P1_R2144_U197
g28179 nand P1_U2765 P1_R2144_U12 ; P1_R2144_U198
g28180 nand P1_R2144_U198 P1_R2144_U197 ; P1_R2144_U199
g28181 nand P1_U2355 P1_R2144_U71 ; P1_R2144_U200
g28182 nand P1_U2764 P1_R2144_U12 ; P1_R2144_U201
g28183 nand P1_U2355 P1_R2144_U76 ; P1_R2144_U202
g28184 nand P1_U2760 P1_R2144_U12 ; P1_R2144_U203
g28185 not P1_R2144_U29 ; P1_R2144_U204
g28186 nand P1_U2355 P1_R2144_U77 ; P1_R2144_U205
g28187 nand P1_U2759 P1_R2144_U12 ; P1_R2144_U206
g28188 not P1_R2144_U27 ; P1_R2144_U207
g28189 nand P1_R2144_U122 P1_R2144_U207 ; P1_R2144_U208
g28190 nand P1_R2144_U27 P1_R2144_U78 ; P1_R2144_U209
g28191 nand P1_R2144_U121 P1_R2144_U204 ; P1_R2144_U210
g28192 nand P1_R2144_U29 P1_R2144_U79 ; P1_R2144_U211
g28193 nand P1_R2144_U57 P1_R2144_U124 P1_R2144_U23 ; P1_R2144_U212
g28194 nand P1_R2144_U5 P1_R2144_U108 ; P1_R2144_U213
g28195 nand P1_R2144_U102 P1_R2144_U156 ; P1_R2144_U214
g28196 nand P1_R2144_U59 P1_R2144_U160 P1_R2144_U81 ; P1_R2144_U215
g28197 nand P1_R2144_U149 P1_R2144_U83 ; P1_R2144_U216
g28198 nand P1_R2144_U44 P1_R2144_U123 ; P1_R2144_U217
g28199 nand P1_R2144_U150 P1_R2144_U84 ; P1_R2144_U218
g28200 nand P1_R2144_U46 P1_R2144_U119 ; P1_R2144_U219
g28201 nand P1_U2355 P1_R2144_U85 ; P1_R2144_U220
g28202 nand P1_U2754 P1_R2144_U12 ; P1_R2144_U221
g28203 not P1_R2144_U32 ; P1_R2144_U222
g28204 nand P1_U2355 P1_R2144_U86 ; P1_R2144_U223
g28205 nand P1_U2753 P1_R2144_U12 ; P1_R2144_U224
g28206 not P1_R2144_U31 ; P1_R2144_U225
g28207 nand P1_U2355 P1_R2144_U87 ; P1_R2144_U226
g28208 nand P1_U2755 P1_R2144_U12 ; P1_R2144_U227
g28209 not P1_R2144_U33 ; P1_R2144_U228
g28210 nand P1_U2355 P1_R2144_U88 ; P1_R2144_U229
g28211 nand P1_U2756 P1_R2144_U12 ; P1_R2144_U230
g28212 not P1_R2144_U34 ; P1_R2144_U231
g28213 nand P1_U2355 P1_R2144_U89 ; P1_R2144_U232
g28214 nand P1_U2757 P1_R2144_U12 ; P1_R2144_U233
g28215 not P1_R2144_U35 ; P1_R2144_U234
g28216 nand P1_U2355 P1_R2144_U90 ; P1_R2144_U235
g28217 nand P1_U2758 P1_R2144_U12 ; P1_R2144_U236
g28218 not P1_R2144_U36 ; P1_R2144_U237
g28219 nand P1_R2144_U163 P1_R2144_U91 ; P1_R2144_U238
g28220 nand P1_R2144_U48 P1_R2144_U133 ; P1_R2144_U239
g28221 nand P1_R2144_U187 P1_U2751 ; P1_R2144_U240
g28222 nand P1_R2144_U28 P1_R2144_U14 ; P1_R2144_U241
g28223 nand P1_R2144_U187 P1_U2751 ; P1_R2144_U242
g28224 nand P1_R2144_U28 P1_R2144_U14 ; P1_R2144_U243
g28225 nand P1_R2144_U243 P1_R2144_U242 ; P1_R2144_U244
g28226 nand P1_R2144_U92 P1_R2144_U93 ; P1_R2144_U245
g28227 nand P1_R2144_U130 P1_R2144_U244 ; P1_R2144_U246
g28228 nand P1_R2144_U147 P1_R2144_U225 ; P1_R2144_U247
g28229 nand P1_R2144_U31 P1_R2144_U94 ; P1_R2144_U248
g28230 nand P1_R2144_U222 P1_R2144_U143 ; P1_R2144_U249
g28231 nand P1_R2144_U32 P1_R2144_U26 ; P1_R2144_U250
g28232 nand P1_R2144_U142 P1_R2144_U228 ; P1_R2144_U251
g28233 nand P1_R2144_U33 P1_R2144_U95 ; P1_R2144_U252
g28234 nand P1_R2144_U231 P1_R2144_U141 ; P1_R2144_U253
g28235 nand P1_R2144_U34 P1_R2144_U25 ; P1_R2144_U254
g28236 nand P1_R2144_U140 P1_R2144_U234 ; P1_R2144_U255
g28237 nand P1_R2144_U35 P1_R2144_U96 ; P1_R2144_U256
g28238 nand P1_R2144_U139 P1_R2144_U237 ; P1_R2144_U257
g28239 nand P1_R2144_U36 P1_R2144_U97 ; P1_R2144_U258
g28240 nand P1_U2355 P1_R2144_U98 ; P1_R2144_U259
g28241 nand P1_R2144_U148 P1_R2144_U12 ; P1_R2144_U260
g28242 and P1_R2278_U466 P1_R2278_U327 ; P1_R2278_U5
g28243 and P1_R2278_U292 P1_R2278_U288 ; P1_R2278_U6
g28244 and P1_R2278_U6 P1_R2278_U295 ; P1_R2278_U7
g28245 and P1_R2278_U302 P1_R2278_U298 P1_R2278_U305 ; P1_R2278_U8
g28246 and P1_R2278_U8 P1_R2278_U308 ; P1_R2278_U9
g28247 and P1_R2278_U313 P1_R2278_U311 P1_R2278_U315 ; P1_R2278_U10
g28248 and P1_R2278_U134 P1_R2278_U10 ; P1_R2278_U11
g28249 and P1_R2278_U295 P1_R2278_U292 ; P1_R2278_U12
g28250 and P1_R2278_U9 P1_R2278_U321 ; P1_R2278_U13
g28251 and P1_R2278_U463 P1_R2278_U462 ; P1_R2278_U14
g28252 and P1_R2278_U344 P1_R2278_U342 ; P1_R2278_U15
g28253 and P1_R2278_U188 P1_R2278_U375 P1_R2278_U468 P1_R2278_U467 ; P1_R2278_U16
g28254 and P1_R2278_U272 P1_R2278_U270 ; P1_R2278_U17
g28255 and P1_R2278_U268 P1_R2278_U266 ; P1_R2278_U18
g28256 nand P1_R2278_U214 P1_R2278_U429 ; P1_R2278_U19
g28257 and P1_R2278_U414 P1_R2278_U335 ; P1_R2278_U20
g28258 not P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2278_U21
g28259 not P1_U2792 ; P1_R2278_U22
g28260 not P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2278_U23
g28261 not P1_U2793 ; P1_R2278_U24
g28262 not P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2278_U25
g28263 not P1_U2794 ; P1_R2278_U26
g28264 not P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2278_U27
g28265 not P1_U2795 ; P1_R2278_U28
g28266 not P1_U2800 ; P1_R2278_U29
g28267 not P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_R2278_U30
g28268 not P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2278_U31
g28269 nand P1_U2800 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_R2278_U32
g28270 not P1_U2799 ; P1_R2278_U33
g28271 not P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2278_U34
g28272 not P1_U2798 ; P1_R2278_U35
g28273 not P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2278_U36
g28274 not P1_U2797 ; P1_R2278_U37
g28275 not P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2278_U38
g28276 not P1_U2796 ; P1_R2278_U39
g28277 nand P1_R2278_U43 P1_R2278_U250 ; P1_R2278_U40
g28278 nand P1_R2278_U254 P1_R2278_U252 P1_R2278_U253 ; P1_R2278_U41
g28279 nand P1_R2278_U246 P1_R2278_U245 ; P1_R2278_U42
g28280 nand P1_R2278_U42 P1_R2278_U248 ; P1_R2278_U43
g28281 not P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2278_U44
g28282 not P1_U2775 ; P1_R2278_U45
g28283 not P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2278_U46
g28284 not P1_U2774 ; P1_R2278_U47
g28285 not P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2278_U48
g28286 not P1_U2776 ; P1_R2278_U49
g28287 not P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2278_U50
g28288 not P1_U2777 ; P1_R2278_U51
g28289 not P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2278_U52
g28290 not P1_U2779 ; P1_R2278_U53
g28291 not P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2278_U54
g28292 not P1_U2780 ; P1_R2278_U55
g28293 not P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2278_U56
g28294 not P1_U2781 ; P1_R2278_U57
g28295 not P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2278_U58
g28296 not P1_U2789 ; P1_R2278_U59
g28297 not P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2278_U60
g28298 not P1_U2790 ; P1_R2278_U61
g28299 not P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2278_U62
g28300 not P1_U2785 ; P1_R2278_U63
g28301 not P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2278_U64
g28302 not P1_U2787 ; P1_R2278_U65
g28303 not P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2278_U66
g28304 not P1_U2786 ; P1_R2278_U67
g28305 nand P1_U2788 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_R2278_U68
g28306 not P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2278_U69
g28307 not P1_U2784 ; P1_R2278_U70
g28308 not P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2278_U71
g28309 not P1_U2783 ; P1_R2278_U72
g28310 nand P1_R2278_U12 P1_R2278_U8 P1_R2278_U359 P1_R2278_U308 ; P1_R2278_U73
g28311 not P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2278_U74
g28312 not P1_U2778 ; P1_R2278_U75
g28313 nand P1_U2778 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2278_U76
g28314 not P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2278_U77
g28315 not P1_U2782 ; P1_R2278_U78
g28316 nand P1_U2782 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2278_U79
g28317 nand P1_R2278_U144 P1_R2278_U8 ; P1_R2278_U80
g28318 not P1_U2772 ; P1_R2278_U81
g28319 not P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2278_U82
g28320 not P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2278_U83
g28321 not P1_U2773 ; P1_R2278_U84
g28322 nand P1_U2773 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2278_U85
g28323 nand P1_R2278_U379 P1_R2278_U322 ; P1_R2278_U86
g28324 nand P1_R2278_U392 P1_R2278_U92 P1_R2278_U93 ; P1_R2278_U87
g28325 not P1_U2770 ; P1_R2278_U88
g28326 not P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2278_U89
g28327 not P1_U2771 ; P1_R2278_U90
g28328 not P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2278_U91
g28329 nand P1_R2278_U143 P1_R2278_U11 ; P1_R2278_U92
g28330 nand P1_R2278_U11 P1_R2278_U321 P1_R2278_U377 ; P1_R2278_U93
g28331 nand P1_R2278_U132 P1_R2278_U372 ; P1_R2278_U94
g28332 nand P1_R2278_U136 P1_R2278_U368 ; P1_R2278_U95
g28333 nand P1_R2278_U11 P1_R2278_U321 P1_R2278_U378 ; P1_R2278_U96
g28334 nand P1_R2278_U229 P1_R2278_U331 ; P1_R2278_U97
g28335 nand P1_R2278_U138 P1_R2278_U354 ; P1_R2278_U98
g28336 nand P1_R2278_U610 P1_R2278_U609 ; P1_R2278_U99
g28337 and P1_R2278_U262 P1_R2278_U261 ; P1_R2278_U100
g28338 nand P1_R2278_U431 P1_R2278_U430 ; P1_R2278_U101
g28339 nand P1_R2278_U438 P1_R2278_U437 ; P1_R2278_U102
g28340 nand P1_R2278_U445 P1_R2278_U444 ; P1_R2278_U103
g28341 nand P1_R2278_U454 P1_R2278_U453 ; P1_R2278_U104
g28342 nand P1_R2278_U461 P1_R2278_U460 ; P1_R2278_U105
g28343 nand P1_R2278_U477 P1_R2278_U476 ; P1_R2278_U106
g28344 nand P1_R2278_U484 P1_R2278_U483 ; P1_R2278_U107
g28345 nand P1_R2278_U491 P1_R2278_U490 ; P1_R2278_U108
g28346 nand P1_R2278_U498 P1_R2278_U497 ; P1_R2278_U109
g28347 nand P1_R2278_U505 P1_R2278_U504 ; P1_R2278_U110
g28348 nand P1_R2278_U512 P1_R2278_U511 ; P1_R2278_U111
g28349 nand P1_R2278_U519 P1_R2278_U518 ; P1_R2278_U112
g28350 nand P1_R2278_U526 P1_R2278_U525 ; P1_R2278_U113
g28351 nand P1_R2278_U533 P1_R2278_U532 ; P1_R2278_U114
g28352 nand P1_R2278_U540 P1_R2278_U539 ; P1_R2278_U115
g28353 nand P1_R2278_U547 P1_R2278_U546 ; P1_R2278_U116
g28354 nand P1_R2278_U554 P1_R2278_U553 ; P1_R2278_U117
g28355 nand P1_R2278_U566 P1_R2278_U565 ; P1_R2278_U118
g28356 nand P1_R2278_U573 P1_R2278_U572 ; P1_R2278_U119
g28357 nand P1_R2278_U580 P1_R2278_U579 ; P1_R2278_U120
g28358 nand P1_R2278_U587 P1_R2278_U586 ; P1_R2278_U121
g28359 nand P1_R2278_U594 P1_R2278_U593 ; P1_R2278_U122
g28360 nand P1_R2278_U599 P1_R2278_U598 ; P1_R2278_U123
g28361 and P1_R2278_U68 P1_R2278_U281 ; P1_R2278_U124
g28362 nand P1_R2278_U601 P1_R2278_U600 ; P1_R2278_U125
g28363 nand P1_R2278_U608 P1_R2278_U607 ; P1_R2278_U126
g28364 and P1_U2793 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2278_U127
g28365 and P1_R2278_U258 P1_R2278_U254 ; P1_R2278_U128
g28366 and P1_R2278_U352 P1_R2278_U259 ; P1_R2278_U129
g28367 and P1_U2777 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2278_U130
g28368 and P1_R2278_U318 P1_R2278_U316 ; P1_R2278_U131
g28369 and P1_R2278_U319 P1_R2278_U317 P1_R2278_U321 ; P1_R2278_U132
g28370 and P1_U2781 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2278_U133
g28371 and P1_R2278_U319 P1_R2278_U317 ; P1_R2278_U134
g28372 and P1_R2278_U321 P1_R2278_U308 ; P1_R2278_U135
g28373 and P1_R2278_U11 P1_R2278_U135 ; P1_R2278_U136
g28374 and P1_R2278_U259 P1_R2278_U228 P1_R2278_U273 ; P1_R2278_U137
g28375 and P1_R2278_U389 P1_R2278_U276 ; P1_R2278_U138
g28376 and P1_R2278_U357 P1_R2278_U140 ; P1_R2278_U139
g28377 and P1_R2278_U281 P1_R2278_U283 P1_R2278_U284 ; P1_R2278_U140
g28378 and P1_R2278_U286 P1_R2278_U410 ; P1_R2278_U141
g28379 and P1_R2278_U7 P1_R2278_U13 ; P1_R2278_U142
g28380 and P1_R2278_U309 P1_R2278_U321 ; P1_R2278_U143
g28381 and P1_R2278_U296 P1_R2278_U308 ; P1_R2278_U144
g28382 and P1_R2278_U95 P1_R2278_U94 ; P1_R2278_U145
g28383 and P1_R2278_U401 P1_R2278_U96 ; P1_R2278_U146
g28384 and P1_R2278_U324 P1_R2278_U5 ; P1_R2278_U147
g28385 and P1_R2278_U324 P1_R2278_U321 P1_R2278_U319 P1_R2278_U317 ; P1_R2278_U148
g28386 and P1_R2278_U321 P1_R2278_U308 P1_R2278_U324 ; P1_R2278_U149
g28387 and P1_R2278_U11 P1_R2278_U149 ; P1_R2278_U150
g28388 and P1_R2278_U286 P1_R2278_U412 ; P1_R2278_U151
g28389 and P1_R2278_U11 P1_R2278_U324 ; P1_R2278_U152
g28390 and P1_R2278_U7 P1_R2278_U13 ; P1_R2278_U153
g28391 and P1_R2278_U324 P1_R2278_U321 ; P1_R2278_U154
g28392 and P1_R2278_U394 P1_R2278_U393 P1_R2278_U395 P1_R2278_U398 P1_R2278_U156 ; P1_R2278_U155
g28393 and P1_R2278_U14 P1_R2278_U400 P1_R2278_U399 ; P1_R2278_U156
g28394 and P1_R2278_U11 P1_R2278_U324 ; P1_R2278_U157
g28395 and P1_R2278_U7 P1_R2278_U13 ; P1_R2278_U158
g28396 and P1_R2278_U403 P1_R2278_U187 P1_R2278_U404 ; P1_R2278_U159
g28397 and P1_R2278_U286 P1_R2278_U417 ; P1_R2278_U160
g28398 and P1_R2278_U9 P1_R2278_U7 ; P1_R2278_U161
g28399 and P1_R2278_U369 P1_R2278_U76 ; P1_R2278_U162
g28400 and P1_R2278_U73 P1_R2278_U80 ; P1_R2278_U163
g28401 and P1_R2278_U317 P1_R2278_U10 ; P1_R2278_U164
g28402 and P1_R2278_U371 P1_R2278_U316 ; P1_R2278_U165
g28403 and P1_R2278_U311 P1_R2278_U313 ; P1_R2278_U166
g28404 and P1_R2278_U370 P1_R2278_U314 ; P1_R2278_U167
g28405 and P1_R2278_U286 P1_R2278_U415 ; P1_R2278_U168
g28406 and P1_R2278_U362 P1_R2278_U79 ; P1_R2278_U169
g28407 and P1_R2278_U367 P1_R2278_U306 ; P1_R2278_U170
g28408 and P1_R2278_U298 P1_R2278_U302 ; P1_R2278_U171
g28409 and P1_R2278_U364 P1_R2278_U303 ; P1_R2278_U172
g28410 and P1_R2278_U589 P1_R2278_U588 P1_R2278_U285 ; P1_R2278_U173
g28411 and P1_R2278_U337 P1_R2278_U227 ; P1_R2278_U174
g28412 and P1_R2278_U603 P1_R2278_U602 P1_R2278_U228 ; P1_R2278_U175
g28413 nand P1_R2278_U129 P1_R2278_U353 ; P1_R2278_U176
g28414 and P1_R2278_U433 P1_R2278_U432 ; P1_R2278_U177
g28415 nand P1_R2278_U41 P1_R2278_U256 ; P1_R2278_U178
g28416 and P1_R2278_U440 P1_R2278_U439 ; P1_R2278_U179
g28417 and P1_R2278_U447 P1_R2278_U446 ; P1_R2278_U180
g28418 and P1_R2278_U449 P1_R2278_U448 ; P1_R2278_U181
g28419 nand P1_R2278_U242 P1_R2278_U241 ; P1_R2278_U182
g28420 and P1_R2278_U456 P1_R2278_U455 ; P1_R2278_U183
g28421 nand P1_R2278_U238 P1_R2278_U237 ; P1_R2278_U184
g28422 not P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_R2278_U185
g28423 not P1_U2769 ; P1_R2278_U186
g28424 nand P1_U2771 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2278_U187
g28425 and P1_R2278_U470 P1_R2278_U469 ; P1_R2278_U188
g28426 and P1_R2278_U472 P1_R2278_U471 ; P1_R2278_U189
g28427 nand P1_R2278_U406 P1_R2278_U405 P1_R2278_U407 P1_R2278_U159 ; P1_R2278_U190
g28428 and P1_R2278_U479 P1_R2278_U478 ; P1_R2278_U191
g28429 nand P1_R2278_U213 P1_R2278_U234 ; P1_R2278_U192
g28430 and P1_R2278_U486 P1_R2278_U485 ; P1_R2278_U193
g28431 nand P1_R2278_U145 P1_R2278_U385 P1_R2278_U146 ; P1_R2278_U194
g28432 and P1_R2278_U493 P1_R2278_U492 ; P1_R2278_U195
g28433 nand P1_R2278_U419 P1_R2278_U409 ; P1_R2278_U196
g28434 and P1_R2278_U500 P1_R2278_U499 ; P1_R2278_U197
g28435 nand P1_R2278_U425 P1_R2278_U373 ; P1_R2278_U198
g28436 and P1_R2278_U507 P1_R2278_U506 ; P1_R2278_U199
g28437 nand P1_R2278_U165 P1_R2278_U423 ; P1_R2278_U200
g28438 and P1_R2278_U514 P1_R2278_U513 ; P1_R2278_U201
g28439 nand P1_R2278_U167 P1_R2278_U427 ; P1_R2278_U202
g28440 and P1_R2278_U521 P1_R2278_U520 ; P1_R2278_U203
g28441 nand P1_R2278_U421 P1_R2278_U312 ; P1_R2278_U204
g28442 and P1_R2278_U528 P1_R2278_U527 ; P1_R2278_U205
g28443 nand P1_R2278_U163 P1_R2278_U376 P1_R2278_U162 ; P1_R2278_U206
g28444 and P1_R2278_U535 P1_R2278_U534 ; P1_R2278_U207
g28445 nand P1_R2278_U170 P1_R2278_U365 ; P1_R2278_U208
g28446 and P1_R2278_U542 P1_R2278_U541 ; P1_R2278_U209
g28447 nand P1_R2278_U172 P1_R2278_U363 ; P1_R2278_U210
g28448 and P1_R2278_U549 P1_R2278_U548 ; P1_R2278_U211
g28449 nand P1_R2278_U300 P1_R2278_U299 ; P1_R2278_U212
g28450 nand P1_U2799 P1_R2278_U232 ; P1_R2278_U213
g28451 and P1_R2278_U559 P1_R2278_U558 ; P1_R2278_U214
g28452 and P1_R2278_U561 P1_R2278_U560 ; P1_R2278_U215
g28453 nand P1_R2278_U169 P1_R2278_U361 ; P1_R2278_U216
g28454 and P1_R2278_U568 P1_R2278_U567 ; P1_R2278_U217
g28455 nand P1_R2278_U360 P1_R2278_U358 ; P1_R2278_U218
g28456 and P1_R2278_U575 P1_R2278_U574 ; P1_R2278_U219
g28457 nand P1_R2278_U290 P1_R2278_U289 ; P1_R2278_U220
g28458 and P1_R2278_U582 P1_R2278_U581 ; P1_R2278_U221
g28459 nand P1_R2278_U168 P1_R2278_U226 ; P1_R2278_U222
g28460 nand P1_R2278_U68 P1_R2278_U328 ; P1_R2278_U223
g28461 nand P1_R2278_U98 P1_R2278_U279 ; P1_R2278_U224
g28462 nand P1_R2278_U274 P1_R2278_U273 ; P1_R2278_U225
g28463 nand P1_R2278_U224 P1_R2278_U139 ; P1_R2278_U226
g28464 nand P1_R2278_U356 P1_R2278_U355 ; P1_R2278_U227
g28465 nand P1_U2790 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2278_U228
g28466 nand P1_U2787 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2278_U229
g28467 not P1_R2278_U213 ; P1_R2278_U230
g28468 nand P1_U2794 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2278_U231
g28469 not P1_R2278_U32 ; P1_R2278_U232
g28470 nand P1_R2278_U33 P1_R2278_U32 ; P1_R2278_U233
g28471 nand P1_R2278_U233 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2278_U234
g28472 not P1_R2278_U192 ; P1_R2278_U235
g28473 or P1_U2798 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2278_U236
g28474 nand P1_R2278_U236 P1_R2278_U192 ; P1_R2278_U237
g28475 nand P1_U2798 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2278_U238
g28476 not P1_R2278_U184 ; P1_R2278_U239
g28477 or P1_U2797 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2278_U240
g28478 nand P1_R2278_U240 P1_R2278_U184 ; P1_R2278_U241
g28479 nand P1_U2797 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2278_U242
g28480 not P1_R2278_U182 ; P1_R2278_U243
g28481 or P1_U2796 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2278_U244
g28482 nand P1_R2278_U244 P1_R2278_U182 ; P1_R2278_U245
g28483 nand P1_U2796 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2278_U246
g28484 not P1_R2278_U42 ; P1_R2278_U247
g28485 or P1_U2795 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2278_U248
g28486 not P1_R2278_U43 ; P1_R2278_U249
g28487 nand P1_U2795 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2278_U250
g28488 not P1_R2278_U40 ; P1_R2278_U251
g28489 nand P1_R2278_U251 P1_R2278_U231 ; P1_R2278_U252
g28490 or P1_U2793 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2278_U253
g28491 or P1_U2794 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2278_U254
g28492 not P1_R2278_U41 ; P1_R2278_U255
g28493 nand P1_U2793 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2278_U256
g28494 not P1_R2278_U178 ; P1_R2278_U257
g28495 or P1_U2792 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2278_U258
g28496 nand P1_U2792 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2278_U259
g28497 not P1_R2278_U176 ; P1_R2278_U260
g28498 or P1_U2791 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2278_U261
g28499 nand P1_U2791 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2278_U262
g28500 nand P1_U2791 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2278_U263
g28501 or P1_U2794 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2278_U264
g28502 nand P1_R2278_U264 P1_R2278_U40 ; P1_R2278_U265
g28503 nand P1_R2278_U265 P1_R2278_U231 P1_R2278_U179 ; P1_R2278_U266
g28504 nand P1_U2793 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2278_U267
g28505 nand P1_R2278_U255 P1_R2278_U267 ; P1_R2278_U268
g28506 or P1_U2794 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2278_U269
g28507 nand P1_R2278_U180 P1_R2278_U247 ; P1_R2278_U270
g28508 nand P1_U2795 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2278_U271
g28509 nand P1_R2278_U249 P1_R2278_U271 ; P1_R2278_U272
g28510 nand P1_U2791 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_R2278_U273
g28511 nand P1_R2278_U261 P1_R2278_U176 ; P1_R2278_U274
g28512 not P1_R2278_U225 ; P1_R2278_U275
g28513 or P1_U2789 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2278_U276
g28514 or P1_U2790 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2278_U277
g28515 not P1_R2278_U98 ; P1_R2278_U278
g28516 nand P1_U2789 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2278_U279
g28517 not P1_R2278_U224 ; P1_R2278_U280
g28518 or P1_U2788 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_R2278_U281
g28519 not P1_R2278_U68 ; P1_R2278_U282
g28520 or P1_U2787 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2278_U283
g28521 or P1_U2786 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2278_U284
g28522 nand P1_U2786 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2278_U285
g28523 nand P1_U2785 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2278_U286
g28524 nand P1_R2278_U391 P1_R2278_U229 P1_R2278_U285 ; P1_R2278_U287
g28525 or P1_U2784 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2278_U288
g28526 nand P1_R2278_U288 P1_R2278_U222 ; P1_R2278_U289
g28527 nand P1_U2784 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2278_U290
g28528 not P1_R2278_U220 ; P1_R2278_U291
g28529 or P1_U2783 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2278_U292
g28530 nand P1_U2783 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2278_U293
g28531 not P1_R2278_U218 ; P1_R2278_U294
g28532 or P1_U2782 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2278_U295
g28533 not P1_R2278_U79 ; P1_R2278_U296
g28534 not P1_R2278_U216 ; P1_R2278_U297
g28535 or P1_U2781 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2278_U298
g28536 nand P1_R2278_U298 P1_R2278_U216 ; P1_R2278_U299
g28537 nand P1_U2781 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2278_U300
g28538 not P1_R2278_U212 ; P1_R2278_U301
g28539 or P1_U2780 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2278_U302
g28540 nand P1_U2780 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2278_U303
g28541 not P1_R2278_U210 ; P1_R2278_U304
g28542 or P1_U2779 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2278_U305
g28543 nand P1_U2779 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2278_U306
g28544 not P1_R2278_U208 ; P1_R2278_U307
g28545 or P1_U2778 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2278_U308
g28546 not P1_R2278_U76 ; P1_R2278_U309
g28547 not P1_R2278_U206 ; P1_R2278_U310
g28548 or P1_U2777 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2278_U311
g28549 nand P1_U2777 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2278_U312
g28550 or P1_U2776 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2278_U313
g28551 nand P1_U2776 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2278_U314
g28552 or P1_U2775 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2278_U315
g28553 nand P1_U2775 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2278_U316
g28554 or P1_U2774 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2278_U317
g28555 nand P1_U2774 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2278_U318
g28556 or P1_U2773 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2278_U319
g28557 not P1_R2278_U85 ; P1_R2278_U320
g28558 or P1_U2772 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2278_U321
g28559 nand P1_U2772 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2278_U322
g28560 not P1_R2278_U194 ; P1_R2278_U323
g28561 or P1_U2771 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2278_U324
g28562 not P1_R2278_U187 ; P1_R2278_U325
g28563 not P1_R2278_U190 ; P1_R2278_U326
g28564 or P1_U2770 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2278_U327
g28565 nand P1_R2278_U281 P1_R2278_U224 ; P1_R2278_U328
g28566 not P1_R2278_U223 ; P1_R2278_U329
g28567 or P1_U2787 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2278_U330
g28568 nand P1_R2278_U330 P1_R2278_U223 ; P1_R2278_U331
g28569 not P1_R2278_U97 ; P1_R2278_U332
g28570 or P1_U2786 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2278_U333
g28571 nand P1_R2278_U333 P1_R2278_U97 ; P1_R2278_U334
g28572 nand P1_R2278_U173 P1_R2278_U334 ; P1_R2278_U335
g28573 nand P1_R2278_U332 P1_R2278_U285 ; P1_R2278_U336
g28574 nand P1_U2785 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2278_U337
g28575 or P1_U2786 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2278_U338
g28576 or P1_U2787 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2278_U339
g28577 or P1_U2790 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2278_U340
g28578 nand P1_R2278_U340 P1_R2278_U225 ; P1_R2278_U341
g28579 nand P1_R2278_U175 P1_R2278_U341 ; P1_R2278_U342
g28580 nand P1_U2789 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2278_U343
g28581 nand P1_R2278_U278 P1_R2278_U343 ; P1_R2278_U344
g28582 or P1_U2790 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2278_U345
g28583 nand P1_R2278_U263 P1_R2278_U261 ; P1_R2278_U346
g28584 nand P1_R2278_U269 P1_R2278_U231 ; P1_R2278_U347
g28585 nand P1_R2278_U338 P1_R2278_U285 ; P1_R2278_U348
g28586 nand P1_R2278_U339 P1_R2278_U229 ; P1_R2278_U349
g28587 nand P1_R2278_U68 P1_R2278_U281 ; P1_R2278_U350
g28588 nand P1_R2278_U345 P1_R2278_U228 ; P1_R2278_U351
g28589 nand P1_R2278_U127 P1_R2278_U258 ; P1_R2278_U352
g28590 nand P1_R2278_U253 P1_R2278_U252 P1_R2278_U128 ; P1_R2278_U353
g28591 nand P1_R2278_U353 P1_R2278_U352 P1_R2278_U137 ; P1_R2278_U354
g28592 nand P1_U2785 P1_R2278_U284 ; P1_R2278_U355
g28593 nand P1_R2278_U284 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2278_U356
g28594 nand P1_R2278_U356 P1_R2278_U63 ; P1_R2278_U357
g28595 nand P1_R2278_U6 P1_R2278_U222 ; P1_R2278_U358
g28596 nand P1_R2278_U293 P1_R2278_U290 ; P1_R2278_U359
g28597 nand P1_R2278_U359 P1_R2278_U292 ; P1_R2278_U360
g28598 nand P1_R2278_U7 P1_R2278_U222 ; P1_R2278_U361
g28599 nand P1_R2278_U12 P1_R2278_U359 ; P1_R2278_U362
g28600 nand P1_R2278_U171 P1_R2278_U216 ; P1_R2278_U363
g28601 nand P1_R2278_U133 P1_R2278_U302 ; P1_R2278_U364
g28602 nand P1_R2278_U8 P1_R2278_U216 ; P1_R2278_U365
g28603 nand P1_R2278_U364 P1_R2278_U303 ; P1_R2278_U366
g28604 nand P1_R2278_U366 P1_R2278_U305 ; P1_R2278_U367
g28605 nand P1_R2278_U367 P1_R2278_U306 ; P1_R2278_U368
g28606 nand P1_R2278_U368 P1_R2278_U308 ; P1_R2278_U369
g28607 nand P1_R2278_U130 P1_R2278_U313 ; P1_R2278_U370
g28608 nand P1_R2278_U381 P1_R2278_U315 ; P1_R2278_U371
g28609 nand P1_R2278_U131 P1_R2278_U371 ; P1_R2278_U372
g28610 nand P1_R2278_U372 P1_R2278_U317 ; P1_R2278_U373
g28611 nand P1_R2278_U372 P1_R2278_U317 ; P1_R2278_U374
g28612 nand P1_R2278_U147 P1_R2278_U194 ; P1_R2278_U375
g28613 nand P1_R2278_U161 P1_R2278_U418 ; P1_R2278_U376
g28614 not P1_R2278_U80 ; P1_R2278_U377
g28615 not P1_R2278_U73 ; P1_R2278_U378
g28616 nand P1_R2278_U320 P1_R2278_U321 ; P1_R2278_U379
g28617 not P1_R2278_U94 ; P1_R2278_U380
g28618 nand P1_R2278_U370 P1_R2278_U314 ; P1_R2278_U381
g28619 nand P1_R2278_U391 P1_R2278_U229 P1_R2278_U285 ; P1_R2278_U382
g28620 not P1_R2278_U92 ; P1_R2278_U383
g28621 not P1_R2278_U95 ; P1_R2278_U384
g28622 nand P1_R2278_U11 P1_R2278_U411 P1_R2278_U142 ; P1_R2278_U385
g28623 not P1_R2278_U93 ; P1_R2278_U386
g28624 not P1_R2278_U96 ; P1_R2278_U387
g28625 nand P1_R2278_U277 P1_R2278_U261 ; P1_R2278_U388
g28626 nand P1_R2278_U388 P1_R2278_U228 ; P1_R2278_U389
g28627 nand P1_R2278_U391 P1_R2278_U229 P1_R2278_U285 ; P1_R2278_U390
g28628 nand P1_R2278_U282 P1_R2278_U283 ; P1_R2278_U391
g28629 not P1_R2278_U86 ; P1_R2278_U392
g28630 nand P1_U2770 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2278_U393
g28631 nand P1_R2278_U148 P1_R2278_U372 ; P1_R2278_U394
g28632 nand P1_R2278_U383 P1_R2278_U324 ; P1_R2278_U395
g28633 nand P1_R2278_U150 P1_R2278_U368 ; P1_R2278_U396
g28634 nand P1_R2278_U152 P1_R2278_U413 P1_R2278_U153 ; P1_R2278_U397
g28635 nand P1_R2278_U386 P1_R2278_U324 ; P1_R2278_U398
g28636 nand P1_R2278_U154 P1_R2278_U11 P1_R2278_U378 ; P1_R2278_U399
g28637 nand P1_R2278_U86 P1_R2278_U324 ; P1_R2278_U400
g28638 not P1_R2278_U87 ; P1_R2278_U401
g28639 nand P1_R2278_U391 P1_R2278_U229 P1_R2278_U285 ; P1_R2278_U402
g28640 nand P1_R2278_U380 P1_R2278_U324 ; P1_R2278_U403
g28641 nand P1_R2278_U384 P1_R2278_U324 ; P1_R2278_U404
g28642 nand P1_R2278_U157 P1_R2278_U411 P1_R2278_U158 ; P1_R2278_U405
g28643 nand P1_R2278_U387 P1_R2278_U324 ; P1_R2278_U406
g28644 nand P1_R2278_U87 P1_R2278_U324 ; P1_R2278_U407
g28645 nand P1_R2278_U374 P1_R2278_U85 ; P1_R2278_U408
g28646 nand P1_R2278_U408 P1_R2278_U319 ; P1_R2278_U409
g28647 nand P1_R2278_U402 P1_R2278_U227 ; P1_R2278_U410
g28648 nand P1_R2278_U141 P1_R2278_U226 ; P1_R2278_U411
g28649 nand P1_R2278_U390 P1_R2278_U227 ; P1_R2278_U412
g28650 nand P1_R2278_U151 P1_R2278_U226 ; P1_R2278_U413
g28651 nand P1_R2278_U174 P1_R2278_U336 ; P1_R2278_U414
g28652 nand P1_R2278_U287 P1_R2278_U227 ; P1_R2278_U415
g28653 not P1_R2278_U222 ; P1_R2278_U416
g28654 nand P1_R2278_U382 P1_R2278_U227 ; P1_R2278_U417
g28655 nand P1_R2278_U160 P1_R2278_U226 ; P1_R2278_U418
g28656 nand P1_R2278_U11 P1_R2278_U206 ; P1_R2278_U419
g28657 not P1_R2278_U196 ; P1_R2278_U420
g28658 nand P1_R2278_U311 P1_R2278_U206 ; P1_R2278_U421
g28659 not P1_R2278_U204 ; P1_R2278_U422
g28660 nand P1_R2278_U10 P1_R2278_U206 ; P1_R2278_U423
g28661 not P1_R2278_U200 ; P1_R2278_U424
g28662 nand P1_R2278_U164 P1_R2278_U206 ; P1_R2278_U425
g28663 not P1_R2278_U198 ; P1_R2278_U426
g28664 nand P1_R2278_U166 P1_R2278_U206 ; P1_R2278_U427
g28665 not P1_R2278_U202 ; P1_R2278_U428
g28666 nand P1_R2278_U557 P1_R2278_U33 ; P1_R2278_U429
g28667 nand P1_R2278_U346 P1_R2278_U176 ; P1_R2278_U430
g28668 nand P1_R2278_U100 P1_R2278_U260 ; P1_R2278_U431
g28669 nand P1_U2792 P1_R2278_U21 ; P1_R2278_U432
g28670 nand P1_R2278_U22 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2278_U433
g28671 nand P1_U2792 P1_R2278_U21 ; P1_R2278_U434
g28672 nand P1_R2278_U22 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_R2278_U435
g28673 nand P1_R2278_U435 P1_R2278_U434 ; P1_R2278_U436
g28674 nand P1_R2278_U177 P1_R2278_U178 ; P1_R2278_U437
g28675 nand P1_R2278_U257 P1_R2278_U436 ; P1_R2278_U438
g28676 nand P1_U2793 P1_R2278_U23 ; P1_R2278_U439
g28677 nand P1_R2278_U24 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_R2278_U440
g28678 nand P1_U2794 P1_R2278_U25 ; P1_R2278_U441
g28679 nand P1_R2278_U26 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_R2278_U442
g28680 nand P1_R2278_U442 P1_R2278_U441 ; P1_R2278_U443
g28681 nand P1_R2278_U347 P1_R2278_U40 ; P1_R2278_U444
g28682 nand P1_R2278_U443 P1_R2278_U251 ; P1_R2278_U445
g28683 nand P1_U2795 P1_R2278_U27 ; P1_R2278_U446
g28684 nand P1_R2278_U28 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_R2278_U447
g28685 nand P1_U2796 P1_R2278_U38 ; P1_R2278_U448
g28686 nand P1_R2278_U39 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2278_U449
g28687 nand P1_U2796 P1_R2278_U38 ; P1_R2278_U450
g28688 nand P1_R2278_U39 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_R2278_U451
g28689 nand P1_R2278_U451 P1_R2278_U450 ; P1_R2278_U452
g28690 nand P1_R2278_U181 P1_R2278_U182 ; P1_R2278_U453
g28691 nand P1_R2278_U243 P1_R2278_U452 ; P1_R2278_U454
g28692 nand P1_U2797 P1_R2278_U36 ; P1_R2278_U455
g28693 nand P1_R2278_U37 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2278_U456
g28694 nand P1_U2797 P1_R2278_U36 ; P1_R2278_U457
g28695 nand P1_R2278_U37 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_R2278_U458
g28696 nand P1_R2278_U458 P1_R2278_U457 ; P1_R2278_U459
g28697 nand P1_R2278_U183 P1_R2278_U184 ; P1_R2278_U460
g28698 nand P1_R2278_U239 P1_R2278_U459 ; P1_R2278_U461
g28699 nand P1_R2278_U186 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_R2278_U462
g28700 nand P1_U2769 P1_R2278_U185 ; P1_R2278_U463
g28701 nand P1_R2278_U186 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_R2278_U464
g28702 nand P1_U2769 P1_R2278_U185 ; P1_R2278_U465
g28703 nand P1_R2278_U465 P1_R2278_U464 ; P1_R2278_U466
g28704 nand P1_R2278_U397 P1_R2278_U396 P1_R2278_U155 P1_R2278_U187 ; P1_R2278_U467
g28705 nand P1_R2278_U325 P1_R2278_U5 ; P1_R2278_U468
g28706 nand P1_R2278_U14 P1_R2278_U88 P1_R2278_U89 ; P1_R2278_U469
g28707 nand P1_U2770 P1_R2278_U466 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2278_U470
g28708 nand P1_R2278_U88 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2278_U471
g28709 nand P1_U2770 P1_R2278_U89 ; P1_R2278_U472
g28710 nand P1_R2278_U88 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_R2278_U473
g28711 nand P1_U2770 P1_R2278_U89 ; P1_R2278_U474
g28712 nand P1_R2278_U474 P1_R2278_U473 ; P1_R2278_U475
g28713 nand P1_R2278_U189 P1_R2278_U190 ; P1_R2278_U476
g28714 nand P1_R2278_U326 P1_R2278_U475 ; P1_R2278_U477
g28715 nand P1_U2798 P1_R2278_U34 ; P1_R2278_U478
g28716 nand P1_R2278_U35 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2278_U479
g28717 nand P1_U2798 P1_R2278_U34 ; P1_R2278_U480
g28718 nand P1_R2278_U35 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_R2278_U481
g28719 nand P1_R2278_U481 P1_R2278_U480 ; P1_R2278_U482
g28720 nand P1_R2278_U191 P1_R2278_U192 ; P1_R2278_U483
g28721 nand P1_R2278_U235 P1_R2278_U482 ; P1_R2278_U484
g28722 nand P1_R2278_U90 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2278_U485
g28723 nand P1_U2771 P1_R2278_U91 ; P1_R2278_U486
g28724 nand P1_R2278_U90 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_R2278_U487
g28725 nand P1_U2771 P1_R2278_U91 ; P1_R2278_U488
g28726 nand P1_R2278_U488 P1_R2278_U487 ; P1_R2278_U489
g28727 nand P1_R2278_U193 P1_R2278_U194 ; P1_R2278_U490
g28728 nand P1_R2278_U323 P1_R2278_U489 ; P1_R2278_U491
g28729 nand P1_R2278_U81 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2278_U492
g28730 nand P1_U2772 P1_R2278_U82 ; P1_R2278_U493
g28731 nand P1_R2278_U81 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_R2278_U494
g28732 nand P1_U2772 P1_R2278_U82 ; P1_R2278_U495
g28733 nand P1_R2278_U495 P1_R2278_U494 ; P1_R2278_U496
g28734 nand P1_R2278_U195 P1_R2278_U196 ; P1_R2278_U497
g28735 nand P1_R2278_U420 P1_R2278_U496 ; P1_R2278_U498
g28736 nand P1_U2773 P1_R2278_U83 ; P1_R2278_U499
g28737 nand P1_R2278_U84 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2278_U500
g28738 nand P1_U2773 P1_R2278_U83 ; P1_R2278_U501
g28739 nand P1_R2278_U84 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_R2278_U502
g28740 nand P1_R2278_U502 P1_R2278_U501 ; P1_R2278_U503
g28741 nand P1_R2278_U197 P1_R2278_U198 ; P1_R2278_U504
g28742 nand P1_R2278_U426 P1_R2278_U503 ; P1_R2278_U505
g28743 nand P1_U2774 P1_R2278_U46 ; P1_R2278_U506
g28744 nand P1_R2278_U47 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2278_U507
g28745 nand P1_U2774 P1_R2278_U46 ; P1_R2278_U508
g28746 nand P1_R2278_U47 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_R2278_U509
g28747 nand P1_R2278_U509 P1_R2278_U508 ; P1_R2278_U510
g28748 nand P1_R2278_U199 P1_R2278_U200 ; P1_R2278_U511
g28749 nand P1_R2278_U424 P1_R2278_U510 ; P1_R2278_U512
g28750 nand P1_U2775 P1_R2278_U44 ; P1_R2278_U513
g28751 nand P1_R2278_U45 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2278_U514
g28752 nand P1_U2775 P1_R2278_U44 ; P1_R2278_U515
g28753 nand P1_R2278_U45 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_R2278_U516
g28754 nand P1_R2278_U516 P1_R2278_U515 ; P1_R2278_U517
g28755 nand P1_R2278_U201 P1_R2278_U202 ; P1_R2278_U518
g28756 nand P1_R2278_U428 P1_R2278_U517 ; P1_R2278_U519
g28757 nand P1_U2776 P1_R2278_U48 ; P1_R2278_U520
g28758 nand P1_R2278_U49 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2278_U521
g28759 nand P1_U2776 P1_R2278_U48 ; P1_R2278_U522
g28760 nand P1_R2278_U49 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_R2278_U523
g28761 nand P1_R2278_U523 P1_R2278_U522 ; P1_R2278_U524
g28762 nand P1_R2278_U203 P1_R2278_U204 ; P1_R2278_U525
g28763 nand P1_R2278_U422 P1_R2278_U524 ; P1_R2278_U526
g28764 nand P1_U2777 P1_R2278_U50 ; P1_R2278_U527
g28765 nand P1_R2278_U51 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2278_U528
g28766 nand P1_U2777 P1_R2278_U50 ; P1_R2278_U529
g28767 nand P1_R2278_U51 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_R2278_U530
g28768 nand P1_R2278_U530 P1_R2278_U529 ; P1_R2278_U531
g28769 nand P1_R2278_U205 P1_R2278_U206 ; P1_R2278_U532
g28770 nand P1_R2278_U310 P1_R2278_U531 ; P1_R2278_U533
g28771 nand P1_U2778 P1_R2278_U74 ; P1_R2278_U534
g28772 nand P1_R2278_U75 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2278_U535
g28773 nand P1_U2778 P1_R2278_U74 ; P1_R2278_U536
g28774 nand P1_R2278_U75 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_R2278_U537
g28775 nand P1_R2278_U537 P1_R2278_U536 ; P1_R2278_U538
g28776 nand P1_R2278_U207 P1_R2278_U208 ; P1_R2278_U539
g28777 nand P1_R2278_U307 P1_R2278_U538 ; P1_R2278_U540
g28778 nand P1_U2779 P1_R2278_U52 ; P1_R2278_U541
g28779 nand P1_R2278_U53 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2278_U542
g28780 nand P1_U2779 P1_R2278_U52 ; P1_R2278_U543
g28781 nand P1_R2278_U53 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_R2278_U544
g28782 nand P1_R2278_U544 P1_R2278_U543 ; P1_R2278_U545
g28783 nand P1_R2278_U209 P1_R2278_U210 ; P1_R2278_U546
g28784 nand P1_R2278_U304 P1_R2278_U545 ; P1_R2278_U547
g28785 nand P1_U2780 P1_R2278_U54 ; P1_R2278_U548
g28786 nand P1_R2278_U55 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2278_U549
g28787 nand P1_U2780 P1_R2278_U54 ; P1_R2278_U550
g28788 nand P1_R2278_U55 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_R2278_U551
g28789 nand P1_R2278_U551 P1_R2278_U550 ; P1_R2278_U552
g28790 nand P1_R2278_U211 P1_R2278_U212 ; P1_R2278_U553
g28791 nand P1_R2278_U301 P1_R2278_U552 ; P1_R2278_U554
g28792 nand P1_R2278_U32 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2278_U555
g28793 nand P1_R2278_U232 P1_R2278_U31 ; P1_R2278_U556
g28794 nand P1_R2278_U556 P1_R2278_U555 ; P1_R2278_U557
g28795 nand P1_U2799 P1_R2278_U32 P1_R2278_U31 ; P1_R2278_U558
g28796 nand P1_R2278_U230 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_R2278_U559
g28797 nand P1_U2781 P1_R2278_U56 ; P1_R2278_U560
g28798 nand P1_R2278_U57 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2278_U561
g28799 nand P1_U2781 P1_R2278_U56 ; P1_R2278_U562
g28800 nand P1_R2278_U57 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_R2278_U563
g28801 nand P1_R2278_U563 P1_R2278_U562 ; P1_R2278_U564
g28802 nand P1_R2278_U215 P1_R2278_U216 ; P1_R2278_U565
g28803 nand P1_R2278_U297 P1_R2278_U564 ; P1_R2278_U566
g28804 nand P1_U2782 P1_R2278_U77 ; P1_R2278_U567
g28805 nand P1_R2278_U78 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2278_U568
g28806 nand P1_U2782 P1_R2278_U77 ; P1_R2278_U569
g28807 nand P1_R2278_U78 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_R2278_U570
g28808 nand P1_R2278_U570 P1_R2278_U569 ; P1_R2278_U571
g28809 nand P1_R2278_U217 P1_R2278_U218 ; P1_R2278_U572
g28810 nand P1_R2278_U294 P1_R2278_U571 ; P1_R2278_U573
g28811 nand P1_U2783 P1_R2278_U71 ; P1_R2278_U574
g28812 nand P1_R2278_U72 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2278_U575
g28813 nand P1_U2783 P1_R2278_U71 ; P1_R2278_U576
g28814 nand P1_R2278_U72 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_R2278_U577
g28815 nand P1_R2278_U577 P1_R2278_U576 ; P1_R2278_U578
g28816 nand P1_R2278_U219 P1_R2278_U220 ; P1_R2278_U579
g28817 nand P1_R2278_U291 P1_R2278_U578 ; P1_R2278_U580
g28818 nand P1_U2784 P1_R2278_U69 ; P1_R2278_U581
g28819 nand P1_R2278_U70 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2278_U582
g28820 nand P1_U2784 P1_R2278_U69 ; P1_R2278_U583
g28821 nand P1_R2278_U70 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_R2278_U584
g28822 nand P1_R2278_U584 P1_R2278_U583 ; P1_R2278_U585
g28823 nand P1_R2278_U221 P1_R2278_U222 ; P1_R2278_U586
g28824 nand P1_R2278_U416 P1_R2278_U585 ; P1_R2278_U587
g28825 nand P1_U2785 P1_R2278_U62 ; P1_R2278_U588
g28826 nand P1_R2278_U63 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_R2278_U589
g28827 nand P1_U2786 P1_R2278_U66 ; P1_R2278_U590
g28828 nand P1_R2278_U67 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_R2278_U591
g28829 nand P1_R2278_U591 P1_R2278_U590 ; P1_R2278_U592
g28830 nand P1_R2278_U348 P1_R2278_U97 ; P1_R2278_U593
g28831 nand P1_R2278_U592 P1_R2278_U332 ; P1_R2278_U594
g28832 nand P1_U2787 P1_R2278_U64 ; P1_R2278_U595
g28833 nand P1_R2278_U65 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_R2278_U596
g28834 nand P1_R2278_U596 P1_R2278_U595 ; P1_R2278_U597
g28835 nand P1_R2278_U349 P1_R2278_U223 ; P1_R2278_U598
g28836 nand P1_R2278_U329 P1_R2278_U597 ; P1_R2278_U599
g28837 nand P1_R2278_U350 P1_R2278_U224 ; P1_R2278_U600
g28838 nand P1_R2278_U124 P1_R2278_U280 ; P1_R2278_U601
g28839 nand P1_U2789 P1_R2278_U58 ; P1_R2278_U602
g28840 nand P1_R2278_U59 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_R2278_U603
g28841 nand P1_U2790 P1_R2278_U60 ; P1_R2278_U604
g28842 nand P1_R2278_U61 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_R2278_U605
g28843 nand P1_R2278_U605 P1_R2278_U604 ; P1_R2278_U606
g28844 nand P1_R2278_U351 P1_R2278_U225 ; P1_R2278_U607
g28845 nand P1_R2278_U275 P1_R2278_U606 ; P1_R2278_U608
g28846 nand P1_R2278_U29 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_R2278_U609
g28847 nand P1_U2800 P1_R2278_U30 ; P1_R2278_U610
g28848 and P1_R2358_U274 P1_R2358_U272 ; P1_R2358_U5
g28849 and P1_R2358_U280 P1_R2358_U278 ; P1_R2358_U6
g28850 and P1_R2358_U6 P1_R2358_U282 ; P1_R2358_U7
g28851 and P1_R2358_U288 P1_R2358_U286 ; P1_R2358_U8
g28852 and P1_R2358_U8 P1_R2358_U290 ; P1_R2358_U9
g28853 and P1_R2358_U9 P1_R2358_U292 ; P1_R2358_U10
g28854 and P1_R2358_U458 P1_R2358_U457 ; P1_R2358_U11
g28855 and P1_R2358_U481 P1_R2358_U480 ; P1_R2358_U12
g28856 and P1_R2358_U555 P1_R2358_U554 ; P1_R2358_U13
g28857 and P1_R2358_U330 P1_R2358_U329 ; P1_R2358_U14
g28858 and P1_R2358_U327 P1_R2358_U325 ; P1_R2358_U15
g28859 and P1_R2358_U320 P1_R2358_U319 ; P1_R2358_U16
g28860 and P1_R2358_U317 P1_R2358_U315 ; P1_R2358_U17
g28861 and P1_R2358_U308 P1_R2358_U307 ; P1_R2358_U18
g28862 and P1_R2358_U254 P1_R2358_U252 ; P1_R2358_U19
g28863 and P1_R2358_U245 P1_R2358_U244 ; P1_R2358_U20
g28864 and P1_R2358_U242 P1_R2358_U240 ; P1_R2358_U21
g28865 and P1_R2358_U566 P1_R2358_U565 P1_R2358_U136 ; P1_R2358_U22
g28866 not P1_U2352 ; P1_R2358_U23
g28867 not P1_U2643 ; P1_R2358_U24
g28868 not P1_U2644 ; P1_R2358_U25
g28869 not P1_U2645 ; P1_R2358_U26
g28870 not P1_U2646 ; P1_R2358_U27
g28871 nand P1_U2646 P1_R2358_U413 ; P1_R2358_U28
g28872 not P1_U2649 ; P1_R2358_U29
g28873 not P1_U2648 ; P1_R2358_U30
g28874 not P1_U2650 ; P1_R2358_U31
g28875 not P1_U2647 ; P1_R2358_U32
g28876 not P1_U2642 ; P1_R2358_U33
g28877 not P1_U2641 ; P1_R2358_U34
g28878 nand P1_R2358_U236 P1_R2358_U220 ; P1_R2358_U35
g28879 nand P1_R2358_U35 P1_R2358_U218 ; P1_R2358_U36
g28880 not P1_U2623 ; P1_R2358_U37
g28881 not P1_U2624 ; P1_R2358_U38
g28882 not P1_U2625 ; P1_R2358_U39
g28883 not P1_U2626 ; P1_R2358_U40
g28884 not P1_U2627 ; P1_R2358_U41
g28885 nand P1_U2627 P1_R2358_U546 ; P1_R2358_U42
g28886 not P1_U2628 ; P1_R2358_U43
g28887 not P1_U2629 ; P1_R2358_U44
g28888 not P1_U2630 ; P1_R2358_U45
g28889 not P1_U2631 ; P1_R2358_U46
g28890 nand P1_U2631 P1_R2358_U521 ; P1_R2358_U47
g28891 not P1_U2632 ; P1_R2358_U48
g28892 not P1_U2633 ; P1_R2358_U49
g28893 not P1_U2634 ; P1_R2358_U50
g28894 nand P1_U2634 P1_R2358_U501 ; P1_R2358_U51
g28895 not P1_U2639 ; P1_R2358_U52
g28896 not P1_U2640 ; P1_R2358_U53
g28897 nand P1_R2358_U400 P1_R2358_U399 P1_R2358_U34 ; P1_R2358_U54
g28898 not P1_U2635 ; P1_R2358_U55
g28899 not P1_U2638 ; P1_R2358_U56
g28900 nand P1_U2638 P1_R2358_U471 ; P1_R2358_U57
g28901 not P1_U2637 ; P1_R2358_U58
g28902 nand P1_U2637 P1_R2358_U463 ; P1_R2358_U59
g28903 not P1_U2636 ; P1_R2358_U60
g28904 nand P1_U2636 P1_R2358_U466 ; P1_R2358_U61
g28905 not P1_U2622 ; P1_R2358_U62
g28906 not P1_U2620 ; P1_R2358_U63
g28907 not P1_U2621 ; P1_R2358_U64
g28908 nand P1_R2358_U206 P1_R2358_U248 ; P1_R2358_U65
g28909 nand P1_R2358_U65 P1_R2358_U202 ; P1_R2358_U66
g28910 nand P1_R2358_U371 P1_R2358_U293 ; P1_R2358_U67
g28911 nand P1_R2358_U369 P1_R2358_U291 ; P1_R2358_U68
g28912 nand P1_R2358_U364 P1_R2358_U283 ; P1_R2358_U69
g28913 nand P1_R2358_U358 P1_R2358_U275 ; P1_R2358_U70
g28914 nand P1_R2358_U59 P1_R2358_U311 ; P1_R2358_U71
g28915 nand P1_R2358_U71 P1_R2358_U255 ; P1_R2358_U72
g28916 nand P1_R2358_U233 P1_R2358_U321 ; P1_R2358_U73
g28917 nand P1_R2358_U73 P1_R2358_U262 ; P1_R2358_U74
g28918 nand P1_R2358_U557 P1_R2358_U556 ; P1_R2358_U75
g28919 nand P1_R2358_U611 P1_R2358_U610 ; P1_R2358_U76
g28920 and P1_R2358_U233 P1_R2358_U54 ; P1_R2358_U77
g28921 nand P1_R2358_U450 P1_R2358_U449 ; P1_R2358_U78
g28922 and P1_R2358_U229 P1_R2358_U228 ; P1_R2358_U79
g28923 nand P1_R2358_U452 P1_R2358_U451 ; P1_R2358_U80
g28924 and P1_R2358_U220 P1_R2358_U219 ; P1_R2358_U81
g28925 nand P1_R2358_U454 P1_R2358_U453 ; P1_R2358_U82
g28926 and P1_R2358_U225 P1_R2358_U28 ; P1_R2358_U83
g28927 nand P1_R2358_U456 P1_R2358_U455 ; P1_R2358_U84
g28928 nand P1_R2358_U575 P1_R2358_U574 ; P1_R2358_U85
g28929 and P1_R2358_U179 P1_R2358_U300 ; P1_R2358_U86
g28930 nand P1_R2358_U577 P1_R2358_U576 ; P1_R2358_U87
g28931 and P1_R2358_U297 P1_R2358_U296 ; P1_R2358_U88
g28932 nand P1_R2358_U579 P1_R2358_U578 ; P1_R2358_U89
g28933 and P1_R2358_U295 P1_R2358_U294 ; P1_R2358_U90
g28934 nand P1_R2358_U581 P1_R2358_U580 ; P1_R2358_U91
g28935 and P1_R2358_U293 P1_R2358_U292 ; P1_R2358_U92
g28936 nand P1_R2358_U583 P1_R2358_U582 ; P1_R2358_U93
g28937 and P1_R2358_U291 P1_R2358_U290 ; P1_R2358_U94
g28938 nand P1_R2358_U585 P1_R2358_U584 ; P1_R2358_U95
g28939 and P1_R2358_U289 P1_R2358_U288 ; P1_R2358_U96
g28940 nand P1_R2358_U587 P1_R2358_U586 ; P1_R2358_U97
g28941 and P1_R2358_U42 P1_R2358_U286 ; P1_R2358_U98
g28942 nand P1_R2358_U589 P1_R2358_U588 ; P1_R2358_U99
g28943 and P1_R2358_U285 P1_R2358_U284 ; P1_R2358_U100
g28944 nand P1_R2358_U591 P1_R2358_U590 ; P1_R2358_U101
g28945 and P1_R2358_U283 P1_R2358_U282 ; P1_R2358_U102
g28946 nand P1_R2358_U593 P1_R2358_U592 ; P1_R2358_U103
g28947 and P1_R2358_U281 P1_R2358_U280 ; P1_R2358_U104
g28948 nand P1_R2358_U595 P1_R2358_U594 ; P1_R2358_U105
g28949 and P1_R2358_U206 P1_R2358_U205 ; P1_R2358_U106
g28950 nand P1_R2358_U597 P1_R2358_U596 ; P1_R2358_U107
g28951 and P1_R2358_U47 P1_R2358_U278 ; P1_R2358_U108
g28952 nand P1_R2358_U599 P1_R2358_U598 ; P1_R2358_U109
g28953 and P1_R2358_U277 P1_R2358_U276 ; P1_R2358_U110
g28954 nand P1_R2358_U601 P1_R2358_U600 ; P1_R2358_U111
g28955 and P1_R2358_U275 P1_R2358_U274 ; P1_R2358_U112
g28956 nand P1_R2358_U603 P1_R2358_U602 ; P1_R2358_U113
g28957 and P1_R2358_U51 P1_R2358_U272 ; P1_R2358_U114
g28958 nand P1_R2358_U605 P1_R2358_U604 ; P1_R2358_U115
g28959 and P1_R2358_U59 P1_R2358_U258 ; P1_R2358_U116
g28960 nand P1_R2358_U607 P1_R2358_U606 ; P1_R2358_U117
g28961 and P1_R2358_U57 P1_R2358_U259 ; P1_R2358_U118
g28962 nand P1_R2358_U609 P1_R2358_U608 ; P1_R2358_U119
g28963 and P1_R2358_U208 P1_R2358_U205 ; P1_R2358_U120
g28964 and P1_R2358_U204 P1_R2358_U202 ; P1_R2358_U121
g28965 and P1_R2358_U217 P1_R2358_U216 ; P1_R2358_U122
g28966 and P1_R2358_U204 P1_R2358_U203 ; P1_R2358_U123
g28967 and P1_R2358_U229 P1_R2358_U54 ; P1_R2358_U124
g28968 and P1_R2358_U265 P1_R2358_U262 ; P1_R2358_U125
g28969 and P1_R2358_U258 P1_R2358_U259 P1_R2358_U255 P1_R2358_U356 ; P1_R2358_U126
g28970 and P1_R2358_U256 P1_R2358_U353 P1_R2358_U355 P1_R2358_U354 ; P1_R2358_U127
g28971 and P1_R2358_U276 P1_R2358_U5 ; P1_R2358_U128
g28972 and P1_R2358_U361 P1_R2358_U277 ; P1_R2358_U129
g28973 and P1_R2358_U7 P1_R2358_U284 ; P1_R2358_U130
g28974 and P1_R2358_U366 P1_R2358_U285 ; P1_R2358_U131
g28975 and P1_R2358_U10 P1_R2358_U294 ; P1_R2358_U132
g28976 and P1_R2358_U373 P1_R2358_U295 ; P1_R2358_U133
g28977 and P1_R2358_U561 P1_R2358_U305 ; P1_R2358_U134
g28978 and P1_R2358_U304 P1_R2358_U13 ; P1_R2358_U135
g28979 and P1_R2358_U180 P1_R2358_U374 ; P1_R2358_U136
g28980 and P1_R2358_U367 P1_R2358_U289 ; P1_R2358_U137
g28981 and P1_R2358_U362 P1_R2358_U281 ; P1_R2358_U138
g28982 and P1_R2358_U257 P1_R2358_U256 ; P1_R2358_U139
g28983 and P1_R2358_U316 P1_R2358_U61 ; P1_R2358_U140
g28984 and P1_R2358_U265 P1_R2358_U264 ; P1_R2358_U141
g28985 and P1_R2358_U326 P1_R2358_U263 ; P1_R2358_U142
g28986 not P1_U2618 ; P1_R2358_U143
g28987 not P1_U2615 ; P1_R2358_U144
g28988 not P1_U2614 ; P1_R2358_U145
g28989 not P1_U2667 ; P1_R2358_U146
g28990 not P1_U2668 ; P1_R2358_U147
g28991 not P1_U2670 ; P1_R2358_U148
g28992 not P1_U2671 ; P1_R2358_U149
g28993 not P1_U2672 ; P1_R2358_U150
g28994 not P1_U2669 ; P1_R2358_U151
g28995 not P1_U2617 ; P1_R2358_U152
g28996 nand P1_R2358_U228 P1_R2358_U230 ; P1_R2358_U153
g28997 nand P1_R2358_U226 P1_R2358_U216 P1_R2358_U224 ; P1_R2358_U154
g28998 nand P1_R2358_U28 P1_R2358_U234 ; P1_R2358_U155
g28999 nand P1_R2358_U203 P1_R2358_U213 ; P1_R2358_U156
g29000 not P1_U2611 ; P1_R2358_U157
g29001 not P1_U2612 ; P1_R2358_U158
g29002 not P1_U2613 ; P1_R2358_U159
g29003 not P1_U2616 ; P1_R2358_U160
g29004 not P1_U2610 ; P1_R2358_U161
g29005 not P1_U2609 ; P1_R2358_U162
g29006 not P1_U2666 ; P1_R2358_U163
g29007 not P1_U2665 ; P1_R2358_U164
g29008 not P1_U2664 ; P1_R2358_U165
g29009 not P1_U2660 ; P1_R2358_U166
g29010 not P1_U2661 ; P1_R2358_U167
g29011 not P1_U2663 ; P1_R2358_U168
g29012 not P1_U2662 ; P1_R2358_U169
g29013 not P1_U2655 ; P1_R2358_U170
g29014 not P1_U2656 ; P1_R2358_U171
g29015 not P1_U2657 ; P1_R2358_U172
g29016 not P1_U2659 ; P1_R2358_U173
g29017 not P1_U2658 ; P1_R2358_U174
g29018 not P1_U2654 ; P1_R2358_U175
g29019 not P1_U2653 ; P1_R2358_U176
g29020 not P1_U2651 ; P1_R2358_U177
g29021 not P1_U2652 ; P1_R2358_U178
g29022 nand P1_U2621 P1_R2358_U564 ; P1_R2358_U179
g29023 and P1_R2358_U568 P1_R2358_U567 ; P1_R2358_U180
g29024 and P1_R2358_U570 P1_R2358_U569 ; P1_R2358_U181
g29025 nand P1_R2358_U179 P1_R2358_U302 ; P1_R2358_U182
g29026 nand P1_R2358_U297 P1_R2358_U298 ; P1_R2358_U183
g29027 nand P1_R2358_U133 P1_R2358_U383 ; P1_R2358_U184
g29028 nand P1_R2358_U372 P1_R2358_U381 ; P1_R2358_U185
g29029 nand P1_R2358_U370 P1_R2358_U379 ; P1_R2358_U186
g29030 nand P1_R2358_U137 P1_R2358_U377 ; P1_R2358_U187
g29031 nand P1_R2358_U375 P1_R2358_U42 ; P1_R2358_U188
g29032 nand P1_R2358_U131 P1_R2358_U385 ; P1_R2358_U189
g29033 nand P1_R2358_U365 P1_R2358_U387 ; P1_R2358_U190
g29034 nand P1_R2358_U138 P1_R2358_U389 ; P1_R2358_U191
g29035 nand P1_R2358_U391 P1_R2358_U47 ; P1_R2358_U192
g29036 nand P1_R2358_U209 P1_R2358_U246 ; P1_R2358_U193
g29037 nand P1_R2358_U129 P1_R2358_U393 ; P1_R2358_U194
g29038 nand P1_R2358_U359 P1_R2358_U395 ; P1_R2358_U195
g29039 nand P1_R2358_U397 P1_R2358_U51 ; P1_R2358_U196
g29040 nand P1_R2358_U201 P1_R2358_U127 ; P1_R2358_U197
g29041 nand P1_R2358_U57 P1_R2358_U309 ; P1_R2358_U198
g29042 nand P1_R2358_U268 P1_R2358_U264 P1_R2358_U267 ; P1_R2358_U199
g29043 nand P1_R2358_U209 P1_R2358_U208 ; P1_R2358_U200
g29044 nand P1_R2358_U126 P1_R2358_U199 ; P1_R2358_U201
g29045 nand P1_R2358_U436 P1_R2358_U435 P1_R2358_U30 ; P1_R2358_U202
g29046 nand P1_U2647 P1_R2358_U441 ; P1_R2358_U203
g29047 nand P1_R2358_U438 P1_R2358_U437 P1_R2358_U32 ; P1_R2358_U204
g29048 nand P1_R2358_U432 P1_R2358_U431 P1_R2358_U29 ; P1_R2358_U205
g29049 nand P1_U2649 P1_R2358_U427 ; P1_R2358_U206
g29050 nand P1_U2648 P1_R2358_U424 ; P1_R2358_U207
g29051 nand P1_R2358_U434 P1_R2358_U433 P1_R2358_U31 ; P1_R2358_U208
g29052 nand P1_U2650 P1_R2358_U430 ; P1_R2358_U209
g29053 nand P1_R2358_U209 P1_R2358_U23 ; P1_R2358_U210
g29054 nand P1_R2358_U120 P1_R2358_U210 ; P1_R2358_U211
g29055 nand P1_R2358_U211 P1_R2358_U206 P1_R2358_U207 ; P1_R2358_U212
g29056 nand P1_R2358_U121 P1_R2358_U212 ; P1_R2358_U213
g29057 not P1_R2358_U156 ; P1_R2358_U214
g29058 nand P1_U2644 P1_R2358_U408 ; P1_R2358_U215
g29059 nand P1_U2643 P1_R2358_U421 ; P1_R2358_U216
g29060 nand P1_R2358_U405 P1_R2358_U404 P1_R2358_U24 ; P1_R2358_U217
g29061 nand P1_R2358_U418 P1_R2358_U417 P1_R2358_U25 ; P1_R2358_U218
g29062 nand P1_R2358_U410 P1_R2358_U409 P1_R2358_U26 ; P1_R2358_U219
g29063 nand P1_U2645 P1_R2358_U416 ; P1_R2358_U220
g29064 not P1_R2358_U28 ; P1_R2358_U221
g29065 nand P1_R2358_U221 P1_R2358_U219 ; P1_R2358_U222
g29066 nand P1_R2358_U220 P1_R2358_U222 P1_R2358_U215 ; P1_R2358_U223
g29067 nand P1_R2358_U218 P1_R2358_U223 P1_R2358_U217 ; P1_R2358_U224
g29068 nand P1_R2358_U443 P1_R2358_U442 P1_R2358_U27 ; P1_R2358_U225
g29069 nand P1_R2358_U225 P1_R2358_U156 P1_R2358_U219 P1_R2358_U218 P1_R2358_U217 ; P1_R2358_U226
g29070 not P1_R2358_U154 ; P1_R2358_U227
g29071 nand P1_U2642 P1_R2358_U448 ; P1_R2358_U228
g29072 nand P1_R2358_U445 P1_R2358_U444 P1_R2358_U33 ; P1_R2358_U229
g29073 nand P1_R2358_U229 P1_R2358_U154 ; P1_R2358_U230
g29074 not P1_R2358_U153 ; P1_R2358_U231
g29075 not P1_R2358_U54 ; P1_R2358_U232
g29076 nand P1_U2641 P1_R2358_U403 ; P1_R2358_U233
g29077 nand P1_R2358_U225 P1_R2358_U156 ; P1_R2358_U234
g29078 not P1_R2358_U155 ; P1_R2358_U235
g29079 nand P1_R2358_U155 P1_R2358_U219 ; P1_R2358_U236
g29080 not P1_R2358_U35 ; P1_R2358_U237
g29081 not P1_R2358_U36 ; P1_R2358_U238
g29082 nand P1_R2358_U36 P1_R2358_U215 ; P1_R2358_U239
g29083 nand P1_R2358_U122 P1_R2358_U239 ; P1_R2358_U240
g29084 nand P1_R2358_U217 P1_R2358_U216 ; P1_R2358_U241
g29085 nand P1_R2358_U36 P1_R2358_U215 P1_R2358_U241 ; P1_R2358_U242
g29086 nand P1_R2358_U218 P1_R2358_U215 ; P1_R2358_U243
g29087 nand P1_R2358_U237 P1_R2358_U243 ; P1_R2358_U244
g29088 nand P1_R2358_U238 P1_R2358_U215 ; P1_R2358_U245
g29089 nand P1_U2352 P1_R2358_U208 ; P1_R2358_U246
g29090 not P1_R2358_U193 ; P1_R2358_U247
g29091 nand P1_R2358_U193 P1_R2358_U205 ; P1_R2358_U248
g29092 not P1_R2358_U65 ; P1_R2358_U249
g29093 not P1_R2358_U66 ; P1_R2358_U250
g29094 nand P1_R2358_U66 P1_R2358_U207 ; P1_R2358_U251
g29095 nand P1_R2358_U123 P1_R2358_U251 ; P1_R2358_U252
g29096 nand P1_R2358_U204 P1_R2358_U203 ; P1_R2358_U253
g29097 nand P1_R2358_U66 P1_R2358_U207 P1_R2358_U253 ; P1_R2358_U254
g29098 nand P1_R2358_U460 P1_R2358_U459 P1_R2358_U60 ; P1_R2358_U255
g29099 nand P1_U2635 P1_R2358_U474 ; P1_R2358_U256
g29100 nand P1_R2358_U11 P1_R2358_U55 ; P1_R2358_U257
g29101 nand P1_R2358_U468 P1_R2358_U467 P1_R2358_U58 ; P1_R2358_U258
g29102 nand P1_R2358_U486 P1_R2358_U485 P1_R2358_U56 ; P1_R2358_U259
g29103 not P1_R2358_U59 ; P1_R2358_U260
g29104 not P1_R2358_U61 ; P1_R2358_U261
g29105 nand P1_R2358_U476 P1_R2358_U475 P1_R2358_U53 ; P1_R2358_U262
g29106 nand P1_U2640 P1_R2358_U479 ; P1_R2358_U263
g29107 nand P1_U2639 P1_R2358_U484 ; P1_R2358_U264
g29108 nand P1_R2358_U12 P1_R2358_U52 ; P1_R2358_U265
g29109 nand P1_R2358_U233 P1_R2358_U228 P1_R2358_U263 ; P1_R2358_U266
g29110 nand P1_R2358_U360 P1_R2358_U357 P1_R2358_U266 P1_R2358_U262 ; P1_R2358_U267
g29111 nand P1_R2358_U124 P1_R2358_U154 P1_R2358_U125 ; P1_R2358_U268
g29112 not P1_R2358_U199 ; P1_R2358_U269
g29113 not P1_R2358_U57 ; P1_R2358_U270
g29114 not P1_R2358_U197 ; P1_R2358_U271
g29115 nand P1_R2358_U488 P1_R2358_U487 P1_R2358_U50 ; P1_R2358_U272
g29116 not P1_R2358_U51 ; P1_R2358_U273
g29117 nand P1_R2358_U490 P1_R2358_U489 P1_R2358_U49 ; P1_R2358_U274
g29118 nand P1_U2633 P1_R2358_U498 ; P1_R2358_U275
g29119 nand P1_R2358_U492 P1_R2358_U491 P1_R2358_U48 ; P1_R2358_U276
g29120 nand P1_U2632 P1_R2358_U495 ; P1_R2358_U277
g29121 nand P1_R2358_U507 P1_R2358_U506 P1_R2358_U46 ; P1_R2358_U278
g29122 not P1_R2358_U47 ; P1_R2358_U279
g29123 nand P1_R2358_U509 P1_R2358_U508 P1_R2358_U45 ; P1_R2358_U280
g29124 nand P1_U2630 P1_R2358_U518 ; P1_R2358_U281
g29125 nand P1_R2358_U505 P1_R2358_U504 P1_R2358_U44 ; P1_R2358_U282
g29126 nand P1_U2629 P1_R2358_U515 ; P1_R2358_U283
g29127 nand P1_R2358_U503 P1_R2358_U502 P1_R2358_U43 ; P1_R2358_U284
g29128 nand P1_U2628 P1_R2358_U512 ; P1_R2358_U285
g29129 nand P1_R2358_U529 P1_R2358_U528 P1_R2358_U41 ; P1_R2358_U286
g29130 not P1_R2358_U42 ; P1_R2358_U287
g29131 nand P1_R2358_U531 P1_R2358_U530 P1_R2358_U40 ; P1_R2358_U288
g29132 nand P1_U2626 P1_R2358_U543 ; P1_R2358_U289
g29133 nand P1_R2358_U527 P1_R2358_U526 P1_R2358_U39 ; P1_R2358_U290
g29134 nand P1_U2625 P1_R2358_U540 ; P1_R2358_U291
g29135 nand P1_R2358_U525 P1_R2358_U524 P1_R2358_U38 ; P1_R2358_U292
g29136 nand P1_U2624 P1_R2358_U537 ; P1_R2358_U293
g29137 nand P1_R2358_U523 P1_R2358_U522 P1_R2358_U37 ; P1_R2358_U294
g29138 nand P1_U2623 P1_R2358_U534 ; P1_R2358_U295
g29139 nand P1_R2358_U548 P1_R2358_U547 P1_R2358_U62 ; P1_R2358_U296
g29140 nand P1_U2622 P1_R2358_U551 ; P1_R2358_U297
g29141 nand P1_R2358_U296 P1_R2358_U184 ; P1_R2358_U298
g29142 not P1_R2358_U183 ; P1_R2358_U299
g29143 nand P1_R2358_U553 P1_R2358_U552 P1_R2358_U64 ; P1_R2358_U300
g29144 not P1_R2358_U179 ; P1_R2358_U301
g29145 nand P1_R2358_U300 P1_R2358_U183 ; P1_R2358_U302
g29146 not P1_R2358_U182 ; P1_R2358_U303
g29147 nand P1_U2620 P1_R2358_U75 ; P1_R2358_U304
g29148 nand P1_R2358_U558 P1_R2358_U63 ; P1_R2358_U305
g29149 nand P1_R2358_U207 P1_R2358_U202 ; P1_R2358_U306
g29150 nand P1_R2358_U249 P1_R2358_U306 ; P1_R2358_U307
g29151 nand P1_R2358_U250 P1_R2358_U207 ; P1_R2358_U308
g29152 nand P1_R2358_U199 P1_R2358_U259 ; P1_R2358_U309
g29153 not P1_R2358_U198 ; P1_R2358_U310
g29154 nand P1_R2358_U198 P1_R2358_U258 ; P1_R2358_U311
g29155 not P1_R2358_U71 ; P1_R2358_U312
g29156 not P1_R2358_U72 ; P1_R2358_U313
g29157 nand P1_R2358_U72 P1_R2358_U61 ; P1_R2358_U314
g29158 nand P1_R2358_U139 P1_R2358_U314 ; P1_R2358_U315
g29159 nand P1_R2358_U257 P1_R2358_U256 ; P1_R2358_U316
g29160 nand P1_R2358_U140 P1_R2358_U72 ; P1_R2358_U317
g29161 nand P1_R2358_U61 P1_R2358_U255 ; P1_R2358_U318
g29162 nand P1_R2358_U312 P1_R2358_U318 ; P1_R2358_U319
g29163 nand P1_R2358_U313 P1_R2358_U61 ; P1_R2358_U320
g29164 nand P1_R2358_U54 P1_R2358_U153 ; P1_R2358_U321
g29165 not P1_R2358_U73 ; P1_R2358_U322
g29166 not P1_R2358_U74 ; P1_R2358_U323
g29167 nand P1_R2358_U74 P1_R2358_U263 ; P1_R2358_U324
g29168 nand P1_R2358_U141 P1_R2358_U324 ; P1_R2358_U325
g29169 nand P1_R2358_U265 P1_R2358_U264 ; P1_R2358_U326
g29170 nand P1_R2358_U142 P1_R2358_U74 ; P1_R2358_U327
g29171 nand P1_R2358_U263 P1_R2358_U262 ; P1_R2358_U328
g29172 nand P1_R2358_U322 P1_R2358_U328 ; P1_R2358_U329
g29173 nand P1_R2358_U323 P1_R2358_U263 ; P1_R2358_U330
g29174 not P1_R2358_U200 ; P1_R2358_U331
g29175 nand P1_R2358_U233 P1_R2358_U54 ; P1_R2358_U332
g29176 nand P1_R2358_U229 P1_R2358_U228 ; P1_R2358_U333
g29177 nand P1_R2358_U220 P1_R2358_U219 ; P1_R2358_U334
g29178 nand P1_R2358_U225 P1_R2358_U28 ; P1_R2358_U335
g29179 nand P1_R2358_U179 P1_R2358_U300 ; P1_R2358_U336
g29180 nand P1_R2358_U297 P1_R2358_U296 ; P1_R2358_U337
g29181 nand P1_R2358_U295 P1_R2358_U294 ; P1_R2358_U338
g29182 nand P1_R2358_U293 P1_R2358_U292 ; P1_R2358_U339
g29183 nand P1_R2358_U291 P1_R2358_U290 ; P1_R2358_U340
g29184 nand P1_R2358_U289 P1_R2358_U288 ; P1_R2358_U341
g29185 nand P1_R2358_U42 P1_R2358_U286 ; P1_R2358_U342
g29186 nand P1_R2358_U285 P1_R2358_U284 ; P1_R2358_U343
g29187 nand P1_R2358_U283 P1_R2358_U282 ; P1_R2358_U344
g29188 nand P1_R2358_U281 P1_R2358_U280 ; P1_R2358_U345
g29189 nand P1_R2358_U206 P1_R2358_U205 ; P1_R2358_U346
g29190 nand P1_R2358_U47 P1_R2358_U278 ; P1_R2358_U347
g29191 nand P1_R2358_U277 P1_R2358_U276 ; P1_R2358_U348
g29192 nand P1_R2358_U275 P1_R2358_U274 ; P1_R2358_U349
g29193 nand P1_R2358_U51 P1_R2358_U272 ; P1_R2358_U350
g29194 nand P1_R2358_U59 P1_R2358_U258 ; P1_R2358_U351
g29195 nand P1_R2358_U57 P1_R2358_U259 ; P1_R2358_U352
g29196 nand P1_R2358_U270 P1_R2358_U258 P1_R2358_U255 P1_R2358_U257 ; P1_R2358_U353
g29197 nand P1_R2358_U260 P1_R2358_U255 P1_R2358_U257 ; P1_R2358_U354
g29198 nand P1_R2358_U261 P1_R2358_U257 ; P1_R2358_U355
g29199 nand P1_R2358_U11 P1_R2358_U55 ; P1_R2358_U356
g29200 nand P1_R2358_U232 P1_R2358_U263 ; P1_R2358_U357
g29201 nand P1_R2358_U273 P1_R2358_U274 ; P1_R2358_U358
g29202 not P1_R2358_U70 ; P1_R2358_U359
g29203 nand P1_R2358_U12 P1_R2358_U52 ; P1_R2358_U360
g29204 nand P1_R2358_U70 P1_R2358_U276 ; P1_R2358_U361
g29205 nand P1_R2358_U279 P1_R2358_U280 ; P1_R2358_U362
g29206 nand P1_R2358_U362 P1_R2358_U281 ; P1_R2358_U363
g29207 nand P1_R2358_U363 P1_R2358_U282 ; P1_R2358_U364
g29208 not P1_R2358_U69 ; P1_R2358_U365
g29209 nand P1_R2358_U69 P1_R2358_U284 ; P1_R2358_U366
g29210 nand P1_R2358_U287 P1_R2358_U288 ; P1_R2358_U367
g29211 nand P1_R2358_U367 P1_R2358_U289 ; P1_R2358_U368
g29212 nand P1_R2358_U368 P1_R2358_U290 ; P1_R2358_U369
g29213 not P1_R2358_U68 ; P1_R2358_U370
g29214 nand P1_R2358_U68 P1_R2358_U292 ; P1_R2358_U371
g29215 not P1_R2358_U67 ; P1_R2358_U372
g29216 nand P1_R2358_U67 P1_R2358_U294 ; P1_R2358_U373
g29217 nand P1_R2358_U300 P1_R2358_U183 P1_R2358_U134 ; P1_R2358_U374
g29218 nand P1_R2358_U286 P1_R2358_U189 ; P1_R2358_U375
g29219 not P1_R2358_U188 ; P1_R2358_U376
g29220 nand P1_R2358_U8 P1_R2358_U189 ; P1_R2358_U377
g29221 not P1_R2358_U187 ; P1_R2358_U378
g29222 nand P1_R2358_U9 P1_R2358_U189 ; P1_R2358_U379
g29223 not P1_R2358_U186 ; P1_R2358_U380
g29224 nand P1_R2358_U10 P1_R2358_U189 ; P1_R2358_U381
g29225 not P1_R2358_U185 ; P1_R2358_U382
g29226 nand P1_R2358_U132 P1_R2358_U189 ; P1_R2358_U383
g29227 not P1_R2358_U184 ; P1_R2358_U384
g29228 nand P1_R2358_U130 P1_R2358_U194 ; P1_R2358_U385
g29229 not P1_R2358_U189 ; P1_R2358_U386
g29230 nand P1_R2358_U7 P1_R2358_U194 ; P1_R2358_U387
g29231 not P1_R2358_U190 ; P1_R2358_U388
g29232 nand P1_R2358_U6 P1_R2358_U194 ; P1_R2358_U389
g29233 not P1_R2358_U191 ; P1_R2358_U390
g29234 nand P1_R2358_U278 P1_R2358_U194 ; P1_R2358_U391
g29235 not P1_R2358_U192 ; P1_R2358_U392
g29236 nand P1_R2358_U128 P1_R2358_U197 ; P1_R2358_U393
g29237 not P1_R2358_U194 ; P1_R2358_U394
g29238 nand P1_R2358_U5 P1_R2358_U197 ; P1_R2358_U395
g29239 not P1_R2358_U195 ; P1_R2358_U396
g29240 nand P1_R2358_U272 P1_R2358_U197 ; P1_R2358_U397
g29241 not P1_R2358_U196 ; P1_R2358_U398
g29242 nand P1_U2352 P1_R2358_U143 ; P1_R2358_U399
g29243 nand P1_U2618 P1_R2358_U23 ; P1_R2358_U400
g29244 nand P1_U2352 P1_R2358_U143 ; P1_R2358_U401
g29245 nand P1_U2618 P1_R2358_U23 ; P1_R2358_U402
g29246 nand P1_R2358_U402 P1_R2358_U401 ; P1_R2358_U403
g29247 nand P1_U2352 P1_R2358_U144 ; P1_R2358_U404
g29248 nand P1_U2615 P1_R2358_U23 ; P1_R2358_U405
g29249 nand P1_U2352 P1_R2358_U145 ; P1_R2358_U406
g29250 nand P1_U2614 P1_R2358_U23 ; P1_R2358_U407
g29251 nand P1_R2358_U407 P1_R2358_U406 ; P1_R2358_U408
g29252 nand P1_U2352 P1_R2358_U146 ; P1_R2358_U409
g29253 nand P1_U2667 P1_R2358_U23 ; P1_R2358_U410
g29254 nand P1_U2352 P1_R2358_U147 ; P1_R2358_U411
g29255 nand P1_U2668 P1_R2358_U23 ; P1_R2358_U412
g29256 nand P1_R2358_U412 P1_R2358_U411 ; P1_R2358_U413
g29257 nand P1_U2352 P1_R2358_U146 ; P1_R2358_U414
g29258 nand P1_U2667 P1_R2358_U23 ; P1_R2358_U415
g29259 nand P1_R2358_U415 P1_R2358_U414 ; P1_R2358_U416
g29260 nand P1_U2352 P1_R2358_U145 ; P1_R2358_U417
g29261 nand P1_U2614 P1_R2358_U23 ; P1_R2358_U418
g29262 nand P1_U2352 P1_R2358_U144 ; P1_R2358_U419
g29263 nand P1_U2615 P1_R2358_U23 ; P1_R2358_U420
g29264 nand P1_R2358_U420 P1_R2358_U419 ; P1_R2358_U421
g29265 nand P1_U2352 P1_R2358_U148 ; P1_R2358_U422
g29266 nand P1_U2670 P1_R2358_U23 ; P1_R2358_U423
g29267 nand P1_R2358_U423 P1_R2358_U422 ; P1_R2358_U424
g29268 nand P1_U2352 P1_R2358_U149 ; P1_R2358_U425
g29269 nand P1_U2671 P1_R2358_U23 ; P1_R2358_U426
g29270 nand P1_R2358_U426 P1_R2358_U425 ; P1_R2358_U427
g29271 nand P1_U2352 P1_R2358_U150 ; P1_R2358_U428
g29272 nand P1_U2672 P1_R2358_U23 ; P1_R2358_U429
g29273 nand P1_R2358_U429 P1_R2358_U428 ; P1_R2358_U430
g29274 nand P1_U2352 P1_R2358_U149 ; P1_R2358_U431
g29275 nand P1_U2671 P1_R2358_U23 ; P1_R2358_U432
g29276 nand P1_U2352 P1_R2358_U150 ; P1_R2358_U433
g29277 nand P1_U2672 P1_R2358_U23 ; P1_R2358_U434
g29278 nand P1_U2352 P1_R2358_U148 ; P1_R2358_U435
g29279 nand P1_U2670 P1_R2358_U23 ; P1_R2358_U436
g29280 nand P1_U2352 P1_R2358_U151 ; P1_R2358_U437
g29281 nand P1_U2669 P1_R2358_U23 ; P1_R2358_U438
g29282 nand P1_U2352 P1_R2358_U151 ; P1_R2358_U439
g29283 nand P1_U2669 P1_R2358_U23 ; P1_R2358_U440
g29284 nand P1_R2358_U440 P1_R2358_U439 ; P1_R2358_U441
g29285 nand P1_U2352 P1_R2358_U147 ; P1_R2358_U442
g29286 nand P1_U2668 P1_R2358_U23 ; P1_R2358_U443
g29287 nand P1_U2352 P1_R2358_U152 ; P1_R2358_U444
g29288 nand P1_U2617 P1_R2358_U23 ; P1_R2358_U445
g29289 nand P1_U2352 P1_R2358_U152 ; P1_R2358_U446
g29290 nand P1_U2617 P1_R2358_U23 ; P1_R2358_U447
g29291 nand P1_R2358_U447 P1_R2358_U446 ; P1_R2358_U448
g29292 nand P1_R2358_U332 P1_R2358_U153 ; P1_R2358_U449
g29293 nand P1_R2358_U77 P1_R2358_U231 ; P1_R2358_U450
g29294 nand P1_R2358_U333 P1_R2358_U154 ; P1_R2358_U451
g29295 nand P1_R2358_U79 P1_R2358_U227 ; P1_R2358_U452
g29296 nand P1_R2358_U334 P1_R2358_U155 ; P1_R2358_U453
g29297 nand P1_R2358_U81 P1_R2358_U235 ; P1_R2358_U454
g29298 nand P1_R2358_U335 P1_R2358_U156 ; P1_R2358_U455
g29299 nand P1_R2358_U83 P1_R2358_U214 ; P1_R2358_U456
g29300 nand P1_U2352 P1_R2358_U157 ; P1_R2358_U457
g29301 nand P1_U2611 P1_R2358_U23 ; P1_R2358_U458
g29302 nand P1_U2352 P1_R2358_U158 ; P1_R2358_U459
g29303 nand P1_U2612 P1_R2358_U23 ; P1_R2358_U460
g29304 nand P1_U2352 P1_R2358_U159 ; P1_R2358_U461
g29305 nand P1_U2613 P1_R2358_U23 ; P1_R2358_U462
g29306 nand P1_R2358_U462 P1_R2358_U461 ; P1_R2358_U463
g29307 nand P1_U2352 P1_R2358_U158 ; P1_R2358_U464
g29308 nand P1_U2612 P1_R2358_U23 ; P1_R2358_U465
g29309 nand P1_R2358_U465 P1_R2358_U464 ; P1_R2358_U466
g29310 nand P1_U2352 P1_R2358_U159 ; P1_R2358_U467
g29311 nand P1_U2613 P1_R2358_U23 ; P1_R2358_U468
g29312 nand P1_U2352 P1_R2358_U160 ; P1_R2358_U469
g29313 nand P1_U2616 P1_R2358_U23 ; P1_R2358_U470
g29314 nand P1_R2358_U470 P1_R2358_U469 ; P1_R2358_U471
g29315 nand P1_U2352 P1_R2358_U157 ; P1_R2358_U472
g29316 nand P1_U2611 P1_R2358_U23 ; P1_R2358_U473
g29317 nand P1_R2358_U473 P1_R2358_U472 ; P1_R2358_U474
g29318 nand P1_U2352 P1_R2358_U161 ; P1_R2358_U475
g29319 nand P1_U2610 P1_R2358_U23 ; P1_R2358_U476
g29320 nand P1_U2352 P1_R2358_U161 ; P1_R2358_U477
g29321 nand P1_U2610 P1_R2358_U23 ; P1_R2358_U478
g29322 nand P1_R2358_U478 P1_R2358_U477 ; P1_R2358_U479
g29323 nand P1_U2352 P1_R2358_U162 ; P1_R2358_U480
g29324 nand P1_U2609 P1_R2358_U23 ; P1_R2358_U481
g29325 nand P1_U2352 P1_R2358_U162 ; P1_R2358_U482
g29326 nand P1_U2609 P1_R2358_U23 ; P1_R2358_U483
g29327 nand P1_R2358_U483 P1_R2358_U482 ; P1_R2358_U484
g29328 nand P1_U2352 P1_R2358_U160 ; P1_R2358_U485
g29329 nand P1_U2616 P1_R2358_U23 ; P1_R2358_U486
g29330 nand P1_U2352 P1_R2358_U163 ; P1_R2358_U487
g29331 nand P1_U2666 P1_R2358_U23 ; P1_R2358_U488
g29332 nand P1_U2352 P1_R2358_U164 ; P1_R2358_U489
g29333 nand P1_U2665 P1_R2358_U23 ; P1_R2358_U490
g29334 nand P1_U2352 P1_R2358_U165 ; P1_R2358_U491
g29335 nand P1_U2664 P1_R2358_U23 ; P1_R2358_U492
g29336 nand P1_U2352 P1_R2358_U165 ; P1_R2358_U493
g29337 nand P1_U2664 P1_R2358_U23 ; P1_R2358_U494
g29338 nand P1_R2358_U494 P1_R2358_U493 ; P1_R2358_U495
g29339 nand P1_U2352 P1_R2358_U164 ; P1_R2358_U496
g29340 nand P1_U2665 P1_R2358_U23 ; P1_R2358_U497
g29341 nand P1_R2358_U497 P1_R2358_U496 ; P1_R2358_U498
g29342 nand P1_U2352 P1_R2358_U163 ; P1_R2358_U499
g29343 nand P1_U2666 P1_R2358_U23 ; P1_R2358_U500
g29344 nand P1_R2358_U500 P1_R2358_U499 ; P1_R2358_U501
g29345 nand P1_U2352 P1_R2358_U166 ; P1_R2358_U502
g29346 nand P1_U2660 P1_R2358_U23 ; P1_R2358_U503
g29347 nand P1_U2352 P1_R2358_U167 ; P1_R2358_U504
g29348 nand P1_U2661 P1_R2358_U23 ; P1_R2358_U505
g29349 nand P1_U2352 P1_R2358_U168 ; P1_R2358_U506
g29350 nand P1_U2663 P1_R2358_U23 ; P1_R2358_U507
g29351 nand P1_U2352 P1_R2358_U169 ; P1_R2358_U508
g29352 nand P1_U2662 P1_R2358_U23 ; P1_R2358_U509
g29353 nand P1_U2352 P1_R2358_U166 ; P1_R2358_U510
g29354 nand P1_U2660 P1_R2358_U23 ; P1_R2358_U511
g29355 nand P1_R2358_U511 P1_R2358_U510 ; P1_R2358_U512
g29356 nand P1_U2352 P1_R2358_U167 ; P1_R2358_U513
g29357 nand P1_U2661 P1_R2358_U23 ; P1_R2358_U514
g29358 nand P1_R2358_U514 P1_R2358_U513 ; P1_R2358_U515
g29359 nand P1_U2352 P1_R2358_U169 ; P1_R2358_U516
g29360 nand P1_U2662 P1_R2358_U23 ; P1_R2358_U517
g29361 nand P1_R2358_U517 P1_R2358_U516 ; P1_R2358_U518
g29362 nand P1_U2352 P1_R2358_U168 ; P1_R2358_U519
g29363 nand P1_U2663 P1_R2358_U23 ; P1_R2358_U520
g29364 nand P1_R2358_U520 P1_R2358_U519 ; P1_R2358_U521
g29365 nand P1_U2352 P1_R2358_U170 ; P1_R2358_U522
g29366 nand P1_U2655 P1_R2358_U23 ; P1_R2358_U523
g29367 nand P1_U2352 P1_R2358_U171 ; P1_R2358_U524
g29368 nand P1_U2656 P1_R2358_U23 ; P1_R2358_U525
g29369 nand P1_U2352 P1_R2358_U172 ; P1_R2358_U526
g29370 nand P1_U2657 P1_R2358_U23 ; P1_R2358_U527
g29371 nand P1_U2352 P1_R2358_U173 ; P1_R2358_U528
g29372 nand P1_U2659 P1_R2358_U23 ; P1_R2358_U529
g29373 nand P1_U2352 P1_R2358_U174 ; P1_R2358_U530
g29374 nand P1_U2658 P1_R2358_U23 ; P1_R2358_U531
g29375 nand P1_U2352 P1_R2358_U170 ; P1_R2358_U532
g29376 nand P1_U2655 P1_R2358_U23 ; P1_R2358_U533
g29377 nand P1_R2358_U533 P1_R2358_U532 ; P1_R2358_U534
g29378 nand P1_U2352 P1_R2358_U171 ; P1_R2358_U535
g29379 nand P1_U2656 P1_R2358_U23 ; P1_R2358_U536
g29380 nand P1_R2358_U536 P1_R2358_U535 ; P1_R2358_U537
g29381 nand P1_U2352 P1_R2358_U172 ; P1_R2358_U538
g29382 nand P1_U2657 P1_R2358_U23 ; P1_R2358_U539
g29383 nand P1_R2358_U539 P1_R2358_U538 ; P1_R2358_U540
g29384 nand P1_U2352 P1_R2358_U174 ; P1_R2358_U541
g29385 nand P1_U2658 P1_R2358_U23 ; P1_R2358_U542
g29386 nand P1_R2358_U542 P1_R2358_U541 ; P1_R2358_U543
g29387 nand P1_U2352 P1_R2358_U173 ; P1_R2358_U544
g29388 nand P1_U2659 P1_R2358_U23 ; P1_R2358_U545
g29389 nand P1_R2358_U545 P1_R2358_U544 ; P1_R2358_U546
g29390 nand P1_U2352 P1_R2358_U175 ; P1_R2358_U547
g29391 nand P1_U2654 P1_R2358_U23 ; P1_R2358_U548
g29392 nand P1_U2352 P1_R2358_U175 ; P1_R2358_U549
g29393 nand P1_U2654 P1_R2358_U23 ; P1_R2358_U550
g29394 nand P1_R2358_U550 P1_R2358_U549 ; P1_R2358_U551
g29395 nand P1_U2352 P1_R2358_U176 ; P1_R2358_U552
g29396 nand P1_U2653 P1_R2358_U23 ; P1_R2358_U553
g29397 nand P1_U2352 P1_R2358_U177 ; P1_R2358_U554
g29398 nand P1_U2651 P1_R2358_U23 ; P1_R2358_U555
g29399 nand P1_U2352 P1_R2358_U178 ; P1_R2358_U556
g29400 nand P1_U2652 P1_R2358_U23 ; P1_R2358_U557
g29401 not P1_R2358_U75 ; P1_R2358_U558
g29402 nand P1_U2352 P1_R2358_U177 ; P1_R2358_U559
g29403 nand P1_U2651 P1_R2358_U23 ; P1_R2358_U560
g29404 nand P1_R2358_U560 P1_R2358_U559 ; P1_R2358_U561
g29405 nand P1_U2352 P1_R2358_U176 ; P1_R2358_U562
g29406 nand P1_U2653 P1_R2358_U23 ; P1_R2358_U563
g29407 nand P1_R2358_U563 P1_R2358_U562 ; P1_R2358_U564
g29408 nand P1_R2358_U135 P1_R2358_U302 P1_R2358_U179 ; P1_R2358_U565
g29409 nand P1_R2358_U561 P1_R2358_U305 P1_R2358_U301 ; P1_R2358_U566
g29410 nand P1_R2358_U13 P1_R2358_U558 P1_R2358_U63 ; P1_R2358_U567
g29411 nand P1_R2358_U561 P1_R2358_U75 P1_U2620 ; P1_R2358_U568
g29412 nand P1_R2358_U558 P1_U2620 ; P1_R2358_U569
g29413 nand P1_R2358_U75 P1_R2358_U63 ; P1_R2358_U570
g29414 nand P1_R2358_U558 P1_U2620 ; P1_R2358_U571
g29415 nand P1_R2358_U75 P1_R2358_U63 ; P1_R2358_U572
g29416 nand P1_R2358_U572 P1_R2358_U571 ; P1_R2358_U573
g29417 nand P1_R2358_U181 P1_R2358_U182 ; P1_R2358_U574
g29418 nand P1_R2358_U303 P1_R2358_U573 ; P1_R2358_U575
g29419 nand P1_R2358_U336 P1_R2358_U183 ; P1_R2358_U576
g29420 nand P1_R2358_U86 P1_R2358_U299 ; P1_R2358_U577
g29421 nand P1_R2358_U184 P1_R2358_U337 ; P1_R2358_U578
g29422 nand P1_R2358_U88 P1_R2358_U384 ; P1_R2358_U579
g29423 nand P1_R2358_U185 P1_R2358_U338 ; P1_R2358_U580
g29424 nand P1_R2358_U90 P1_R2358_U382 ; P1_R2358_U581
g29425 nand P1_R2358_U186 P1_R2358_U339 ; P1_R2358_U582
g29426 nand P1_R2358_U92 P1_R2358_U380 ; P1_R2358_U583
g29427 nand P1_R2358_U187 P1_R2358_U340 ; P1_R2358_U584
g29428 nand P1_R2358_U94 P1_R2358_U378 ; P1_R2358_U585
g29429 nand P1_R2358_U188 P1_R2358_U341 ; P1_R2358_U586
g29430 nand P1_R2358_U96 P1_R2358_U376 ; P1_R2358_U587
g29431 nand P1_R2358_U189 P1_R2358_U342 ; P1_R2358_U588
g29432 nand P1_R2358_U98 P1_R2358_U386 ; P1_R2358_U589
g29433 nand P1_R2358_U190 P1_R2358_U343 ; P1_R2358_U590
g29434 nand P1_R2358_U100 P1_R2358_U388 ; P1_R2358_U591
g29435 nand P1_R2358_U191 P1_R2358_U344 ; P1_R2358_U592
g29436 nand P1_R2358_U102 P1_R2358_U390 ; P1_R2358_U593
g29437 nand P1_R2358_U192 P1_R2358_U345 ; P1_R2358_U594
g29438 nand P1_R2358_U104 P1_R2358_U392 ; P1_R2358_U595
g29439 nand P1_R2358_U346 P1_R2358_U193 ; P1_R2358_U596
g29440 nand P1_R2358_U106 P1_R2358_U247 ; P1_R2358_U597
g29441 nand P1_R2358_U194 P1_R2358_U347 ; P1_R2358_U598
g29442 nand P1_R2358_U108 P1_R2358_U394 ; P1_R2358_U599
g29443 nand P1_R2358_U195 P1_R2358_U348 ; P1_R2358_U600
g29444 nand P1_R2358_U110 P1_R2358_U396 ; P1_R2358_U601
g29445 nand P1_R2358_U196 P1_R2358_U349 ; P1_R2358_U602
g29446 nand P1_R2358_U112 P1_R2358_U398 ; P1_R2358_U603
g29447 nand P1_R2358_U350 P1_R2358_U197 ; P1_R2358_U604
g29448 nand P1_R2358_U114 P1_R2358_U271 ; P1_R2358_U605
g29449 nand P1_R2358_U351 P1_R2358_U198 ; P1_R2358_U606
g29450 nand P1_R2358_U116 P1_R2358_U310 ; P1_R2358_U607
g29451 nand P1_R2358_U352 P1_R2358_U199 ; P1_R2358_U608
g29452 nand P1_R2358_U118 P1_R2358_U269 ; P1_R2358_U609
g29453 nand P1_U2352 P1_R2358_U200 ; P1_R2358_U610
g29454 nand P1_R2358_U331 P1_R2358_U23 ; P1_R2358_U611
g29455 or P1_LT_589_U8 P1_U2673 ; P1_LT_589_U6
g29456 and P1_R584_U7 P1_R584_U6 ; P1_LT_589_U7
g29457 nor P1_LT_589_U7 P1_R584_U9 P1_R584_U8 ; P1_LT_589_U8
g29458 not P1_U2676 ; P1_R584_U6
g29459 not P1_U2677 ; P1_R584_U7
g29460 not P1_U2674 ; P1_R584_U8
g29461 not P1_U2675 ; P1_R584_U9
g29462 not P1_U4190 ; P1_R2099_U4
g29463 not P1_U4189 ; P1_R2099_U5
g29464 not P1_U2678 ; P1_R2099_U6
g29465 nand P1_R2099_U88 P1_R2099_U137 ; P1_R2099_U7
g29466 nand P1_R2099_U89 P1_R2099_U155 ; P1_R2099_U8
g29467 nand P1_R2099_U90 P1_R2099_U157 ; P1_R2099_U9
g29468 nand P1_R2099_U91 P1_R2099_U159 ; P1_R2099_U10
g29469 nand P1_R2099_U92 P1_R2099_U161 ; P1_R2099_U11
g29470 nand P1_R2099_U93 P1_R2099_U163 ; P1_R2099_U12
g29471 nand P1_R2099_U94 P1_R2099_U165 ; P1_R2099_U13
g29472 nand P1_R2099_U95 P1_R2099_U167 ; P1_R2099_U14
g29473 nand P1_R2099_U169 P1_R2099_U55 ; P1_R2099_U15
g29474 nand P1_R2099_U170 P1_R2099_U54 ; P1_R2099_U16
g29475 nand P1_R2099_U171 P1_R2099_U53 ; P1_R2099_U17
g29476 nand P1_R2099_U172 P1_R2099_U52 ; P1_R2099_U18
g29477 nand P1_R2099_U173 P1_R2099_U51 ; P1_R2099_U19
g29478 nand P1_R2099_U174 P1_R2099_U50 ; P1_R2099_U20
g29479 nand P1_R2099_U175 P1_R2099_U49 ; P1_R2099_U21
g29480 nand P1_R2099_U176 P1_R2099_U48 ; P1_R2099_U22
g29481 nand P1_R2099_U177 P1_R2099_U47 ; P1_R2099_U23
g29482 nand P1_R2099_U178 P1_R2099_U46 ; P1_R2099_U24
g29483 nand P1_R2099_U179 P1_R2099_U45 ; P1_R2099_U25
g29484 nand P1_R2099_U210 P1_R2099_U209 ; P1_R2099_U26
g29485 nand P1_R2099_U183 P1_R2099_U182 ; P1_R2099_U27
g29486 nand P1_R2099_U204 P1_R2099_U203 ; P1_R2099_U28
g29487 nand P1_R2099_U207 P1_R2099_U206 ; P1_R2099_U29
g29488 nand P1_R2099_U198 P1_R2099_U197 ; P1_R2099_U30
g29489 nand P1_R2099_U201 P1_R2099_U200 ; P1_R2099_U31
g29490 nand P1_R2099_U186 P1_R2099_U185 ; P1_R2099_U32
g29491 nand P1_R2099_U189 P1_R2099_U188 ; P1_R2099_U33
g29492 nand P1_R2099_U195 P1_R2099_U194 ; P1_R2099_U34
g29493 nand P1_R2099_U192 P1_R2099_U191 ; P1_R2099_U35
g29494 nand P1_R2099_U213 P1_R2099_U212 ; P1_R2099_U36
g29495 nand P1_R2099_U215 P1_R2099_U214 ; P1_R2099_U37
g29496 nand P1_R2099_U217 P1_R2099_U216 ; P1_R2099_U38
g29497 nand P1_R2099_U219 P1_R2099_U218 ; P1_R2099_U39
g29498 nand P1_R2099_U221 P1_R2099_U220 ; P1_R2099_U40
g29499 nand P1_R2099_U223 P1_R2099_U222 ; P1_R2099_U41
g29500 nand P1_R2099_U225 P1_R2099_U224 ; P1_R2099_U42
g29501 nand P1_R2099_U284 P1_R2099_U283 ; P1_R2099_U43
g29502 nand P1_R2099_U287 P1_R2099_U286 ; P1_R2099_U44
g29503 nand P1_R2099_U227 P1_R2099_U226 ; P1_R2099_U45
g29504 nand P1_R2099_U230 P1_R2099_U229 ; P1_R2099_U46
g29505 nand P1_R2099_U233 P1_R2099_U232 ; P1_R2099_U47
g29506 nand P1_R2099_U236 P1_R2099_U235 ; P1_R2099_U48
g29507 nand P1_R2099_U239 P1_R2099_U238 ; P1_R2099_U49
g29508 nand P1_R2099_U242 P1_R2099_U241 ; P1_R2099_U50
g29509 nand P1_R2099_U245 P1_R2099_U244 ; P1_R2099_U51
g29510 nand P1_R2099_U248 P1_R2099_U247 ; P1_R2099_U52
g29511 nand P1_R2099_U251 P1_R2099_U250 ; P1_R2099_U53
g29512 nand P1_R2099_U254 P1_R2099_U253 ; P1_R2099_U54
g29513 nand P1_R2099_U257 P1_R2099_U256 ; P1_R2099_U55
g29514 nand P1_R2099_U278 P1_R2099_U277 ; P1_R2099_U56
g29515 nand P1_R2099_U281 P1_R2099_U280 ; P1_R2099_U57
g29516 nand P1_R2099_U272 P1_R2099_U271 ; P1_R2099_U58
g29517 nand P1_R2099_U275 P1_R2099_U274 ; P1_R2099_U59
g29518 nand P1_R2099_U266 P1_R2099_U265 ; P1_R2099_U60
g29519 nand P1_R2099_U269 P1_R2099_U268 ; P1_R2099_U61
g29520 nand P1_R2099_U260 P1_R2099_U259 ; P1_R2099_U62
g29521 nand P1_R2099_U263 P1_R2099_U262 ; P1_R2099_U63
g29522 nand P1_R2099_U293 P1_R2099_U292 ; P1_R2099_U64
g29523 nand P1_R2099_U295 P1_R2099_U294 ; P1_R2099_U65
g29524 nand P1_R2099_U299 P1_R2099_U298 ; P1_R2099_U66
g29525 nand P1_R2099_U301 P1_R2099_U300 ; P1_R2099_U67
g29526 nand P1_R2099_U303 P1_R2099_U302 ; P1_R2099_U68
g29527 nand P1_R2099_U305 P1_R2099_U304 ; P1_R2099_U69
g29528 nand P1_R2099_U307 P1_R2099_U306 ; P1_R2099_U70
g29529 nand P1_R2099_U309 P1_R2099_U308 ; P1_R2099_U71
g29530 nand P1_R2099_U311 P1_R2099_U310 ; P1_R2099_U72
g29531 nand P1_R2099_U313 P1_R2099_U312 ; P1_R2099_U73
g29532 nand P1_R2099_U315 P1_R2099_U314 ; P1_R2099_U74
g29533 nand P1_R2099_U317 P1_R2099_U316 ; P1_R2099_U75
g29534 nand P1_R2099_U326 P1_R2099_U325 ; P1_R2099_U76
g29535 nand P1_R2099_U328 P1_R2099_U327 ; P1_R2099_U77
g29536 nand P1_R2099_U330 P1_R2099_U329 ; P1_R2099_U78
g29537 nand P1_R2099_U332 P1_R2099_U331 ; P1_R2099_U79
g29538 nand P1_R2099_U334 P1_R2099_U333 ; P1_R2099_U80
g29539 nand P1_R2099_U336 P1_R2099_U335 ; P1_R2099_U81
g29540 nand P1_R2099_U338 P1_R2099_U337 ; P1_R2099_U82
g29541 nand P1_R2099_U340 P1_R2099_U339 ; P1_R2099_U83
g29542 nand P1_R2099_U342 P1_R2099_U341 ; P1_R2099_U84
g29543 nand P1_R2099_U344 P1_R2099_U343 ; P1_R2099_U85
g29544 nand P1_R2099_U349 P1_R2099_U348 ; P1_R2099_U86
g29545 nand P1_R2099_U324 P1_R2099_U323 ; P1_R2099_U87
g29546 and P1_R2099_U34 P1_R2099_U35 ; P1_R2099_U88
g29547 and P1_R2099_U31 P1_R2099_U30 ; P1_R2099_U89
g29548 and P1_R2099_U29 P1_R2099_U28 ; P1_R2099_U90
g29549 and P1_R2099_U26 P1_R2099_U27 ; P1_R2099_U91
g29550 and P1_R2099_U63 P1_R2099_U62 ; P1_R2099_U92
g29551 and P1_R2099_U61 P1_R2099_U60 ; P1_R2099_U93
g29552 and P1_R2099_U59 P1_R2099_U58 ; P1_R2099_U94
g29553 and P1_R2099_U57 P1_R2099_U56 ; P1_R2099_U95
g29554 and P1_R2099_U44 P1_R2099_U43 ; P1_R2099_U96
g29555 nand P1_R2099_U290 P1_R2099_U289 ; P1_R2099_U97
g29556 nand P1_R2099_U346 P1_R2099_U345 ; P1_R2099_U98
g29557 not P1_U2702 ; P1_R2099_U99
g29558 not P1_U2710 ; P1_R2099_U100
g29559 not P1_U2709 ; P1_R2099_U101
g29560 not P1_U2708 ; P1_R2099_U102
g29561 not P1_U2707 ; P1_R2099_U103
g29562 not P1_U2706 ; P1_R2099_U104
g29563 not P1_U2705 ; P1_R2099_U105
g29564 not P1_U2704 ; P1_R2099_U106
g29565 not P1_U2703 ; P1_R2099_U107
g29566 not P1_U2701 ; P1_R2099_U108
g29567 nand P1_R2099_U159 P1_R2099_U27 ; P1_R2099_U109
g29568 nand P1_R2099_U157 P1_R2099_U28 ; P1_R2099_U110
g29569 nand P1_R2099_U155 P1_R2099_U30 ; P1_R2099_U111
g29570 nand P1_R2099_U35 P1_R2099_U137 ; P1_R2099_U112
g29571 not P1_U2682 ; P1_R2099_U113
g29572 not P1_U2683 ; P1_R2099_U114
g29573 not P1_U2684 ; P1_R2099_U115
g29574 not P1_U2685 ; P1_R2099_U116
g29575 not P1_U2686 ; P1_R2099_U117
g29576 not P1_U2687 ; P1_R2099_U118
g29577 not P1_U2688 ; P1_R2099_U119
g29578 not P1_U2689 ; P1_R2099_U120
g29579 not P1_U2690 ; P1_R2099_U121
g29580 not P1_U2691 ; P1_R2099_U122
g29581 not P1_U2692 ; P1_R2099_U123
g29582 not P1_U2700 ; P1_R2099_U124
g29583 not P1_U2699 ; P1_R2099_U125
g29584 not P1_U2698 ; P1_R2099_U126
g29585 not P1_U2697 ; P1_R2099_U127
g29586 not P1_U2696 ; P1_R2099_U128
g29587 not P1_U2695 ; P1_R2099_U129
g29588 not P1_U2694 ; P1_R2099_U130
g29589 not P1_U2693 ; P1_R2099_U131
g29590 not P1_U2680 ; P1_R2099_U132
g29591 not P1_U2681 ; P1_R2099_U133
g29592 not P1_U2679 ; P1_R2099_U134
g29593 nand P1_R2099_U96 P1_R2099_U180 ; P1_R2099_U135
g29594 nand P1_R2099_U180 P1_R2099_U44 ; P1_R2099_U136
g29595 nand P1_R2099_U152 P1_R2099_U151 ; P1_R2099_U137
g29596 and P1_R2099_U297 P1_R2099_U296 ; P1_R2099_U138
g29597 and P1_R2099_U319 P1_R2099_U318 ; P1_R2099_U139
g29598 nand P1_R2099_U148 P1_R2099_U147 ; P1_R2099_U140
g29599 nand P1_R2099_U167 P1_R2099_U56 ; P1_R2099_U141
g29600 nand P1_R2099_U165 P1_R2099_U58 ; P1_R2099_U142
g29601 nand P1_R2099_U163 P1_R2099_U60 ; P1_R2099_U143
g29602 nand P1_R2099_U161 P1_R2099_U62 ; P1_R2099_U144
g29603 not P1_R2099_U135 ; P1_R2099_U145
g29604 or P1_U4190 P1_U4189 ; P1_R2099_U146
g29605 nand P1_R2099_U32 P1_R2099_U146 ; P1_R2099_U147
g29606 nand P1_U4189 P1_U4190 ; P1_R2099_U148
g29607 not P1_R2099_U140 ; P1_R2099_U149
g29608 nand P1_R2099_U190 P1_R2099_U6 ; P1_R2099_U150
g29609 nand P1_R2099_U150 P1_R2099_U140 ; P1_R2099_U151
g29610 nand P1_U2678 P1_R2099_U33 ; P1_R2099_U152
g29611 not P1_R2099_U137 ; P1_R2099_U153
g29612 not P1_R2099_U112 ; P1_R2099_U154
g29613 not P1_R2099_U7 ; P1_R2099_U155
g29614 not P1_R2099_U111 ; P1_R2099_U156
g29615 not P1_R2099_U8 ; P1_R2099_U157
g29616 not P1_R2099_U110 ; P1_R2099_U158
g29617 not P1_R2099_U9 ; P1_R2099_U159
g29618 not P1_R2099_U109 ; P1_R2099_U160
g29619 not P1_R2099_U10 ; P1_R2099_U161
g29620 not P1_R2099_U144 ; P1_R2099_U162
g29621 not P1_R2099_U11 ; P1_R2099_U163
g29622 not P1_R2099_U143 ; P1_R2099_U164
g29623 not P1_R2099_U12 ; P1_R2099_U165
g29624 not P1_R2099_U142 ; P1_R2099_U166
g29625 not P1_R2099_U13 ; P1_R2099_U167
g29626 not P1_R2099_U141 ; P1_R2099_U168
g29627 not P1_R2099_U14 ; P1_R2099_U169
g29628 not P1_R2099_U15 ; P1_R2099_U170
g29629 not P1_R2099_U16 ; P1_R2099_U171
g29630 not P1_R2099_U17 ; P1_R2099_U172
g29631 not P1_R2099_U18 ; P1_R2099_U173
g29632 not P1_R2099_U19 ; P1_R2099_U174
g29633 not P1_R2099_U20 ; P1_R2099_U175
g29634 not P1_R2099_U21 ; P1_R2099_U176
g29635 not P1_R2099_U22 ; P1_R2099_U177
g29636 not P1_R2099_U23 ; P1_R2099_U178
g29637 not P1_R2099_U24 ; P1_R2099_U179
g29638 not P1_R2099_U25 ; P1_R2099_U180
g29639 not P1_R2099_U136 ; P1_R2099_U181
g29640 nand P1_U4190 P1_R2099_U99 ; P1_R2099_U182
g29641 nand P1_U2702 P1_R2099_U4 ; P1_R2099_U183
g29642 not P1_R2099_U27 ; P1_R2099_U184
g29643 nand P1_U4190 P1_R2099_U100 ; P1_R2099_U185
g29644 nand P1_U2710 P1_R2099_U4 ; P1_R2099_U186
g29645 not P1_R2099_U32 ; P1_R2099_U187
g29646 nand P1_U4190 P1_R2099_U101 ; P1_R2099_U188
g29647 nand P1_U2709 P1_R2099_U4 ; P1_R2099_U189
g29648 not P1_R2099_U33 ; P1_R2099_U190
g29649 nand P1_U4190 P1_R2099_U102 ; P1_R2099_U191
g29650 nand P1_U2708 P1_R2099_U4 ; P1_R2099_U192
g29651 not P1_R2099_U35 ; P1_R2099_U193
g29652 nand P1_U4190 P1_R2099_U103 ; P1_R2099_U194
g29653 nand P1_U2707 P1_R2099_U4 ; P1_R2099_U195
g29654 not P1_R2099_U34 ; P1_R2099_U196
g29655 nand P1_U4190 P1_R2099_U104 ; P1_R2099_U197
g29656 nand P1_U2706 P1_R2099_U4 ; P1_R2099_U198
g29657 not P1_R2099_U30 ; P1_R2099_U199
g29658 nand P1_U4190 P1_R2099_U105 ; P1_R2099_U200
g29659 nand P1_U2705 P1_R2099_U4 ; P1_R2099_U201
g29660 not P1_R2099_U31 ; P1_R2099_U202
g29661 nand P1_U4190 P1_R2099_U106 ; P1_R2099_U203
g29662 nand P1_U2704 P1_R2099_U4 ; P1_R2099_U204
g29663 not P1_R2099_U28 ; P1_R2099_U205
g29664 nand P1_U4190 P1_R2099_U107 ; P1_R2099_U206
g29665 nand P1_U2703 P1_R2099_U4 ; P1_R2099_U207
g29666 not P1_R2099_U29 ; P1_R2099_U208
g29667 nand P1_U4190 P1_R2099_U108 ; P1_R2099_U209
g29668 nand P1_U2701 P1_R2099_U4 ; P1_R2099_U210
g29669 not P1_R2099_U26 ; P1_R2099_U211
g29670 nand P1_R2099_U160 P1_R2099_U211 ; P1_R2099_U212
g29671 nand P1_R2099_U26 P1_R2099_U109 ; P1_R2099_U213
g29672 nand P1_R2099_U184 P1_R2099_U159 ; P1_R2099_U214
g29673 nand P1_R2099_U27 P1_R2099_U9 ; P1_R2099_U215
g29674 nand P1_R2099_U158 P1_R2099_U208 ; P1_R2099_U216
g29675 nand P1_R2099_U29 P1_R2099_U110 ; P1_R2099_U217
g29676 nand P1_R2099_U205 P1_R2099_U157 ; P1_R2099_U218
g29677 nand P1_R2099_U28 P1_R2099_U8 ; P1_R2099_U219
g29678 nand P1_R2099_U156 P1_R2099_U202 ; P1_R2099_U220
g29679 nand P1_R2099_U31 P1_R2099_U111 ; P1_R2099_U221
g29680 nand P1_R2099_U199 P1_R2099_U155 ; P1_R2099_U222
g29681 nand P1_R2099_U30 P1_R2099_U7 ; P1_R2099_U223
g29682 nand P1_R2099_U154 P1_R2099_U196 ; P1_R2099_U224
g29683 nand P1_R2099_U34 P1_R2099_U112 ; P1_R2099_U225
g29684 nand P1_U4190 P1_R2099_U113 ; P1_R2099_U226
g29685 nand P1_U2682 P1_R2099_U4 ; P1_R2099_U227
g29686 not P1_R2099_U45 ; P1_R2099_U228
g29687 nand P1_U4190 P1_R2099_U114 ; P1_R2099_U229
g29688 nand P1_U2683 P1_R2099_U4 ; P1_R2099_U230
g29689 not P1_R2099_U46 ; P1_R2099_U231
g29690 nand P1_U4190 P1_R2099_U115 ; P1_R2099_U232
g29691 nand P1_U2684 P1_R2099_U4 ; P1_R2099_U233
g29692 not P1_R2099_U47 ; P1_R2099_U234
g29693 nand P1_U4190 P1_R2099_U116 ; P1_R2099_U235
g29694 nand P1_U2685 P1_R2099_U4 ; P1_R2099_U236
g29695 not P1_R2099_U48 ; P1_R2099_U237
g29696 nand P1_U4190 P1_R2099_U117 ; P1_R2099_U238
g29697 nand P1_U2686 P1_R2099_U4 ; P1_R2099_U239
g29698 not P1_R2099_U49 ; P1_R2099_U240
g29699 nand P1_U4190 P1_R2099_U118 ; P1_R2099_U241
g29700 nand P1_U2687 P1_R2099_U4 ; P1_R2099_U242
g29701 not P1_R2099_U50 ; P1_R2099_U243
g29702 nand P1_U4190 P1_R2099_U119 ; P1_R2099_U244
g29703 nand P1_U2688 P1_R2099_U4 ; P1_R2099_U245
g29704 not P1_R2099_U51 ; P1_R2099_U246
g29705 nand P1_U4190 P1_R2099_U120 ; P1_R2099_U247
g29706 nand P1_U2689 P1_R2099_U4 ; P1_R2099_U248
g29707 not P1_R2099_U52 ; P1_R2099_U249
g29708 nand P1_U4190 P1_R2099_U121 ; P1_R2099_U250
g29709 nand P1_U2690 P1_R2099_U4 ; P1_R2099_U251
g29710 not P1_R2099_U53 ; P1_R2099_U252
g29711 nand P1_U4190 P1_R2099_U122 ; P1_R2099_U253
g29712 nand P1_U2691 P1_R2099_U4 ; P1_R2099_U254
g29713 not P1_R2099_U54 ; P1_R2099_U255
g29714 nand P1_U4190 P1_R2099_U123 ; P1_R2099_U256
g29715 nand P1_U2692 P1_R2099_U4 ; P1_R2099_U257
g29716 not P1_R2099_U55 ; P1_R2099_U258
g29717 nand P1_U4190 P1_R2099_U124 ; P1_R2099_U259
g29718 nand P1_U2700 P1_R2099_U4 ; P1_R2099_U260
g29719 not P1_R2099_U62 ; P1_R2099_U261
g29720 nand P1_U4190 P1_R2099_U125 ; P1_R2099_U262
g29721 nand P1_U2699 P1_R2099_U4 ; P1_R2099_U263
g29722 not P1_R2099_U63 ; P1_R2099_U264
g29723 nand P1_U4190 P1_R2099_U126 ; P1_R2099_U265
g29724 nand P1_U2698 P1_R2099_U4 ; P1_R2099_U266
g29725 not P1_R2099_U60 ; P1_R2099_U267
g29726 nand P1_U4190 P1_R2099_U127 ; P1_R2099_U268
g29727 nand P1_U2697 P1_R2099_U4 ; P1_R2099_U269
g29728 not P1_R2099_U61 ; P1_R2099_U270
g29729 nand P1_U4190 P1_R2099_U128 ; P1_R2099_U271
g29730 nand P1_U2696 P1_R2099_U4 ; P1_R2099_U272
g29731 not P1_R2099_U58 ; P1_R2099_U273
g29732 nand P1_U4190 P1_R2099_U129 ; P1_R2099_U274
g29733 nand P1_U2695 P1_R2099_U4 ; P1_R2099_U275
g29734 not P1_R2099_U59 ; P1_R2099_U276
g29735 nand P1_U4190 P1_R2099_U130 ; P1_R2099_U277
g29736 nand P1_U2694 P1_R2099_U4 ; P1_R2099_U278
g29737 not P1_R2099_U56 ; P1_R2099_U279
g29738 nand P1_U4190 P1_R2099_U131 ; P1_R2099_U280
g29739 nand P1_U2693 P1_R2099_U4 ; P1_R2099_U281
g29740 not P1_R2099_U57 ; P1_R2099_U282
g29741 nand P1_U4190 P1_R2099_U132 ; P1_R2099_U283
g29742 nand P1_U2680 P1_R2099_U4 ; P1_R2099_U284
g29743 not P1_R2099_U43 ; P1_R2099_U285
g29744 nand P1_U4190 P1_R2099_U133 ; P1_R2099_U286
g29745 nand P1_U2681 P1_R2099_U4 ; P1_R2099_U287
g29746 not P1_R2099_U44 ; P1_R2099_U288
g29747 nand P1_U4190 P1_R2099_U134 ; P1_R2099_U289
g29748 nand P1_U2679 P1_R2099_U4 ; P1_R2099_U290
g29749 not P1_R2099_U97 ; P1_R2099_U291
g29750 nand P1_R2099_U145 P1_R2099_U291 ; P1_R2099_U292
g29751 nand P1_R2099_U97 P1_R2099_U135 ; P1_R2099_U293
g29752 nand P1_R2099_U181 P1_R2099_U285 ; P1_R2099_U294
g29753 nand P1_R2099_U43 P1_R2099_U136 ; P1_R2099_U295
g29754 nand P1_R2099_U153 P1_R2099_U193 ; P1_R2099_U296
g29755 nand P1_R2099_U35 P1_R2099_U137 ; P1_R2099_U297
g29756 nand P1_R2099_U288 P1_R2099_U180 ; P1_R2099_U298
g29757 nand P1_R2099_U44 P1_R2099_U25 ; P1_R2099_U299
g29758 nand P1_R2099_U228 P1_R2099_U179 ; P1_R2099_U300
g29759 nand P1_R2099_U45 P1_R2099_U24 ; P1_R2099_U301
g29760 nand P1_R2099_U231 P1_R2099_U178 ; P1_R2099_U302
g29761 nand P1_R2099_U46 P1_R2099_U23 ; P1_R2099_U303
g29762 nand P1_R2099_U234 P1_R2099_U177 ; P1_R2099_U304
g29763 nand P1_R2099_U47 P1_R2099_U22 ; P1_R2099_U305
g29764 nand P1_R2099_U237 P1_R2099_U176 ; P1_R2099_U306
g29765 nand P1_R2099_U48 P1_R2099_U21 ; P1_R2099_U307
g29766 nand P1_R2099_U240 P1_R2099_U175 ; P1_R2099_U308
g29767 nand P1_R2099_U49 P1_R2099_U20 ; P1_R2099_U309
g29768 nand P1_R2099_U243 P1_R2099_U174 ; P1_R2099_U310
g29769 nand P1_R2099_U50 P1_R2099_U19 ; P1_R2099_U311
g29770 nand P1_R2099_U246 P1_R2099_U173 ; P1_R2099_U312
g29771 nand P1_R2099_U51 P1_R2099_U18 ; P1_R2099_U313
g29772 nand P1_R2099_U249 P1_R2099_U172 ; P1_R2099_U314
g29773 nand P1_R2099_U52 P1_R2099_U17 ; P1_R2099_U315
g29774 nand P1_R2099_U252 P1_R2099_U171 ; P1_R2099_U316
g29775 nand P1_R2099_U53 P1_R2099_U16 ; P1_R2099_U317
g29776 nand P1_R2099_U190 P1_U2678 ; P1_R2099_U318
g29777 nand P1_R2099_U33 P1_R2099_U6 ; P1_R2099_U319
g29778 nand P1_R2099_U190 P1_U2678 ; P1_R2099_U320
g29779 nand P1_R2099_U33 P1_R2099_U6 ; P1_R2099_U321
g29780 nand P1_R2099_U321 P1_R2099_U320 ; P1_R2099_U322
g29781 nand P1_R2099_U139 P1_R2099_U140 ; P1_R2099_U323
g29782 nand P1_R2099_U149 P1_R2099_U322 ; P1_R2099_U324
g29783 nand P1_R2099_U255 P1_R2099_U170 ; P1_R2099_U325
g29784 nand P1_R2099_U54 P1_R2099_U15 ; P1_R2099_U326
g29785 nand P1_R2099_U258 P1_R2099_U169 ; P1_R2099_U327
g29786 nand P1_R2099_U55 P1_R2099_U14 ; P1_R2099_U328
g29787 nand P1_R2099_U168 P1_R2099_U282 ; P1_R2099_U329
g29788 nand P1_R2099_U57 P1_R2099_U141 ; P1_R2099_U330
g29789 nand P1_R2099_U279 P1_R2099_U167 ; P1_R2099_U331
g29790 nand P1_R2099_U56 P1_R2099_U13 ; P1_R2099_U332
g29791 nand P1_R2099_U166 P1_R2099_U276 ; P1_R2099_U333
g29792 nand P1_R2099_U59 P1_R2099_U142 ; P1_R2099_U334
g29793 nand P1_R2099_U273 P1_R2099_U165 ; P1_R2099_U335
g29794 nand P1_R2099_U58 P1_R2099_U12 ; P1_R2099_U336
g29795 nand P1_R2099_U164 P1_R2099_U270 ; P1_R2099_U337
g29796 nand P1_R2099_U61 P1_R2099_U143 ; P1_R2099_U338
g29797 nand P1_R2099_U267 P1_R2099_U163 ; P1_R2099_U339
g29798 nand P1_R2099_U60 P1_R2099_U11 ; P1_R2099_U340
g29799 nand P1_R2099_U162 P1_R2099_U264 ; P1_R2099_U341
g29800 nand P1_R2099_U63 P1_R2099_U144 ; P1_R2099_U342
g29801 nand P1_R2099_U261 P1_R2099_U161 ; P1_R2099_U343
g29802 nand P1_R2099_U62 P1_R2099_U10 ; P1_R2099_U344
g29803 nand P1_U4189 P1_R2099_U4 ; P1_R2099_U345
g29804 nand P1_U4190 P1_R2099_U5 ; P1_R2099_U346
g29805 not P1_R2099_U98 ; P1_R2099_U347
g29806 nand P1_R2099_U32 P1_R2099_U347 ; P1_R2099_U348
g29807 nand P1_R2099_U98 P1_R2099_U187 ; P1_R2099_U349
g29808 not P1_U2716 ; P1_R2167_U6
g29809 not P1_U2714 ; P1_R2167_U7
g29810 not P1_U2720 ; P1_R2167_U8
g29811 not P1_U2719 ; P1_R2167_U9
g29812 not P1_U2713 ; P1_R2167_U10
g29813 not P1_U2712 ; P1_R2167_U11
g29814 not P1_U2718 ; P1_R2167_U12
g29815 not P1_U2717 ; P1_R2167_U13
g29816 not P1_U2711 ; P1_R2167_U14
g29817 not P1_U2356 ; P1_R2167_U15
g29818 not P1_STATE2_REG_0__SCAN_IN ; P1_R2167_U16
g29819 nand P1_R2167_U50 P1_R2167_U49 ; P1_R2167_U17
g29820 and P1_R2167_U29 P1_R2167_U30 ; P1_R2167_U18
g29821 and P1_R2167_U32 P1_R2167_U33 ; P1_R2167_U19
g29822 and P1_R2167_U35 P1_R2167_U36 ; P1_R2167_U20
g29823 and P1_R2167_U38 P1_R2167_U39 ; P1_R2167_U21
g29824 not P1_U2721 ; P1_R2167_U22
g29825 not P1_U2722 ; P1_R2167_U23
g29826 nand P1_U2715 P1_R2167_U23 ; P1_R2167_U24
g29827 nand P1_U2715 P1_R2167_U22 ; P1_R2167_U25
g29828 or P1_U2721 P1_U2722 ; P1_R2167_U26
g29829 nand P1_U2714 P1_R2167_U8 ; P1_R2167_U27
g29830 nand P1_R2167_U27 P1_R2167_U26 P1_R2167_U25 P1_R2167_U24 ; P1_R2167_U28
g29831 nand P1_U2720 P1_R2167_U7 ; P1_R2167_U29
g29832 nand P1_U2719 P1_R2167_U10 ; P1_R2167_U30
g29833 nand P1_R2167_U18 P1_R2167_U28 ; P1_R2167_U31
g29834 nand P1_U2713 P1_R2167_U9 ; P1_R2167_U32
g29835 nand P1_U2712 P1_R2167_U12 ; P1_R2167_U33
g29836 nand P1_R2167_U19 P1_R2167_U31 ; P1_R2167_U34
g29837 nand P1_U2718 P1_R2167_U11 ; P1_R2167_U35
g29838 nand P1_U2717 P1_R2167_U14 ; P1_R2167_U36
g29839 nand P1_R2167_U20 P1_R2167_U34 ; P1_R2167_U37
g29840 nand P1_U2711 P1_R2167_U13 ; P1_R2167_U38
g29841 nand P1_U2356 P1_R2167_U6 ; P1_R2167_U39
g29842 nand P1_R2167_U21 P1_R2167_U37 ; P1_R2167_U40
g29843 nand P1_U2716 P1_R2167_U15 ; P1_R2167_U41
g29844 nand P1_R2167_U40 P1_R2167_U41 ; P1_R2167_U42
g29845 nand P1_U2716 P1_R2167_U16 ; P1_R2167_U43
g29846 nand P1_R2167_U42 P1_R2167_U6 ; P1_R2167_U44
g29847 nand P1_R2167_U44 P1_R2167_U43 ; P1_R2167_U45
g29848 nand P1_R2167_U6 P1_STATE2_REG_0__SCAN_IN ; P1_R2167_U46
g29849 nand P1_U2716 P1_R2167_U42 ; P1_R2167_U47
g29850 nand P1_R2167_U47 P1_R2167_U46 ; P1_R2167_U48
g29851 nand P1_R2167_U45 P1_R2167_U15 ; P1_R2167_U49
g29852 nand P1_U2356 P1_R2167_U48 ; P1_R2167_U50
g29853 not P1_PHYADDRPOINTER_REG_1__SCAN_IN ; P1_R2337_U4
g29854 not P1_PHYADDRPOINTER_REG_2__SCAN_IN ; P1_R2337_U5
g29855 nand P1_PHYADDRPOINTER_REG_1__SCAN_IN P1_PHYADDRPOINTER_REG_2__SCAN_IN ; P1_R2337_U6
g29856 not P1_PHYADDRPOINTER_REG_3__SCAN_IN ; P1_R2337_U7
g29857 nand P1_R2337_U94 P1_PHYADDRPOINTER_REG_3__SCAN_IN ; P1_R2337_U8
g29858 not P1_PHYADDRPOINTER_REG_4__SCAN_IN ; P1_R2337_U9
g29859 nand P1_R2337_U95 P1_PHYADDRPOINTER_REG_4__SCAN_IN ; P1_R2337_U10
g29860 not P1_PHYADDRPOINTER_REG_5__SCAN_IN ; P1_R2337_U11
g29861 nand P1_R2337_U96 P1_PHYADDRPOINTER_REG_5__SCAN_IN ; P1_R2337_U12
g29862 not P1_PHYADDRPOINTER_REG_6__SCAN_IN ; P1_R2337_U13
g29863 nand P1_R2337_U97 P1_PHYADDRPOINTER_REG_6__SCAN_IN ; P1_R2337_U14
g29864 not P1_PHYADDRPOINTER_REG_7__SCAN_IN ; P1_R2337_U15
g29865 nand P1_R2337_U98 P1_PHYADDRPOINTER_REG_7__SCAN_IN ; P1_R2337_U16
g29866 not P1_PHYADDRPOINTER_REG_8__SCAN_IN ; P1_R2337_U17
g29867 not P1_PHYADDRPOINTER_REG_9__SCAN_IN ; P1_R2337_U18
g29868 nand P1_R2337_U99 P1_PHYADDRPOINTER_REG_8__SCAN_IN ; P1_R2337_U19
g29869 nand P1_R2337_U100 P1_PHYADDRPOINTER_REG_9__SCAN_IN ; P1_R2337_U20
g29870 not P1_PHYADDRPOINTER_REG_10__SCAN_IN ; P1_R2337_U21
g29871 nand P1_R2337_U101 P1_PHYADDRPOINTER_REG_10__SCAN_IN ; P1_R2337_U22
g29872 not P1_PHYADDRPOINTER_REG_11__SCAN_IN ; P1_R2337_U23
g29873 nand P1_R2337_U102 P1_PHYADDRPOINTER_REG_11__SCAN_IN ; P1_R2337_U24
g29874 not P1_PHYADDRPOINTER_REG_12__SCAN_IN ; P1_R2337_U25
g29875 nand P1_R2337_U103 P1_PHYADDRPOINTER_REG_12__SCAN_IN ; P1_R2337_U26
g29876 not P1_PHYADDRPOINTER_REG_13__SCAN_IN ; P1_R2337_U27
g29877 nand P1_R2337_U104 P1_PHYADDRPOINTER_REG_13__SCAN_IN ; P1_R2337_U28
g29878 not P1_PHYADDRPOINTER_REG_14__SCAN_IN ; P1_R2337_U29
g29879 nand P1_R2337_U105 P1_PHYADDRPOINTER_REG_14__SCAN_IN ; P1_R2337_U30
g29880 not P1_PHYADDRPOINTER_REG_15__SCAN_IN ; P1_R2337_U31
g29881 nand P1_R2337_U106 P1_PHYADDRPOINTER_REG_15__SCAN_IN ; P1_R2337_U32
g29882 not P1_PHYADDRPOINTER_REG_16__SCAN_IN ; P1_R2337_U33
g29883 nand P1_R2337_U107 P1_PHYADDRPOINTER_REG_16__SCAN_IN ; P1_R2337_U34
g29884 not P1_PHYADDRPOINTER_REG_17__SCAN_IN ; P1_R2337_U35
g29885 nand P1_R2337_U108 P1_PHYADDRPOINTER_REG_17__SCAN_IN ; P1_R2337_U36
g29886 not P1_PHYADDRPOINTER_REG_18__SCAN_IN ; P1_R2337_U37
g29887 nand P1_R2337_U109 P1_PHYADDRPOINTER_REG_18__SCAN_IN ; P1_R2337_U38
g29888 not P1_PHYADDRPOINTER_REG_19__SCAN_IN ; P1_R2337_U39
g29889 nand P1_R2337_U110 P1_PHYADDRPOINTER_REG_19__SCAN_IN ; P1_R2337_U40
g29890 not P1_PHYADDRPOINTER_REG_20__SCAN_IN ; P1_R2337_U41
g29891 nand P1_R2337_U111 P1_PHYADDRPOINTER_REG_20__SCAN_IN ; P1_R2337_U42
g29892 not P1_PHYADDRPOINTER_REG_21__SCAN_IN ; P1_R2337_U43
g29893 nand P1_R2337_U112 P1_PHYADDRPOINTER_REG_21__SCAN_IN ; P1_R2337_U44
g29894 not P1_PHYADDRPOINTER_REG_22__SCAN_IN ; P1_R2337_U45
g29895 nand P1_R2337_U113 P1_PHYADDRPOINTER_REG_22__SCAN_IN ; P1_R2337_U46
g29896 not P1_PHYADDRPOINTER_REG_23__SCAN_IN ; P1_R2337_U47
g29897 nand P1_R2337_U114 P1_PHYADDRPOINTER_REG_23__SCAN_IN ; P1_R2337_U48
g29898 not P1_PHYADDRPOINTER_REG_24__SCAN_IN ; P1_R2337_U49
g29899 nand P1_R2337_U115 P1_PHYADDRPOINTER_REG_24__SCAN_IN ; P1_R2337_U50
g29900 not P1_PHYADDRPOINTER_REG_25__SCAN_IN ; P1_R2337_U51
g29901 nand P1_R2337_U116 P1_PHYADDRPOINTER_REG_25__SCAN_IN ; P1_R2337_U52
g29902 not P1_PHYADDRPOINTER_REG_26__SCAN_IN ; P1_R2337_U53
g29903 nand P1_R2337_U117 P1_PHYADDRPOINTER_REG_26__SCAN_IN ; P1_R2337_U54
g29904 not P1_PHYADDRPOINTER_REG_27__SCAN_IN ; P1_R2337_U55
g29905 nand P1_R2337_U118 P1_PHYADDRPOINTER_REG_27__SCAN_IN ; P1_R2337_U56
g29906 not P1_PHYADDRPOINTER_REG_28__SCAN_IN ; P1_R2337_U57
g29907 nand P1_R2337_U119 P1_PHYADDRPOINTER_REG_28__SCAN_IN ; P1_R2337_U58
g29908 not P1_PHYADDRPOINTER_REG_29__SCAN_IN ; P1_R2337_U59
g29909 nand P1_R2337_U120 P1_PHYADDRPOINTER_REG_29__SCAN_IN ; P1_R2337_U60
g29910 not P1_PHYADDRPOINTER_REG_30__SCAN_IN ; P1_R2337_U61
g29911 nand P1_R2337_U124 P1_R2337_U123 ; P1_R2337_U62
g29912 nand P1_R2337_U126 P1_R2337_U125 ; P1_R2337_U63
g29913 nand P1_R2337_U128 P1_R2337_U127 ; P1_R2337_U64
g29914 nand P1_R2337_U130 P1_R2337_U129 ; P1_R2337_U65
g29915 nand P1_R2337_U132 P1_R2337_U131 ; P1_R2337_U66
g29916 nand P1_R2337_U134 P1_R2337_U133 ; P1_R2337_U67
g29917 nand P1_R2337_U136 P1_R2337_U135 ; P1_R2337_U68
g29918 nand P1_R2337_U138 P1_R2337_U137 ; P1_R2337_U69
g29919 nand P1_R2337_U140 P1_R2337_U139 ; P1_R2337_U70
g29920 nand P1_R2337_U142 P1_R2337_U141 ; P1_R2337_U71
g29921 nand P1_R2337_U144 P1_R2337_U143 ; P1_R2337_U72
g29922 nand P1_R2337_U146 P1_R2337_U145 ; P1_R2337_U73
g29923 nand P1_R2337_U148 P1_R2337_U147 ; P1_R2337_U74
g29924 nand P1_R2337_U150 P1_R2337_U149 ; P1_R2337_U75
g29925 nand P1_R2337_U152 P1_R2337_U151 ; P1_R2337_U76
g29926 nand P1_R2337_U154 P1_R2337_U153 ; P1_R2337_U77
g29927 nand P1_R2337_U156 P1_R2337_U155 ; P1_R2337_U78
g29928 nand P1_R2337_U158 P1_R2337_U157 ; P1_R2337_U79
g29929 nand P1_R2337_U160 P1_R2337_U159 ; P1_R2337_U80
g29930 nand P1_R2337_U162 P1_R2337_U161 ; P1_R2337_U81
g29931 nand P1_R2337_U164 P1_R2337_U163 ; P1_R2337_U82
g29932 nand P1_R2337_U166 P1_R2337_U165 ; P1_R2337_U83
g29933 nand P1_R2337_U168 P1_R2337_U167 ; P1_R2337_U84
g29934 nand P1_R2337_U170 P1_R2337_U169 ; P1_R2337_U85
g29935 nand P1_R2337_U172 P1_R2337_U171 ; P1_R2337_U86
g29936 nand P1_R2337_U174 P1_R2337_U173 ; P1_R2337_U87
g29937 nand P1_R2337_U176 P1_R2337_U175 ; P1_R2337_U88
g29938 nand P1_R2337_U178 P1_R2337_U177 ; P1_R2337_U89
g29939 nand P1_R2337_U180 P1_R2337_U179 ; P1_R2337_U90
g29940 nand P1_R2337_U182 P1_R2337_U181 ; P1_R2337_U91
g29941 not P1_PHYADDRPOINTER_REG_31__SCAN_IN ; P1_R2337_U92
g29942 nand P1_R2337_U121 P1_PHYADDRPOINTER_REG_30__SCAN_IN ; P1_R2337_U93
g29943 not P1_R2337_U6 ; P1_R2337_U94
g29944 not P1_R2337_U8 ; P1_R2337_U95
g29945 not P1_R2337_U10 ; P1_R2337_U96
g29946 not P1_R2337_U12 ; P1_R2337_U97
g29947 not P1_R2337_U14 ; P1_R2337_U98
g29948 not P1_R2337_U16 ; P1_R2337_U99
g29949 not P1_R2337_U19 ; P1_R2337_U100
g29950 not P1_R2337_U20 ; P1_R2337_U101
g29951 not P1_R2337_U22 ; P1_R2337_U102
g29952 not P1_R2337_U24 ; P1_R2337_U103
g29953 not P1_R2337_U26 ; P1_R2337_U104
g29954 not P1_R2337_U28 ; P1_R2337_U105
g29955 not P1_R2337_U30 ; P1_R2337_U106
g29956 not P1_R2337_U32 ; P1_R2337_U107
g29957 not P1_R2337_U34 ; P1_R2337_U108
g29958 not P1_R2337_U36 ; P1_R2337_U109
g29959 not P1_R2337_U38 ; P1_R2337_U110
g29960 not P1_R2337_U40 ; P1_R2337_U111
g29961 not P1_R2337_U42 ; P1_R2337_U112
g29962 not P1_R2337_U44 ; P1_R2337_U113
g29963 not P1_R2337_U46 ; P1_R2337_U114
g29964 not P1_R2337_U48 ; P1_R2337_U115
g29965 not P1_R2337_U50 ; P1_R2337_U116
g29966 not P1_R2337_U52 ; P1_R2337_U117
g29967 not P1_R2337_U54 ; P1_R2337_U118
g29968 not P1_R2337_U56 ; P1_R2337_U119
g29969 not P1_R2337_U58 ; P1_R2337_U120
g29970 not P1_R2337_U60 ; P1_R2337_U121
g29971 not P1_R2337_U93 ; P1_R2337_U122
g29972 nand P1_R2337_U19 P1_PHYADDRPOINTER_REG_9__SCAN_IN ; P1_R2337_U123
g29973 nand P1_R2337_U100 P1_R2337_U18 ; P1_R2337_U124
g29974 nand P1_R2337_U16 P1_PHYADDRPOINTER_REG_8__SCAN_IN ; P1_R2337_U125
g29975 nand P1_R2337_U99 P1_R2337_U17 ; P1_R2337_U126
g29976 nand P1_R2337_U14 P1_PHYADDRPOINTER_REG_7__SCAN_IN ; P1_R2337_U127
g29977 nand P1_R2337_U98 P1_R2337_U15 ; P1_R2337_U128
g29978 nand P1_R2337_U12 P1_PHYADDRPOINTER_REG_6__SCAN_IN ; P1_R2337_U129
g29979 nand P1_R2337_U97 P1_R2337_U13 ; P1_R2337_U130
g29980 nand P1_R2337_U10 P1_PHYADDRPOINTER_REG_5__SCAN_IN ; P1_R2337_U131
g29981 nand P1_R2337_U96 P1_R2337_U11 ; P1_R2337_U132
g29982 nand P1_R2337_U8 P1_PHYADDRPOINTER_REG_4__SCAN_IN ; P1_R2337_U133
g29983 nand P1_R2337_U95 P1_R2337_U9 ; P1_R2337_U134
g29984 nand P1_R2337_U6 P1_PHYADDRPOINTER_REG_3__SCAN_IN ; P1_R2337_U135
g29985 nand P1_R2337_U94 P1_R2337_U7 ; P1_R2337_U136
g29986 nand P1_R2337_U93 P1_PHYADDRPOINTER_REG_31__SCAN_IN ; P1_R2337_U137
g29987 nand P1_R2337_U122 P1_R2337_U92 ; P1_R2337_U138
g29988 nand P1_R2337_U60 P1_PHYADDRPOINTER_REG_30__SCAN_IN ; P1_R2337_U139
g29989 nand P1_R2337_U121 P1_R2337_U61 ; P1_R2337_U140
g29990 nand P1_R2337_U4 P1_PHYADDRPOINTER_REG_2__SCAN_IN ; P1_R2337_U141
g29991 nand P1_R2337_U5 P1_PHYADDRPOINTER_REG_1__SCAN_IN ; P1_R2337_U142
g29992 nand P1_R2337_U58 P1_PHYADDRPOINTER_REG_29__SCAN_IN ; P1_R2337_U143
g29993 nand P1_R2337_U120 P1_R2337_U59 ; P1_R2337_U144
g29994 nand P1_R2337_U56 P1_PHYADDRPOINTER_REG_28__SCAN_IN ; P1_R2337_U145
g29995 nand P1_R2337_U119 P1_R2337_U57 ; P1_R2337_U146
g29996 nand P1_R2337_U54 P1_PHYADDRPOINTER_REG_27__SCAN_IN ; P1_R2337_U147
g29997 nand P1_R2337_U118 P1_R2337_U55 ; P1_R2337_U148
g29998 nand P1_R2337_U52 P1_PHYADDRPOINTER_REG_26__SCAN_IN ; P1_R2337_U149
g29999 nand P1_R2337_U117 P1_R2337_U53 ; P1_R2337_U150
g30000 nand P1_R2337_U50 P1_PHYADDRPOINTER_REG_25__SCAN_IN ; P1_R2337_U151
g30001 nand P1_R2337_U116 P1_R2337_U51 ; P1_R2337_U152
g30002 nand P1_R2337_U48 P1_PHYADDRPOINTER_REG_24__SCAN_IN ; P1_R2337_U153
g30003 nand P1_R2337_U115 P1_R2337_U49 ; P1_R2337_U154
g30004 nand P1_R2337_U46 P1_PHYADDRPOINTER_REG_23__SCAN_IN ; P1_R2337_U155
g30005 nand P1_R2337_U114 P1_R2337_U47 ; P1_R2337_U156
g30006 nand P1_R2337_U44 P1_PHYADDRPOINTER_REG_22__SCAN_IN ; P1_R2337_U157
g30007 nand P1_R2337_U113 P1_R2337_U45 ; P1_R2337_U158
g30008 nand P1_R2337_U42 P1_PHYADDRPOINTER_REG_21__SCAN_IN ; P1_R2337_U159
g30009 nand P1_R2337_U112 P1_R2337_U43 ; P1_R2337_U160
g30010 nand P1_R2337_U40 P1_PHYADDRPOINTER_REG_20__SCAN_IN ; P1_R2337_U161
g30011 nand P1_R2337_U111 P1_R2337_U41 ; P1_R2337_U162
g30012 nand P1_R2337_U38 P1_PHYADDRPOINTER_REG_19__SCAN_IN ; P1_R2337_U163
g30013 nand P1_R2337_U110 P1_R2337_U39 ; P1_R2337_U164
g30014 nand P1_R2337_U36 P1_PHYADDRPOINTER_REG_18__SCAN_IN ; P1_R2337_U165
g30015 nand P1_R2337_U109 P1_R2337_U37 ; P1_R2337_U166
g30016 nand P1_R2337_U34 P1_PHYADDRPOINTER_REG_17__SCAN_IN ; P1_R2337_U167
g30017 nand P1_R2337_U108 P1_R2337_U35 ; P1_R2337_U168
g30018 nand P1_R2337_U32 P1_PHYADDRPOINTER_REG_16__SCAN_IN ; P1_R2337_U169
g30019 nand P1_R2337_U107 P1_R2337_U33 ; P1_R2337_U170
g30020 nand P1_R2337_U30 P1_PHYADDRPOINTER_REG_15__SCAN_IN ; P1_R2337_U171
g30021 nand P1_R2337_U106 P1_R2337_U31 ; P1_R2337_U172
g30022 nand P1_R2337_U28 P1_PHYADDRPOINTER_REG_14__SCAN_IN ; P1_R2337_U173
g30023 nand P1_R2337_U105 P1_R2337_U29 ; P1_R2337_U174
g30024 nand P1_R2337_U26 P1_PHYADDRPOINTER_REG_13__SCAN_IN ; P1_R2337_U175
g30025 nand P1_R2337_U104 P1_R2337_U27 ; P1_R2337_U176
g30026 nand P1_R2337_U24 P1_PHYADDRPOINTER_REG_12__SCAN_IN ; P1_R2337_U177
g30027 nand P1_R2337_U103 P1_R2337_U25 ; P1_R2337_U178
g30028 nand P1_R2337_U22 P1_PHYADDRPOINTER_REG_11__SCAN_IN ; P1_R2337_U179
g30029 nand P1_R2337_U102 P1_R2337_U23 ; P1_R2337_U180
g30030 nand P1_R2337_U20 P1_PHYADDRPOINTER_REG_10__SCAN_IN ; P1_R2337_U181
g30031 nand P1_R2337_U101 P1_R2337_U21 ; P1_R2337_U182
g30032 not P1_U3233 ; P1_SUB_357_U6
g30033 not P1_U3228 ; P1_SUB_357_U7
g30034 not P1_U3234 ; P1_SUB_357_U8
g30035 not P1_U3232 ; P1_SUB_357_U9
g30036 not P1_U3227 ; P1_SUB_357_U10
g30037 not P1_U3230 ; P1_SUB_357_U11
g30038 not P1_U3229 ; P1_SUB_357_U12
g30039 not P1_U3231 ; P1_SUB_357_U13
g30040 and P1_LT_563_1260_U9 P1_LT_563_1260_U8 ; P1_LT_563_1260_U6
g30041 not P1_U2673 ; P1_LT_563_1260_U7
g30042 nand P1_R584_U8 P1_LT_563_1260_U7 ; P1_LT_563_1260_U8
g30043 nand P1_R584_U9 P1_LT_563_1260_U7 ; P1_LT_563_1260_U9
g30044 nand P1_SUB_580_U10 P1_SUB_580_U9 ; P1_SUB_580_U6
g30045 not P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_SUB_580_U7
g30046 not P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_SUB_580_U8
g30047 nand P1_SUB_580_U8 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_SUB_580_U9
g30048 nand P1_SUB_580_U7 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_SUB_580_U10
g30049 not P1_REIP_REG_1__SCAN_IN ; P1_R2096_U4
g30050 not P1_REIP_REG_2__SCAN_IN ; P1_R2096_U5
g30051 nand P1_REIP_REG_1__SCAN_IN P1_REIP_REG_2__SCAN_IN ; P1_R2096_U6
g30052 not P1_REIP_REG_3__SCAN_IN ; P1_R2096_U7
g30053 nand P1_R2096_U94 P1_REIP_REG_3__SCAN_IN ; P1_R2096_U8
g30054 not P1_REIP_REG_4__SCAN_IN ; P1_R2096_U9
g30055 nand P1_R2096_U95 P1_REIP_REG_4__SCAN_IN ; P1_R2096_U10
g30056 not P1_REIP_REG_5__SCAN_IN ; P1_R2096_U11
g30057 nand P1_R2096_U96 P1_REIP_REG_5__SCAN_IN ; P1_R2096_U12
g30058 not P1_REIP_REG_6__SCAN_IN ; P1_R2096_U13
g30059 nand P1_R2096_U97 P1_REIP_REG_6__SCAN_IN ; P1_R2096_U14
g30060 not P1_REIP_REG_7__SCAN_IN ; P1_R2096_U15
g30061 nand P1_R2096_U98 P1_REIP_REG_7__SCAN_IN ; P1_R2096_U16
g30062 not P1_REIP_REG_8__SCAN_IN ; P1_R2096_U17
g30063 not P1_REIP_REG_9__SCAN_IN ; P1_R2096_U18
g30064 nand P1_R2096_U99 P1_REIP_REG_8__SCAN_IN ; P1_R2096_U19
g30065 nand P1_R2096_U100 P1_REIP_REG_9__SCAN_IN ; P1_R2096_U20
g30066 not P1_REIP_REG_10__SCAN_IN ; P1_R2096_U21
g30067 nand P1_R2096_U101 P1_REIP_REG_10__SCAN_IN ; P1_R2096_U22
g30068 not P1_REIP_REG_11__SCAN_IN ; P1_R2096_U23
g30069 nand P1_R2096_U102 P1_REIP_REG_11__SCAN_IN ; P1_R2096_U24
g30070 not P1_REIP_REG_12__SCAN_IN ; P1_R2096_U25
g30071 nand P1_R2096_U103 P1_REIP_REG_12__SCAN_IN ; P1_R2096_U26
g30072 not P1_REIP_REG_13__SCAN_IN ; P1_R2096_U27
g30073 nand P1_R2096_U104 P1_REIP_REG_13__SCAN_IN ; P1_R2096_U28
g30074 not P1_REIP_REG_14__SCAN_IN ; P1_R2096_U29
g30075 nand P1_R2096_U105 P1_REIP_REG_14__SCAN_IN ; P1_R2096_U30
g30076 not P1_REIP_REG_15__SCAN_IN ; P1_R2096_U31
g30077 nand P1_R2096_U106 P1_REIP_REG_15__SCAN_IN ; P1_R2096_U32
g30078 not P1_REIP_REG_16__SCAN_IN ; P1_R2096_U33
g30079 nand P1_R2096_U107 P1_REIP_REG_16__SCAN_IN ; P1_R2096_U34
g30080 not P1_REIP_REG_17__SCAN_IN ; P1_R2096_U35
g30081 nand P1_R2096_U108 P1_REIP_REG_17__SCAN_IN ; P1_R2096_U36
g30082 not P1_REIP_REG_18__SCAN_IN ; P1_R2096_U37
g30083 nand P1_R2096_U109 P1_REIP_REG_18__SCAN_IN ; P1_R2096_U38
g30084 not P1_REIP_REG_19__SCAN_IN ; P1_R2096_U39
g30085 nand P1_R2096_U110 P1_REIP_REG_19__SCAN_IN ; P1_R2096_U40
g30086 not P1_REIP_REG_20__SCAN_IN ; P1_R2096_U41
g30087 nand P1_R2096_U111 P1_REIP_REG_20__SCAN_IN ; P1_R2096_U42
g30088 not P1_REIP_REG_21__SCAN_IN ; P1_R2096_U43
g30089 nand P1_R2096_U112 P1_REIP_REG_21__SCAN_IN ; P1_R2096_U44
g30090 not P1_REIP_REG_22__SCAN_IN ; P1_R2096_U45
g30091 nand P1_R2096_U113 P1_REIP_REG_22__SCAN_IN ; P1_R2096_U46
g30092 not P1_REIP_REG_23__SCAN_IN ; P1_R2096_U47
g30093 nand P1_R2096_U114 P1_REIP_REG_23__SCAN_IN ; P1_R2096_U48
g30094 not P1_REIP_REG_24__SCAN_IN ; P1_R2096_U49
g30095 nand P1_R2096_U115 P1_REIP_REG_24__SCAN_IN ; P1_R2096_U50
g30096 not P1_REIP_REG_25__SCAN_IN ; P1_R2096_U51
g30097 nand P1_R2096_U116 P1_REIP_REG_25__SCAN_IN ; P1_R2096_U52
g30098 not P1_REIP_REG_26__SCAN_IN ; P1_R2096_U53
g30099 nand P1_R2096_U117 P1_REIP_REG_26__SCAN_IN ; P1_R2096_U54
g30100 not P1_REIP_REG_27__SCAN_IN ; P1_R2096_U55
g30101 nand P1_R2096_U118 P1_REIP_REG_27__SCAN_IN ; P1_R2096_U56
g30102 not P1_REIP_REG_28__SCAN_IN ; P1_R2096_U57
g30103 nand P1_R2096_U119 P1_REIP_REG_28__SCAN_IN ; P1_R2096_U58
g30104 not P1_REIP_REG_29__SCAN_IN ; P1_R2096_U59
g30105 nand P1_R2096_U120 P1_REIP_REG_29__SCAN_IN ; P1_R2096_U60
g30106 not P1_REIP_REG_30__SCAN_IN ; P1_R2096_U61
g30107 nand P1_R2096_U124 P1_R2096_U123 ; P1_R2096_U62
g30108 nand P1_R2096_U126 P1_R2096_U125 ; P1_R2096_U63
g30109 nand P1_R2096_U128 P1_R2096_U127 ; P1_R2096_U64
g30110 nand P1_R2096_U130 P1_R2096_U129 ; P1_R2096_U65
g30111 nand P1_R2096_U132 P1_R2096_U131 ; P1_R2096_U66
g30112 nand P1_R2096_U134 P1_R2096_U133 ; P1_R2096_U67
g30113 nand P1_R2096_U136 P1_R2096_U135 ; P1_R2096_U68
g30114 nand P1_R2096_U138 P1_R2096_U137 ; P1_R2096_U69
g30115 nand P1_R2096_U140 P1_R2096_U139 ; P1_R2096_U70
g30116 nand P1_R2096_U142 P1_R2096_U141 ; P1_R2096_U71
g30117 nand P1_R2096_U144 P1_R2096_U143 ; P1_R2096_U72
g30118 nand P1_R2096_U146 P1_R2096_U145 ; P1_R2096_U73
g30119 nand P1_R2096_U148 P1_R2096_U147 ; P1_R2096_U74
g30120 nand P1_R2096_U150 P1_R2096_U149 ; P1_R2096_U75
g30121 nand P1_R2096_U152 P1_R2096_U151 ; P1_R2096_U76
g30122 nand P1_R2096_U154 P1_R2096_U153 ; P1_R2096_U77
g30123 nand P1_R2096_U156 P1_R2096_U155 ; P1_R2096_U78
g30124 nand P1_R2096_U158 P1_R2096_U157 ; P1_R2096_U79
g30125 nand P1_R2096_U160 P1_R2096_U159 ; P1_R2096_U80
g30126 nand P1_R2096_U162 P1_R2096_U161 ; P1_R2096_U81
g30127 nand P1_R2096_U164 P1_R2096_U163 ; P1_R2096_U82
g30128 nand P1_R2096_U166 P1_R2096_U165 ; P1_R2096_U83
g30129 nand P1_R2096_U168 P1_R2096_U167 ; P1_R2096_U84
g30130 nand P1_R2096_U170 P1_R2096_U169 ; P1_R2096_U85
g30131 nand P1_R2096_U172 P1_R2096_U171 ; P1_R2096_U86
g30132 nand P1_R2096_U174 P1_R2096_U173 ; P1_R2096_U87
g30133 nand P1_R2096_U176 P1_R2096_U175 ; P1_R2096_U88
g30134 nand P1_R2096_U178 P1_R2096_U177 ; P1_R2096_U89
g30135 nand P1_R2096_U180 P1_R2096_U179 ; P1_R2096_U90
g30136 nand P1_R2096_U182 P1_R2096_U181 ; P1_R2096_U91
g30137 not P1_REIP_REG_31__SCAN_IN ; P1_R2096_U92
g30138 nand P1_R2096_U121 P1_REIP_REG_30__SCAN_IN ; P1_R2096_U93
g30139 not P1_R2096_U6 ; P1_R2096_U94
g30140 not P1_R2096_U8 ; P1_R2096_U95
g30141 not P1_R2096_U10 ; P1_R2096_U96
g30142 not P1_R2096_U12 ; P1_R2096_U97
g30143 not P1_R2096_U14 ; P1_R2096_U98
g30144 not P1_R2096_U16 ; P1_R2096_U99
g30145 not P1_R2096_U19 ; P1_R2096_U100
g30146 not P1_R2096_U20 ; P1_R2096_U101
g30147 not P1_R2096_U22 ; P1_R2096_U102
g30148 not P1_R2096_U24 ; P1_R2096_U103
g30149 not P1_R2096_U26 ; P1_R2096_U104
g30150 not P1_R2096_U28 ; P1_R2096_U105
g30151 not P1_R2096_U30 ; P1_R2096_U106
g30152 not P1_R2096_U32 ; P1_R2096_U107
g30153 not P1_R2096_U34 ; P1_R2096_U108
g30154 not P1_R2096_U36 ; P1_R2096_U109
g30155 not P1_R2096_U38 ; P1_R2096_U110
g30156 not P1_R2096_U40 ; P1_R2096_U111
g30157 not P1_R2096_U42 ; P1_R2096_U112
g30158 not P1_R2096_U44 ; P1_R2096_U113
g30159 not P1_R2096_U46 ; P1_R2096_U114
g30160 not P1_R2096_U48 ; P1_R2096_U115
g30161 not P1_R2096_U50 ; P1_R2096_U116
g30162 not P1_R2096_U52 ; P1_R2096_U117
g30163 not P1_R2096_U54 ; P1_R2096_U118
g30164 not P1_R2096_U56 ; P1_R2096_U119
g30165 not P1_R2096_U58 ; P1_R2096_U120
g30166 not P1_R2096_U60 ; P1_R2096_U121
g30167 not P1_R2096_U93 ; P1_R2096_U122
g30168 nand P1_R2096_U19 P1_REIP_REG_9__SCAN_IN ; P1_R2096_U123
g30169 nand P1_R2096_U100 P1_R2096_U18 ; P1_R2096_U124
g30170 nand P1_R2096_U16 P1_REIP_REG_8__SCAN_IN ; P1_R2096_U125
g30171 nand P1_R2096_U99 P1_R2096_U17 ; P1_R2096_U126
g30172 nand P1_R2096_U14 P1_REIP_REG_7__SCAN_IN ; P1_R2096_U127
g30173 nand P1_R2096_U98 P1_R2096_U15 ; P1_R2096_U128
g30174 nand P1_R2096_U12 P1_REIP_REG_6__SCAN_IN ; P1_R2096_U129
g30175 nand P1_R2096_U97 P1_R2096_U13 ; P1_R2096_U130
g30176 nand P1_R2096_U10 P1_REIP_REG_5__SCAN_IN ; P1_R2096_U131
g30177 nand P1_R2096_U96 P1_R2096_U11 ; P1_R2096_U132
g30178 nand P1_R2096_U8 P1_REIP_REG_4__SCAN_IN ; P1_R2096_U133
g30179 nand P1_R2096_U95 P1_R2096_U9 ; P1_R2096_U134
g30180 nand P1_R2096_U6 P1_REIP_REG_3__SCAN_IN ; P1_R2096_U135
g30181 nand P1_R2096_U94 P1_R2096_U7 ; P1_R2096_U136
g30182 nand P1_R2096_U93 P1_REIP_REG_31__SCAN_IN ; P1_R2096_U137
g30183 nand P1_R2096_U122 P1_R2096_U92 ; P1_R2096_U138
g30184 nand P1_R2096_U60 P1_REIP_REG_30__SCAN_IN ; P1_R2096_U139
g30185 nand P1_R2096_U121 P1_R2096_U61 ; P1_R2096_U140
g30186 nand P1_R2096_U4 P1_REIP_REG_2__SCAN_IN ; P1_R2096_U141
g30187 nand P1_R2096_U5 P1_REIP_REG_1__SCAN_IN ; P1_R2096_U142
g30188 nand P1_R2096_U58 P1_REIP_REG_29__SCAN_IN ; P1_R2096_U143
g30189 nand P1_R2096_U120 P1_R2096_U59 ; P1_R2096_U144
g30190 nand P1_R2096_U56 P1_REIP_REG_28__SCAN_IN ; P1_R2096_U145
g30191 nand P1_R2096_U119 P1_R2096_U57 ; P1_R2096_U146
g30192 nand P1_R2096_U54 P1_REIP_REG_27__SCAN_IN ; P1_R2096_U147
g30193 nand P1_R2096_U118 P1_R2096_U55 ; P1_R2096_U148
g30194 nand P1_R2096_U52 P1_REIP_REG_26__SCAN_IN ; P1_R2096_U149
g30195 nand P1_R2096_U117 P1_R2096_U53 ; P1_R2096_U150
g30196 nand P1_R2096_U50 P1_REIP_REG_25__SCAN_IN ; P1_R2096_U151
g30197 nand P1_R2096_U116 P1_R2096_U51 ; P1_R2096_U152
g30198 nand P1_R2096_U48 P1_REIP_REG_24__SCAN_IN ; P1_R2096_U153
g30199 nand P1_R2096_U115 P1_R2096_U49 ; P1_R2096_U154
g30200 nand P1_R2096_U46 P1_REIP_REG_23__SCAN_IN ; P1_R2096_U155
g30201 nand P1_R2096_U114 P1_R2096_U47 ; P1_R2096_U156
g30202 nand P1_R2096_U44 P1_REIP_REG_22__SCAN_IN ; P1_R2096_U157
g30203 nand P1_R2096_U113 P1_R2096_U45 ; P1_R2096_U158
g30204 nand P1_R2096_U42 P1_REIP_REG_21__SCAN_IN ; P1_R2096_U159
g30205 nand P1_R2096_U112 P1_R2096_U43 ; P1_R2096_U160
g30206 nand P1_R2096_U40 P1_REIP_REG_20__SCAN_IN ; P1_R2096_U161
g30207 nand P1_R2096_U111 P1_R2096_U41 ; P1_R2096_U162
g30208 nand P1_R2096_U38 P1_REIP_REG_19__SCAN_IN ; P1_R2096_U163
g30209 nand P1_R2096_U110 P1_R2096_U39 ; P1_R2096_U164
g30210 nand P1_R2096_U36 P1_REIP_REG_18__SCAN_IN ; P1_R2096_U165
g30211 nand P1_R2096_U109 P1_R2096_U37 ; P1_R2096_U166
g30212 nand P1_R2096_U34 P1_REIP_REG_17__SCAN_IN ; P1_R2096_U167
g30213 nand P1_R2096_U108 P1_R2096_U35 ; P1_R2096_U168
g30214 nand P1_R2096_U32 P1_REIP_REG_16__SCAN_IN ; P1_R2096_U169
g30215 nand P1_R2096_U107 P1_R2096_U33 ; P1_R2096_U170
g30216 nand P1_R2096_U30 P1_REIP_REG_15__SCAN_IN ; P1_R2096_U171
g30217 nand P1_R2096_U106 P1_R2096_U31 ; P1_R2096_U172
g30218 nand P1_R2096_U28 P1_REIP_REG_14__SCAN_IN ; P1_R2096_U173
g30219 nand P1_R2096_U105 P1_R2096_U29 ; P1_R2096_U174
g30220 nand P1_R2096_U26 P1_REIP_REG_13__SCAN_IN ; P1_R2096_U175
g30221 nand P1_R2096_U104 P1_R2096_U27 ; P1_R2096_U176
g30222 nand P1_R2096_U24 P1_REIP_REG_12__SCAN_IN ; P1_R2096_U177
g30223 nand P1_R2096_U103 P1_R2096_U25 ; P1_R2096_U178
g30224 nand P1_R2096_U22 P1_REIP_REG_11__SCAN_IN ; P1_R2096_U179
g30225 nand P1_R2096_U102 P1_R2096_U23 ; P1_R2096_U180
g30226 nand P1_R2096_U20 P1_REIP_REG_10__SCAN_IN ; P1_R2096_U181
g30227 nand P1_R2096_U101 P1_R2096_U21 ; P1_R2096_U182
g30228 and P1_LT_563_U27 P1_LT_563_U26 ; P1_LT_563_U6
g30229 not P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_LT_563_U7
g30230 not P1_U3491 ; P1_LT_563_U8
g30231 not P1_U3490 ; P1_LT_563_U9
g30232 not P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_LT_563_U10
g30233 not P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_LT_563_U11
g30234 not P1_U3489 ; P1_LT_563_U12
g30235 and P1_LT_563_U21 P1_LT_563_U22 ; P1_LT_563_U13
g30236 and P1_LT_563_U24 P1_LT_563_U25 ; P1_LT_563_U14
g30237 not P1_U3492 ; P1_LT_563_U15
g30238 not P1_U3493 ; P1_LT_563_U16
g30239 nand P1_LT_563_U16 P1_LT_563_U15 P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_LT_563_U17
g30240 nand P1_LT_563_U15 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_LT_563_U18
g30241 nand P1_LT_563_U8 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_LT_563_U19
g30242 nand P1_LT_563_U28 P1_LT_563_U19 P1_LT_563_U18 P1_LT_563_U17 ; P1_LT_563_U20
g30243 nand P1_U3491 P1_LT_563_U7 ; P1_LT_563_U21
g30244 nand P1_U3490 P1_LT_563_U10 ; P1_LT_563_U22
g30245 nand P1_LT_563_U13 P1_LT_563_U20 ; P1_LT_563_U23
g30246 nand P1_LT_563_U9 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_LT_563_U24
g30247 nand P1_LT_563_U12 P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_LT_563_U25
g30248 nand P1_LT_563_U14 P1_LT_563_U23 ; P1_LT_563_U26
g30249 nand P1_U3489 P1_LT_563_U11 ; P1_LT_563_U27
g30250 nand P1_LT_563_U16 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_LT_563_U28
g30251 nand P1_R2238_U45 P1_R2238_U44 ; P1_R2238_U6
g30252 nand P1_R2238_U9 P1_R2238_U46 ; P1_R2238_U7
g30253 not P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_R2238_U8
g30254 nand P1_R2238_U18 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_R2238_U9
g30255 not P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_R2238_U10
g30256 not P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_R2238_U11
g30257 not P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_R2238_U12
g30258 not P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_R2238_U13
g30259 not P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_R2238_U14
g30260 not P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_R2238_U15
g30261 nand P1_R2238_U41 P1_R2238_U40 ; P1_R2238_U16
g30262 not P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_R2238_U17
g30263 not P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_R2238_U18
g30264 nand P1_R2238_U51 P1_R2238_U50 ; P1_R2238_U19
g30265 nand P1_R2238_U56 P1_R2238_U55 ; P1_R2238_U20
g30266 nand P1_R2238_U61 P1_R2238_U60 ; P1_R2238_U21
g30267 nand P1_R2238_U66 P1_R2238_U65 ; P1_R2238_U22
g30268 nand P1_R2238_U48 P1_R2238_U47 ; P1_R2238_U23
g30269 nand P1_R2238_U53 P1_R2238_U52 ; P1_R2238_U24
g30270 nand P1_R2238_U58 P1_R2238_U57 ; P1_R2238_U25
g30271 nand P1_R2238_U63 P1_R2238_U62 ; P1_R2238_U26
g30272 nand P1_R2238_U37 P1_R2238_U36 ; P1_R2238_U27
g30273 nand P1_R2238_U33 P1_R2238_U32 ; P1_R2238_U28
g30274 not P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_R2238_U29
g30275 not P1_R2238_U9 ; P1_R2238_U30
g30276 nand P1_R2238_U30 P1_R2238_U10 ; P1_R2238_U31
g30277 nand P1_R2238_U31 P1_R2238_U29 ; P1_R2238_U32
g30278 nand P1_R2238_U9 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_R2238_U33
g30279 not P1_R2238_U28 ; P1_R2238_U34
g30280 nand P1_R2238_U12 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_R2238_U35
g30281 nand P1_R2238_U35 P1_R2238_U28 ; P1_R2238_U36
g30282 nand P1_R2238_U11 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_R2238_U37
g30283 not P1_R2238_U27 ; P1_R2238_U38
g30284 nand P1_R2238_U14 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_R2238_U39
g30285 nand P1_R2238_U39 P1_R2238_U27 ; P1_R2238_U40
g30286 nand P1_R2238_U13 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_R2238_U41
g30287 not P1_R2238_U16 ; P1_R2238_U42
g30288 nand P1_R2238_U17 P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_R2238_U43
g30289 nand P1_R2238_U42 P1_R2238_U43 ; P1_R2238_U44
g30290 nand P1_R2238_U15 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_R2238_U45
g30291 nand P1_R2238_U8 P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_R2238_U46
g30292 nand P1_R2238_U15 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_R2238_U47
g30293 nand P1_R2238_U17 P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_R2238_U48
g30294 not P1_R2238_U23 ; P1_R2238_U49
g30295 nand P1_R2238_U49 P1_R2238_U42 ; P1_R2238_U50
g30296 nand P1_R2238_U23 P1_R2238_U16 ; P1_R2238_U51
g30297 nand P1_R2238_U14 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_R2238_U52
g30298 nand P1_R2238_U13 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_R2238_U53
g30299 not P1_R2238_U24 ; P1_R2238_U54
g30300 nand P1_R2238_U38 P1_R2238_U54 ; P1_R2238_U55
g30301 nand P1_R2238_U24 P1_R2238_U27 ; P1_R2238_U56
g30302 nand P1_R2238_U12 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_R2238_U57
g30303 nand P1_R2238_U11 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_R2238_U58
g30304 not P1_R2238_U25 ; P1_R2238_U59
g30305 nand P1_R2238_U34 P1_R2238_U59 ; P1_R2238_U60
g30306 nand P1_R2238_U25 P1_R2238_U28 ; P1_R2238_U61
g30307 nand P1_R2238_U10 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_R2238_U62
g30308 nand P1_R2238_U29 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_R2238_U63
g30309 not P1_R2238_U26 ; P1_R2238_U64
g30310 nand P1_R2238_U64 P1_R2238_U30 ; P1_R2238_U65
g30311 nand P1_R2238_U26 P1_R2238_U9 ; P1_R2238_U66
g30312 nand P1_SUB_450_U45 P1_SUB_450_U44 ; P1_SUB_450_U6
g30313 nand P1_SUB_450_U9 P1_SUB_450_U46 ; P1_SUB_450_U7
g30314 not P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_SUB_450_U8
g30315 nand P1_SUB_450_U18 P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN ; P1_SUB_450_U9
g30316 not P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_SUB_450_U10
g30317 not P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_SUB_450_U11
g30318 not P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_SUB_450_U12
g30319 not P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_SUB_450_U13
g30320 not P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_SUB_450_U14
g30321 not P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_SUB_450_U15
g30322 nand P1_SUB_450_U41 P1_SUB_450_U40 ; P1_SUB_450_U16
g30323 not P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_SUB_450_U17
g30324 not P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_SUB_450_U18
g30325 nand P1_SUB_450_U51 P1_SUB_450_U50 ; P1_SUB_450_U19
g30326 nand P1_SUB_450_U56 P1_SUB_450_U55 ; P1_SUB_450_U20
g30327 nand P1_SUB_450_U61 P1_SUB_450_U60 ; P1_SUB_450_U21
g30328 nand P1_SUB_450_U66 P1_SUB_450_U65 ; P1_SUB_450_U22
g30329 nand P1_SUB_450_U48 P1_SUB_450_U47 ; P1_SUB_450_U23
g30330 nand P1_SUB_450_U53 P1_SUB_450_U52 ; P1_SUB_450_U24
g30331 nand P1_SUB_450_U58 P1_SUB_450_U57 ; P1_SUB_450_U25
g30332 nand P1_SUB_450_U63 P1_SUB_450_U62 ; P1_SUB_450_U26
g30333 nand P1_SUB_450_U37 P1_SUB_450_U36 ; P1_SUB_450_U27
g30334 nand P1_SUB_450_U33 P1_SUB_450_U32 ; P1_SUB_450_U28
g30335 not P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_SUB_450_U29
g30336 not P1_SUB_450_U9 ; P1_SUB_450_U30
g30337 nand P1_SUB_450_U30 P1_SUB_450_U10 ; P1_SUB_450_U31
g30338 nand P1_SUB_450_U31 P1_SUB_450_U29 ; P1_SUB_450_U32
g30339 nand P1_SUB_450_U9 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_SUB_450_U33
g30340 not P1_SUB_450_U28 ; P1_SUB_450_U34
g30341 nand P1_SUB_450_U12 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_SUB_450_U35
g30342 nand P1_SUB_450_U35 P1_SUB_450_U28 ; P1_SUB_450_U36
g30343 nand P1_SUB_450_U11 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_SUB_450_U37
g30344 not P1_SUB_450_U27 ; P1_SUB_450_U38
g30345 nand P1_SUB_450_U14 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_SUB_450_U39
g30346 nand P1_SUB_450_U39 P1_SUB_450_U27 ; P1_SUB_450_U40
g30347 nand P1_SUB_450_U13 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_SUB_450_U41
g30348 not P1_SUB_450_U16 ; P1_SUB_450_U42
g30349 nand P1_SUB_450_U17 P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_SUB_450_U43
g30350 nand P1_SUB_450_U42 P1_SUB_450_U43 ; P1_SUB_450_U44
g30351 nand P1_SUB_450_U15 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_SUB_450_U45
g30352 nand P1_SUB_450_U8 P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; P1_SUB_450_U46
g30353 nand P1_SUB_450_U15 P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN ; P1_SUB_450_U47
g30354 nand P1_SUB_450_U17 P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; P1_SUB_450_U48
g30355 not P1_SUB_450_U23 ; P1_SUB_450_U49
g30356 nand P1_SUB_450_U49 P1_SUB_450_U42 ; P1_SUB_450_U50
g30357 nand P1_SUB_450_U23 P1_SUB_450_U16 ; P1_SUB_450_U51
g30358 nand P1_SUB_450_U14 P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN ; P1_SUB_450_U52
g30359 nand P1_SUB_450_U13 P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; P1_SUB_450_U53
g30360 not P1_SUB_450_U24 ; P1_SUB_450_U54
g30361 nand P1_SUB_450_U38 P1_SUB_450_U54 ; P1_SUB_450_U55
g30362 nand P1_SUB_450_U24 P1_SUB_450_U27 ; P1_SUB_450_U56
g30363 nand P1_SUB_450_U12 P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN ; P1_SUB_450_U57
g30364 nand P1_SUB_450_U11 P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; P1_SUB_450_U58
g30365 not P1_SUB_450_U25 ; P1_SUB_450_U59
g30366 nand P1_SUB_450_U34 P1_SUB_450_U59 ; P1_SUB_450_U60
g30367 nand P1_SUB_450_U25 P1_SUB_450_U28 ; P1_SUB_450_U61
g30368 nand P1_SUB_450_U10 P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN ; P1_SUB_450_U62
g30369 nand P1_SUB_450_U29 P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; P1_SUB_450_U63
g30370 not P1_SUB_450_U26 ; P1_SUB_450_U64
g30371 nand P1_SUB_450_U64 P1_SUB_450_U30 ; P1_SUB_450_U65
g30372 nand P1_SUB_450_U26 P1_SUB_450_U9 ; P1_SUB_450_U66
g30373 not P1_U3227 ; P1_ADD_371_U4
g30374 nand P1_ADD_371_U23 P1_ADD_371_U31 ; P1_ADD_371_U5
g30375 and P1_ADD_371_U22 P1_ADD_371_U30 ; P1_ADD_371_U6
g30376 not P1_U3228 ; P1_ADD_371_U7
g30377 not P1_U3230 ; P1_ADD_371_U8
g30378 nand P1_U3230 P1_ADD_371_U23 ; P1_ADD_371_U9
g30379 not P1_U3231 ; P1_ADD_371_U10
g30380 nand P1_U3231 P1_ADD_371_U28 ; P1_ADD_371_U11
g30381 not P1_U3232 ; P1_ADD_371_U12
g30382 not P1_U3233 ; P1_ADD_371_U13
g30383 nand P1_U3232 P1_ADD_371_U29 ; P1_ADD_371_U14
g30384 not P1_U3229 ; P1_ADD_371_U15
g30385 not P1_U3234 ; P1_ADD_371_U16
g30386 nand P1_ADD_371_U34 P1_ADD_371_U33 ; P1_ADD_371_U17
g30387 nand P1_ADD_371_U36 P1_ADD_371_U35 ; P1_ADD_371_U18
g30388 nand P1_ADD_371_U38 P1_ADD_371_U37 ; P1_ADD_371_U19
g30389 nand P1_ADD_371_U42 P1_ADD_371_U41 ; P1_ADD_371_U20
g30390 nand P1_ADD_371_U44 P1_ADD_371_U43 ; P1_ADD_371_U21
g30391 and P1_U3234 P1_U3233 ; P1_ADD_371_U22
g30392 nand P1_ADD_371_U15 P1_ADD_371_U26 ; P1_ADD_371_U23
g30393 and P1_ADD_371_U40 P1_ADD_371_U39 ; P1_ADD_371_U24
g30394 nand P1_ADD_371_U30 P1_U3233 ; P1_ADD_371_U25
g30395 nand P1_U3228 P1_U3227 ; P1_ADD_371_U26
g30396 not P1_ADD_371_U23 ; P1_ADD_371_U27
g30397 not P1_ADD_371_U9 ; P1_ADD_371_U28
g30398 not P1_ADD_371_U11 ; P1_ADD_371_U29
g30399 not P1_ADD_371_U14 ; P1_ADD_371_U30
g30400 nand P1_U3228 P1_U3227 P1_U3229 ; P1_ADD_371_U31
g30401 not P1_ADD_371_U25 ; P1_ADD_371_U32
g30402 nand P1_U3233 P1_ADD_371_U14 ; P1_ADD_371_U33
g30403 nand P1_ADD_371_U30 P1_ADD_371_U13 ; P1_ADD_371_U34
g30404 nand P1_U3231 P1_ADD_371_U9 ; P1_ADD_371_U35
g30405 nand P1_ADD_371_U28 P1_ADD_371_U10 ; P1_ADD_371_U36
g30406 nand P1_U3232 P1_ADD_371_U11 ; P1_ADD_371_U37
g30407 nand P1_ADD_371_U29 P1_ADD_371_U12 ; P1_ADD_371_U38
g30408 nand P1_U3230 P1_ADD_371_U23 ; P1_ADD_371_U39
g30409 nand P1_ADD_371_U27 P1_ADD_371_U8 ; P1_ADD_371_U40
g30410 nand P1_U3228 P1_ADD_371_U4 ; P1_ADD_371_U41
g30411 nand P1_U3227 P1_ADD_371_U7 ; P1_ADD_371_U42
g30412 nand P1_U3234 P1_ADD_371_U25 ; P1_ADD_371_U43
g30413 nand P1_ADD_371_U32 P1_ADD_371_U16 ; P1_ADD_371_U44
g30414 not P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_ADD_405_U4
g30415 nand P1_ADD_405_U94 P1_ADD_405_U125 ; P1_ADD_405_U5
g30416 not P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_ADD_405_U6
g30417 not P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_ADD_405_U7
g30418 nand P1_ADD_405_U94 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_ADD_405_U8
g30419 not P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_ADD_405_U9
g30420 nand P1_ADD_405_U98 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_ADD_405_U10
g30421 not P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_ADD_405_U11
g30422 not P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_ADD_405_U12
g30423 nand P1_ADD_405_U99 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_ADD_405_U13
g30424 nand P1_ADD_405_U100 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_ADD_405_U14
g30425 not P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_ADD_405_U15
g30426 nand P1_ADD_405_U101 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_ADD_405_U16
g30427 not P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_ADD_405_U17
g30428 nand P1_ADD_405_U102 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_ADD_405_U18
g30429 not P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_ADD_405_U19
g30430 nand P1_ADD_405_U103 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_ADD_405_U20
g30431 not P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_ADD_405_U21
g30432 nand P1_ADD_405_U104 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_ADD_405_U22
g30433 not P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_ADD_405_U23
g30434 nand P1_ADD_405_U105 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_ADD_405_U24
g30435 not P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_ADD_405_U25
g30436 nand P1_ADD_405_U106 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_ADD_405_U26
g30437 not P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_ADD_405_U27
g30438 nand P1_ADD_405_U107 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_ADD_405_U28
g30439 not P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_ADD_405_U29
g30440 nand P1_ADD_405_U108 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_ADD_405_U30
g30441 not P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_ADD_405_U31
g30442 nand P1_ADD_405_U109 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_ADD_405_U32
g30443 not P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_ADD_405_U33
g30444 nand P1_ADD_405_U110 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_ADD_405_U34
g30445 not P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_ADD_405_U35
g30446 nand P1_ADD_405_U111 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_ADD_405_U36
g30447 not P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_ADD_405_U37
g30448 nand P1_ADD_405_U112 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_ADD_405_U38
g30449 not P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_ADD_405_U39
g30450 nand P1_ADD_405_U113 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_ADD_405_U40
g30451 not P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_ADD_405_U41
g30452 nand P1_ADD_405_U114 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_ADD_405_U42
g30453 not P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_ADD_405_U43
g30454 nand P1_ADD_405_U115 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_ADD_405_U44
g30455 not P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_ADD_405_U45
g30456 nand P1_ADD_405_U116 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_ADD_405_U46
g30457 not P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_ADD_405_U47
g30458 nand P1_ADD_405_U117 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_ADD_405_U48
g30459 not P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_ADD_405_U49
g30460 nand P1_ADD_405_U118 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_ADD_405_U50
g30461 not P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_ADD_405_U51
g30462 nand P1_ADD_405_U119 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_ADD_405_U52
g30463 not P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_ADD_405_U53
g30464 nand P1_ADD_405_U120 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_ADD_405_U54
g30465 not P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_ADD_405_U55
g30466 nand P1_ADD_405_U121 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_ADD_405_U56
g30467 not P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_ADD_405_U57
g30468 nand P1_ADD_405_U122 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_ADD_405_U58
g30469 not P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_ADD_405_U59
g30470 not P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_ADD_405_U60
g30471 nand P1_ADD_405_U123 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_ADD_405_U61
g30472 not P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_ADD_405_U62
g30473 nand P1_ADD_405_U128 P1_ADD_405_U127 ; P1_ADD_405_U63
g30474 nand P1_ADD_405_U130 P1_ADD_405_U129 ; P1_ADD_405_U64
g30475 nand P1_ADD_405_U132 P1_ADD_405_U131 ; P1_ADD_405_U65
g30476 nand P1_ADD_405_U134 P1_ADD_405_U133 ; P1_ADD_405_U66
g30477 nand P1_ADD_405_U136 P1_ADD_405_U135 ; P1_ADD_405_U67
g30478 nand P1_ADD_405_U138 P1_ADD_405_U137 ; P1_ADD_405_U68
g30479 nand P1_ADD_405_U140 P1_ADD_405_U139 ; P1_ADD_405_U69
g30480 nand P1_ADD_405_U142 P1_ADD_405_U141 ; P1_ADD_405_U70
g30481 nand P1_ADD_405_U144 P1_ADD_405_U143 ; P1_ADD_405_U71
g30482 nand P1_ADD_405_U146 P1_ADD_405_U145 ; P1_ADD_405_U72
g30483 nand P1_ADD_405_U148 P1_ADD_405_U147 ; P1_ADD_405_U73
g30484 nand P1_ADD_405_U150 P1_ADD_405_U149 ; P1_ADD_405_U74
g30485 nand P1_ADD_405_U152 P1_ADD_405_U151 ; P1_ADD_405_U75
g30486 nand P1_ADD_405_U154 P1_ADD_405_U153 ; P1_ADD_405_U76
g30487 nand P1_ADD_405_U156 P1_ADD_405_U155 ; P1_ADD_405_U77
g30488 nand P1_ADD_405_U158 P1_ADD_405_U157 ; P1_ADD_405_U78
g30489 nand P1_ADD_405_U160 P1_ADD_405_U159 ; P1_ADD_405_U79
g30490 nand P1_ADD_405_U162 P1_ADD_405_U161 ; P1_ADD_405_U80
g30491 nand P1_ADD_405_U164 P1_ADD_405_U163 ; P1_ADD_405_U81
g30492 nand P1_ADD_405_U166 P1_ADD_405_U165 ; P1_ADD_405_U82
g30493 nand P1_ADD_405_U168 P1_ADD_405_U167 ; P1_ADD_405_U83
g30494 nand P1_ADD_405_U170 P1_ADD_405_U169 ; P1_ADD_405_U84
g30495 nand P1_ADD_405_U174 P1_ADD_405_U173 ; P1_ADD_405_U85
g30496 nand P1_ADD_405_U176 P1_ADD_405_U175 ; P1_ADD_405_U86
g30497 nand P1_ADD_405_U178 P1_ADD_405_U177 ; P1_ADD_405_U87
g30498 nand P1_ADD_405_U180 P1_ADD_405_U179 ; P1_ADD_405_U88
g30499 nand P1_ADD_405_U182 P1_ADD_405_U181 ; P1_ADD_405_U89
g30500 nand P1_ADD_405_U184 P1_ADD_405_U183 ; P1_ADD_405_U90
g30501 nand P1_ADD_405_U186 P1_ADD_405_U185 ; P1_ADD_405_U91
g30502 not P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_ADD_405_U92
g30503 nand P1_ADD_405_U124 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_ADD_405_U93
g30504 nand P1_ADD_405_U62 P1_ADD_405_U96 ; P1_ADD_405_U94
g30505 and P1_ADD_405_U172 P1_ADD_405_U171 ; P1_ADD_405_U95
g30506 nand P1_INSTADDRPOINTER_REG_0__SCAN_IN P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_ADD_405_U96
g30507 not P1_ADD_405_U94 ; P1_ADD_405_U97
g30508 not P1_ADD_405_U8 ; P1_ADD_405_U98
g30509 not P1_ADD_405_U10 ; P1_ADD_405_U99
g30510 not P1_ADD_405_U13 ; P1_ADD_405_U100
g30511 not P1_ADD_405_U14 ; P1_ADD_405_U101
g30512 not P1_ADD_405_U16 ; P1_ADD_405_U102
g30513 not P1_ADD_405_U18 ; P1_ADD_405_U103
g30514 not P1_ADD_405_U20 ; P1_ADD_405_U104
g30515 not P1_ADD_405_U22 ; P1_ADD_405_U105
g30516 not P1_ADD_405_U24 ; P1_ADD_405_U106
g30517 not P1_ADD_405_U26 ; P1_ADD_405_U107
g30518 not P1_ADD_405_U28 ; P1_ADD_405_U108
g30519 not P1_ADD_405_U30 ; P1_ADD_405_U109
g30520 not P1_ADD_405_U32 ; P1_ADD_405_U110
g30521 not P1_ADD_405_U34 ; P1_ADD_405_U111
g30522 not P1_ADD_405_U36 ; P1_ADD_405_U112
g30523 not P1_ADD_405_U38 ; P1_ADD_405_U113
g30524 not P1_ADD_405_U40 ; P1_ADD_405_U114
g30525 not P1_ADD_405_U42 ; P1_ADD_405_U115
g30526 not P1_ADD_405_U44 ; P1_ADD_405_U116
g30527 not P1_ADD_405_U46 ; P1_ADD_405_U117
g30528 not P1_ADD_405_U48 ; P1_ADD_405_U118
g30529 not P1_ADD_405_U50 ; P1_ADD_405_U119
g30530 not P1_ADD_405_U52 ; P1_ADD_405_U120
g30531 not P1_ADD_405_U54 ; P1_ADD_405_U121
g30532 not P1_ADD_405_U56 ; P1_ADD_405_U122
g30533 not P1_ADD_405_U58 ; P1_ADD_405_U123
g30534 not P1_ADD_405_U61 ; P1_ADD_405_U124
g30535 nand P1_INSTADDRPOINTER_REG_0__SCAN_IN P1_INSTADDRPOINTER_REG_1__SCAN_IN P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_ADD_405_U125
g30536 not P1_ADD_405_U93 ; P1_ADD_405_U126
g30537 nand P1_ADD_405_U13 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_ADD_405_U127
g30538 nand P1_ADD_405_U100 P1_ADD_405_U12 ; P1_ADD_405_U128
g30539 nand P1_ADD_405_U61 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_ADD_405_U129
g30540 nand P1_ADD_405_U124 P1_ADD_405_U60 ; P1_ADD_405_U130
g30541 nand P1_ADD_405_U58 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_ADD_405_U131
g30542 nand P1_ADD_405_U123 P1_ADD_405_U59 ; P1_ADD_405_U132
g30543 nand P1_ADD_405_U48 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_ADD_405_U133
g30544 nand P1_ADD_405_U118 P1_ADD_405_U49 ; P1_ADD_405_U134
g30545 nand P1_ADD_405_U34 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_ADD_405_U135
g30546 nand P1_ADD_405_U111 P1_ADD_405_U35 ; P1_ADD_405_U136
g30547 nand P1_ADD_405_U40 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_ADD_405_U137
g30548 nand P1_ADD_405_U114 P1_ADD_405_U41 ; P1_ADD_405_U138
g30549 nand P1_ADD_405_U26 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_ADD_405_U139
g30550 nand P1_ADD_405_U107 P1_ADD_405_U27 ; P1_ADD_405_U140
g30551 nand P1_ADD_405_U18 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_ADD_405_U141
g30552 nand P1_ADD_405_U103 P1_ADD_405_U19 ; P1_ADD_405_U142
g30553 nand P1_ADD_405_U44 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_ADD_405_U143
g30554 nand P1_ADD_405_U116 P1_ADD_405_U45 ; P1_ADD_405_U144
g30555 nand P1_ADD_405_U36 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_ADD_405_U145
g30556 nand P1_ADD_405_U112 P1_ADD_405_U37 ; P1_ADD_405_U146
g30557 nand P1_ADD_405_U22 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_ADD_405_U147
g30558 nand P1_ADD_405_U105 P1_ADD_405_U23 ; P1_ADD_405_U148
g30559 nand P1_ADD_405_U52 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_ADD_405_U149
g30560 nand P1_ADD_405_U120 P1_ADD_405_U53 ; P1_ADD_405_U150
g30561 nand P1_ADD_405_U30 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_ADD_405_U151
g30562 nand P1_ADD_405_U109 P1_ADD_405_U31 ; P1_ADD_405_U152
g30563 nand P1_ADD_405_U8 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_ADD_405_U153
g30564 nand P1_ADD_405_U98 P1_ADD_405_U9 ; P1_ADD_405_U154
g30565 nand P1_ADD_405_U54 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_ADD_405_U155
g30566 nand P1_ADD_405_U121 P1_ADD_405_U55 ; P1_ADD_405_U156
g30567 nand P1_ADD_405_U28 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_ADD_405_U157
g30568 nand P1_ADD_405_U108 P1_ADD_405_U29 ; P1_ADD_405_U158
g30569 nand P1_ADD_405_U10 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_ADD_405_U159
g30570 nand P1_ADD_405_U99 P1_ADD_405_U11 ; P1_ADD_405_U160
g30571 nand P1_ADD_405_U16 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_ADD_405_U161
g30572 nand P1_ADD_405_U102 P1_ADD_405_U17 ; P1_ADD_405_U162
g30573 nand P1_ADD_405_U46 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_ADD_405_U163
g30574 nand P1_ADD_405_U117 P1_ADD_405_U47 ; P1_ADD_405_U164
g30575 nand P1_ADD_405_U38 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_ADD_405_U165
g30576 nand P1_ADD_405_U113 P1_ADD_405_U39 ; P1_ADD_405_U166
g30577 nand P1_ADD_405_U20 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_ADD_405_U167
g30578 nand P1_ADD_405_U104 P1_ADD_405_U21 ; P1_ADD_405_U168
g30579 nand P1_ADD_405_U93 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_ADD_405_U169
g30580 nand P1_ADD_405_U126 P1_ADD_405_U92 ; P1_ADD_405_U170
g30581 nand P1_ADD_405_U94 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_ADD_405_U171
g30582 nand P1_ADD_405_U97 P1_ADD_405_U7 ; P1_ADD_405_U172
g30583 nand P1_ADD_405_U4 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_ADD_405_U173
g30584 nand P1_ADD_405_U6 P1_INSTADDRPOINTER_REG_0__SCAN_IN ; P1_ADD_405_U174
g30585 nand P1_ADD_405_U56 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_ADD_405_U175
g30586 nand P1_ADD_405_U122 P1_ADD_405_U57 ; P1_ADD_405_U176
g30587 nand P1_ADD_405_U42 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_ADD_405_U177
g30588 nand P1_ADD_405_U115 P1_ADD_405_U43 ; P1_ADD_405_U178
g30589 nand P1_ADD_405_U24 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_ADD_405_U179
g30590 nand P1_ADD_405_U106 P1_ADD_405_U25 ; P1_ADD_405_U180
g30591 nand P1_ADD_405_U14 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_ADD_405_U181
g30592 nand P1_ADD_405_U101 P1_ADD_405_U15 ; P1_ADD_405_U182
g30593 nand P1_ADD_405_U50 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_ADD_405_U183
g30594 nand P1_ADD_405_U119 P1_ADD_405_U51 ; P1_ADD_405_U184
g30595 nand P1_ADD_405_U32 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_ADD_405_U185
g30596 nand P1_ADD_405_U110 P1_ADD_405_U33 ; P1_ADD_405_U186
g30597 nor P1_R2238_U6 P1_GTE_485_U7 ; P1_GTE_485_U6
g30598 nor P1_R2238_U19 P1_R2238_U20 P1_R2238_U22 P1_R2238_U21 ; P1_GTE_485_U7
g30599 not P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_ADD_515_U4
g30600 not P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_ADD_515_U5
g30601 nand P1_INSTADDRPOINTER_REG_1__SCAN_IN P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_ADD_515_U6
g30602 not P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_ADD_515_U7
g30603 nand P1_ADD_515_U94 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_ADD_515_U8
g30604 not P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_ADD_515_U9
g30605 nand P1_ADD_515_U95 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_ADD_515_U10
g30606 not P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_ADD_515_U11
g30607 not P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_ADD_515_U12
g30608 nand P1_ADD_515_U96 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_ADD_515_U13
g30609 nand P1_ADD_515_U97 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_ADD_515_U14
g30610 not P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_ADD_515_U15
g30611 nand P1_ADD_515_U98 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_ADD_515_U16
g30612 not P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_ADD_515_U17
g30613 nand P1_ADD_515_U99 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_ADD_515_U18
g30614 not P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_ADD_515_U19
g30615 nand P1_ADD_515_U100 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_ADD_515_U20
g30616 not P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_ADD_515_U21
g30617 nand P1_ADD_515_U101 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_ADD_515_U22
g30618 not P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_ADD_515_U23
g30619 nand P1_ADD_515_U102 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_ADD_515_U24
g30620 not P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_ADD_515_U25
g30621 nand P1_ADD_515_U103 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_ADD_515_U26
g30622 not P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_ADD_515_U27
g30623 nand P1_ADD_515_U104 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_ADD_515_U28
g30624 not P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_ADD_515_U29
g30625 nand P1_ADD_515_U105 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_ADD_515_U30
g30626 not P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_ADD_515_U31
g30627 nand P1_ADD_515_U106 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_ADD_515_U32
g30628 not P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_ADD_515_U33
g30629 nand P1_ADD_515_U107 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_ADD_515_U34
g30630 not P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_ADD_515_U35
g30631 nand P1_ADD_515_U108 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_ADD_515_U36
g30632 not P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_ADD_515_U37
g30633 nand P1_ADD_515_U109 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_ADD_515_U38
g30634 not P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_ADD_515_U39
g30635 nand P1_ADD_515_U110 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_ADD_515_U40
g30636 not P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_ADD_515_U41
g30637 nand P1_ADD_515_U111 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_ADD_515_U42
g30638 not P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_ADD_515_U43
g30639 nand P1_ADD_515_U112 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_ADD_515_U44
g30640 not P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_ADD_515_U45
g30641 nand P1_ADD_515_U113 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_ADD_515_U46
g30642 not P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_ADD_515_U47
g30643 nand P1_ADD_515_U114 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_ADD_515_U48
g30644 not P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_ADD_515_U49
g30645 nand P1_ADD_515_U115 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_ADD_515_U50
g30646 not P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_ADD_515_U51
g30647 nand P1_ADD_515_U116 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_ADD_515_U52
g30648 not P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_ADD_515_U53
g30649 nand P1_ADD_515_U117 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_ADD_515_U54
g30650 not P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_ADD_515_U55
g30651 nand P1_ADD_515_U118 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_ADD_515_U56
g30652 not P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_ADD_515_U57
g30653 nand P1_ADD_515_U119 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_ADD_515_U58
g30654 not P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_ADD_515_U59
g30655 not P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_ADD_515_U60
g30656 nand P1_ADD_515_U120 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_ADD_515_U61
g30657 nand P1_ADD_515_U124 P1_ADD_515_U123 ; P1_ADD_515_U62
g30658 nand P1_ADD_515_U126 P1_ADD_515_U125 ; P1_ADD_515_U63
g30659 nand P1_ADD_515_U128 P1_ADD_515_U127 ; P1_ADD_515_U64
g30660 nand P1_ADD_515_U130 P1_ADD_515_U129 ; P1_ADD_515_U65
g30661 nand P1_ADD_515_U132 P1_ADD_515_U131 ; P1_ADD_515_U66
g30662 nand P1_ADD_515_U134 P1_ADD_515_U133 ; P1_ADD_515_U67
g30663 nand P1_ADD_515_U136 P1_ADD_515_U135 ; P1_ADD_515_U68
g30664 nand P1_ADD_515_U138 P1_ADD_515_U137 ; P1_ADD_515_U69
g30665 nand P1_ADD_515_U140 P1_ADD_515_U139 ; P1_ADD_515_U70
g30666 nand P1_ADD_515_U142 P1_ADD_515_U141 ; P1_ADD_515_U71
g30667 nand P1_ADD_515_U144 P1_ADD_515_U143 ; P1_ADD_515_U72
g30668 nand P1_ADD_515_U146 P1_ADD_515_U145 ; P1_ADD_515_U73
g30669 nand P1_ADD_515_U148 P1_ADD_515_U147 ; P1_ADD_515_U74
g30670 nand P1_ADD_515_U150 P1_ADD_515_U149 ; P1_ADD_515_U75
g30671 nand P1_ADD_515_U152 P1_ADD_515_U151 ; P1_ADD_515_U76
g30672 nand P1_ADD_515_U154 P1_ADD_515_U153 ; P1_ADD_515_U77
g30673 nand P1_ADD_515_U156 P1_ADD_515_U155 ; P1_ADD_515_U78
g30674 nand P1_ADD_515_U158 P1_ADD_515_U157 ; P1_ADD_515_U79
g30675 nand P1_ADD_515_U160 P1_ADD_515_U159 ; P1_ADD_515_U80
g30676 nand P1_ADD_515_U162 P1_ADD_515_U161 ; P1_ADD_515_U81
g30677 nand P1_ADD_515_U164 P1_ADD_515_U163 ; P1_ADD_515_U82
g30678 nand P1_ADD_515_U166 P1_ADD_515_U165 ; P1_ADD_515_U83
g30679 nand P1_ADD_515_U168 P1_ADD_515_U167 ; P1_ADD_515_U84
g30680 nand P1_ADD_515_U170 P1_ADD_515_U169 ; P1_ADD_515_U85
g30681 nand P1_ADD_515_U172 P1_ADD_515_U171 ; P1_ADD_515_U86
g30682 nand P1_ADD_515_U174 P1_ADD_515_U173 ; P1_ADD_515_U87
g30683 nand P1_ADD_515_U176 P1_ADD_515_U175 ; P1_ADD_515_U88
g30684 nand P1_ADD_515_U178 P1_ADD_515_U177 ; P1_ADD_515_U89
g30685 nand P1_ADD_515_U180 P1_ADD_515_U179 ; P1_ADD_515_U90
g30686 nand P1_ADD_515_U182 P1_ADD_515_U181 ; P1_ADD_515_U91
g30687 not P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_ADD_515_U92
g30688 nand P1_ADD_515_U121 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_ADD_515_U93
g30689 not P1_ADD_515_U6 ; P1_ADD_515_U94
g30690 not P1_ADD_515_U8 ; P1_ADD_515_U95
g30691 not P1_ADD_515_U10 ; P1_ADD_515_U96
g30692 not P1_ADD_515_U13 ; P1_ADD_515_U97
g30693 not P1_ADD_515_U14 ; P1_ADD_515_U98
g30694 not P1_ADD_515_U16 ; P1_ADD_515_U99
g30695 not P1_ADD_515_U18 ; P1_ADD_515_U100
g30696 not P1_ADD_515_U20 ; P1_ADD_515_U101
g30697 not P1_ADD_515_U22 ; P1_ADD_515_U102
g30698 not P1_ADD_515_U24 ; P1_ADD_515_U103
g30699 not P1_ADD_515_U26 ; P1_ADD_515_U104
g30700 not P1_ADD_515_U28 ; P1_ADD_515_U105
g30701 not P1_ADD_515_U30 ; P1_ADD_515_U106
g30702 not P1_ADD_515_U32 ; P1_ADD_515_U107
g30703 not P1_ADD_515_U34 ; P1_ADD_515_U108
g30704 not P1_ADD_515_U36 ; P1_ADD_515_U109
g30705 not P1_ADD_515_U38 ; P1_ADD_515_U110
g30706 not P1_ADD_515_U40 ; P1_ADD_515_U111
g30707 not P1_ADD_515_U42 ; P1_ADD_515_U112
g30708 not P1_ADD_515_U44 ; P1_ADD_515_U113
g30709 not P1_ADD_515_U46 ; P1_ADD_515_U114
g30710 not P1_ADD_515_U48 ; P1_ADD_515_U115
g30711 not P1_ADD_515_U50 ; P1_ADD_515_U116
g30712 not P1_ADD_515_U52 ; P1_ADD_515_U117
g30713 not P1_ADD_515_U54 ; P1_ADD_515_U118
g30714 not P1_ADD_515_U56 ; P1_ADD_515_U119
g30715 not P1_ADD_515_U58 ; P1_ADD_515_U120
g30716 not P1_ADD_515_U61 ; P1_ADD_515_U121
g30717 not P1_ADD_515_U93 ; P1_ADD_515_U122
g30718 nand P1_ADD_515_U13 P1_INSTADDRPOINTER_REG_6__SCAN_IN ; P1_ADD_515_U123
g30719 nand P1_ADD_515_U97 P1_ADD_515_U12 ; P1_ADD_515_U124
g30720 nand P1_ADD_515_U61 P1_INSTADDRPOINTER_REG_30__SCAN_IN ; P1_ADD_515_U125
g30721 nand P1_ADD_515_U121 P1_ADD_515_U60 ; P1_ADD_515_U126
g30722 nand P1_ADD_515_U58 P1_INSTADDRPOINTER_REG_29__SCAN_IN ; P1_ADD_515_U127
g30723 nand P1_ADD_515_U120 P1_ADD_515_U59 ; P1_ADD_515_U128
g30724 nand P1_ADD_515_U48 P1_INSTADDRPOINTER_REG_24__SCAN_IN ; P1_ADD_515_U129
g30725 nand P1_ADD_515_U115 P1_ADD_515_U49 ; P1_ADD_515_U130
g30726 nand P1_ADD_515_U34 P1_INSTADDRPOINTER_REG_17__SCAN_IN ; P1_ADD_515_U131
g30727 nand P1_ADD_515_U108 P1_ADD_515_U35 ; P1_ADD_515_U132
g30728 nand P1_ADD_515_U4 P1_INSTADDRPOINTER_REG_2__SCAN_IN ; P1_ADD_515_U133
g30729 nand P1_ADD_515_U5 P1_INSTADDRPOINTER_REG_1__SCAN_IN ; P1_ADD_515_U134
g30730 nand P1_ADD_515_U40 P1_INSTADDRPOINTER_REG_20__SCAN_IN ; P1_ADD_515_U135
g30731 nand P1_ADD_515_U111 P1_ADD_515_U41 ; P1_ADD_515_U136
g30732 nand P1_ADD_515_U26 P1_INSTADDRPOINTER_REG_13__SCAN_IN ; P1_ADD_515_U137
g30733 nand P1_ADD_515_U104 P1_ADD_515_U27 ; P1_ADD_515_U138
g30734 nand P1_ADD_515_U18 P1_INSTADDRPOINTER_REG_9__SCAN_IN ; P1_ADD_515_U139
g30735 nand P1_ADD_515_U100 P1_ADD_515_U19 ; P1_ADD_515_U140
g30736 nand P1_ADD_515_U44 P1_INSTADDRPOINTER_REG_22__SCAN_IN ; P1_ADD_515_U141
g30737 nand P1_ADD_515_U113 P1_ADD_515_U45 ; P1_ADD_515_U142
g30738 nand P1_ADD_515_U36 P1_INSTADDRPOINTER_REG_18__SCAN_IN ; P1_ADD_515_U143
g30739 nand P1_ADD_515_U109 P1_ADD_515_U37 ; P1_ADD_515_U144
g30740 nand P1_ADD_515_U22 P1_INSTADDRPOINTER_REG_11__SCAN_IN ; P1_ADD_515_U145
g30741 nand P1_ADD_515_U102 P1_ADD_515_U23 ; P1_ADD_515_U146
g30742 nand P1_ADD_515_U52 P1_INSTADDRPOINTER_REG_26__SCAN_IN ; P1_ADD_515_U147
g30743 nand P1_ADD_515_U117 P1_ADD_515_U53 ; P1_ADD_515_U148
g30744 nand P1_ADD_515_U30 P1_INSTADDRPOINTER_REG_15__SCAN_IN ; P1_ADD_515_U149
g30745 nand P1_ADD_515_U106 P1_ADD_515_U31 ; P1_ADD_515_U150
g30746 nand P1_ADD_515_U8 P1_INSTADDRPOINTER_REG_4__SCAN_IN ; P1_ADD_515_U151
g30747 nand P1_ADD_515_U95 P1_ADD_515_U9 ; P1_ADD_515_U152
g30748 nand P1_ADD_515_U54 P1_INSTADDRPOINTER_REG_27__SCAN_IN ; P1_ADD_515_U153
g30749 nand P1_ADD_515_U118 P1_ADD_515_U55 ; P1_ADD_515_U154
g30750 nand P1_ADD_515_U28 P1_INSTADDRPOINTER_REG_14__SCAN_IN ; P1_ADD_515_U155
g30751 nand P1_ADD_515_U105 P1_ADD_515_U29 ; P1_ADD_515_U156
g30752 nand P1_ADD_515_U10 P1_INSTADDRPOINTER_REG_5__SCAN_IN ; P1_ADD_515_U157
g30753 nand P1_ADD_515_U96 P1_ADD_515_U11 ; P1_ADD_515_U158
g30754 nand P1_ADD_515_U16 P1_INSTADDRPOINTER_REG_8__SCAN_IN ; P1_ADD_515_U159
g30755 nand P1_ADD_515_U99 P1_ADD_515_U17 ; P1_ADD_515_U160
g30756 nand P1_ADD_515_U46 P1_INSTADDRPOINTER_REG_23__SCAN_IN ; P1_ADD_515_U161
g30757 nand P1_ADD_515_U114 P1_ADD_515_U47 ; P1_ADD_515_U162
g30758 nand P1_ADD_515_U38 P1_INSTADDRPOINTER_REG_19__SCAN_IN ; P1_ADD_515_U163
g30759 nand P1_ADD_515_U110 P1_ADD_515_U39 ; P1_ADD_515_U164
g30760 nand P1_ADD_515_U20 P1_INSTADDRPOINTER_REG_10__SCAN_IN ; P1_ADD_515_U165
g30761 nand P1_ADD_515_U101 P1_ADD_515_U21 ; P1_ADD_515_U166
g30762 nand P1_ADD_515_U93 P1_INSTADDRPOINTER_REG_31__SCAN_IN ; P1_ADD_515_U167
g30763 nand P1_ADD_515_U122 P1_ADD_515_U92 ; P1_ADD_515_U168
g30764 nand P1_ADD_515_U6 P1_INSTADDRPOINTER_REG_3__SCAN_IN ; P1_ADD_515_U169
g30765 nand P1_ADD_515_U94 P1_ADD_515_U7 ; P1_ADD_515_U170
g30766 nand P1_ADD_515_U56 P1_INSTADDRPOINTER_REG_28__SCAN_IN ; P1_ADD_515_U171
g30767 nand P1_ADD_515_U119 P1_ADD_515_U57 ; P1_ADD_515_U172
g30768 nand P1_ADD_515_U42 P1_INSTADDRPOINTER_REG_21__SCAN_IN ; P1_ADD_515_U173
g30769 nand P1_ADD_515_U112 P1_ADD_515_U43 ; P1_ADD_515_U174
g30770 nand P1_ADD_515_U24 P1_INSTADDRPOINTER_REG_12__SCAN_IN ; P1_ADD_515_U175
g30771 nand P1_ADD_515_U103 P1_ADD_515_U25 ; P1_ADD_515_U176
g30772 nand P1_ADD_515_U14 P1_INSTADDRPOINTER_REG_7__SCAN_IN ; P1_ADD_515_U177
g30773 nand P1_ADD_515_U98 P1_ADD_515_U15 ; P1_ADD_515_U178
g30774 nand P1_ADD_515_U50 P1_INSTADDRPOINTER_REG_25__SCAN_IN ; P1_ADD_515_U179
g30775 nand P1_ADD_515_U116 P1_ADD_515_U51 ; P1_ADD_515_U180
g30776 nand P1_ADD_515_U32 P1_INSTADDRPOINTER_REG_16__SCAN_IN ; P1_ADD_515_U181
g30777 nand P1_ADD_515_U107 P1_ADD_515_U33 ; P1_ADD_515_U182
