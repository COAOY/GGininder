i P2_WR_REG_SCAN_IN
i SI_31_
i SI_30_
i SI_29_
i SI_28_
i SI_27_
i SI_26_
i SI_25_
i SI_24_
i SI_23_
i SI_22_
i SI_21_
i SI_20_
i SI_19_
i SI_18_
i SI_17_
i SI_16_
i SI_15_
i SI_14_
i SI_13_
i SI_12_
i SI_11_
i SI_10_
i SI_9_
i SI_8_
i SI_7_
i SI_6_
i SI_5_
i SI_4_
i SI_3_
i SI_2_
i SI_1_
i SI_0_
i P2_RD_REG_SCAN_IN
i P2_STATE_REG_SCAN_IN
i P2_REG3_REG_7__SCAN_IN
i P2_REG3_REG_27__SCAN_IN
i P2_REG3_REG_14__SCAN_IN
i P2_REG3_REG_23__SCAN_IN
i P2_REG3_REG_10__SCAN_IN
i P2_REG3_REG_3__SCAN_IN
i P2_REG3_REG_19__SCAN_IN
i P2_REG3_REG_28__SCAN_IN
i P2_REG3_REG_8__SCAN_IN
i P2_REG3_REG_1__SCAN_IN
i P2_REG3_REG_21__SCAN_IN
i P2_REG3_REG_12__SCAN_IN
i P2_REG3_REG_25__SCAN_IN
i P2_REG3_REG_16__SCAN_IN
i P2_REG3_REG_5__SCAN_IN
i P2_REG3_REG_17__SCAN_IN
i P2_REG3_REG_24__SCAN_IN
i P2_REG3_REG_4__SCAN_IN
i P2_REG3_REG_9__SCAN_IN
i P2_REG3_REG_0__SCAN_IN
i P2_REG3_REG_20__SCAN_IN
i P2_REG3_REG_13__SCAN_IN
i P2_REG3_REG_22__SCAN_IN
i P2_REG3_REG_11__SCAN_IN
i P2_REG3_REG_2__SCAN_IN
i P2_REG3_REG_18__SCAN_IN
i P2_REG3_REG_6__SCAN_IN
i P2_REG3_REG_26__SCAN_IN
i P2_REG3_REG_15__SCAN_IN
i P2_B_REG_SCAN_IN
i P2_DATAO_REG_31__SCAN_IN
i P2_DATAO_REG_30__SCAN_IN
i P2_DATAO_REG_29__SCAN_IN
i P2_DATAO_REG_28__SCAN_IN
i P2_DATAO_REG_27__SCAN_IN
i P2_DATAO_REG_26__SCAN_IN
i P2_DATAO_REG_25__SCAN_IN
i P2_DATAO_REG_24__SCAN_IN
i P2_DATAO_REG_23__SCAN_IN
i P2_DATAO_REG_22__SCAN_IN
i P2_DATAO_REG_21__SCAN_IN
i P2_DATAO_REG_20__SCAN_IN
i P2_DATAO_REG_19__SCAN_IN
i P2_DATAO_REG_18__SCAN_IN
i P2_DATAO_REG_17__SCAN_IN
i P2_DATAO_REG_16__SCAN_IN
i P2_DATAO_REG_15__SCAN_IN
i P2_DATAO_REG_14__SCAN_IN
i P2_DATAO_REG_13__SCAN_IN
i P2_DATAO_REG_12__SCAN_IN
i P2_DATAO_REG_11__SCAN_IN
i P2_DATAO_REG_10__SCAN_IN
i P2_DATAO_REG_9__SCAN_IN
i P2_DATAO_REG_8__SCAN_IN
i P2_DATAO_REG_7__SCAN_IN
i P2_DATAO_REG_6__SCAN_IN
i P1_IR_REG_0__SCAN_IN
i P1_IR_REG_1__SCAN_IN
i P1_IR_REG_2__SCAN_IN
i P1_IR_REG_3__SCAN_IN
i P1_IR_REG_4__SCAN_IN
i P1_IR_REG_5__SCAN_IN
i P1_IR_REG_6__SCAN_IN
i P1_IR_REG_7__SCAN_IN
i P1_IR_REG_8__SCAN_IN
i P1_IR_REG_9__SCAN_IN
i P1_IR_REG_10__SCAN_IN
i P1_IR_REG_11__SCAN_IN
i P1_IR_REG_12__SCAN_IN
i P1_IR_REG_13__SCAN_IN
i P1_IR_REG_14__SCAN_IN
i P1_IR_REG_15__SCAN_IN
i P1_IR_REG_16__SCAN_IN
i P1_IR_REG_17__SCAN_IN
i P1_IR_REG_18__SCAN_IN
i P1_IR_REG_19__SCAN_IN
i P1_IR_REG_20__SCAN_IN
i P1_IR_REG_21__SCAN_IN
i P1_IR_REG_22__SCAN_IN
i P1_IR_REG_23__SCAN_IN
i P1_IR_REG_24__SCAN_IN
i P1_IR_REG_25__SCAN_IN
i P1_IR_REG_26__SCAN_IN
i P1_IR_REG_27__SCAN_IN
i P1_IR_REG_28__SCAN_IN
i P1_IR_REG_29__SCAN_IN
i P1_IR_REG_30__SCAN_IN
i P1_IR_REG_31__SCAN_IN
i P1_D_REG_0__SCAN_IN
i P1_D_REG_1__SCAN_IN
i P1_D_REG_2__SCAN_IN
i P1_D_REG_3__SCAN_IN
i P1_D_REG_4__SCAN_IN
i P1_D_REG_5__SCAN_IN
i P1_D_REG_6__SCAN_IN
i P1_D_REG_7__SCAN_IN
i P1_D_REG_8__SCAN_IN
i P1_D_REG_9__SCAN_IN
i P1_D_REG_10__SCAN_IN
i P1_D_REG_11__SCAN_IN
i P1_D_REG_12__SCAN_IN
i P1_D_REG_13__SCAN_IN
i P1_D_REG_14__SCAN_IN
i P1_D_REG_15__SCAN_IN
i P1_D_REG_16__SCAN_IN
i P1_D_REG_17__SCAN_IN
i P1_D_REG_18__SCAN_IN
i P1_D_REG_19__SCAN_IN
i P1_D_REG_20__SCAN_IN
i P1_D_REG_21__SCAN_IN
i P1_D_REG_22__SCAN_IN
i P1_D_REG_23__SCAN_IN
i P1_D_REG_24__SCAN_IN
i P1_D_REG_25__SCAN_IN
i P1_D_REG_26__SCAN_IN
i P1_D_REG_27__SCAN_IN
i P1_D_REG_28__SCAN_IN
i P1_D_REG_29__SCAN_IN
i P1_D_REG_30__SCAN_IN
i P1_D_REG_31__SCAN_IN
i P1_REG0_REG_0__SCAN_IN
i P1_REG0_REG_1__SCAN_IN
i P1_REG0_REG_2__SCAN_IN
i P1_REG0_REG_3__SCAN_IN
i P1_REG0_REG_4__SCAN_IN
i P1_REG0_REG_5__SCAN_IN
i P1_REG0_REG_6__SCAN_IN
i P1_REG0_REG_7__SCAN_IN
i P1_REG0_REG_8__SCAN_IN
i P1_REG0_REG_9__SCAN_IN
i P1_REG0_REG_10__SCAN_IN
i P1_REG0_REG_11__SCAN_IN
i P1_REG0_REG_12__SCAN_IN
i P1_REG0_REG_13__SCAN_IN
i P1_REG0_REG_14__SCAN_IN
i P1_REG0_REG_15__SCAN_IN
i P1_REG0_REG_16__SCAN_IN
i P1_REG0_REG_17__SCAN_IN
i P1_REG0_REG_18__SCAN_IN
i P1_REG0_REG_19__SCAN_IN
i P1_REG0_REG_20__SCAN_IN
i P1_REG0_REG_21__SCAN_IN
i P1_REG0_REG_22__SCAN_IN
i P1_REG0_REG_23__SCAN_IN
i P1_REG0_REG_24__SCAN_IN
i P1_REG0_REG_25__SCAN_IN
i P1_REG0_REG_26__SCAN_IN
i P1_REG0_REG_27__SCAN_IN
i P1_REG0_REG_28__SCAN_IN
i P1_REG0_REG_29__SCAN_IN
i P1_REG0_REG_30__SCAN_IN
i P1_REG0_REG_31__SCAN_IN
i P1_REG1_REG_0__SCAN_IN
i P1_REG1_REG_1__SCAN_IN
i P1_REG1_REG_2__SCAN_IN
i P1_REG1_REG_3__SCAN_IN
i P1_REG1_REG_4__SCAN_IN
i P1_REG1_REG_5__SCAN_IN
i P1_REG1_REG_6__SCAN_IN
i P1_REG1_REG_7__SCAN_IN
i P1_REG1_REG_8__SCAN_IN
i P1_REG1_REG_9__SCAN_IN
i P1_REG1_REG_10__SCAN_IN
i P1_REG1_REG_11__SCAN_IN
i P1_REG1_REG_12__SCAN_IN
i P1_REG1_REG_13__SCAN_IN
i P1_REG1_REG_14__SCAN_IN
i P1_REG1_REG_15__SCAN_IN
i P1_REG1_REG_16__SCAN_IN
i P1_REG1_REG_17__SCAN_IN
i P1_REG1_REG_18__SCAN_IN
i P1_REG1_REG_19__SCAN_IN
i P1_REG1_REG_20__SCAN_IN
i P1_REG1_REG_21__SCAN_IN
i P1_REG1_REG_22__SCAN_IN
i P1_REG1_REG_23__SCAN_IN
i P1_REG1_REG_24__SCAN_IN
i P1_REG1_REG_25__SCAN_IN
i P1_REG1_REG_26__SCAN_IN
i P1_REG1_REG_27__SCAN_IN
i P1_REG1_REG_28__SCAN_IN
i P1_REG1_REG_29__SCAN_IN
i P1_REG1_REG_30__SCAN_IN
i P1_REG1_REG_31__SCAN_IN
i P1_REG2_REG_0__SCAN_IN
i P1_REG2_REG_1__SCAN_IN
i P1_REG2_REG_2__SCAN_IN
i P1_REG2_REG_3__SCAN_IN
i P1_REG2_REG_4__SCAN_IN
i P1_REG2_REG_5__SCAN_IN
i P1_REG2_REG_6__SCAN_IN
i P1_REG2_REG_7__SCAN_IN
i P1_REG2_REG_8__SCAN_IN
i P1_REG2_REG_9__SCAN_IN
i P1_REG2_REG_10__SCAN_IN
i P1_REG2_REG_11__SCAN_IN
i P1_REG2_REG_12__SCAN_IN
i P1_REG2_REG_13__SCAN_IN
i P1_REG2_REG_14__SCAN_IN
i P1_REG2_REG_15__SCAN_IN
i P1_REG2_REG_16__SCAN_IN
i P1_REG2_REG_17__SCAN_IN
i P1_REG2_REG_18__SCAN_IN
i P1_REG2_REG_19__SCAN_IN
i P1_REG2_REG_20__SCAN_IN
i P1_REG2_REG_21__SCAN_IN
i P1_REG2_REG_22__SCAN_IN
i P1_REG2_REG_23__SCAN_IN
i P1_REG2_REG_24__SCAN_IN
i P1_REG2_REG_25__SCAN_IN
i P1_REG2_REG_26__SCAN_IN
i P1_REG2_REG_27__SCAN_IN
i P1_REG2_REG_28__SCAN_IN
i P1_REG2_REG_29__SCAN_IN
i P1_REG2_REG_30__SCAN_IN
i P1_REG2_REG_31__SCAN_IN
i P1_ADDR_REG_19__SCAN_IN
i P1_ADDR_REG_18__SCAN_IN
i P1_ADDR_REG_17__SCAN_IN
i P1_ADDR_REG_16__SCAN_IN
i P1_ADDR_REG_15__SCAN_IN
i P1_ADDR_REG_14__SCAN_IN
i P1_ADDR_REG_13__SCAN_IN
i P1_ADDR_REG_12__SCAN_IN
i P1_ADDR_REG_11__SCAN_IN
i P1_ADDR_REG_10__SCAN_IN
i P1_ADDR_REG_9__SCAN_IN
i P1_ADDR_REG_8__SCAN_IN
i P1_ADDR_REG_7__SCAN_IN
i P1_ADDR_REG_6__SCAN_IN
i P1_ADDR_REG_5__SCAN_IN
i P1_ADDR_REG_4__SCAN_IN
i P1_ADDR_REG_3__SCAN_IN
i P1_ADDR_REG_2__SCAN_IN
i P1_ADDR_REG_1__SCAN_IN
i P1_ADDR_REG_0__SCAN_IN
i P1_DATAO_REG_0__SCAN_IN
i P1_DATAO_REG_1__SCAN_IN
i P1_DATAO_REG_2__SCAN_IN
i P1_DATAO_REG_3__SCAN_IN
i P1_DATAO_REG_4__SCAN_IN
i P1_DATAO_REG_5__SCAN_IN
i P1_DATAO_REG_6__SCAN_IN
i P1_DATAO_REG_7__SCAN_IN
i P1_DATAO_REG_8__SCAN_IN
i P1_DATAO_REG_9__SCAN_IN
i P1_DATAO_REG_10__SCAN_IN
i P1_DATAO_REG_11__SCAN_IN
i P1_DATAO_REG_12__SCAN_IN
i P1_DATAO_REG_13__SCAN_IN
i P1_DATAO_REG_14__SCAN_IN
i P1_DATAO_REG_15__SCAN_IN
i P1_DATAO_REG_16__SCAN_IN
i P1_DATAO_REG_17__SCAN_IN
i P1_DATAO_REG_18__SCAN_IN
i P1_DATAO_REG_19__SCAN_IN
i P1_DATAO_REG_20__SCAN_IN
i P1_DATAO_REG_21__SCAN_IN
i P1_DATAO_REG_22__SCAN_IN
i P1_DATAO_REG_23__SCAN_IN
i P1_DATAO_REG_24__SCAN_IN
i P1_DATAO_REG_25__SCAN_IN
i P1_DATAO_REG_26__SCAN_IN
i P1_DATAO_REG_27__SCAN_IN
i P1_DATAO_REG_28__SCAN_IN
i P1_DATAO_REG_29__SCAN_IN
i P1_DATAO_REG_30__SCAN_IN
i P1_DATAO_REG_31__SCAN_IN
i P1_B_REG_SCAN_IN
i P1_REG3_REG_15__SCAN_IN
i P1_REG3_REG_26__SCAN_IN
i P1_REG3_REG_6__SCAN_IN
i P1_REG3_REG_18__SCAN_IN
i P1_REG3_REG_2__SCAN_IN
i P1_REG3_REG_11__SCAN_IN
i P1_REG3_REG_22__SCAN_IN
i P1_REG3_REG_13__SCAN_IN
i P1_REG3_REG_20__SCAN_IN
i P1_REG3_REG_0__SCAN_IN
i P1_REG3_REG_9__SCAN_IN
i P1_REG3_REG_4__SCAN_IN
i P1_REG3_REG_24__SCAN_IN
i P1_REG3_REG_17__SCAN_IN
i P1_REG3_REG_5__SCAN_IN
i P1_REG3_REG_16__SCAN_IN
i P1_REG3_REG_25__SCAN_IN
i P1_REG3_REG_12__SCAN_IN
i P1_REG3_REG_21__SCAN_IN
i P1_REG3_REG_1__SCAN_IN
i P1_REG3_REG_8__SCAN_IN
i P1_REG3_REG_28__SCAN_IN
i P1_REG3_REG_19__SCAN_IN
i P1_REG3_REG_3__SCAN_IN
i P1_REG3_REG_10__SCAN_IN
i P1_REG3_REG_23__SCAN_IN
i P1_REG3_REG_14__SCAN_IN
i P1_REG3_REG_27__SCAN_IN
i P1_REG3_REG_7__SCAN_IN
i P1_STATE_REG_SCAN_IN
i P1_RD_REG_SCAN_IN
i P1_WR_REG_SCAN_IN
i P2_IR_REG_0__SCAN_IN
i P2_IR_REG_1__SCAN_IN
i P2_IR_REG_2__SCAN_IN
i P2_IR_REG_3__SCAN_IN
i P2_IR_REG_4__SCAN_IN
i P2_IR_REG_5__SCAN_IN
i P2_IR_REG_6__SCAN_IN
i P2_IR_REG_7__SCAN_IN
i P2_IR_REG_8__SCAN_IN
i P2_IR_REG_9__SCAN_IN
i P2_IR_REG_10__SCAN_IN
i P2_IR_REG_11__SCAN_IN
i P2_IR_REG_12__SCAN_IN
i P2_IR_REG_13__SCAN_IN
i P2_IR_REG_14__SCAN_IN
i P2_IR_REG_15__SCAN_IN
i P2_IR_REG_16__SCAN_IN
i P2_IR_REG_17__SCAN_IN
i P2_IR_REG_18__SCAN_IN
i P2_IR_REG_19__SCAN_IN
i P2_IR_REG_20__SCAN_IN
i P2_IR_REG_21__SCAN_IN
i P2_IR_REG_22__SCAN_IN
i P2_IR_REG_23__SCAN_IN
i P2_IR_REG_24__SCAN_IN
i P2_IR_REG_25__SCAN_IN
i P2_IR_REG_26__SCAN_IN
i P2_IR_REG_27__SCAN_IN
i P2_IR_REG_28__SCAN_IN
i P2_IR_REG_29__SCAN_IN
i P2_IR_REG_30__SCAN_IN
i P2_IR_REG_31__SCAN_IN
i P2_D_REG_0__SCAN_IN
i P2_D_REG_1__SCAN_IN
i P2_D_REG_2__SCAN_IN
i P2_D_REG_3__SCAN_IN
i P2_D_REG_4__SCAN_IN
i P2_D_REG_5__SCAN_IN
i P2_D_REG_6__SCAN_IN
i P2_D_REG_7__SCAN_IN
i P2_D_REG_8__SCAN_IN
i P2_D_REG_9__SCAN_IN
i P2_D_REG_10__SCAN_IN
i P2_D_REG_11__SCAN_IN
i P2_D_REG_12__SCAN_IN
i P2_D_REG_13__SCAN_IN
i P2_D_REG_14__SCAN_IN
i P2_D_REG_15__SCAN_IN
i P2_D_REG_16__SCAN_IN
i P2_D_REG_17__SCAN_IN
i P2_D_REG_18__SCAN_IN
i P2_D_REG_19__SCAN_IN
i P2_D_REG_20__SCAN_IN
i P2_D_REG_21__SCAN_IN
i P2_D_REG_22__SCAN_IN
i P2_D_REG_23__SCAN_IN
i P2_D_REG_24__SCAN_IN
i P2_D_REG_25__SCAN_IN
i P2_D_REG_26__SCAN_IN
i P2_D_REG_27__SCAN_IN
i P2_D_REG_28__SCAN_IN
i P2_D_REG_29__SCAN_IN
i P2_D_REG_30__SCAN_IN
i P2_D_REG_31__SCAN_IN
i P2_REG0_REG_0__SCAN_IN
i P2_REG0_REG_1__SCAN_IN
i P2_REG0_REG_2__SCAN_IN
i P2_REG0_REG_3__SCAN_IN
i P2_REG0_REG_4__SCAN_IN
i P2_REG0_REG_5__SCAN_IN
i P2_REG0_REG_6__SCAN_IN
i P2_REG0_REG_7__SCAN_IN
i P2_REG0_REG_8__SCAN_IN
i P2_REG0_REG_9__SCAN_IN
i P2_REG0_REG_10__SCAN_IN
i P2_REG0_REG_11__SCAN_IN
i P2_REG0_REG_12__SCAN_IN
i P2_REG0_REG_13__SCAN_IN
i P2_REG0_REG_14__SCAN_IN
i P2_REG0_REG_15__SCAN_IN
i P2_REG0_REG_16__SCAN_IN
i P2_REG0_REG_17__SCAN_IN
i P2_REG0_REG_18__SCAN_IN
i P2_REG0_REG_19__SCAN_IN
i P2_REG0_REG_20__SCAN_IN
i P2_REG0_REG_21__SCAN_IN
i P2_REG0_REG_22__SCAN_IN
i P2_REG0_REG_23__SCAN_IN
i P2_REG0_REG_24__SCAN_IN
i P2_REG0_REG_25__SCAN_IN
i P2_REG0_REG_26__SCAN_IN
i P2_REG0_REG_27__SCAN_IN
i P2_REG0_REG_28__SCAN_IN
i P2_REG0_REG_29__SCAN_IN
i P2_REG0_REG_30__SCAN_IN
i P2_REG0_REG_31__SCAN_IN
i P2_REG1_REG_0__SCAN_IN
i P2_REG1_REG_1__SCAN_IN
i P2_REG1_REG_2__SCAN_IN
i P2_REG1_REG_3__SCAN_IN
i P2_REG1_REG_4__SCAN_IN
i P2_REG1_REG_5__SCAN_IN
i P2_REG1_REG_6__SCAN_IN
i P2_REG1_REG_7__SCAN_IN
i P2_REG1_REG_8__SCAN_IN
i P2_REG1_REG_9__SCAN_IN
i P2_REG1_REG_10__SCAN_IN
i P2_REG1_REG_11__SCAN_IN
i P2_REG1_REG_12__SCAN_IN
i P2_REG1_REG_13__SCAN_IN
i P2_REG1_REG_14__SCAN_IN
i P2_REG1_REG_15__SCAN_IN
i P2_REG1_REG_16__SCAN_IN
i P2_REG1_REG_17__SCAN_IN
i P2_REG1_REG_18__SCAN_IN
i P2_REG1_REG_19__SCAN_IN
i P2_REG1_REG_20__SCAN_IN
i P2_REG1_REG_21__SCAN_IN
i P2_REG1_REG_22__SCAN_IN
i P2_REG1_REG_23__SCAN_IN
i P2_REG1_REG_24__SCAN_IN
i P2_REG1_REG_25__SCAN_IN
i P2_REG1_REG_26__SCAN_IN
i P2_REG1_REG_27__SCAN_IN
i P2_REG1_REG_28__SCAN_IN
i P2_REG1_REG_29__SCAN_IN
i P2_REG1_REG_30__SCAN_IN
i P2_REG1_REG_31__SCAN_IN
i P2_REG2_REG_0__SCAN_IN
i P2_REG2_REG_1__SCAN_IN
i P2_REG2_REG_2__SCAN_IN
i P2_REG2_REG_3__SCAN_IN
i P2_REG2_REG_4__SCAN_IN
i P2_REG2_REG_5__SCAN_IN
i P2_REG2_REG_6__SCAN_IN
i P2_REG2_REG_7__SCAN_IN
i P2_REG2_REG_8__SCAN_IN
i P2_REG2_REG_9__SCAN_IN
i P2_REG2_REG_10__SCAN_IN
i P2_REG2_REG_11__SCAN_IN
i P2_REG2_REG_12__SCAN_IN
i P2_REG2_REG_13__SCAN_IN
i P2_REG2_REG_14__SCAN_IN
i P2_REG2_REG_15__SCAN_IN
i P2_REG2_REG_16__SCAN_IN
i P2_REG2_REG_17__SCAN_IN
i P2_REG2_REG_18__SCAN_IN
i P2_REG2_REG_19__SCAN_IN
i P2_REG2_REG_20__SCAN_IN
i P2_REG2_REG_21__SCAN_IN
i P2_REG2_REG_22__SCAN_IN
i P2_REG2_REG_23__SCAN_IN
i P2_REG2_REG_24__SCAN_IN
i P2_REG2_REG_25__SCAN_IN
i P2_REG2_REG_26__SCAN_IN
i P2_REG2_REG_27__SCAN_IN
i P2_REG2_REG_28__SCAN_IN
i P2_REG2_REG_29__SCAN_IN
i P2_REG2_REG_30__SCAN_IN
i P2_REG2_REG_31__SCAN_IN
i P2_ADDR_REG_19__SCAN_IN
i P2_ADDR_REG_18__SCAN_IN
i P2_ADDR_REG_17__SCAN_IN
i P2_ADDR_REG_16__SCAN_IN
i P2_ADDR_REG_15__SCAN_IN
i P2_ADDR_REG_14__SCAN_IN
i P2_ADDR_REG_13__SCAN_IN
i P2_ADDR_REG_12__SCAN_IN
i P2_ADDR_REG_11__SCAN_IN
i P2_ADDR_REG_10__SCAN_IN
i P2_ADDR_REG_9__SCAN_IN
i P2_ADDR_REG_8__SCAN_IN
i P2_ADDR_REG_7__SCAN_IN
i P2_ADDR_REG_6__SCAN_IN
i P2_ADDR_REG_5__SCAN_IN
i P2_ADDR_REG_4__SCAN_IN
i P2_ADDR_REG_3__SCAN_IN
i P2_ADDR_REG_2__SCAN_IN
i P2_ADDR_REG_1__SCAN_IN
i P2_ADDR_REG_0__SCAN_IN
i P2_DATAO_REG_0__SCAN_IN
i P2_DATAO_REG_1__SCAN_IN
i P2_DATAO_REG_2__SCAN_IN
i P2_DATAO_REG_3__SCAN_IN
i P2_DATAO_REG_4__SCAN_IN
i P2_DATAO_REG_5__SCAN_IN
o ADD_1071_U4
o ADD_1071_U55
o ADD_1071_U56
o ADD_1071_U57
o ADD_1071_U58
o ADD_1071_U59
o ADD_1071_U60
o ADD_1071_U61
o ADD_1071_U62
o ADD_1071_U63
o ADD_1071_U47
o ADD_1071_U48
o ADD_1071_U49
o ADD_1071_U50
o ADD_1071_U51
o ADD_1071_U52
o ADD_1071_U53
o ADD_1071_U54
o ADD_1071_U5
o ADD_1071_U46
o U126
o U123
o P1_U3353
o P1_U3352
o P1_U3351
o P1_U3350
o P1_U3349
o P1_U3348
o P1_U3347
o P1_U3346
o P1_U3345
o P1_U3344
o P1_U3343
o P1_U3342
o P1_U3341
o P1_U3340
o P1_U3339
o P1_U3338
o P1_U3337
o P1_U3336
o P1_U3335
o P1_U3334
o P1_U3333
o P1_U3332
o P1_U3331
o P1_U3330
o P1_U3329
o P1_U3328
o P1_U3327
o P1_U3326
o P1_U3325
o P1_U3324
o P1_U3323
o P1_U3322
o P1_U3440
o P1_U3441
o P1_U3321
o P1_U3320
o P1_U3319
o P1_U3318
o P1_U3317
o P1_U3316
o P1_U3315
o P1_U3314
o P1_U3313
o P1_U3312
o P1_U3311
o P1_U3310
o P1_U3309
o P1_U3308
o P1_U3307
o P1_U3306
o P1_U3305
o P1_U3304
o P1_U3303
o P1_U3302
o P1_U3301
o P1_U3300
o P1_U3299
o P1_U3298
o P1_U3297
o P1_U3296
o P1_U3295
o P1_U3294
o P1_U3293
o P1_U3292
o P1_U3454
o P1_U3457
o P1_U3460
o P1_U3463
o P1_U3466
o P1_U3469
o P1_U3472
o P1_U3475
o P1_U3478
o P1_U3481
o P1_U3484
o P1_U3487
o P1_U3490
o P1_U3493
o P1_U3496
o P1_U3499
o P1_U3502
o P1_U3505
o P1_U3508
o P1_U3510
o P1_U3511
o P1_U3512
o P1_U3513
o P1_U3514
o P1_U3515
o P1_U3516
o P1_U3517
o P1_U3518
o P1_U3519
o P1_U3520
o P1_U3521
o P1_U3522
o P1_U3523
o P1_U3524
o P1_U3525
o P1_U3526
o P1_U3527
o P1_U3528
o P1_U3529
o P1_U3530
o P1_U3531
o P1_U3532
o P1_U3533
o P1_U3534
o P1_U3535
o P1_U3536
o P1_U3537
o P1_U3538
o P1_U3539
o P1_U3540
o P1_U3541
o P1_U3542
o P1_U3543
o P1_U3544
o P1_U3545
o P1_U3546
o P1_U3547
o P1_U3548
o P1_U3549
o P1_U3550
o P1_U3551
o P1_U3552
o P1_U3553
o P1_U3554
o P1_U3291
o P1_U3290
o P1_U3289
o P1_U3288
o P1_U3287
o P1_U3286
o P1_U3285
o P1_U3284
o P1_U3283
o P1_U3282
o P1_U3281
o P1_U3280
o P1_U3279
o P1_U3278
o P1_U3277
o P1_U3276
o P1_U3275
o P1_U3274
o P1_U3273
o P1_U3272
o P1_U3271
o P1_U3270
o P1_U3269
o P1_U3268
o P1_U3267
o P1_U3266
o P1_U3265
o P1_U3264
o P1_U3263
o P1_U3355
o P1_U3262
o P1_U3261
o P1_U3260
o P1_U3259
o P1_U3258
o P1_U3257
o P1_U3256
o P1_U3255
o P1_U3254
o P1_U3253
o P1_U3252
o P1_U3251
o P1_U3250
o P1_U3249
o P1_U3248
o P1_U3247
o P1_U3246
o P1_U3245
o P1_U3244
o P1_U3243
o P1_U3242
o P1_U3241
o P1_U3555
o P1_U3556
o P1_U3557
o P1_U3558
o P1_U3559
o P1_U3560
o P1_U3561
o P1_U3562
o P1_U3563
o P1_U3564
o P1_U3565
o P1_U3566
o P1_U3567
o P1_U3568
o P1_U3569
o P1_U3570
o P1_U3571
o P1_U3572
o P1_U3573
o P1_U3574
o P1_U3575
o P1_U3576
o P1_U3577
o P1_U3578
o P1_U3579
o P1_U3580
o P1_U3581
o P1_U3582
o P1_U3583
o P1_U3584
o P1_U3585
o P1_U3586
o P1_U3240
o P1_U3239
o P1_U3238
o P1_U3237
o P1_U3236
o P1_U3235
o P1_U3234
o P1_U3233
o P1_U3232
o P1_U3231
o P1_U3230
o P1_U3229
o P1_U3228
o P1_U3227
o P1_U3226
o P1_U3225
o P1_U3224
o P1_U3223
o P1_U3222
o P1_U3221
o P1_U3220
o P1_U3219
o P1_U3218
o P1_U3217
o P1_U3216
o P1_U3215
o P1_U3214
o P1_U3213
o P1_U3212
o P1_U3211
o P1_U3084
o P1_U3083
o P1_U4006
o P2_U3358
o P2_U3357
o P2_U3356
o P2_U3355
o P2_U3354
o P2_U3353
o P2_U3352
o P2_U3351
o P2_U3350
o P2_U3349
o P2_U3348
o P2_U3347
o P2_U3346
o P2_U3345
o P2_U3344
o P2_U3343
o P2_U3342
o P2_U3341
o P2_U3340
o P2_U3339
o P2_U3338
o P2_U3337
o P2_U3336
o P2_U3335
o P2_U3334
o P2_U3333
o P2_U3332
o P2_U3331
o P2_U3330
o P2_U3329
o P2_U3328
o P2_U3327
o P2_U3437
o P2_U3438
o P2_U3326
o P2_U3325
o P2_U3324
o P2_U3323
o P2_U3322
o P2_U3321
o P2_U3320
o P2_U3319
o P2_U3318
o P2_U3317
o P2_U3316
o P2_U3315
o P2_U3314
o P2_U3313
o P2_U3312
o P2_U3311
o P2_U3310
o P2_U3309
o P2_U3308
o P2_U3307
o P2_U3306
o P2_U3305
o P2_U3304
o P2_U3303
o P2_U3302
o P2_U3301
o P2_U3300
o P2_U3299
o P2_U3298
o P2_U3297
o P2_U3451
o P2_U3454
o P2_U3457
o P2_U3460
o P2_U3463
o P2_U3466
o P2_U3469
o P2_U3472
o P2_U3475
o P2_U3478
o P2_U3481
o P2_U3484
o P2_U3487
o P2_U3490
o P2_U3493
o P2_U3496
o P2_U3499
o P2_U3502
o P2_U3505
o P2_U3507
o P2_U3508
o P2_U3509
o P2_U3510
o P2_U3511
o P2_U3512
o P2_U3513
o P2_U3514
o P2_U3515
o P2_U3516
o P2_U3517
o P2_U3518
o P2_U3519
o P2_U3520
o P2_U3521
o P2_U3522
o P2_U3523
o P2_U3524
o P2_U3525
o P2_U3526
o P2_U3527
o P2_U3528
o P2_U3529
o P2_U3530
o P2_U3531
o P2_U3532
o P2_U3533
o P2_U3534
o P2_U3535
o P2_U3536
o P2_U3537
o P2_U3538
o P2_U3539
o P2_U3540
o P2_U3541
o P2_U3542
o P2_U3543
o P2_U3544
o P2_U3545
o P2_U3546
o P2_U3547
o P2_U3548
o P2_U3549
o P2_U3550
o P2_U3551
o P2_U3296
o P2_U3295
o P2_U3294
o P2_U3293
o P2_U3292
o P2_U3291
o P2_U3290
o P2_U3289
o P2_U3288
o P2_U3287
o P2_U3286
o P2_U3285
o P2_U3284
o P2_U3283
o P2_U3282
o P2_U3281
o P2_U3280
o P2_U3279
o P2_U3278
o P2_U3277
o P2_U3276
o P2_U3275
o P2_U3274
o P2_U3273
o P2_U3272
o P2_U3271
o P2_U3270
o P2_U3269
o P2_U3268
o P2_U3267
o P2_U3266
o P2_U3265
o P2_U3264
o P2_U3263
o P2_U3262
o P2_U3261
o P2_U3260
o P2_U3259
o P2_U3258
o P2_U3257
o P2_U3256
o P2_U3255
o P2_U3254
o P2_U3253
o P2_U3252
o P2_U3251
o P2_U3250
o P2_U3249
o P2_U3248
o P2_U3247
o P2_U3246
o P2_U3245
o P2_U3552
o P2_U3553
o P2_U3554
o P2_U3555
o P2_U3556
o P2_U3557
o P2_U3558
o P2_U3559
o P2_U3560
o P2_U3561
o P2_U3562
o P2_U3563
o P2_U3564
o P2_U3565
o P2_U3566
o P2_U3567
o P2_U3568
o P2_U3569
o P2_U3570
o P2_U3571
o P2_U3572
o P2_U3573
o P2_U3574
o P2_U3575
o P2_U3576
o P2_U3577
o P2_U3578
o P2_U3579
o P2_U3580
o P2_U3581
o P2_U3582
o P2_U3583
o P2_U3244
o P2_U3243
o P2_U3242
o P2_U3241
o P2_U3240
o P2_U3239
o P2_U3238
o P2_U3237
o P2_U3236
o P2_U3235
o P2_U3234
o P2_U3233
o P2_U3232
o P2_U3231
o P2_U3230
o P2_U3229
o P2_U3228
o P2_U3227
o P2_U3226
o P2_U3225
o P2_U3224
o P2_U3223
o P2_U3222
o P2_U3221
o P2_U3220
o P2_U3219
o P2_U3218
o P2_U3217
o P2_U3216
o P2_U3215
o P2_U3152
o P2_U3151
o P2_U3966
g1 nand U136 U135 ; U25
g2 nand U138 U137 ; U26
g3 nand U140 U139 ; U27
g4 nand U142 U141 ; U28
g5 nand U144 U143 ; U29
g6 nand U146 U145 ; U30
g7 nand U148 U147 ; U31
g8 nand U150 U149 ; U32
g9 nand U152 U151 ; U33
g10 nand U154 U153 ; U34
g11 nand U156 U155 ; U35
g12 nand U158 U157 ; U36
g13 nand U160 U159 ; U37
g14 nand U162 U161 ; U38
g15 nand U164 U163 ; U39
g16 nand U166 U165 ; U40
g17 nand U168 U167 ; U41
g18 nand U170 U169 ; U42
g19 nand U172 U171 ; U43
g20 nand U174 U173 ; U44
g21 nand U176 U175 ; U45
g22 nand U178 U177 ; U46
g23 nand U180 U179 ; U47
g24 nand U182 U181 ; U48
g25 nand U184 U183 ; U49
g26 nand U186 U185 ; U50
g27 nand U188 U187 ; U51
g28 nand U190 U189 ; U52
g29 nand U192 U191 ; U53
g30 nand U194 U193 ; U54
g31 nand U196 U195 ; U55
g32 nand U198 U197 ; U56
g33 nand U200 U199 ; U57
g34 nand U202 U201 ; U58
g35 nand U204 U203 ; U59
g36 nand U206 U205 ; U60
g37 nand U208 U207 ; U61
g38 nand U210 U209 ; U62
g39 nand U212 U211 ; U63
g40 nand U214 U213 ; U64
g41 nand U216 U215 ; U65
g42 nand U218 U217 ; U66
g43 nand U220 U219 ; U67
g44 nand U222 U221 ; U68
g45 nand U224 U223 ; U69
g46 nand U226 U225 ; U70
g47 nand U228 U227 ; U71
g48 nand U230 U229 ; U72
g49 nand U232 U231 ; U73
g50 nand U234 U233 ; U74
g51 nand U236 U235 ; U75
g52 nand U238 U237 ; U76
g53 nand U240 U239 ; U77
g54 nand U242 U241 ; U78
g55 nand U244 U243 ; U79
g56 nand U246 U245 ; U80
g57 nand U248 U247 ; U81
g58 nand U250 U249 ; U82
g59 nand U252 U251 ; U83
g60 nand U254 U253 ; U84
g61 nand U256 U255 ; U85
g62 nand U258 U257 ; U86
g63 nand U260 U259 ; U87
g64 nand U262 U261 ; U88
g65 nand U264 U263 ; U89
g66 nand U266 U265 ; U90
g67 nand U268 U267 ; U91
g68 nand U270 U269 ; U92
g69 nand U272 U271 ; U93
g70 nand U274 U273 ; U94
g71 nand U276 U275 ; U95
g72 nand U278 U277 ; U96
g73 nand U280 U279 ; U97
g74 nand U282 U281 ; U98
g75 nand U284 U283 ; U99
g76 nand U286 U285 ; U100
g77 nand U288 U287 ; U101
g78 nand U290 U289 ; U102
g79 nand U292 U291 ; U103
g80 nand U294 U293 ; U104
g81 nand U296 U295 ; U105
g82 nand U298 U297 ; U106
g83 nand U300 U299 ; U107
g84 nand U302 U301 ; U108
g85 nand U304 U303 ; U109
g86 nand U306 U305 ; U110
g87 nand U308 U307 ; U111
g88 nand U310 U309 ; U112
g89 nand U312 U311 ; U113
g90 nand U314 U313 ; U114
g91 nand U316 U315 ; U115
g92 nand U318 U317 ; U116
g93 nand U320 U319 ; U117
g94 nand U322 U321 ; U118
g95 nand U324 U323 ; U119
g96 nand U326 U325 ; U120
g97 not P2_WR_REG_SCAN_IN ; U121
g98 not P1_WR_REG_SCAN_IN ; U122
g99 and U132 U131 ; U123
g100 not P2_RD_REG_SCAN_IN ; U124
g101 not P1_RD_REG_SCAN_IN ; U125
g102 and U134 U133 ; U126
g103 nand U129 U128 ; U127
g104 nand LT_1079_U6 U125 LT_1079_19_U6 ; U128
g105 nand U124 P1_ADDR_REG_19__SCAN_IN P2_ADDR_REG_19__SCAN_IN ; U129
g106 not U127 ; U130
g107 nand U122 P2_WR_REG_SCAN_IN ; U131
g108 nand U121 P1_WR_REG_SCAN_IN ; U132
g109 nand U125 P2_RD_REG_SCAN_IN ; U133
g110 nand U124 P1_RD_REG_SCAN_IN ; U134
g111 nand U127 P1_DATAO_REG_9__SCAN_IN ; U135
g112 nand R140_U84 U130 ; U136
g113 nand U127 P1_DATAO_REG_8__SCAN_IN ; U137
g114 nand R140_U85 U130 ; U138
g115 nand U127 P1_DATAO_REG_7__SCAN_IN ; U139
g116 nand R140_U86 U130 ; U140
g117 nand U127 P1_DATAO_REG_6__SCAN_IN ; U141
g118 nand R140_U87 U130 ; U142
g119 nand U127 P1_DATAO_REG_5__SCAN_IN ; U143
g120 nand R140_U88 U130 ; U144
g121 nand U127 P1_DATAO_REG_4__SCAN_IN ; U145
g122 nand R140_U89 U130 ; U146
g123 nand U127 P1_DATAO_REG_3__SCAN_IN ; U147
g124 nand R140_U90 U130 ; U148
g125 nand U127 P1_DATAO_REG_31__SCAN_IN ; U149
g126 nand R140_U11 U130 ; U150
g127 nand U127 P1_DATAO_REG_30__SCAN_IN ; U151
g128 nand R140_U91 U130 ; U152
g129 nand U127 P1_DATAO_REG_2__SCAN_IN ; U153
g130 nand R140_U92 U130 ; U154
g131 nand U127 P1_DATAO_REG_29__SCAN_IN ; U155
g132 nand R140_U93 U130 ; U156
g133 nand U127 P1_DATAO_REG_28__SCAN_IN ; U157
g134 nand R140_U94 U130 ; U158
g135 nand U127 P1_DATAO_REG_27__SCAN_IN ; U159
g136 nand R140_U95 U130 ; U160
g137 nand U127 P1_DATAO_REG_26__SCAN_IN ; U161
g138 nand R140_U96 U130 ; U162
g139 nand U127 P1_DATAO_REG_25__SCAN_IN ; U163
g140 nand R140_U97 U130 ; U164
g141 nand U127 P1_DATAO_REG_24__SCAN_IN ; U165
g142 nand R140_U98 U130 ; U166
g143 nand U127 P1_DATAO_REG_23__SCAN_IN ; U167
g144 nand R140_U99 U130 ; U168
g145 nand U127 P1_DATAO_REG_22__SCAN_IN ; U169
g146 nand R140_U100 U130 ; U170
g147 nand U127 P1_DATAO_REG_21__SCAN_IN ; U171
g148 nand R140_U101 U130 ; U172
g149 nand U127 P1_DATAO_REG_20__SCAN_IN ; U173
g150 nand R140_U102 U130 ; U174
g151 nand U127 P1_DATAO_REG_1__SCAN_IN ; U175
g152 nand R140_U10 U130 ; U176
g153 nand U127 P1_DATAO_REG_19__SCAN_IN ; U177
g154 nand R140_U103 U130 ; U178
g155 nand U127 P1_DATAO_REG_18__SCAN_IN ; U179
g156 nand R140_U104 U130 ; U180
g157 nand U127 P1_DATAO_REG_17__SCAN_IN ; U181
g158 nand R140_U105 U130 ; U182
g159 nand U127 P1_DATAO_REG_16__SCAN_IN ; U183
g160 nand R140_U106 U130 ; U184
g161 nand U127 P1_DATAO_REG_15__SCAN_IN ; U185
g162 nand R140_U107 U130 ; U186
g163 nand U127 P1_DATAO_REG_14__SCAN_IN ; U187
g164 nand R140_U108 U130 ; U188
g165 nand U127 P1_DATAO_REG_13__SCAN_IN ; U189
g166 nand R140_U109 U130 ; U190
g167 nand U127 P1_DATAO_REG_12__SCAN_IN ; U191
g168 nand R140_U110 U130 ; U192
g169 nand U127 P1_DATAO_REG_11__SCAN_IN ; U193
g170 nand R140_U111 U130 ; U194
g171 nand U127 P1_DATAO_REG_10__SCAN_IN ; U195
g172 nand R140_U112 U130 ; U196
g173 nand U127 P1_DATAO_REG_0__SCAN_IN ; U197
g174 nand R140_U83 U130 ; U198
g175 nand R140_U84 U127 ; U199
g176 nand U130 P2_DATAO_REG_9__SCAN_IN ; U200
g177 nand R140_U85 U127 ; U201
g178 nand U130 P2_DATAO_REG_8__SCAN_IN ; U202
g179 nand R140_U86 U127 ; U203
g180 nand U130 P2_DATAO_REG_7__SCAN_IN ; U204
g181 nand R140_U87 U127 ; U205
g182 nand U130 P2_DATAO_REG_6__SCAN_IN ; U206
g183 nand R140_U88 U127 ; U207
g184 nand U130 P2_DATAO_REG_5__SCAN_IN ; U208
g185 nand R140_U89 U127 ; U209
g186 nand U130 P2_DATAO_REG_4__SCAN_IN ; U210
g187 nand R140_U90 U127 ; U211
g188 nand U130 P2_DATAO_REG_3__SCAN_IN ; U212
g189 nand R140_U11 U127 ; U213
g190 nand U130 P2_DATAO_REG_31__SCAN_IN ; U214
g191 nand R140_U91 U127 ; U215
g192 nand U130 P2_DATAO_REG_30__SCAN_IN ; U216
g193 nand R140_U92 U127 ; U217
g194 nand U130 P2_DATAO_REG_2__SCAN_IN ; U218
g195 nand R140_U93 U127 ; U219
g196 nand U130 P2_DATAO_REG_29__SCAN_IN ; U220
g197 nand R140_U94 U127 ; U221
g198 nand U130 P2_DATAO_REG_28__SCAN_IN ; U222
g199 nand R140_U95 U127 ; U223
g200 nand U130 P2_DATAO_REG_27__SCAN_IN ; U224
g201 nand R140_U96 U127 ; U225
g202 nand U130 P2_DATAO_REG_26__SCAN_IN ; U226
g203 nand R140_U97 U127 ; U227
g204 nand U130 P2_DATAO_REG_25__SCAN_IN ; U228
g205 nand R140_U98 U127 ; U229
g206 nand U130 P2_DATAO_REG_24__SCAN_IN ; U230
g207 nand R140_U99 U127 ; U231
g208 nand U130 P2_DATAO_REG_23__SCAN_IN ; U232
g209 nand R140_U100 U127 ; U233
g210 nand U130 P2_DATAO_REG_22__SCAN_IN ; U234
g211 nand R140_U101 U127 ; U235
g212 nand U130 P2_DATAO_REG_21__SCAN_IN ; U236
g213 nand R140_U102 U127 ; U237
g214 nand U130 P2_DATAO_REG_20__SCAN_IN ; U238
g215 nand R140_U10 U127 ; U239
g216 nand U130 P2_DATAO_REG_1__SCAN_IN ; U240
g217 nand R140_U103 U127 ; U241
g218 nand U130 P2_DATAO_REG_19__SCAN_IN ; U242
g219 nand R140_U104 U127 ; U243
g220 nand U130 P2_DATAO_REG_18__SCAN_IN ; U244
g221 nand R140_U105 U127 ; U245
g222 nand U130 P2_DATAO_REG_17__SCAN_IN ; U246
g223 nand R140_U106 U127 ; U247
g224 nand U130 P2_DATAO_REG_16__SCAN_IN ; U248
g225 nand R140_U107 U127 ; U249
g226 nand U130 P2_DATAO_REG_15__SCAN_IN ; U250
g227 nand R140_U108 U127 ; U251
g228 nand U130 P2_DATAO_REG_14__SCAN_IN ; U252
g229 nand R140_U109 U127 ; U253
g230 nand U130 P2_DATAO_REG_13__SCAN_IN ; U254
g231 nand R140_U110 U127 ; U255
g232 nand U130 P2_DATAO_REG_12__SCAN_IN ; U256
g233 nand R140_U111 U127 ; U257
g234 nand U130 P2_DATAO_REG_11__SCAN_IN ; U258
g235 nand R140_U112 U127 ; U259
g236 nand U130 P2_DATAO_REG_10__SCAN_IN ; U260
g237 nand R140_U83 U127 ; U261
g238 nand U130 P2_DATAO_REG_0__SCAN_IN ; U262
g239 nand U127 P2_DATAO_REG_9__SCAN_IN ; U263
g240 nand U130 P1_DATAO_REG_9__SCAN_IN ; U264
g241 nand U127 P2_DATAO_REG_8__SCAN_IN ; U265
g242 nand U130 P1_DATAO_REG_8__SCAN_IN ; U266
g243 nand U127 P2_DATAO_REG_7__SCAN_IN ; U267
g244 nand U130 P1_DATAO_REG_7__SCAN_IN ; U268
g245 nand U127 P2_DATAO_REG_6__SCAN_IN ; U269
g246 nand U130 P1_DATAO_REG_6__SCAN_IN ; U270
g247 nand U127 P2_DATAO_REG_5__SCAN_IN ; U271
g248 nand U130 P1_DATAO_REG_5__SCAN_IN ; U272
g249 nand U127 P2_DATAO_REG_4__SCAN_IN ; U273
g250 nand U130 P1_DATAO_REG_4__SCAN_IN ; U274
g251 nand U127 P2_DATAO_REG_31__SCAN_IN ; U275
g252 nand U130 P1_DATAO_REG_31__SCAN_IN ; U276
g253 nand U127 P2_DATAO_REG_30__SCAN_IN ; U277
g254 nand U130 P1_DATAO_REG_30__SCAN_IN ; U278
g255 nand U127 P2_DATAO_REG_3__SCAN_IN ; U279
g256 nand U130 P1_DATAO_REG_3__SCAN_IN ; U280
g257 nand U127 P2_DATAO_REG_29__SCAN_IN ; U281
g258 nand U130 P1_DATAO_REG_29__SCAN_IN ; U282
g259 nand U127 P2_DATAO_REG_28__SCAN_IN ; U283
g260 nand U130 P1_DATAO_REG_28__SCAN_IN ; U284
g261 nand U127 P2_DATAO_REG_27__SCAN_IN ; U285
g262 nand U130 P1_DATAO_REG_27__SCAN_IN ; U286
g263 nand U127 P2_DATAO_REG_26__SCAN_IN ; U287
g264 nand U130 P1_DATAO_REG_26__SCAN_IN ; U288
g265 nand U127 P2_DATAO_REG_25__SCAN_IN ; U289
g266 nand U130 P1_DATAO_REG_25__SCAN_IN ; U290
g267 nand U127 P2_DATAO_REG_24__SCAN_IN ; U291
g268 nand U130 P1_DATAO_REG_24__SCAN_IN ; U292
g269 nand U127 P2_DATAO_REG_23__SCAN_IN ; U293
g270 nand U130 P1_DATAO_REG_23__SCAN_IN ; U294
g271 nand U127 P2_DATAO_REG_22__SCAN_IN ; U295
g272 nand U130 P1_DATAO_REG_22__SCAN_IN ; U296
g273 nand U127 P2_DATAO_REG_21__SCAN_IN ; U297
g274 nand U130 P1_DATAO_REG_21__SCAN_IN ; U298
g275 nand U127 P2_DATAO_REG_20__SCAN_IN ; U299
g276 nand U130 P1_DATAO_REG_20__SCAN_IN ; U300
g277 nand U127 P2_DATAO_REG_2__SCAN_IN ; U301
g278 nand U130 P1_DATAO_REG_2__SCAN_IN ; U302
g279 nand U127 P2_DATAO_REG_19__SCAN_IN ; U303
g280 nand U130 P1_DATAO_REG_19__SCAN_IN ; U304
g281 nand U127 P2_DATAO_REG_18__SCAN_IN ; U305
g282 nand U130 P1_DATAO_REG_18__SCAN_IN ; U306
g283 nand U127 P2_DATAO_REG_17__SCAN_IN ; U307
g284 nand U130 P1_DATAO_REG_17__SCAN_IN ; U308
g285 nand U127 P2_DATAO_REG_16__SCAN_IN ; U309
g286 nand U130 P1_DATAO_REG_16__SCAN_IN ; U310
g287 nand U127 P2_DATAO_REG_15__SCAN_IN ; U311
g288 nand U130 P1_DATAO_REG_15__SCAN_IN ; U312
g289 nand U127 P2_DATAO_REG_14__SCAN_IN ; U313
g290 nand U130 P1_DATAO_REG_14__SCAN_IN ; U314
g291 nand U127 P2_DATAO_REG_13__SCAN_IN ; U315
g292 nand U130 P1_DATAO_REG_13__SCAN_IN ; U316
g293 nand U127 P2_DATAO_REG_12__SCAN_IN ; U317
g294 nand U130 P1_DATAO_REG_12__SCAN_IN ; U318
g295 nand U127 P2_DATAO_REG_11__SCAN_IN ; U319
g296 nand U130 P1_DATAO_REG_11__SCAN_IN ; U320
g297 nand U127 P2_DATAO_REG_10__SCAN_IN ; U321
g298 nand U130 P1_DATAO_REG_10__SCAN_IN ; U322
g299 nand U127 P2_DATAO_REG_1__SCAN_IN ; U323
g300 nand U130 P1_DATAO_REG_1__SCAN_IN ; U324
g301 nand U127 P2_DATAO_REG_0__SCAN_IN ; U325
g302 nand U130 P1_DATAO_REG_0__SCAN_IN ; U326
g303 and P1_U3989 P1_U3444 ; P1_U3014
g304 and P1_U3450 P1_U3447 ; P1_U3015
g305 and P1_U3632 P1_U3627 ; P1_U3016
g306 and P1_U3445 P1_U3446 ; P1_U3017
g307 and P1_U5725 P1_U3445 ; P1_U3018
g308 and P1_U5722 P1_U3446 ; P1_U3019
g309 and P1_U5722 P1_U5725 ; P1_U3020
g310 and P1_U5400 P1_U3421 ; P1_U3021
g311 and P1_U3046 P1_STATE_REG_SCAN_IN ; P1_U3022
g312 and P1_U3049 P1_U5716 ; P1_U3023
g313 and P1_U3817 P1_U3423 ; P1_U3024
g314 and P1_U4020 P1_U5728 ; P1_U3025
g315 and P1_U3986 P1_U5716 ; P1_U3026
g316 and P1_U3880 P1_U4005 ; P1_U3027
g317 and P1_U3356 P1_STATE_REG_SCAN_IN ; P1_U3028
g318 and P1_U3997 P1_U4022 ; P1_U3029
g319 and P1_U4022 P1_U3422 ; P1_U3030
g320 and P1_U3990 P1_U4022 ; P1_U3031
g321 and P1_U3998 P1_U4022 ; P1_U3032
g322 and P1_U4020 P1_U3447 ; P1_U3033
g323 and P1_U4005 P1_U5728 ; P1_U3034
g324 and P1_U4022 P1_U3025 ; P1_U3035
g325 and P1_U4005 P1_U3447 ; P1_U3036
g326 and P1_U5734 P1_U4913 ; P1_U3037
g327 and P1_U3024 P1_U5734 ; P1_U3038
g328 and P1_U5728 P1_U4913 ; P1_U3039
g329 and P1_U3024 P1_U5728 ; P1_U3040
g330 and P1_U3015 P1_U4913 ; P1_U3041
g331 and P1_U3024 P1_U3015 ; P1_U3042
g332 and P1_U3022 P1_U3423 ; P1_U3043
g333 and P1_U5145 P1_STATE_REG_SCAN_IN ; P1_U3044
g334 and P1_U3022 P1_U5147 ; P1_U3045
g335 and P1_U5703 P1_U3421 ; P1_U3046
g336 and P1_U3633 P1_U3016 ; P1_U3047
g337 and P1_U5716 P1_U3443 ; P1_U3048
g338 and P1_U5710 P1_U5719 ; P1_U3049
g339 and P1_U3436 P1_U3438 ; P1_U3050
g340 nand P1_U4670 P1_U4671 P1_U4669 P1_U4672 ; P1_U3051
g341 nand P1_U4689 P1_U4690 P1_U4688 P1_U4691 ; P1_U3052
g342 nand P1_U4710 P1_U4709 P1_U4708 P1_U4707 ; P1_U3053
g343 nand P1_U4747 P1_U4748 P1_U4746 ; P1_U3054
g344 nand P1_U4651 P1_U4652 P1_U4650 P1_U4653 ; P1_U3055
g345 nand P1_U4632 P1_U4633 P1_U4631 P1_U4634 ; P1_U3056
g346 nand P1_U4727 P1_U4728 P1_U4726 ; P1_U3057
g347 nand P1_U4235 P1_U4234 P1_U4233 P1_U4232 ; P1_U3058
g348 nand P1_U4575 P1_U4576 P1_U4574 P1_U4577 ; P1_U3059
g349 nand P1_U4347 P1_U4348 P1_U4346 P1_U4349 ; P1_U3060
g350 nand P1_U4366 P1_U4367 P1_U4365 P1_U4368 ; P1_U3061
g351 nand P1_U4216 P1_U4215 P1_U4214 P1_U4213 ; P1_U3062
g352 nand P1_U4613 P1_U4614 P1_U4612 P1_U4615 ; P1_U3063
g353 nand P1_U4594 P1_U4595 P1_U4593 P1_U4596 ; P1_U3064
g354 nand P1_U4254 P1_U4253 P1_U4252 P1_U4251 ; P1_U3065
g355 nand P1_U4192 P1_U4191 P1_U4190 P1_U4189 ; P1_U3066
g356 nand P1_U4480 P1_U4481 P1_U4479 P1_U4482 ; P1_U3067
g357 nand P1_U4292 P1_U4291 P1_U4290 P1_U4289 ; P1_U3068
g358 nand P1_U4273 P1_U4272 P1_U4271 P1_U4270 ; P1_U3069
g359 nand P1_U4385 P1_U4386 P1_U4384 P1_U4387 ; P1_U3070
g360 nand P1_U4461 P1_U4462 P1_U4460 P1_U4463 ; P1_U3071
g361 nand P1_U4442 P1_U4443 P1_U4441 P1_U4444 ; P1_U3072
g362 nand P1_U4556 P1_U4557 P1_U4555 P1_U4558 ; P1_U3073
g363 nand P1_U4537 P1_U4538 P1_U4536 P1_U4539 ; P1_U3074
g364 nand P1_U4197 P1_U4196 P1_U4195 P1_U4194 ; P1_U3075
g365 nand P1_U4173 P1_U4172 P1_U4171 P1_U4170 ; P1_U3076
g366 nand P1_U4423 P1_U4424 P1_U4422 P1_U4425 ; P1_U3077
g367 nand P1_U4404 P1_U4405 P1_U4403 P1_U4406 ; P1_U3078
g368 nand P1_U4518 P1_U4519 P1_U4517 P1_U4520 ; P1_U3079
g369 nand P1_U4499 P1_U4500 P1_U4498 P1_U4501 ; P1_U3080
g370 nand P1_U4328 P1_U4329 P1_U4327 P1_U4330 ; P1_U3081
g371 nand P1_U4311 P1_U4310 P1_U4309 P1_U4308 ; P1_U3082
g372 nand P1_U4920 P1_STATE_REG_SCAN_IN ; P1_U3083
g373 not P1_STATE_REG_SCAN_IN ; P1_U3084
g374 nand P1_U5608 P1_U5607 ; P1_U3085
g375 nand P1_U5610 P1_U5609 ; P1_U3086
g376 nand P1_U5615 P1_U5614 P1_U5616 ; P1_U3087
g377 nand P1_U3923 P1_U5618 ; P1_U3088
g378 nand P1_U3924 P1_U5621 ; P1_U3089
g379 nand P1_U3925 P1_U5624 ; P1_U3090
g380 nand P1_U3926 P1_U5627 ; P1_U3091
g381 nand P1_U3927 P1_U5630 ; P1_U3092
g382 nand P1_U3928 P1_U5633 ; P1_U3093
g383 nand P1_U3929 P1_U5636 ; P1_U3094
g384 nand P1_U3930 P1_U5639 ; P1_U3095
g385 nand P1_U3931 P1_U5642 ; P1_U3096
g386 nand P1_U3933 P1_U5648 ; P1_U3097
g387 nand P1_U3934 P1_U5651 ; P1_U3098
g388 nand P1_U3935 P1_U5654 ; P1_U3099
g389 nand P1_U3936 P1_U5657 ; P1_U3100
g390 nand P1_U3937 P1_U5660 ; P1_U3101
g391 nand P1_U3938 P1_U5663 ; P1_U3102
g392 nand P1_U3939 P1_U5666 ; P1_U3103
g393 nand P1_U3940 P1_U5669 ; P1_U3104
g394 nand P1_U3941 P1_U5672 ; P1_U3105
g395 nand P1_U3942 P1_U5675 ; P1_U3106
g396 nand P1_U5590 P1_U5591 P1_U5589 ; P1_U3107
g397 nand P1_U5593 P1_U5594 P1_U5592 ; P1_U3108
g398 nand P1_U5596 P1_U5597 P1_U5595 ; P1_U3109
g399 nand P1_U5599 P1_U5600 P1_U5598 ; P1_U3110
g400 nand P1_U5602 P1_U5603 P1_U5601 ; P1_U3111
g401 nand P1_U3921 P1_U5605 ; P1_U3112
g402 nand P1_U3922 P1_U5612 ; P1_U3113
g403 nand P1_U3932 P1_U5645 ; P1_U3114
g404 nand P1_U3943 P1_U5678 ; P1_U3115
g405 nand P1_U5681 P1_U5680 ; P1_U3116
g406 nand P1_U5538 P1_U5537 ; P1_U3117
g407 nand P1_U5540 P1_U5539 ; P1_U3118
g408 nand P1_U3898 P1_U5543 ; P1_U3119
g409 nand P1_U3899 P1_U5545 ; P1_U3120
g410 nand P1_U3900 P1_U5547 ; P1_U3121
g411 nand P1_U3901 P1_U5549 ; P1_U3122
g412 nand P1_U3902 P1_U5551 ; P1_U3123
g413 nand P1_U3903 P1_U5553 ; P1_U3124
g414 nand P1_U3904 P1_U5555 ; P1_U3125
g415 nand P1_U3905 P1_U5557 ; P1_U3126
g416 nand P1_U3906 P1_U5559 ; P1_U3127
g417 nand P1_U3907 P1_U5561 ; P1_U3128
g418 nand P1_U3909 P1_U5566 ; P1_U3129
g419 nand P1_U3910 P1_U5568 ; P1_U3130
g420 nand P1_U3911 P1_U5570 ; P1_U3131
g421 nand P1_U3912 P1_U5572 ; P1_U3132
g422 nand P1_U3913 P1_U5574 ; P1_U3133
g423 nand P1_U3914 P1_U5576 ; P1_U3134
g424 nand P1_U3915 P1_U5578 ; P1_U3135
g425 nand P1_U3916 P1_U5580 ; P1_U3136
g426 nand P1_U3917 P1_U5582 ; P1_U3137
g427 nand P1_U3918 P1_U5584 ; P1_U3138
g428 nand P1_U5526 P1_U3439 P1_U5525 ; P1_U3139
g429 nand P1_U5528 P1_U3439 P1_U5527 ; P1_U3140
g430 nand P1_U5530 P1_U3439 P1_U5529 ; P1_U3141
g431 nand P1_U5532 P1_U3439 P1_U5531 ; P1_U3142
g432 nand P1_U5534 P1_U3439 P1_U5533 ; P1_U3143
g433 nand P1_U3896 P1_U5536 ; P1_U3144
g434 nand P1_U3897 P1_U5542 ; P1_U3145
g435 nand P1_U3908 P1_U5564 ; P1_U3146
g436 nand P1_U3919 P1_U5586 ; P1_U3147
g437 nand P1_U3920 P1_U5588 ; P1_U3148
g438 nand P1_U3986 P1_U3439 ; P1_U3149
g439 nand P1_U5703 P1_U3371 ; P1_U3150
g440 nand P1_U5480 P1_U5479 ; P1_U3151
g441 nand P1_U5482 P1_U5481 ; P1_U3152
g442 nand P1_U5484 P1_U5483 ; P1_U3153
g443 nand P1_U5486 P1_U5485 ; P1_U3154
g444 nand P1_U5488 P1_U5487 ; P1_U3155
g445 nand P1_U5490 P1_U5489 ; P1_U3156
g446 nand P1_U5492 P1_U5491 ; P1_U3157
g447 nand P1_U5494 P1_U5493 ; P1_U3158
g448 nand P1_U5496 P1_U5495 ; P1_U3159
g449 nand P1_U5500 P1_U5499 ; P1_U3160
g450 nand P1_U5502 P1_U5501 ; P1_U3161
g451 nand P1_U5504 P1_U5503 ; P1_U3162
g452 nand P1_U5506 P1_U5505 ; P1_U3163
g453 nand P1_U5508 P1_U5507 ; P1_U3164
g454 nand P1_U5510 P1_U5509 ; P1_U3165
g455 nand P1_U5512 P1_U5511 ; P1_U3166
g456 nand P1_U5514 P1_U5513 ; P1_U3167
g457 nand P1_U5516 P1_U5515 ; P1_U3168
g458 nand P1_U5518 P1_U5517 ; P1_U3169
g459 nand P1_U5466 P1_U5465 ; P1_U3170
g460 nand P1_U5468 P1_U5467 ; P1_U3171
g461 nand P1_U5470 P1_U5469 ; P1_U3172
g462 nand P1_U5472 P1_U5471 ; P1_U3173
g463 nand P1_U5474 P1_U5473 ; P1_U3174
g464 nand P1_U5476 P1_U5475 ; P1_U3175
g465 nand P1_U5478 P1_U5477 ; P1_U3176
g466 nand P1_U5498 P1_U5497 ; P1_U3177
g467 nand P1_U5520 P1_U5519 ; P1_U3178
g468 nand P1_U3895 P1_U5522 ; P1_U3179
g469 nand P1_U5421 P1_U5420 ; P1_U3180
g470 nand P1_U5423 P1_U5422 ; P1_U3181
g471 nand P1_U5425 P1_U5424 ; P1_U3182
g472 nand P1_U5427 P1_U5426 ; P1_U3183
g473 nand P1_U5429 P1_U5428 ; P1_U3184
g474 nand P1_U5431 P1_U5430 ; P1_U3185
g475 nand P1_U5433 P1_U5432 ; P1_U3186
g476 nand P1_U5435 P1_U5434 ; P1_U3187
g477 nand P1_U5437 P1_U5436 ; P1_U3188
g478 nand P1_U5441 P1_U5440 ; P1_U3189
g479 nand P1_U5443 P1_U5442 ; P1_U3190
g480 nand P1_U5445 P1_U5444 ; P1_U3191
g481 nand P1_U5447 P1_U5446 ; P1_U3192
g482 nand P1_U5449 P1_U5448 ; P1_U3193
g483 nand P1_U5451 P1_U5450 ; P1_U3194
g484 nand P1_U5453 P1_U5452 ; P1_U3195
g485 nand P1_U5455 P1_U5454 ; P1_U3196
g486 nand P1_U5457 P1_U5456 ; P1_U3197
g487 nand P1_U5459 P1_U5458 ; P1_U3198
g488 nand P1_U5407 P1_U5406 ; P1_U3199
g489 nand P1_U5409 P1_U5408 ; P1_U3200
g490 nand P1_U5411 P1_U5410 ; P1_U3201
g491 nand P1_U5413 P1_U5412 ; P1_U3202
g492 nand P1_U5415 P1_U5414 ; P1_U3203
g493 nand P1_U5417 P1_U5416 ; P1_U3204
g494 nand P1_U5419 P1_U5418 ; P1_U3205
g495 nand P1_U5439 P1_U5438 ; P1_U3206
g496 nand P1_U5461 P1_U5460 ; P1_U3207
g497 nand P1_U3894 P1_U5462 ; P1_U3208
g498 and P1_U5399 P1_U3421 ; P1_U3209
g499 nand P1_U6266 P1_U6265 P1_U5397 ; P1_U3210
g500 nand P1_U5391 P1_U5390 P1_U5394 P1_U5392 P1_U5393 ; P1_U3211
g501 nand P1_U5382 P1_U5381 P1_U5385 P1_U5383 P1_U5384 ; P1_U3212
g502 nand P1_U5373 P1_U5372 P1_U5376 P1_U5374 P1_U5375 ; P1_U3213
g503 nand P1_U5364 P1_U5363 P1_U5367 P1_U5365 P1_U5366 ; P1_U3214
g504 nand P1_U5355 P1_U5354 P1_U5358 P1_U5356 P1_U5357 ; P1_U3215
g505 nand P1_U3891 P1_U5346 P1_U5347 ; P1_U3216
g506 nand P1_U5337 P1_U5336 P1_U5340 P1_U5338 P1_U5339 ; P1_U3217
g507 nand P1_U5328 P1_U5327 P1_U5331 P1_U5329 P1_U5330 ; P1_U3218
g508 nand P1_U5319 P1_U5318 P1_U5322 P1_U5320 P1_U5321 ; P1_U3219
g509 nand P1_U3889 P1_U5310 P1_U5311 ; P1_U3220
g510 nand P1_U5301 P1_U5300 P1_U5304 P1_U5302 P1_U5303 ; P1_U3221
g511 nand P1_U5292 P1_U5291 P1_U5295 P1_U5293 P1_U5294 ; P1_U3222
g512 nand P1_U5283 P1_U5282 P1_U5286 P1_U5284 P1_U5285 ; P1_U3223
g513 nand P1_U5274 P1_U5273 P1_U5277 P1_U5275 P1_U5276 ; P1_U3224
g514 nand P1_U5265 P1_U5264 P1_U5266 P1_U3888 ; P1_U3225
g515 nand P1_U5256 P1_U5255 P1_U5259 P1_U5257 P1_U5258 ; P1_U3226
g516 nand P1_U5247 P1_U5246 P1_U5250 P1_U5248 P1_U5249 ; P1_U3227
g517 nand P1_U3886 P1_U5238 P1_U5239 ; P1_U3228
g518 nand P1_U5229 P1_U5228 P1_U5232 P1_U5230 P1_U5231 ; P1_U3229
g519 nand P1_U3885 P1_U5221 P1_U3884 ; P1_U3230
g520 nand P1_U5212 P1_U5211 P1_U5215 P1_U5213 P1_U5214 ; P1_U3231
g521 nand P1_U5203 P1_U5202 P1_U5206 P1_U5204 P1_U5205 ; P1_U3232
g522 nand P1_U5194 P1_U5193 P1_U5197 P1_U5195 P1_U5196 ; P1_U3233
g523 nand P1_U5185 P1_U5184 P1_U5188 P1_U5186 P1_U5187 ; P1_U3234
g524 nand P1_U3881 P1_U5176 P1_U5177 ; P1_U3235
g525 nand P1_U5167 P1_U5166 P1_U5170 P1_U5168 P1_U5169 ; P1_U3236
g526 nand P1_U5158 P1_U5157 P1_U5161 P1_U5159 P1_U5160 ; P1_U3237
g527 nand P1_U5149 P1_U5148 P1_U5152 P1_U5150 P1_U5151 ; P1_U3238
g528 nand P1_U5136 P1_U5135 P1_U5139 P1_U5137 P1_U5138 ; P1_U3239
g529 and P1_U5120 P1_U5682 ; P1_U3240
g530 nand P1_U3859 P1_U3858 ; P1_U3241
g531 nand P1_U3857 P1_U3856 ; P1_U3242
g532 nand P1_U3855 P1_U3854 ; P1_U3243
g533 nand P1_U3852 P1_U3851 ; P1_U3244
g534 nand P1_U3850 P1_U3849 ; P1_U3245
g535 nand P1_U3847 P1_U3846 ; P1_U3246
g536 nand P1_U3845 P1_U3844 ; P1_U3247
g537 nand P1_U3842 P1_U3843 P1_U5043 ; P1_U3248
g538 nand P1_U3840 P1_U3841 P1_U5033 ; P1_U3249
g539 nand P1_U3838 P1_U3839 P1_U5023 ; P1_U3250
g540 nand P1_U3836 P1_U3837 P1_U5013 ; P1_U3251
g541 nand P1_U3834 P1_U3835 P1_U5003 ; P1_U3252
g542 nand P1_U3832 P1_U3833 P1_U4993 ; P1_U3253
g543 nand P1_U3830 P1_U3831 P1_U4983 ; P1_U3254
g544 nand P1_U3828 P1_U3829 P1_U4973 ; P1_U3255
g545 nand P1_U3826 P1_U3827 P1_U4963 ; P1_U3256
g546 nand P1_U3824 P1_U3825 P1_U4953 ; P1_U3257
g547 nand P1_U3822 P1_U3823 P1_U4943 ; P1_U3258
g548 nand P1_U3820 P1_U3821 P1_U4933 ; P1_U3259
g549 nand P1_U3818 P1_U3819 P1_U4923 ; P1_U3260
g550 nand P1_U3981 P1_U4911 P1_U4912 ; P1_U3261
g551 nand P1_U3980 P1_U4909 P1_U4910 ; P1_U3262
g552 nand P1_U3811 P1_U3812 P1_U4902 P1_U3977 ; P1_U3263
g553 nand P1_U3809 P1_U3810 P1_U4897 P1_U3976 ; P1_U3264
g554 nand P1_U3807 P1_U3808 P1_U4892 P1_U3975 ; P1_U3265
g555 nand P1_U3805 P1_U3806 P1_U4887 P1_U3974 ; P1_U3266
g556 nand P1_U3803 P1_U3804 P1_U4882 P1_U3973 ; P1_U3267
g557 nand P1_U3801 P1_U3802 P1_U4877 P1_U3972 ; P1_U3268
g558 nand P1_U3799 P1_U3800 P1_U4872 P1_U3971 ; P1_U3269
g559 nand P1_U3797 P1_U3798 P1_U4867 P1_U3970 ; P1_U3270
g560 nand P1_U3795 P1_U3796 P1_U4862 P1_U3969 ; P1_U3271
g561 nand P1_U3793 P1_U3794 P1_U4857 P1_U3968 ; P1_U3272
g562 nand P1_U3792 P1_U3791 P1_U3967 ; P1_U3273
g563 nand P1_U3790 P1_U3789 P1_U3966 ; P1_U3274
g564 nand P1_U3787 P1_U3788 P1_U4842 P1_U3965 ; P1_U3275
g565 nand P1_U3785 P1_U3786 P1_U4837 P1_U3964 ; P1_U3276
g566 nand P1_U3784 P1_U3783 P1_U3963 ; P1_U3277
g567 nand P1_U3782 P1_U3781 P1_U3962 ; P1_U3278
g568 nand P1_U3780 P1_U3779 P1_U3961 ; P1_U3279
g569 nand P1_U3778 P1_U3777 P1_U3960 ; P1_U3280
g570 nand P1_U3775 P1_U3776 P1_U4812 P1_U3959 ; P1_U3281
g571 nand P1_U3773 P1_U3774 P1_U4807 P1_U3958 ; P1_U3282
g572 nand P1_U3772 P1_U3771 P1_U3957 ; P1_U3283
g573 nand P1_U3770 P1_U3769 P1_U3956 ; P1_U3284
g574 nand P1_U3768 P1_U3767 P1_U3955 ; P1_U3285
g575 nand P1_U3766 P1_U3765 P1_U3954 ; P1_U3286
g576 nand P1_U3764 P1_U3763 ; P1_U3287
g577 nand P1_U3762 P1_U3761 ; P1_U3288
g578 nand P1_U3760 P1_U3759 ; P1_U3289
g579 nand P1_U3758 P1_U3757 ; P1_U3290
g580 nand P1_U3756 P1_U3755 ; P1_U3291
g581 and P1_U3945 P1_D_REG_31__SCAN_IN ; P1_U3292
g582 and P1_U3945 P1_D_REG_30__SCAN_IN ; P1_U3293
g583 and P1_U3945 P1_D_REG_29__SCAN_IN ; P1_U3294
g584 and P1_U3945 P1_D_REG_28__SCAN_IN ; P1_U3295
g585 and P1_U3945 P1_D_REG_27__SCAN_IN ; P1_U3296
g586 and P1_U3945 P1_D_REG_26__SCAN_IN ; P1_U3297
g587 and P1_U3945 P1_D_REG_25__SCAN_IN ; P1_U3298
g588 and P1_U3945 P1_D_REG_24__SCAN_IN ; P1_U3299
g589 and P1_U3945 P1_D_REG_23__SCAN_IN ; P1_U3300
g590 and P1_U3945 P1_D_REG_22__SCAN_IN ; P1_U3301
g591 and P1_U3945 P1_D_REG_21__SCAN_IN ; P1_U3302
g592 and P1_U3945 P1_D_REG_20__SCAN_IN ; P1_U3303
g593 and P1_U3945 P1_D_REG_19__SCAN_IN ; P1_U3304
g594 and P1_U3945 P1_D_REG_18__SCAN_IN ; P1_U3305
g595 and P1_U3945 P1_D_REG_17__SCAN_IN ; P1_U3306
g596 and P1_U3945 P1_D_REG_16__SCAN_IN ; P1_U3307
g597 and P1_U3945 P1_D_REG_15__SCAN_IN ; P1_U3308
g598 and P1_U3945 P1_D_REG_14__SCAN_IN ; P1_U3309
g599 and P1_U3945 P1_D_REG_13__SCAN_IN ; P1_U3310
g600 and P1_U3945 P1_D_REG_12__SCAN_IN ; P1_U3311
g601 and P1_U3945 P1_D_REG_11__SCAN_IN ; P1_U3312
g602 and P1_U3945 P1_D_REG_10__SCAN_IN ; P1_U3313
g603 and P1_U3945 P1_D_REG_9__SCAN_IN ; P1_U3314
g604 and P1_U3945 P1_D_REG_8__SCAN_IN ; P1_U3315
g605 and P1_U3945 P1_D_REG_7__SCAN_IN ; P1_U3316
g606 and P1_U3945 P1_D_REG_6__SCAN_IN ; P1_U3317
g607 and P1_U3945 P1_D_REG_5__SCAN_IN ; P1_U3318
g608 and P1_U3945 P1_D_REG_4__SCAN_IN ; P1_U3319
g609 and P1_U3945 P1_D_REG_3__SCAN_IN ; P1_U3320
g610 and P1_U3945 P1_D_REG_2__SCAN_IN ; P1_U3321
g611 nand P1_U4132 P1_U4133 P1_U4131 ; P1_U3322
g612 nand P1_U4129 P1_U4130 P1_U4128 ; P1_U3323
g613 nand P1_U4126 P1_U4127 P1_U4125 ; P1_U3324
g614 nand P1_U4123 P1_U4124 P1_U4122 ; P1_U3325
g615 nand P1_U4120 P1_U4121 P1_U4119 ; P1_U3326
g616 nand P1_U4117 P1_U4118 P1_U4116 ; P1_U3327
g617 nand P1_U4114 P1_U4115 P1_U4113 ; P1_U3328
g618 nand P1_U4111 P1_U4112 P1_U4110 ; P1_U3329
g619 nand P1_U4108 P1_U4109 P1_U4107 ; P1_U3330
g620 nand P1_U4105 P1_U4106 P1_U4104 ; P1_U3331
g621 nand P1_U4102 P1_U4103 P1_U4101 ; P1_U3332
g622 nand P1_U4099 P1_U4100 P1_U4098 ; P1_U3333
g623 nand P1_U4096 P1_U4097 P1_U4095 ; P1_U3334
g624 nand P1_U4093 P1_U4094 P1_U4092 ; P1_U3335
g625 nand P1_U4090 P1_U4091 P1_U4089 ; P1_U3336
g626 nand P1_U4087 P1_U4088 P1_U4086 ; P1_U3337
g627 nand P1_U4084 P1_U4085 P1_U4083 ; P1_U3338
g628 nand P1_U4081 P1_U4082 P1_U4080 ; P1_U3339
g629 nand P1_U4078 P1_U4079 P1_U4077 ; P1_U3340
g630 nand P1_U4075 P1_U4076 P1_U4074 ; P1_U3341
g631 nand P1_U4072 P1_U4073 P1_U4071 ; P1_U3342
g632 nand P1_U4069 P1_U4070 P1_U4068 ; P1_U3343
g633 nand P1_U4066 P1_U4067 P1_U4065 ; P1_U3344
g634 nand P1_U4063 P1_U4064 P1_U4062 ; P1_U3345
g635 nand P1_U4060 P1_U4061 P1_U4059 ; P1_U3346
g636 nand P1_U4057 P1_U4058 P1_U4056 ; P1_U3347
g637 nand P1_U4054 P1_U4055 P1_U4053 ; P1_U3348
g638 nand P1_U4051 P1_U4052 P1_U4050 ; P1_U3349
g639 nand P1_U4048 P1_U4049 P1_U4047 ; P1_U3350
g640 nand P1_U4045 P1_U4046 P1_U4044 ; P1_U3351
g641 nand P1_U4042 P1_U4043 P1_U4041 ; P1_U3352
g642 nand P1_U4039 P1_U4040 P1_U4038 ; P1_U3353
g643 and P1_U3443 P1_U3439 ; P1_U3354
g644 nand P1_U4907 P1_U4905 P1_U4908 P1_U4906 P1_U3978 ; P1_U3355
g645 nand P1_U3944 P1_STATE_REG_SCAN_IN ; P1_U3356
g646 nand P1_U3438 P1_U5695 ; P1_U3357
g647 not P1_B_REG_SCAN_IN ; P1_U3358
g648 nand P1_U5700 P1_U5699 P1_U3438 ; P1_U3359
g649 nand P1_U3048 P1_U3444 ; P1_U3360
g650 nand P1_U3442 P1_U3443 P1_U3444 ; P1_U3361
g651 nand P1_U3442 P1_U5713 ; P1_U3362
g652 nand P1_U4034 P1_U3444 ; P1_U3363
g653 nand P1_U3442 P1_U3443 P1_U3448 ; P1_U3364
g654 nand P1_U4034 P1_U3448 ; P1_U3365
g655 nand P1_U5716 P1_U5713 ; P1_U3366
g656 nand P1_U4035 P1_U3444 ; P1_U3367
g657 nand P1_U3993 P1_U5719 ; P1_U3368
g658 nand P1_U4035 P1_U3448 ; P1_U3369
g659 nand P1_U3989 P1_U5710 ; P1_U3370
g660 nand P1_U5710 P1_U3443 ; P1_U3371
g661 nand P1_U3444 P1_U3448 ; P1_U3372
g662 nand P1_U4181 P1_U4180 P1_U4182 P1_U3620 P1_U3619 ; P1_U3373
g663 not P1_REG2_REG_0__SCAN_IN ; P1_U3374
g664 nand P1_U4200 P1_U4199 P1_U3635 P1_U3637 ; P1_U3375
g665 nand P1_U4219 P1_U4218 P1_U3639 P1_U3641 ; P1_U3376
g666 nand P1_U4238 P1_U4237 P1_U3643 P1_U3645 ; P1_U3377
g667 nand P1_U4257 P1_U4256 P1_U3647 P1_U3649 ; P1_U3378
g668 nand P1_U4276 P1_U4275 P1_U3651 P1_U3653 ; P1_U3379
g669 nand P1_U4295 P1_U4294 P1_U3655 P1_U3657 ; P1_U3380
g670 nand P1_U4314 P1_U4313 P1_U3659 P1_U3661 ; P1_U3381
g671 nand P1_U4333 P1_U4332 P1_U3663 P1_U3665 ; P1_U3382
g672 nand P1_U4352 P1_U4351 P1_U3667 P1_U3669 ; P1_U3383
g673 nand P1_U4371 P1_U4370 P1_U3671 P1_U3673 ; P1_U3384
g674 nand P1_U4390 P1_U4389 P1_U3675 P1_U3677 ; P1_U3385
g675 nand P1_U4409 P1_U4408 P1_U3679 P1_U3681 ; P1_U3386
g676 nand P1_U4428 P1_U4427 P1_U3683 P1_U3685 ; P1_U3387
g677 nand P1_U4447 P1_U4446 P1_U3687 P1_U3689 ; P1_U3388
g678 nand P1_U4466 P1_U4465 P1_U3691 P1_U3693 ; P1_U3389
g679 nand P1_U4485 P1_U4484 P1_U3695 P1_U3697 ; P1_U3390
g680 nand P1_U4504 P1_U4503 P1_U3699 P1_U3701 ; P1_U3391
g681 nand P1_U4523 P1_U4522 P1_U3703 P1_U3705 ; P1_U3392
g682 nand P1_U4542 P1_U4541 P1_U3707 P1_U3709 ; P1_U3393
g683 nand U76 P1_U3946 ; P1_U3394
g684 nand P1_U4561 P1_U4560 P1_U3711 P1_U3713 ; P1_U3395
g685 nand U75 P1_U3946 ; P1_U3396
g686 nand P1_U4580 P1_U4579 P1_U3715 P1_U3717 ; P1_U3397
g687 nand U74 P1_U3946 ; P1_U3398
g688 nand P1_U4599 P1_U4598 P1_U3719 P1_U3721 ; P1_U3399
g689 nand U73 P1_U3946 ; P1_U3400
g690 nand P1_U4618 P1_U4617 P1_U3723 P1_U3725 ; P1_U3401
g691 nand U72 P1_U3946 ; P1_U3402
g692 nand P1_U4637 P1_U4636 P1_U3727 P1_U3729 ; P1_U3403
g693 nand U71 P1_U3946 ; P1_U3404
g694 nand P1_U4656 P1_U4655 P1_U3731 P1_U3733 ; P1_U3405
g695 nand U70 P1_U3946 ; P1_U3406
g696 nand P1_U4675 P1_U4674 P1_U3735 P1_U3737 ; P1_U3407
g697 nand U69 P1_U3946 ; P1_U3408
g698 nand P1_U4694 P1_U4693 P1_U3739 P1_U3741 ; P1_U3409
g699 nand U68 P1_U3946 ; P1_U3410
g700 nand P1_U4713 P1_U4712 P1_U3743 P1_U3745 ; P1_U3411
g701 nand U67 P1_U3946 ; P1_U3412
g702 nand P1_U3750 P1_U3748 ; P1_U3413
g703 nand U65 P1_U3946 ; P1_U3414
g704 nand U64 P1_U3946 ; P1_U3415
g705 nand P1_U3986 P1_U5719 ; P1_U3416
g706 nand P1_U3022 P1_U4757 ; P1_U3417
g707 nand P1_U4021 P1_U5716 ; P1_U3418
g708 nand P1_U3048 P1_U3448 ; P1_U3419
g709 nand P1_U3023 P1_U5713 ; P1_U3420
g710 nand P1_U3050 P1_U3437 ; P1_U3421
g711 nand P1_U3999 P1_U4758 ; P1_U3422
g712 nand P1_U3424 P1_U4921 ; P1_U3423
g713 nand P1_U4135 P1_U5703 ; P1_U3424
g714 nand P1_U4032 P1_STATE_REG_SCAN_IN ; P1_U3425
g715 nand P1_U3444 P1_U3439 ; P1_U3426
g716 nand P1_U3014 P1_U3015 ; P1_U3427
g717 nand P1_U3439 P1_U5713 ; P1_U3428
g718 not P1_R1375_U14 ; P1_U3429
g719 nand P1_U3022 P1_U3422 ; P1_U3430
g720 nand P1_U3876 P1_U3016 ; P1_U3431
g721 nand P1_U3014 P1_U3022 ; P1_U3432
g722 nand P1_U3879 P1_U5133 ; P1_U3433
g723 nand P1_U3443 P1_U5719 ; P1_U3434
g724 nand P1_U5403 P1_U5402 ; P1_U3435
g725 nand P1_U5691 P1_U5690 ; P1_U3436
g726 nand P1_U5694 P1_U5693 ; P1_U3437
g727 nand P1_U5697 P1_U5696 ; P1_U3438
g728 nand P1_U5702 P1_U5701 ; P1_U3439
g729 nand P1_U5705 P1_U5704 ; P1_U3440
g730 nand P1_U5707 P1_U5706 ; P1_U3441
g731 nand P1_U5715 P1_U5714 ; P1_U3442
g732 nand P1_U5712 P1_U5711 ; P1_U3443
g733 nand P1_U5709 P1_U5708 ; P1_U3444
g734 nand P1_U5721 P1_U5720 ; P1_U3445
g735 nand P1_U5724 P1_U5723 ; P1_U3446
g736 nand P1_U5727 P1_U5726 ; P1_U3447
g737 nand P1_U5718 P1_U5717 ; P1_U3448
g738 nand P1_U5730 P1_U5729 ; P1_U3449
g739 nand P1_U5733 P1_U5732 ; P1_U3450
g740 nand P1_U5736 P1_U5735 ; P1_U3451
g741 nand P1_U5744 P1_U5743 ; P1_U3452
g742 nand P1_U5741 P1_U5740 ; P1_U3453
g743 nand P1_U5747 P1_U5746 ; P1_U3454
g744 nand P1_U5749 P1_U5748 ; P1_U3455
g745 nand P1_U5751 P1_U5750 ; P1_U3456
g746 nand P1_U5754 P1_U5753 ; P1_U3457
g747 nand P1_U5756 P1_U5755 ; P1_U3458
g748 nand P1_U5758 P1_U5757 ; P1_U3459
g749 nand P1_U5761 P1_U5760 ; P1_U3460
g750 nand P1_U5763 P1_U5762 ; P1_U3461
g751 nand P1_U5765 P1_U5764 ; P1_U3462
g752 nand P1_U5768 P1_U5767 ; P1_U3463
g753 nand P1_U5770 P1_U5769 ; P1_U3464
g754 nand P1_U5772 P1_U5771 ; P1_U3465
g755 nand P1_U5775 P1_U5774 ; P1_U3466
g756 nand P1_U5777 P1_U5776 ; P1_U3467
g757 nand P1_U5779 P1_U5778 ; P1_U3468
g758 nand P1_U5782 P1_U5781 ; P1_U3469
g759 nand P1_U5784 P1_U5783 ; P1_U3470
g760 nand P1_U5786 P1_U5785 ; P1_U3471
g761 nand P1_U5789 P1_U5788 ; P1_U3472
g762 nand P1_U5791 P1_U5790 ; P1_U3473
g763 nand P1_U5793 P1_U5792 ; P1_U3474
g764 nand P1_U5796 P1_U5795 ; P1_U3475
g765 nand P1_U5798 P1_U5797 ; P1_U3476
g766 nand P1_U5800 P1_U5799 ; P1_U3477
g767 nand P1_U5803 P1_U5802 ; P1_U3478
g768 nand P1_U5805 P1_U5804 ; P1_U3479
g769 nand P1_U5807 P1_U5806 ; P1_U3480
g770 nand P1_U5810 P1_U5809 ; P1_U3481
g771 nand P1_U5812 P1_U5811 ; P1_U3482
g772 nand P1_U5814 P1_U5813 ; P1_U3483
g773 nand P1_U5817 P1_U5816 ; P1_U3484
g774 nand P1_U5819 P1_U5818 ; P1_U3485
g775 nand P1_U5821 P1_U5820 ; P1_U3486
g776 nand P1_U5824 P1_U5823 ; P1_U3487
g777 nand P1_U5826 P1_U5825 ; P1_U3488
g778 nand P1_U5828 P1_U5827 ; P1_U3489
g779 nand P1_U5831 P1_U5830 ; P1_U3490
g780 nand P1_U5833 P1_U5832 ; P1_U3491
g781 nand P1_U5835 P1_U5834 ; P1_U3492
g782 nand P1_U5838 P1_U5837 ; P1_U3493
g783 nand P1_U5840 P1_U5839 ; P1_U3494
g784 nand P1_U5842 P1_U5841 ; P1_U3495
g785 nand P1_U5845 P1_U5844 ; P1_U3496
g786 nand P1_U5847 P1_U5846 ; P1_U3497
g787 nand P1_U5849 P1_U5848 ; P1_U3498
g788 nand P1_U5852 P1_U5851 ; P1_U3499
g789 nand P1_U5854 P1_U5853 ; P1_U3500
g790 nand P1_U5856 P1_U5855 ; P1_U3501
g791 nand P1_U5859 P1_U5858 ; P1_U3502
g792 nand P1_U5861 P1_U5860 ; P1_U3503
g793 nand P1_U5863 P1_U5862 ; P1_U3504
g794 nand P1_U5866 P1_U5865 ; P1_U3505
g795 nand P1_U5868 P1_U5867 ; P1_U3506
g796 nand P1_U5870 P1_U5869 ; P1_U3507
g797 nand P1_U5873 P1_U5872 ; P1_U3508
g798 nand P1_U5875 P1_U5874 ; P1_U3509
g799 nand P1_U5878 P1_U5877 ; P1_U3510
g800 nand P1_U5880 P1_U5879 ; P1_U3511
g801 nand P1_U5882 P1_U5881 ; P1_U3512
g802 nand P1_U5884 P1_U5883 ; P1_U3513
g803 nand P1_U5886 P1_U5885 ; P1_U3514
g804 nand P1_U5888 P1_U5887 ; P1_U3515
g805 nand P1_U5890 P1_U5889 ; P1_U3516
g806 nand P1_U5892 P1_U5891 ; P1_U3517
g807 nand P1_U5894 P1_U5893 ; P1_U3518
g808 nand P1_U5896 P1_U5895 ; P1_U3519
g809 nand P1_U5898 P1_U5897 ; P1_U3520
g810 nand P1_U5900 P1_U5899 ; P1_U3521
g811 nand P1_U5902 P1_U5901 ; P1_U3522
g812 nand P1_U5904 P1_U5903 ; P1_U3523
g813 nand P1_U5906 P1_U5905 ; P1_U3524
g814 nand P1_U5908 P1_U5907 ; P1_U3525
g815 nand P1_U5910 P1_U5909 ; P1_U3526
g816 nand P1_U5912 P1_U5911 ; P1_U3527
g817 nand P1_U5914 P1_U5913 ; P1_U3528
g818 nand P1_U5916 P1_U5915 ; P1_U3529
g819 nand P1_U5918 P1_U5917 ; P1_U3530
g820 nand P1_U5920 P1_U5919 ; P1_U3531
g821 nand P1_U5922 P1_U5921 ; P1_U3532
g822 nand P1_U5924 P1_U5923 ; P1_U3533
g823 nand P1_U5926 P1_U5925 ; P1_U3534
g824 nand P1_U5928 P1_U5927 ; P1_U3535
g825 nand P1_U5930 P1_U5929 ; P1_U3536
g826 nand P1_U5932 P1_U5931 ; P1_U3537
g827 nand P1_U5934 P1_U5933 ; P1_U3538
g828 nand P1_U5936 P1_U5935 ; P1_U3539
g829 nand P1_U5938 P1_U5937 ; P1_U3540
g830 nand P1_U5940 P1_U5939 ; P1_U3541
g831 nand P1_U5942 P1_U5941 ; P1_U3542
g832 nand P1_U5944 P1_U5943 ; P1_U3543
g833 nand P1_U5946 P1_U5945 ; P1_U3544
g834 nand P1_U5948 P1_U5947 ; P1_U3545
g835 nand P1_U5950 P1_U5949 ; P1_U3546
g836 nand P1_U5952 P1_U5951 ; P1_U3547
g837 nand P1_U5954 P1_U5953 ; P1_U3548
g838 nand P1_U5956 P1_U5955 ; P1_U3549
g839 nand P1_U5958 P1_U5957 ; P1_U3550
g840 nand P1_U5960 P1_U5959 ; P1_U3551
g841 nand P1_U5962 P1_U5961 ; P1_U3552
g842 nand P1_U5964 P1_U5963 ; P1_U3553
g843 nand P1_U5966 P1_U5965 ; P1_U3554
g844 nand P1_U6032 P1_U6031 ; P1_U3555
g845 nand P1_U6034 P1_U6033 ; P1_U3556
g846 nand P1_U6036 P1_U6035 ; P1_U3557
g847 nand P1_U6038 P1_U6037 ; P1_U3558
g848 nand P1_U6040 P1_U6039 ; P1_U3559
g849 nand P1_U6042 P1_U6041 ; P1_U3560
g850 nand P1_U6044 P1_U6043 ; P1_U3561
g851 nand P1_U6046 P1_U6045 ; P1_U3562
g852 nand P1_U6048 P1_U6047 ; P1_U3563
g853 nand P1_U6050 P1_U6049 ; P1_U3564
g854 nand P1_U6052 P1_U6051 ; P1_U3565
g855 nand P1_U6054 P1_U6053 ; P1_U3566
g856 nand P1_U6056 P1_U6055 ; P1_U3567
g857 nand P1_U6058 P1_U6057 ; P1_U3568
g858 nand P1_U6060 P1_U6059 ; P1_U3569
g859 nand P1_U6062 P1_U6061 ; P1_U3570
g860 nand P1_U6064 P1_U6063 ; P1_U3571
g861 nand P1_U6066 P1_U6065 ; P1_U3572
g862 nand P1_U6068 P1_U6067 ; P1_U3573
g863 nand P1_U6070 P1_U6069 ; P1_U3574
g864 nand P1_U6072 P1_U6071 ; P1_U3575
g865 nand P1_U6074 P1_U6073 ; P1_U3576
g866 nand P1_U6076 P1_U6075 ; P1_U3577
g867 nand P1_U6078 P1_U6077 ; P1_U3578
g868 nand P1_U6080 P1_U6079 ; P1_U3579
g869 nand P1_U6082 P1_U6081 ; P1_U3580
g870 nand P1_U6084 P1_U6083 ; P1_U3581
g871 nand P1_U6086 P1_U6085 ; P1_U3582
g872 nand P1_U6088 P1_U6087 ; P1_U3583
g873 nand P1_U6090 P1_U6089 ; P1_U3584
g874 nand P1_U6092 P1_U6091 ; P1_U3585
g875 nand P1_U6094 P1_U6093 ; P1_U3586
g876 nand P1_U6202 P1_U6201 ; P1_U3587
g877 nand P1_U6204 P1_U6203 ; P1_U3588
g878 nand P1_U6206 P1_U6205 ; P1_U3589
g879 nand P1_U6208 P1_U6207 ; P1_U3590
g880 nand P1_U6210 P1_U6209 ; P1_U3591
g881 nand P1_U6212 P1_U6211 ; P1_U3592
g882 nand P1_U6214 P1_U6213 ; P1_U3593
g883 nand P1_U6216 P1_U6215 ; P1_U3594
g884 nand P1_U6218 P1_U6217 ; P1_U3595
g885 nand P1_U6220 P1_U6219 ; P1_U3596
g886 nand P1_U6222 P1_U6221 ; P1_U3597
g887 nand P1_U6224 P1_U6223 ; P1_U3598
g888 nand P1_U6226 P1_U6225 ; P1_U3599
g889 nand P1_U6228 P1_U6227 ; P1_U3600
g890 nand P1_U6230 P1_U6229 ; P1_U3601
g891 nand P1_U6232 P1_U6231 ; P1_U3602
g892 nand P1_U6234 P1_U6233 ; P1_U3603
g893 nand P1_U6236 P1_U6235 ; P1_U3604
g894 nand P1_U6238 P1_U6237 ; P1_U3605
g895 nand P1_U6240 P1_U6239 ; P1_U3606
g896 nand P1_U6242 P1_U6241 ; P1_U3607
g897 nand P1_U6244 P1_U6243 ; P1_U3608
g898 nand P1_U6246 P1_U6245 ; P1_U3609
g899 nand P1_U6248 P1_U6247 ; P1_U3610
g900 nand P1_U6250 P1_U6249 ; P1_U3611
g901 nand P1_U6252 P1_U6251 ; P1_U3612
g902 nand P1_U6254 P1_U6253 ; P1_U3613
g903 nand P1_U6256 P1_U6255 ; P1_U3614
g904 nand P1_U6258 P1_U6257 ; P1_U3615
g905 nand P1_U6260 P1_U6259 ; P1_U3616
g906 nand P1_U6262 P1_U6261 ; P1_U3617
g907 nand P1_U6264 P1_U6263 ; P1_U3618
g908 and P1_U4177 P1_U4176 ; P1_U3619
g909 and P1_U4179 P1_U4178 ; P1_U3620
g910 and P1_U4186 P1_U4184 ; P1_U3621
g911 and P1_U4187 P1_U4185 P1_U3621 ; P1_U3622
g912 and P1_U4141 P1_U4140 P1_U4139 P1_U4138 ; P1_U3623
g913 and P1_U4145 P1_U4144 P1_U4143 P1_U4142 ; P1_U3624
g914 and P1_U4149 P1_U4148 P1_U4147 P1_U4146 ; P1_U3625
g915 and P1_U4151 P1_U4150 P1_U4152 ; P1_U3626
g916 and P1_U3626 P1_U3625 P1_U3624 P1_U3623 ; P1_U3627
g917 and P1_U4156 P1_U4155 P1_U4154 P1_U4153 ; P1_U3628
g918 and P1_U4160 P1_U4159 P1_U4158 P1_U4157 ; P1_U3629
g919 and P1_U4164 P1_U4163 P1_U4162 P1_U4161 ; P1_U3630
g920 and P1_U4166 P1_U4165 P1_U4167 ; P1_U3631
g921 and P1_U3631 P1_U3630 P1_U3629 P1_U3628 ; P1_U3632
g922 and P1_U5742 P1_U4169 ; P1_U3633
g923 and P1_U5745 P1_U3022 ; P1_U3634
g924 and P1_U4202 P1_U4201 ; P1_U3635
g925 and P1_U4204 P1_U4203 ; P1_U3636
g926 and P1_U4206 P1_U4205 P1_U3636 ; P1_U3637
g927 and P1_U4209 P1_U4210 P1_U4211 P1_U4208 ; P1_U3638
g928 and P1_U4221 P1_U4220 ; P1_U3639
g929 and P1_U4223 P1_U4222 ; P1_U3640
g930 and P1_U4225 P1_U4224 P1_U3640 ; P1_U3641
g931 and P1_U4228 P1_U4229 P1_U4230 P1_U4227 ; P1_U3642
g932 and P1_U4240 P1_U4239 ; P1_U3643
g933 and P1_U4242 P1_U4241 ; P1_U3644
g934 and P1_U4244 P1_U4243 P1_U3644 ; P1_U3645
g935 and P1_U4247 P1_U4248 P1_U4249 P1_U4246 ; P1_U3646
g936 and P1_U4259 P1_U4258 ; P1_U3647
g937 and P1_U4261 P1_U4260 ; P1_U3648
g938 and P1_U4263 P1_U4262 P1_U3648 ; P1_U3649
g939 and P1_U4266 P1_U4267 P1_U4268 P1_U4265 ; P1_U3650
g940 and P1_U4278 P1_U4277 ; P1_U3651
g941 and P1_U4280 P1_U4279 ; P1_U3652
g942 and P1_U4282 P1_U4281 P1_U3652 ; P1_U3653
g943 and P1_U4285 P1_U4286 P1_U4287 P1_U4284 ; P1_U3654
g944 and P1_U4297 P1_U4296 ; P1_U3655
g945 and P1_U4299 P1_U4298 ; P1_U3656
g946 and P1_U4301 P1_U4300 P1_U3656 ; P1_U3657
g947 and P1_U4304 P1_U4305 P1_U4306 P1_U4303 ; P1_U3658
g948 and P1_U4316 P1_U4315 ; P1_U3659
g949 and P1_U4318 P1_U4317 ; P1_U3660
g950 and P1_U4320 P1_U4319 P1_U3660 ; P1_U3661
g951 and P1_U4323 P1_U4324 P1_U4325 P1_U4322 ; P1_U3662
g952 and P1_U4335 P1_U4334 ; P1_U3663
g953 and P1_U4337 P1_U4336 ; P1_U3664
g954 and P1_U4339 P1_U4338 P1_U3664 ; P1_U3665
g955 and P1_U4342 P1_U4343 P1_U4344 P1_U4341 ; P1_U3666
g956 and P1_U4354 P1_U4353 ; P1_U3667
g957 and P1_U4356 P1_U4355 ; P1_U3668
g958 and P1_U4358 P1_U4357 P1_U3668 ; P1_U3669
g959 and P1_U4361 P1_U4362 P1_U4363 P1_U4360 ; P1_U3670
g960 and P1_U4373 P1_U4372 ; P1_U3671
g961 and P1_U4375 P1_U4374 ; P1_U3672
g962 and P1_U4377 P1_U4376 P1_U3672 ; P1_U3673
g963 and P1_U4380 P1_U4381 P1_U4382 P1_U4379 ; P1_U3674
g964 and P1_U4392 P1_U4391 ; P1_U3675
g965 and P1_U4394 P1_U4393 ; P1_U3676
g966 and P1_U4396 P1_U4395 P1_U3676 ; P1_U3677
g967 and P1_U4401 P1_U4400 P1_U4399 P1_U4398 ; P1_U3678
g968 and P1_U4411 P1_U4410 ; P1_U3679
g969 and P1_U4413 P1_U4412 ; P1_U3680
g970 and P1_U4415 P1_U4414 P1_U3680 ; P1_U3681
g971 and P1_U4420 P1_U4419 P1_U4418 P1_U4417 ; P1_U3682
g972 and P1_U4430 P1_U4429 ; P1_U3683
g973 and P1_U4432 P1_U4431 ; P1_U3684
g974 and P1_U4434 P1_U4433 P1_U3684 ; P1_U3685
g975 and P1_U4439 P1_U4438 P1_U4437 P1_U4436 ; P1_U3686
g976 and P1_U4449 P1_U4448 ; P1_U3687
g977 and P1_U4451 P1_U4450 ; P1_U3688
g978 and P1_U4453 P1_U4452 P1_U3688 ; P1_U3689
g979 and P1_U4458 P1_U4455 P1_U4456 P1_U4457 ; P1_U3690
g980 and P1_U4468 P1_U4467 ; P1_U3691
g981 and P1_U4470 P1_U4469 ; P1_U3692
g982 and P1_U4472 P1_U4471 P1_U3692 ; P1_U3693
g983 and P1_U4475 P1_U4476 P1_U4477 P1_U4474 ; P1_U3694
g984 and P1_U4487 P1_U4486 ; P1_U3695
g985 and P1_U4489 P1_U4488 ; P1_U3696
g986 and P1_U4491 P1_U4490 P1_U3696 ; P1_U3697
g987 and P1_U4494 P1_U4495 P1_U4496 P1_U4493 ; P1_U3698
g988 and P1_U4506 P1_U4505 ; P1_U3699
g989 and P1_U4508 P1_U4507 ; P1_U3700
g990 and P1_U4510 P1_U4509 P1_U3700 ; P1_U3701
g991 and P1_U4515 P1_U4512 P1_U4513 P1_U4514 ; P1_U3702
g992 and P1_U4525 P1_U4524 ; P1_U3703
g993 and P1_U4527 P1_U4526 ; P1_U3704
g994 and P1_U4529 P1_U4528 P1_U3704 ; P1_U3705
g995 and P1_U4534 P1_U4531 P1_U4532 P1_U4533 ; P1_U3706
g996 and P1_U4544 P1_U4543 ; P1_U3707
g997 and P1_U4546 P1_U4545 ; P1_U3708
g998 and P1_U4548 P1_U4547 P1_U3708 ; P1_U3709
g999 and P1_U4551 P1_U4552 P1_U4553 P1_U4550 ; P1_U3710
g1000 and P1_U4563 P1_U4562 ; P1_U3711
g1001 and P1_U4565 P1_U4564 ; P1_U3712
g1002 and P1_U4567 P1_U4566 P1_U3712 ; P1_U3713
g1003 and P1_U4570 P1_U4571 P1_U4572 P1_U4569 ; P1_U3714
g1004 and P1_U4582 P1_U4581 ; P1_U3715
g1005 and P1_U4584 P1_U4583 ; P1_U3716
g1006 and P1_U4586 P1_U4585 P1_U3716 ; P1_U3717
g1007 and P1_U4589 P1_U4590 P1_U4591 P1_U4588 ; P1_U3718
g1008 and P1_U4601 P1_U4600 ; P1_U3719
g1009 and P1_U4603 P1_U4602 ; P1_U3720
g1010 and P1_U4605 P1_U4604 P1_U3720 ; P1_U3721
g1011 and P1_U4608 P1_U4609 P1_U4610 P1_U4607 ; P1_U3722
g1012 and P1_U4620 P1_U4619 ; P1_U3723
g1013 and P1_U4622 P1_U4621 ; P1_U3724
g1014 and P1_U4624 P1_U4623 P1_U3724 ; P1_U3725
g1015 and P1_U4627 P1_U4628 P1_U4629 P1_U4626 ; P1_U3726
g1016 and P1_U4639 P1_U4638 ; P1_U3727
g1017 and P1_U4641 P1_U4640 ; P1_U3728
g1018 and P1_U4643 P1_U4642 P1_U3728 ; P1_U3729
g1019 and P1_U4646 P1_U4647 P1_U4648 P1_U4645 ; P1_U3730
g1020 and P1_U4658 P1_U4657 ; P1_U3731
g1021 and P1_U4660 P1_U4659 ; P1_U3732
g1022 and P1_U4662 P1_U4661 P1_U3732 ; P1_U3733
g1023 and P1_U4665 P1_U4666 P1_U4667 P1_U4664 ; P1_U3734
g1024 and P1_U4677 P1_U4676 ; P1_U3735
g1025 and P1_U4679 P1_U4678 ; P1_U3736
g1026 and P1_U4681 P1_U4680 P1_U3736 ; P1_U3737
g1027 and P1_U4684 P1_U4685 P1_U4686 P1_U4683 ; P1_U3738
g1028 and P1_U4696 P1_U4695 ; P1_U3739
g1029 and P1_U4698 P1_U4697 ; P1_U3740
g1030 and P1_U4700 P1_U4699 P1_U3740 ; P1_U3741
g1031 and P1_U4703 P1_U4704 P1_U4705 P1_U4702 ; P1_U3742
g1032 and P1_U4715 P1_U4714 ; P1_U3743
g1033 and P1_U4717 P1_U4716 ; P1_U3744
g1034 and P1_U4719 P1_U4718 P1_U3744 ; P1_U3745
g1035 and P1_U4722 P1_U4723 P1_U4724 P1_U4721 ; P1_U3746
g1036 and P1_U4731 P1_U4020 ; P1_U3747
g1037 and P1_U4733 P1_U4732 P1_U4734 P1_U4735 P1_U4736 ; P1_U3748
g1038 and P1_U4738 P1_U4737 ; P1_U3749
g1039 and P1_U4740 P1_U4739 P1_U3749 ; P1_U3750
g1040 and P1_U4743 P1_U4744 P1_U4742 ; P1_U3751
g1041 and P1_U4020 P1_U4731 ; P1_U3752
g1042 and P1_U3022 P1_U3452 ; P1_U3753
g1043 and P1_U5745 P1_U4002 P1_U3453 ; P1_U3754
g1044 and P1_U4761 P1_U4760 P1_U4762 ; P1_U3755
g1045 and P1_U4764 P1_U4763 P1_U3949 ; P1_U3756
g1046 and P1_U4766 P1_U4765 P1_U4767 ; P1_U3757
g1047 and P1_U4769 P1_U4768 P1_U3950 ; P1_U3758
g1048 and P1_U4771 P1_U4770 P1_U4772 ; P1_U3759
g1049 and P1_U4774 P1_U4773 P1_U3951 ; P1_U3760
g1050 and P1_U4776 P1_U4775 P1_U4777 ; P1_U3761
g1051 and P1_U4779 P1_U4778 P1_U3952 ; P1_U3762
g1052 and P1_U4781 P1_U4780 P1_U4782 ; P1_U3763
g1053 and P1_U4784 P1_U4783 P1_U3953 ; P1_U3764
g1054 and P1_U4786 P1_U4785 P1_U4787 ; P1_U3765
g1055 and P1_U4789 P1_U4788 ; P1_U3766
g1056 and P1_U4791 P1_U4790 P1_U4792 ; P1_U3767
g1057 and P1_U4794 P1_U4793 ; P1_U3768
g1058 and P1_U4796 P1_U4795 P1_U4797 ; P1_U3769
g1059 and P1_U4799 P1_U4798 ; P1_U3770
g1060 and P1_U4801 P1_U4800 P1_U4802 ; P1_U3771
g1061 and P1_U4804 P1_U4803 ; P1_U3772
g1062 and P1_U4806 P1_U4805 ; P1_U3773
g1063 and P1_U4809 P1_U4808 ; P1_U3774
g1064 and P1_U4811 P1_U4810 ; P1_U3775
g1065 and P1_U4814 P1_U4813 ; P1_U3776
g1066 and P1_U4816 P1_U4815 P1_U4817 ; P1_U3777
g1067 and P1_U4819 P1_U4818 ; P1_U3778
g1068 and P1_U4821 P1_U4820 P1_U4822 ; P1_U3779
g1069 and P1_U4824 P1_U4823 ; P1_U3780
g1070 and P1_U4826 P1_U4825 P1_U4827 ; P1_U3781
g1071 and P1_U4829 P1_U4828 ; P1_U3782
g1072 and P1_U4831 P1_U4830 P1_U4832 ; P1_U3783
g1073 and P1_U4834 P1_U4833 ; P1_U3784
g1074 and P1_U4836 P1_U4835 ; P1_U3785
g1075 and P1_U4839 P1_U4838 ; P1_U3786
g1076 and P1_U4841 P1_U4840 ; P1_U3787
g1077 and P1_U4844 P1_U4843 ; P1_U3788
g1078 and P1_U4846 P1_U4845 P1_U4847 ; P1_U3789
g1079 and P1_U4849 P1_U4848 ; P1_U3790
g1080 and P1_U4851 P1_U4850 P1_U4852 ; P1_U3791
g1081 and P1_U4854 P1_U4853 ; P1_U3792
g1082 and P1_U4856 P1_U4855 ; P1_U3793
g1083 and P1_U4859 P1_U4858 ; P1_U3794
g1084 and P1_U4861 P1_U4860 ; P1_U3795
g1085 and P1_U4864 P1_U4863 ; P1_U3796
g1086 and P1_U4866 P1_U4865 ; P1_U3797
g1087 and P1_U4869 P1_U4868 ; P1_U3798
g1088 and P1_U4871 P1_U4870 ; P1_U3799
g1089 and P1_U4874 P1_U4873 ; P1_U3800
g1090 and P1_U4876 P1_U4875 ; P1_U3801
g1091 and P1_U4879 P1_U4878 ; P1_U3802
g1092 and P1_U4881 P1_U4880 ; P1_U3803
g1093 and P1_U4884 P1_U4883 ; P1_U3804
g1094 and P1_U4886 P1_U4885 ; P1_U3805
g1095 and P1_U4889 P1_U4888 ; P1_U3806
g1096 and P1_U4891 P1_U4890 ; P1_U3807
g1097 and P1_U4894 P1_U4893 ; P1_U3808
g1098 and P1_U4896 P1_U4895 ; P1_U3809
g1099 and P1_U4899 P1_U4898 ; P1_U3810
g1100 and P1_U4901 P1_U4900 ; P1_U3811
g1101 and P1_U4904 P1_U4903 ; P1_U3812
g1102 and P1_U3419 P1_U3369 P1_U3365 ; P1_U3813
g1103 and P1_U3367 P1_U3364 P1_U3360 ; P1_U3814
g1104 and P1_U3361 P1_U3363 ; P1_U3815
g1105 and P1_U3815 P1_U3420 ; P1_U3816
g1106 and P1_U3439 P1_STATE_REG_SCAN_IN ; P1_U3817
g1107 and P1_U4924 P1_U4925 ; P1_U3818
g1108 and P1_U4928 P1_U4926 P1_U4927 ; P1_U3819
g1109 and P1_U4934 P1_U4935 ; P1_U3820
g1110 and P1_U4938 P1_U4936 P1_U4937 ; P1_U3821
g1111 and P1_U4944 P1_U4945 ; P1_U3822
g1112 and P1_U4948 P1_U4946 P1_U4947 ; P1_U3823
g1113 and P1_U4954 P1_U4955 ; P1_U3824
g1114 and P1_U4958 P1_U4956 P1_U4957 ; P1_U3825
g1115 and P1_U4964 P1_U4965 ; P1_U3826
g1116 and P1_U4968 P1_U4966 P1_U4967 ; P1_U3827
g1117 and P1_U4974 P1_U4975 ; P1_U3828
g1118 and P1_U4978 P1_U4976 P1_U4977 ; P1_U3829
g1119 and P1_U4984 P1_U4985 ; P1_U3830
g1120 and P1_U4988 P1_U4986 P1_U4987 ; P1_U3831
g1121 and P1_U4994 P1_U4995 ; P1_U3832
g1122 and P1_U4998 P1_U4996 P1_U4997 ; P1_U3833
g1123 and P1_U5004 P1_U5005 ; P1_U3834
g1124 and P1_U5008 P1_U5006 P1_U5007 ; P1_U3835
g1125 and P1_U5014 P1_U5015 ; P1_U3836
g1126 and P1_U5018 P1_U5016 P1_U5017 ; P1_U3837
g1127 and P1_U5024 P1_U5025 ; P1_U3838
g1128 and P1_U5028 P1_U5026 P1_U5027 ; P1_U3839
g1129 and P1_U5034 P1_U5035 ; P1_U3840
g1130 and P1_U5038 P1_U5036 P1_U5037 ; P1_U3841
g1131 and P1_U5044 P1_U5045 ; P1_U3842
g1132 and P1_U5047 P1_U5046 P1_U5048 ; P1_U3843
g1133 and P1_U5054 P1_U5055 P1_U5053 ; P1_U3844
g1134 and P1_U5057 P1_U5056 P1_U5058 ; P1_U3845
g1135 and P1_U5064 P1_U5065 P1_U5063 ; P1_U3846
g1136 and P1_U5067 P1_U5066 P1_U5068 ; P1_U3847
g1137 and P1_U5073 P1_U4031 ; P1_U3848
g1138 and P1_U5075 P1_U5074 P1_U3848 ; P1_U3849
g1139 and P1_U5077 P1_U5076 P1_U5078 ; P1_U3850
g1140 and P1_U5084 P1_U5085 P1_U5083 ; P1_U3851
g1141 and P1_U5087 P1_U5086 P1_U5088 ; P1_U3852
g1142 and P1_U5093 P1_U4031 ; P1_U3853
g1143 and P1_U5095 P1_U5094 P1_U3853 ; P1_U3854
g1144 and P1_U5097 P1_U5096 P1_U5098 ; P1_U3855
g1145 and P1_U5104 P1_U5105 P1_U5103 ; P1_U3856
g1146 and P1_U5107 P1_U5106 P1_U5108 ; P1_U3857
g1147 and P1_U5114 P1_U5115 P1_U5113 ; P1_U3858
g1148 and P1_U5117 P1_U5116 P1_U5118 ; P1_U3859
g1149 and P1_U3426 P1_STATE_REG_SCAN_IN ; P1_U3860
g1150 and P1_U3860 P1_U3424 ; P1_U3861
g1151 and P1_U6127 P1_U6124 P1_U6130 ; P1_U3862
g1152 and P1_U3864 P1_U3862 P1_U6142 ; P1_U3863
g1153 and P1_U6139 P1_U6136 P1_U6133 ; P1_U3864
g1154 and P1_U6151 P1_U6148 P1_U6154 ; P1_U3865
g1155 and P1_U6160 P1_U6157 P1_U6163 ; P1_U3866
g1156 and P1_U3866 P1_U3865 P1_U6145 ; P1_U3867
g1157 and P1_U3867 P1_U3863 P1_U6121 P1_U6166 ; P1_U3868
g1158 and P1_U6190 P1_U6187 ; P1_U3869
g1159 and P1_U6181 P1_U6178 P1_U6175 P1_U6172 P1_U6184 ; P1_U3870
g1160 and P1_U3870 P1_U6169 ; P1_U3871
g1161 and P1_U6112 P1_U6109 P1_U6106 P1_U6103 ; P1_U3872
g1162 and P1_U6118 P1_U6115 ; P1_U3873
g1163 and P1_U3873 P1_U3872 P1_U6100 P1_U6097 ; P1_U3874
g1164 and P1_U5689 P1_U5123 P1_U3984 P1_U5687 ; P1_U3875
g1165 and P1_U3452 P1_U3453 ; P1_U3876
g1166 and P1_U3370 P1_U3368 P1_U3420 ; P1_U3877
g1167 and P1_U5703 P1_U4002 ; P1_U3878
g1168 and P1_U3424 P1_U3878 ; P1_U3879
g1169 and P1_U3022 P1_U5132 ; P1_U3880
g1170 and P1_U3882 P1_U5175 ; P1_U3881
g1171 and P1_U5179 P1_U5178 ; P1_U3882
g1172 and P1_U4027 P1_U3076 ; P1_U3883
g1173 and P1_U5220 P1_U5219 ; P1_U3884
g1174 and P1_U5223 P1_U5222 ; P1_U3885
g1175 and P1_U3887 P1_U5237 ; P1_U3886
g1176 and P1_U5241 P1_U5240 ; P1_U3887
g1177 and P1_U5268 P1_U5267 ; P1_U3888
g1178 and P1_U3890 P1_U5309 ; P1_U3889
g1179 and P1_U5313 P1_U5312 ; P1_U3890
g1180 and P1_U3892 P1_U5345 ; P1_U3891
g1181 and P1_U5349 P1_U5348 ; P1_U3892
g1182 and P1_U3434 P1_U5398 ; P1_U3893
g1183 and P1_U5463 P1_U5464 ; P1_U3894
g1184 and P1_U5523 P1_U5521 ; P1_U3895
g1185 and P1_U3439 P1_U5535 ; P1_U3896
g1186 and P1_U3439 P1_U5541 ; P1_U3897
g1187 and P1_U5544 P1_U3439 ; P1_U3898
g1188 and P1_U5546 P1_U3439 ; P1_U3899
g1189 and P1_U5548 P1_U3439 ; P1_U3900
g1190 and P1_U5550 P1_U3439 ; P1_U3901
g1191 and P1_U5552 P1_U3439 ; P1_U3902
g1192 and P1_U5554 P1_U3439 ; P1_U3903
g1193 and P1_U5556 P1_U3439 ; P1_U3904
g1194 and P1_U5558 P1_U3439 ; P1_U3905
g1195 and P1_U5560 P1_U3439 ; P1_U3906
g1196 and P1_U5562 P1_U3439 ; P1_U3907
g1197 and P1_U3439 P1_U5563 ; P1_U3908
g1198 and P1_U3439 P1_U5565 ; P1_U3909
g1199 and P1_U3439 P1_U5567 ; P1_U3910
g1200 and P1_U3439 P1_U5569 ; P1_U3911
g1201 and P1_U3439 P1_U5571 ; P1_U3912
g1202 and P1_U3439 P1_U5573 ; P1_U3913
g1203 and P1_U3439 P1_U5575 ; P1_U3914
g1204 and P1_U3439 P1_U5577 ; P1_U3915
g1205 and P1_U3439 P1_U5579 ; P1_U3916
g1206 and P1_U3439 P1_U5581 ; P1_U3917
g1207 and P1_U3439 P1_U5583 ; P1_U3918
g1208 and P1_U3439 P1_U5585 ; P1_U3919
g1209 and P1_U3439 P1_U5587 ; P1_U3920
g1210 and P1_U5606 P1_U5604 ; P1_U3921
g1211 and P1_U5613 P1_U5611 ; P1_U3922
g1212 and P1_U5619 P1_U5617 ; P1_U3923
g1213 and P1_U5622 P1_U5620 ; P1_U3924
g1214 and P1_U5625 P1_U5623 ; P1_U3925
g1215 and P1_U5628 P1_U5626 ; P1_U3926
g1216 and P1_U5631 P1_U5629 ; P1_U3927
g1217 and P1_U5634 P1_U5632 ; P1_U3928
g1218 and P1_U5637 P1_U5635 ; P1_U3929
g1219 and P1_U5640 P1_U5638 ; P1_U3930
g1220 and P1_U5643 P1_U5641 ; P1_U3931
g1221 and P1_U5646 P1_U5644 ; P1_U3932
g1222 and P1_U5649 P1_U5647 ; P1_U3933
g1223 and P1_U5652 P1_U5650 ; P1_U3934
g1224 and P1_U5655 P1_U5653 ; P1_U3935
g1225 and P1_U5658 P1_U5656 ; P1_U3936
g1226 and P1_U5661 P1_U5659 ; P1_U3937
g1227 and P1_U5664 P1_U5662 ; P1_U3938
g1228 and P1_U5667 P1_U5665 ; P1_U3939
g1229 and P1_U5670 P1_U5668 ; P1_U3940
g1230 and P1_U5673 P1_U5671 ; P1_U3941
g1231 and P1_U5676 P1_U5674 ; P1_U3942
g1232 and P1_U5679 P1_U5677 ; P1_U3943
g1233 not P1_IR_REG_31__SCAN_IN ; P1_U3944
g1234 nand P1_U3022 P1_U3359 ; P1_U3945
g1235 nand P1_U5734 P1_U5728 ; P1_U3946
g1236 nand P1_U3634 P1_U3047 ; P1_U3947
g1237 nand P1_U3753 P1_U3047 ; P1_U3948
g1238 and P1_U5968 P1_U5967 ; P1_U3949
g1239 and P1_U5970 P1_U5969 ; P1_U3950
g1240 and P1_U5972 P1_U5971 ; P1_U3951
g1241 and P1_U5974 P1_U5973 ; P1_U3952
g1242 and P1_U5976 P1_U5975 ; P1_U3953
g1243 and P1_U5978 P1_U5977 ; P1_U3954
g1244 and P1_U5980 P1_U5979 ; P1_U3955
g1245 and P1_U5982 P1_U5981 ; P1_U3956
g1246 and P1_U5984 P1_U5983 ; P1_U3957
g1247 and P1_U5986 P1_U5985 ; P1_U3958
g1248 and P1_U5988 P1_U5987 ; P1_U3959
g1249 and P1_U5990 P1_U5989 ; P1_U3960
g1250 and P1_U5992 P1_U5991 ; P1_U3961
g1251 and P1_U5994 P1_U5993 ; P1_U3962
g1252 and P1_U5996 P1_U5995 ; P1_U3963
g1253 and P1_U5998 P1_U5997 ; P1_U3964
g1254 and P1_U6000 P1_U5999 ; P1_U3965
g1255 and P1_U6002 P1_U6001 ; P1_U3966
g1256 and P1_U6004 P1_U6003 ; P1_U3967
g1257 and P1_U6006 P1_U6005 ; P1_U3968
g1258 and P1_U6008 P1_U6007 ; P1_U3969
g1259 and P1_U6010 P1_U6009 ; P1_U3970
g1260 and P1_U6012 P1_U6011 ; P1_U3971
g1261 and P1_U6014 P1_U6013 ; P1_U3972
g1262 and P1_U6016 P1_U6015 ; P1_U3973
g1263 and P1_U6018 P1_U6017 ; P1_U3974
g1264 and P1_U6020 P1_U6019 ; P1_U3975
g1265 and P1_U6022 P1_U6021 ; P1_U3976
g1266 and P1_U6024 P1_U6023 ; P1_U3977
g1267 and P1_U6026 P1_U6025 ; P1_U3978
g1268 nand P1_U3752 P1_U3054 ; P1_U3979
g1269 and P1_U6028 P1_U6027 ; P1_U3980
g1270 and P1_U6030 P1_U6029 ; P1_U3981
g1271 nand P1_U3871 P1_U3868 P1_U3869 P1_U3874 ; P1_U3982
g1272 not P1_R1360_U14 ; P1_U3983
g1273 and P1_U6200 P1_U6199 ; P1_U3984
g1274 not P1_R1352_U6 ; P1_U3985
g1275 not P1_U3371 ; P1_U3986
g1276 not P1_U3428 ; P1_U3987
g1277 not P1_U3426 ; P1_U3988
g1278 not P1_U3369 ; P1_U3989
g1279 not P1_U3419 ; P1_U3990
g1280 not P1_U3365 ; P1_U3991
g1281 not P1_U3364 ; P1_U3992
g1282 not P1_U3367 ; P1_U3993
g1283 not P1_U3360 ; P1_U3994
g1284 not P1_U3363 ; P1_U3995
g1285 not P1_U3361 ; P1_U3996
g1286 not P1_U3420 ; P1_U3997
g1287 not P1_U3418 ; P1_U3998
g1288 nand P1_U3049 P1_U4034 ; P1_U3999
g1289 not P1_U3370 ; P1_U4000
g1290 not P1_U3368 ; P1_U4001
g1291 nand P1_U4020 P1_U3366 ; P1_U4002
g1292 nand P1_U3049 P1_U3421 ; P1_U4003
g1293 not P1_U3946 ; P1_U4004
g1294 not P1_U3431 ; P1_U4005
g1295 not P1_U3425 ; P1_U4006
g1296 not P1_U3410 ; P1_U4007
g1297 not P1_U3408 ; P1_U4008
g1298 not P1_U3406 ; P1_U4009
g1299 not P1_U3404 ; P1_U4010
g1300 not P1_U3402 ; P1_U4011
g1301 not P1_U3400 ; P1_U4012
g1302 not P1_U3398 ; P1_U4013
g1303 not P1_U3396 ; P1_U4014
g1304 not P1_U3394 ; P1_U4015
g1305 not P1_U3415 ; P1_U4016
g1306 not P1_U3414 ; P1_U4017
g1307 not P1_U3412 ; P1_U4018
g1308 not P1_U3427 ; P1_U4019
g1309 not P1_U3372 ; P1_U4020
g1310 not P1_U3416 ; P1_U4021
g1311 not P1_U3417 ; P1_U4022
g1312 not P1_U3948 ; P1_U4023
g1313 not P1_U3947 ; P1_U4024
g1314 not P1_U3945 ; P1_U4025
g1315 not P1_U3979 ; P1_U4026
g1316 not P1_U3432 ; P1_U4027
g1317 nand P1_U3433 P1_STATE_REG_SCAN_IN ; P1_U4028
g1318 nand P1_U3998 P1_U3022 ; P1_U4029
g1319 not P1_U3430 ; P1_U4030
g1320 nand P1_U4006 P1_U3210 ; P1_U4031
g1321 not P1_U3424 ; P1_U4032
g1322 not P1_U3434 ; P1_U4033
g1323 not P1_U3362 ; P1_U4034
g1324 not P1_U3366 ; P1_U4035
g1325 not P1_U3357 ; P1_U4036
g1326 not P1_U3356 ; P1_U4037
g1327 nand U88 P1_U3084 ; P1_U4038
g1328 nand P1_U3028 P1_IR_REG_0__SCAN_IN ; P1_U4039
g1329 nand P1_U4037 P1_IR_REG_0__SCAN_IN ; P1_U4040
g1330 nand U77 P1_U3084 ; P1_U4041
g1331 nand P1_SUB_88_U40 P1_U3028 ; P1_U4042
g1332 nand P1_U4037 P1_IR_REG_1__SCAN_IN ; P1_U4043
g1333 nand U66 P1_U3084 ; P1_U4044
g1334 nand P1_SUB_88_U21 P1_U3028 ; P1_U4045
g1335 nand P1_U4037 P1_IR_REG_2__SCAN_IN ; P1_U4046
g1336 nand U63 P1_U3084 ; P1_U4047
g1337 nand P1_SUB_88_U22 P1_U3028 ; P1_U4048
g1338 nand P1_U4037 P1_IR_REG_3__SCAN_IN ; P1_U4049
g1339 nand U62 P1_U3084 ; P1_U4050
g1340 nand P1_SUB_88_U23 P1_U3028 ; P1_U4051
g1341 nand P1_U4037 P1_IR_REG_4__SCAN_IN ; P1_U4052
g1342 nand U61 P1_U3084 ; P1_U4053
g1343 nand P1_SUB_88_U162 P1_U3028 ; P1_U4054
g1344 nand P1_U4037 P1_IR_REG_5__SCAN_IN ; P1_U4055
g1345 nand U60 P1_U3084 ; P1_U4056
g1346 nand P1_SUB_88_U24 P1_U3028 ; P1_U4057
g1347 nand P1_U4037 P1_IR_REG_6__SCAN_IN ; P1_U4058
g1348 nand U59 P1_U3084 ; P1_U4059
g1349 nand P1_SUB_88_U25 P1_U3028 ; P1_U4060
g1350 nand P1_U4037 P1_IR_REG_7__SCAN_IN ; P1_U4061
g1351 nand U58 P1_U3084 ; P1_U4062
g1352 nand P1_SUB_88_U26 P1_U3028 ; P1_U4063
g1353 nand P1_U4037 P1_IR_REG_8__SCAN_IN ; P1_U4064
g1354 nand U57 P1_U3084 ; P1_U4065
g1355 nand P1_SUB_88_U160 P1_U3028 ; P1_U4066
g1356 nand P1_U4037 P1_IR_REG_9__SCAN_IN ; P1_U4067
g1357 nand U87 P1_U3084 ; P1_U4068
g1358 nand P1_SUB_88_U6 P1_U3028 ; P1_U4069
g1359 nand P1_U4037 P1_IR_REG_10__SCAN_IN ; P1_U4070
g1360 nand U86 P1_U3084 ; P1_U4071
g1361 nand P1_SUB_88_U7 P1_U3028 ; P1_U4072
g1362 nand P1_U4037 P1_IR_REG_11__SCAN_IN ; P1_U4073
g1363 nand U85 P1_U3084 ; P1_U4074
g1364 nand P1_SUB_88_U8 P1_U3028 ; P1_U4075
g1365 nand P1_U4037 P1_IR_REG_12__SCAN_IN ; P1_U4076
g1366 nand U84 P1_U3084 ; P1_U4077
g1367 nand P1_SUB_88_U179 P1_U3028 ; P1_U4078
g1368 nand P1_U4037 P1_IR_REG_13__SCAN_IN ; P1_U4079
g1369 nand U83 P1_U3084 ; P1_U4080
g1370 nand P1_SUB_88_U9 P1_U3028 ; P1_U4081
g1371 nand P1_U4037 P1_IR_REG_14__SCAN_IN ; P1_U4082
g1372 nand U82 P1_U3084 ; P1_U4083
g1373 nand P1_SUB_88_U10 P1_U3028 ; P1_U4084
g1374 nand P1_U4037 P1_IR_REG_15__SCAN_IN ; P1_U4085
g1375 nand U81 P1_U3084 ; P1_U4086
g1376 nand P1_SUB_88_U11 P1_U3028 ; P1_U4087
g1377 nand P1_U4037 P1_IR_REG_16__SCAN_IN ; P1_U4088
g1378 nand U80 P1_U3084 ; P1_U4089
g1379 nand P1_SUB_88_U177 P1_U3028 ; P1_U4090
g1380 nand P1_U4037 P1_IR_REG_17__SCAN_IN ; P1_U4091
g1381 nand U79 P1_U3084 ; P1_U4092
g1382 nand P1_SUB_88_U12 P1_U3028 ; P1_U4093
g1383 nand P1_U4037 P1_IR_REG_18__SCAN_IN ; P1_U4094
g1384 nand U78 P1_U3084 ; P1_U4095
g1385 nand P1_SUB_88_U13 P1_U3028 ; P1_U4096
g1386 nand P1_U4037 P1_IR_REG_19__SCAN_IN ; P1_U4097
g1387 nand U76 P1_U3084 ; P1_U4098
g1388 nand P1_SUB_88_U14 P1_U3028 ; P1_U4099
g1389 nand P1_U4037 P1_IR_REG_20__SCAN_IN ; P1_U4100
g1390 nand U75 P1_U3084 ; P1_U4101
g1391 nand P1_SUB_88_U173 P1_U3028 ; P1_U4102
g1392 nand P1_U4037 P1_IR_REG_21__SCAN_IN ; P1_U4103
g1393 nand U74 P1_U3084 ; P1_U4104
g1394 nand P1_SUB_88_U15 P1_U3028 ; P1_U4105
g1395 nand P1_U4037 P1_IR_REG_22__SCAN_IN ; P1_U4106
g1396 nand U73 P1_U3084 ; P1_U4107
g1397 nand P1_SUB_88_U16 P1_U3028 ; P1_U4108
g1398 nand P1_U4037 P1_IR_REG_23__SCAN_IN ; P1_U4109
g1399 nand U72 P1_U3084 ; P1_U4110
g1400 nand P1_SUB_88_U17 P1_U3028 ; P1_U4111
g1401 nand P1_U4037 P1_IR_REG_24__SCAN_IN ; P1_U4112
g1402 nand U71 P1_U3084 ; P1_U4113
g1403 nand P1_SUB_88_U170 P1_U3028 ; P1_U4114
g1404 nand P1_U4037 P1_IR_REG_25__SCAN_IN ; P1_U4115
g1405 nand U70 P1_U3084 ; P1_U4116
g1406 nand P1_SUB_88_U18 P1_U3028 ; P1_U4117
g1407 nand P1_U4037 P1_IR_REG_26__SCAN_IN ; P1_U4118
g1408 nand U69 P1_U3084 ; P1_U4119
g1409 nand P1_SUB_88_U42 P1_U3028 ; P1_U4120
g1410 nand P1_U4037 P1_IR_REG_27__SCAN_IN ; P1_U4121
g1411 nand U68 P1_U3084 ; P1_U4122
g1412 nand P1_SUB_88_U19 P1_U3028 ; P1_U4123
g1413 nand P1_U4037 P1_IR_REG_28__SCAN_IN ; P1_U4124
g1414 nand U67 P1_U3084 ; P1_U4125
g1415 nand P1_SUB_88_U20 P1_U3028 ; P1_U4126
g1416 nand P1_U4037 P1_IR_REG_29__SCAN_IN ; P1_U4127
g1417 nand U65 P1_U3084 ; P1_U4128
g1418 nand P1_SUB_88_U165 P1_U3028 ; P1_U4129
g1419 nand P1_U4037 P1_IR_REG_30__SCAN_IN ; P1_U4130
g1420 nand U64 P1_U3084 ; P1_U4131
g1421 nand P1_SUB_88_U41 P1_U3028 ; P1_U4132
g1422 nand P1_U4037 P1_IR_REG_31__SCAN_IN ; P1_U4133
g1423 not P1_U3359 ; P1_U4134
g1424 not P1_U3421 ; P1_U4135
g1425 nand P1_U3357 P1_U5692 ; P1_U4136
g1426 nand P1_U3357 P1_U5695 ; P1_U4137
g1427 nand P1_U4134 P1_D_REG_10__SCAN_IN ; P1_U4138
g1428 nand P1_U4134 P1_D_REG_11__SCAN_IN ; P1_U4139
g1429 nand P1_U4134 P1_D_REG_12__SCAN_IN ; P1_U4140
g1430 nand P1_U4134 P1_D_REG_13__SCAN_IN ; P1_U4141
g1431 nand P1_U4134 P1_D_REG_14__SCAN_IN ; P1_U4142
g1432 nand P1_U4134 P1_D_REG_15__SCAN_IN ; P1_U4143
g1433 nand P1_U4134 P1_D_REG_16__SCAN_IN ; P1_U4144
g1434 nand P1_U4134 P1_D_REG_17__SCAN_IN ; P1_U4145
g1435 nand P1_U4134 P1_D_REG_18__SCAN_IN ; P1_U4146
g1436 nand P1_U4134 P1_D_REG_19__SCAN_IN ; P1_U4147
g1437 nand P1_U4134 P1_D_REG_20__SCAN_IN ; P1_U4148
g1438 nand P1_U4134 P1_D_REG_21__SCAN_IN ; P1_U4149
g1439 nand P1_U4134 P1_D_REG_22__SCAN_IN ; P1_U4150
g1440 nand P1_U4134 P1_D_REG_23__SCAN_IN ; P1_U4151
g1441 nand P1_U4134 P1_D_REG_24__SCAN_IN ; P1_U4152
g1442 nand P1_U4134 P1_D_REG_25__SCAN_IN ; P1_U4153
g1443 nand P1_U4134 P1_D_REG_26__SCAN_IN ; P1_U4154
g1444 nand P1_U4134 P1_D_REG_27__SCAN_IN ; P1_U4155
g1445 nand P1_U4134 P1_D_REG_28__SCAN_IN ; P1_U4156
g1446 nand P1_U4134 P1_D_REG_29__SCAN_IN ; P1_U4157
g1447 nand P1_U4134 P1_D_REG_2__SCAN_IN ; P1_U4158
g1448 nand P1_U4134 P1_D_REG_30__SCAN_IN ; P1_U4159
g1449 nand P1_U4134 P1_D_REG_31__SCAN_IN ; P1_U4160
g1450 nand P1_U4134 P1_D_REG_3__SCAN_IN ; P1_U4161
g1451 nand P1_U4134 P1_D_REG_4__SCAN_IN ; P1_U4162
g1452 nand P1_U4134 P1_D_REG_5__SCAN_IN ; P1_U4163
g1453 nand P1_U4134 P1_D_REG_6__SCAN_IN ; P1_U4164
g1454 nand P1_U4134 P1_D_REG_7__SCAN_IN ; P1_U4165
g1455 nand P1_U4134 P1_D_REG_8__SCAN_IN ; P1_U4166
g1456 nand P1_U4134 P1_D_REG_9__SCAN_IN ; P1_U4167
g1457 nand P1_U5716 P1_U5719 ; P1_U4168
g1458 nand P1_U5739 P1_U5738 P1_U3366 ; P1_U4169
g1459 nand P1_U3018 P1_REG2_REG_1__SCAN_IN ; P1_U4170
g1460 nand P1_U3019 P1_REG1_REG_1__SCAN_IN ; P1_U4171
g1461 nand P1_U3020 P1_REG0_REG_1__SCAN_IN ; P1_U4172
g1462 nand P1_U3017 P1_REG3_REG_1__SCAN_IN ; P1_U4173
g1463 not P1_U3076 ; P1_U4174
g1464 nand P1_U3999 P1_U3416 ; P1_U4175
g1465 nand P1_U3994 P1_R1150_U21 ; P1_U4176
g1466 nand P1_U3996 P1_R1117_U21 ; P1_U4177
g1467 nand P1_U3995 P1_R1138_U96 ; P1_U4178
g1468 nand P1_U3992 P1_R1192_U21 ; P1_U4179
g1469 nand P1_U3991 P1_R1207_U21 ; P1_U4180
g1470 nand P1_U4001 P1_R1171_U96 ; P1_U4181
g1471 nand P1_U4000 P1_R1240_U96 ; P1_U4182
g1472 not P1_U3373 ; P1_U4183
g1473 nand P1_R1222_U96 P1_U3026 ; P1_U4184
g1474 nand P1_U3025 P1_U3076 ; P1_U4185
g1475 nand P1_U3451 P1_U3023 ; P1_U4186
g1476 nand P1_U3451 P1_U4175 ; P1_U4187
g1477 nand P1_U3622 P1_U4183 ; P1_U4188
g1478 nand P1_U3018 P1_REG2_REG_2__SCAN_IN ; P1_U4189
g1479 nand P1_U3019 P1_REG1_REG_2__SCAN_IN ; P1_U4190
g1480 nand P1_U3020 P1_REG0_REG_2__SCAN_IN ; P1_U4191
g1481 nand P1_U3017 P1_REG3_REG_2__SCAN_IN ; P1_U4192
g1482 not P1_U3066 ; P1_U4193
g1483 nand P1_U3020 P1_REG0_REG_0__SCAN_IN ; P1_U4194
g1484 nand P1_U3019 P1_REG1_REG_0__SCAN_IN ; P1_U4195
g1485 nand P1_U3018 P1_REG2_REG_0__SCAN_IN ; P1_U4196
g1486 nand P1_U3017 P1_REG3_REG_0__SCAN_IN ; P1_U4197
g1487 not P1_U3075 ; P1_U4198
g1488 nand P1_U3033 P1_U3075 ; P1_U4199
g1489 nand P1_R1150_U98 P1_U3994 ; P1_U4200
g1490 nand P1_R1117_U98 P1_U3996 ; P1_U4201
g1491 nand P1_R1138_U95 P1_U3995 ; P1_U4202
g1492 nand P1_R1192_U98 P1_U3992 ; P1_U4203
g1493 nand P1_R1207_U98 P1_U3991 ; P1_U4204
g1494 nand P1_R1171_U95 P1_U4001 ; P1_U4205
g1495 nand P1_R1240_U95 P1_U4000 ; P1_U4206
g1496 not P1_U3375 ; P1_U4207
g1497 nand P1_R1222_U95 P1_U3026 ; P1_U4208
g1498 nand P1_U3025 P1_U3066 ; P1_U4209
g1499 nand P1_R1282_U57 P1_U3023 ; P1_U4210
g1500 nand P1_U3456 P1_U4175 ; P1_U4211
g1501 nand P1_U3638 P1_U4207 ; P1_U4212
g1502 nand P1_U3018 P1_REG2_REG_3__SCAN_IN ; P1_U4213
g1503 nand P1_U3019 P1_REG1_REG_3__SCAN_IN ; P1_U4214
g1504 nand P1_U3020 P1_REG0_REG_3__SCAN_IN ; P1_U4215
g1505 nand P1_ADD_99_U4 P1_U3017 ; P1_U4216
g1506 not P1_U3062 ; P1_U4217
g1507 nand P1_U3033 P1_U3076 ; P1_U4218
g1508 nand P1_R1150_U108 P1_U3994 ; P1_U4219
g1509 nand P1_R1117_U108 P1_U3996 ; P1_U4220
g1510 nand P1_R1138_U17 P1_U3995 ; P1_U4221
g1511 nand P1_R1192_U108 P1_U3992 ; P1_U4222
g1512 nand P1_R1207_U108 P1_U3991 ; P1_U4223
g1513 nand P1_R1171_U17 P1_U4001 ; P1_U4224
g1514 nand P1_R1240_U17 P1_U4000 ; P1_U4225
g1515 not P1_U3376 ; P1_U4226
g1516 nand P1_R1222_U17 P1_U3026 ; P1_U4227
g1517 nand P1_U3025 P1_U3062 ; P1_U4228
g1518 nand P1_R1282_U18 P1_U3023 ; P1_U4229
g1519 nand P1_U3459 P1_U4175 ; P1_U4230
g1520 nand P1_U3642 P1_U4226 ; P1_U4231
g1521 nand P1_U3018 P1_REG2_REG_4__SCAN_IN ; P1_U4232
g1522 nand P1_U3019 P1_REG1_REG_4__SCAN_IN ; P1_U4233
g1523 nand P1_U3020 P1_REG0_REG_4__SCAN_IN ; P1_U4234
g1524 nand P1_ADD_99_U59 P1_U3017 ; P1_U4235
g1525 not P1_U3058 ; P1_U4236
g1526 nand P1_U3033 P1_U3066 ; P1_U4237
g1527 nand P1_R1150_U18 P1_U3994 ; P1_U4238
g1528 nand P1_R1117_U18 P1_U3996 ; P1_U4239
g1529 nand P1_R1138_U101 P1_U3995 ; P1_U4240
g1530 nand P1_R1192_U18 P1_U3992 ; P1_U4241
g1531 nand P1_R1207_U18 P1_U3991 ; P1_U4242
g1532 nand P1_R1171_U101 P1_U4001 ; P1_U4243
g1533 nand P1_R1240_U101 P1_U4000 ; P1_U4244
g1534 not P1_U3377 ; P1_U4245
g1535 nand P1_R1222_U101 P1_U3026 ; P1_U4246
g1536 nand P1_U3025 P1_U3058 ; P1_U4247
g1537 nand P1_R1282_U20 P1_U3023 ; P1_U4248
g1538 nand P1_U3462 P1_U4175 ; P1_U4249
g1539 nand P1_U3646 P1_U4245 ; P1_U4250
g1540 nand P1_U3018 P1_REG2_REG_5__SCAN_IN ; P1_U4251
g1541 nand P1_U3019 P1_REG1_REG_5__SCAN_IN ; P1_U4252
g1542 nand P1_U3020 P1_REG0_REG_5__SCAN_IN ; P1_U4253
g1543 nand P1_ADD_99_U58 P1_U3017 ; P1_U4254
g1544 not P1_U3065 ; P1_U4255
g1545 nand P1_U3033 P1_U3062 ; P1_U4256
g1546 nand P1_R1150_U107 P1_U3994 ; P1_U4257
g1547 nand P1_R1117_U107 P1_U3996 ; P1_U4258
g1548 nand P1_R1138_U100 P1_U3995 ; P1_U4259
g1549 nand P1_R1192_U107 P1_U3992 ; P1_U4260
g1550 nand P1_R1207_U107 P1_U3991 ; P1_U4261
g1551 nand P1_R1171_U100 P1_U4001 ; P1_U4262
g1552 nand P1_R1240_U100 P1_U4000 ; P1_U4263
g1553 not P1_U3378 ; P1_U4264
g1554 nand P1_R1222_U100 P1_U3026 ; P1_U4265
g1555 nand P1_U3025 P1_U3065 ; P1_U4266
g1556 nand P1_R1282_U21 P1_U3023 ; P1_U4267
g1557 nand P1_U3465 P1_U4175 ; P1_U4268
g1558 nand P1_U3650 P1_U4264 ; P1_U4269
g1559 nand P1_U3018 P1_REG2_REG_6__SCAN_IN ; P1_U4270
g1560 nand P1_U3019 P1_REG1_REG_6__SCAN_IN ; P1_U4271
g1561 nand P1_U3020 P1_REG0_REG_6__SCAN_IN ; P1_U4272
g1562 nand P1_ADD_99_U57 P1_U3017 ; P1_U4273
g1563 not P1_U3069 ; P1_U4274
g1564 nand P1_U3033 P1_U3058 ; P1_U4275
g1565 nand P1_R1150_U106 P1_U3994 ; P1_U4276
g1566 nand P1_R1117_U106 P1_U3996 ; P1_U4277
g1567 nand P1_R1138_U18 P1_U3995 ; P1_U4278
g1568 nand P1_R1192_U106 P1_U3992 ; P1_U4279
g1569 nand P1_R1207_U106 P1_U3991 ; P1_U4280
g1570 nand P1_R1171_U18 P1_U4001 ; P1_U4281
g1571 nand P1_R1240_U18 P1_U4000 ; P1_U4282
g1572 not P1_U3379 ; P1_U4283
g1573 nand P1_R1222_U18 P1_U3026 ; P1_U4284
g1574 nand P1_U3025 P1_U3069 ; P1_U4285
g1575 nand P1_R1282_U65 P1_U3023 ; P1_U4286
g1576 nand P1_U3468 P1_U4175 ; P1_U4287
g1577 nand P1_U3654 P1_U4283 ; P1_U4288
g1578 nand P1_U3018 P1_REG2_REG_7__SCAN_IN ; P1_U4289
g1579 nand P1_U3019 P1_REG1_REG_7__SCAN_IN ; P1_U4290
g1580 nand P1_U3020 P1_REG0_REG_7__SCAN_IN ; P1_U4291
g1581 nand P1_ADD_99_U56 P1_U3017 ; P1_U4292
g1582 not P1_U3068 ; P1_U4293
g1583 nand P1_U3033 P1_U3065 ; P1_U4294
g1584 nand P1_R1150_U19 P1_U3994 ; P1_U4295
g1585 nand P1_R1117_U19 P1_U3996 ; P1_U4296
g1586 nand P1_R1138_U99 P1_U3995 ; P1_U4297
g1587 nand P1_R1192_U19 P1_U3992 ; P1_U4298
g1588 nand P1_R1207_U19 P1_U3991 ; P1_U4299
g1589 nand P1_R1171_U99 P1_U4001 ; P1_U4300
g1590 nand P1_R1240_U99 P1_U4000 ; P1_U4301
g1591 not P1_U3380 ; P1_U4302
g1592 nand P1_R1222_U99 P1_U3026 ; P1_U4303
g1593 nand P1_U3025 P1_U3068 ; P1_U4304
g1594 nand P1_R1282_U22 P1_U3023 ; P1_U4305
g1595 nand P1_U3471 P1_U4175 ; P1_U4306
g1596 nand P1_U3658 P1_U4302 ; P1_U4307
g1597 nand P1_U3018 P1_REG2_REG_8__SCAN_IN ; P1_U4308
g1598 nand P1_U3019 P1_REG1_REG_8__SCAN_IN ; P1_U4309
g1599 nand P1_U3020 P1_REG0_REG_8__SCAN_IN ; P1_U4310
g1600 nand P1_ADD_99_U55 P1_U3017 ; P1_U4311
g1601 not P1_U3082 ; P1_U4312
g1602 nand P1_U3033 P1_U3069 ; P1_U4313
g1603 nand P1_R1150_U105 P1_U3994 ; P1_U4314
g1604 nand P1_R1117_U105 P1_U3996 ; P1_U4315
g1605 nand P1_R1138_U19 P1_U3995 ; P1_U4316
g1606 nand P1_R1192_U105 P1_U3992 ; P1_U4317
g1607 nand P1_R1207_U105 P1_U3991 ; P1_U4318
g1608 nand P1_R1171_U19 P1_U4001 ; P1_U4319
g1609 nand P1_R1240_U19 P1_U4000 ; P1_U4320
g1610 not P1_U3381 ; P1_U4321
g1611 nand P1_R1222_U19 P1_U3026 ; P1_U4322
g1612 nand P1_U3025 P1_U3082 ; P1_U4323
g1613 nand P1_R1282_U23 P1_U3023 ; P1_U4324
g1614 nand P1_U3474 P1_U4175 ; P1_U4325
g1615 nand P1_U3662 P1_U4321 ; P1_U4326
g1616 nand P1_U3018 P1_REG2_REG_9__SCAN_IN ; P1_U4327
g1617 nand P1_U3019 P1_REG1_REG_9__SCAN_IN ; P1_U4328
g1618 nand P1_U3020 P1_REG0_REG_9__SCAN_IN ; P1_U4329
g1619 nand P1_ADD_99_U54 P1_U3017 ; P1_U4330
g1620 not P1_U3081 ; P1_U4331
g1621 nand P1_U3033 P1_U3068 ; P1_U4332
g1622 nand P1_R1150_U20 P1_U3994 ; P1_U4333
g1623 nand P1_R1117_U20 P1_U3996 ; P1_U4334
g1624 nand P1_R1138_U98 P1_U3995 ; P1_U4335
g1625 nand P1_R1192_U20 P1_U3992 ; P1_U4336
g1626 nand P1_R1207_U20 P1_U3991 ; P1_U4337
g1627 nand P1_R1171_U98 P1_U4001 ; P1_U4338
g1628 nand P1_R1240_U98 P1_U4000 ; P1_U4339
g1629 not P1_U3382 ; P1_U4340
g1630 nand P1_R1222_U98 P1_U3026 ; P1_U4341
g1631 nand P1_U3025 P1_U3081 ; P1_U4342
g1632 nand P1_R1282_U24 P1_U3023 ; P1_U4343
g1633 nand P1_U3477 P1_U4175 ; P1_U4344
g1634 nand P1_U3666 P1_U4340 ; P1_U4345
g1635 nand P1_U3018 P1_REG2_REG_10__SCAN_IN ; P1_U4346
g1636 nand P1_U3019 P1_REG1_REG_10__SCAN_IN ; P1_U4347
g1637 nand P1_U3020 P1_REG0_REG_10__SCAN_IN ; P1_U4348
g1638 nand P1_ADD_99_U78 P1_U3017 ; P1_U4349
g1639 not P1_U3060 ; P1_U4350
g1640 nand P1_U3033 P1_U3082 ; P1_U4351
g1641 nand P1_R1150_U104 P1_U3994 ; P1_U4352
g1642 nand P1_R1117_U104 P1_U3996 ; P1_U4353
g1643 nand P1_R1138_U97 P1_U3995 ; P1_U4354
g1644 nand P1_R1192_U104 P1_U3992 ; P1_U4355
g1645 nand P1_R1207_U104 P1_U3991 ; P1_U4356
g1646 nand P1_R1171_U97 P1_U4001 ; P1_U4357
g1647 nand P1_R1240_U97 P1_U4000 ; P1_U4358
g1648 not P1_U3383 ; P1_U4359
g1649 nand P1_R1222_U97 P1_U3026 ; P1_U4360
g1650 nand P1_U3025 P1_U3060 ; P1_U4361
g1651 nand P1_R1282_U63 P1_U3023 ; P1_U4362
g1652 nand P1_U3480 P1_U4175 ; P1_U4363
g1653 nand P1_U3670 P1_U4359 ; P1_U4364
g1654 nand P1_U3018 P1_REG2_REG_11__SCAN_IN ; P1_U4365
g1655 nand P1_U3019 P1_REG1_REG_11__SCAN_IN ; P1_U4366
g1656 nand P1_U3020 P1_REG0_REG_11__SCAN_IN ; P1_U4367
g1657 nand P1_ADD_99_U77 P1_U3017 ; P1_U4368
g1658 not P1_U3061 ; P1_U4369
g1659 nand P1_U3033 P1_U3081 ; P1_U4370
g1660 nand P1_R1150_U114 P1_U3994 ; P1_U4371
g1661 nand P1_R1117_U114 P1_U3996 ; P1_U4372
g1662 nand P1_R1138_U11 P1_U3995 ; P1_U4373
g1663 nand P1_R1192_U114 P1_U3992 ; P1_U4374
g1664 nand P1_R1207_U114 P1_U3991 ; P1_U4375
g1665 nand P1_R1171_U11 P1_U4001 ; P1_U4376
g1666 nand P1_R1240_U11 P1_U4000 ; P1_U4377
g1667 not P1_U3384 ; P1_U4378
g1668 nand P1_R1222_U11 P1_U3026 ; P1_U4379
g1669 nand P1_U3025 P1_U3061 ; P1_U4380
g1670 nand P1_R1282_U6 P1_U3023 ; P1_U4381
g1671 nand P1_U3483 P1_U4175 ; P1_U4382
g1672 nand P1_U3674 P1_U4378 ; P1_U4383
g1673 nand P1_U3018 P1_REG2_REG_12__SCAN_IN ; P1_U4384
g1674 nand P1_U3019 P1_REG1_REG_12__SCAN_IN ; P1_U4385
g1675 nand P1_U3020 P1_REG0_REG_12__SCAN_IN ; P1_U4386
g1676 nand P1_ADD_99_U76 P1_U3017 ; P1_U4387
g1677 not P1_U3070 ; P1_U4388
g1678 nand P1_U3033 P1_U3060 ; P1_U4389
g1679 nand P1_R1150_U13 P1_U3994 ; P1_U4390
g1680 nand P1_R1117_U13 P1_U3996 ; P1_U4391
g1681 nand P1_R1138_U115 P1_U3995 ; P1_U4392
g1682 nand P1_R1192_U13 P1_U3992 ; P1_U4393
g1683 nand P1_R1207_U13 P1_U3991 ; P1_U4394
g1684 nand P1_R1171_U115 P1_U4001 ; P1_U4395
g1685 nand P1_R1240_U115 P1_U4000 ; P1_U4396
g1686 not P1_U3385 ; P1_U4397
g1687 nand P1_R1222_U115 P1_U3026 ; P1_U4398
g1688 nand P1_U3025 P1_U3070 ; P1_U4399
g1689 nand P1_R1282_U7 P1_U3023 ; P1_U4400
g1690 nand P1_U3486 P1_U4175 ; P1_U4401
g1691 nand P1_U3678 P1_U4397 ; P1_U4402
g1692 nand P1_U3018 P1_REG2_REG_13__SCAN_IN ; P1_U4403
g1693 nand P1_U3019 P1_REG1_REG_13__SCAN_IN ; P1_U4404
g1694 nand P1_U3020 P1_REG0_REG_13__SCAN_IN ; P1_U4405
g1695 nand P1_ADD_99_U75 P1_U3017 ; P1_U4406
g1696 not P1_U3078 ; P1_U4407
g1697 nand P1_U3033 P1_U3061 ; P1_U4408
g1698 nand P1_R1150_U103 P1_U3994 ; P1_U4409
g1699 nand P1_R1117_U103 P1_U3996 ; P1_U4410
g1700 nand P1_R1138_U114 P1_U3995 ; P1_U4411
g1701 nand P1_R1192_U103 P1_U3992 ; P1_U4412
g1702 nand P1_R1207_U103 P1_U3991 ; P1_U4413
g1703 nand P1_R1171_U114 P1_U4001 ; P1_U4414
g1704 nand P1_R1240_U114 P1_U4000 ; P1_U4415
g1705 not P1_U3386 ; P1_U4416
g1706 nand P1_R1222_U114 P1_U3026 ; P1_U4417
g1707 nand P1_U3025 P1_U3078 ; P1_U4418
g1708 nand P1_R1282_U8 P1_U3023 ; P1_U4419
g1709 nand P1_U3489 P1_U4175 ; P1_U4420
g1710 nand P1_U3682 P1_U4416 ; P1_U4421
g1711 nand P1_U3018 P1_REG2_REG_14__SCAN_IN ; P1_U4422
g1712 nand P1_U3019 P1_REG1_REG_14__SCAN_IN ; P1_U4423
g1713 nand P1_U3020 P1_REG0_REG_14__SCAN_IN ; P1_U4424
g1714 nand P1_ADD_99_U74 P1_U3017 ; P1_U4425
g1715 not P1_U3077 ; P1_U4426
g1716 nand P1_U3033 P1_U3070 ; P1_U4427
g1717 nand P1_R1150_U102 P1_U3994 ; P1_U4428
g1718 nand P1_R1117_U102 P1_U3996 ; P1_U4429
g1719 nand P1_R1138_U12 P1_U3995 ; P1_U4430
g1720 nand P1_R1192_U102 P1_U3992 ; P1_U4431
g1721 nand P1_R1207_U102 P1_U3991 ; P1_U4432
g1722 nand P1_R1171_U12 P1_U4001 ; P1_U4433
g1723 nand P1_R1240_U12 P1_U4000 ; P1_U4434
g1724 not P1_U3387 ; P1_U4435
g1725 nand P1_R1222_U12 P1_U3026 ; P1_U4436
g1726 nand P1_U3025 P1_U3077 ; P1_U4437
g1727 nand P1_R1282_U86 P1_U3023 ; P1_U4438
g1728 nand P1_U3492 P1_U4175 ; P1_U4439
g1729 nand P1_U3686 P1_U4435 ; P1_U4440
g1730 nand P1_U3018 P1_REG2_REG_15__SCAN_IN ; P1_U4441
g1731 nand P1_U3019 P1_REG1_REG_15__SCAN_IN ; P1_U4442
g1732 nand P1_U3020 P1_REG0_REG_15__SCAN_IN ; P1_U4443
g1733 nand P1_ADD_99_U73 P1_U3017 ; P1_U4444
g1734 not P1_U3072 ; P1_U4445
g1735 nand P1_U3033 P1_U3078 ; P1_U4446
g1736 nand P1_R1150_U113 P1_U3994 ; P1_U4447
g1737 nand P1_R1117_U113 P1_U3996 ; P1_U4448
g1738 nand P1_R1138_U113 P1_U3995 ; P1_U4449
g1739 nand P1_R1192_U113 P1_U3992 ; P1_U4450
g1740 nand P1_R1207_U113 P1_U3991 ; P1_U4451
g1741 nand P1_R1171_U113 P1_U4001 ; P1_U4452
g1742 nand P1_R1240_U113 P1_U4000 ; P1_U4453
g1743 not P1_U3388 ; P1_U4454
g1744 nand P1_R1222_U113 P1_U3026 ; P1_U4455
g1745 nand P1_U3025 P1_U3072 ; P1_U4456
g1746 nand P1_R1282_U9 P1_U3023 ; P1_U4457
g1747 nand P1_U3495 P1_U4175 ; P1_U4458
g1748 nand P1_U3690 P1_U4454 ; P1_U4459
g1749 nand P1_U3018 P1_REG2_REG_16__SCAN_IN ; P1_U4460
g1750 nand P1_U3019 P1_REG1_REG_16__SCAN_IN ; P1_U4461
g1751 nand P1_U3020 P1_REG0_REG_16__SCAN_IN ; P1_U4462
g1752 nand P1_ADD_99_U72 P1_U3017 ; P1_U4463
g1753 not P1_U3071 ; P1_U4464
g1754 nand P1_U3033 P1_U3077 ; P1_U4465
g1755 nand P1_R1150_U112 P1_U3994 ; P1_U4466
g1756 nand P1_R1117_U112 P1_U3996 ; P1_U4467
g1757 nand P1_R1138_U112 P1_U3995 ; P1_U4468
g1758 nand P1_R1192_U112 P1_U3992 ; P1_U4469
g1759 nand P1_R1207_U112 P1_U3991 ; P1_U4470
g1760 nand P1_R1171_U112 P1_U4001 ; P1_U4471
g1761 nand P1_R1240_U112 P1_U4000 ; P1_U4472
g1762 not P1_U3389 ; P1_U4473
g1763 nand P1_R1222_U112 P1_U3026 ; P1_U4474
g1764 nand P1_U3025 P1_U3071 ; P1_U4475
g1765 nand P1_R1282_U10 P1_U3023 ; P1_U4476
g1766 nand P1_U3498 P1_U4175 ; P1_U4477
g1767 nand P1_U3694 P1_U4473 ; P1_U4478
g1768 nand P1_U3018 P1_REG2_REG_17__SCAN_IN ; P1_U4479
g1769 nand P1_U3019 P1_REG1_REG_17__SCAN_IN ; P1_U4480
g1770 nand P1_U3020 P1_REG0_REG_17__SCAN_IN ; P1_U4481
g1771 nand P1_ADD_99_U71 P1_U3017 ; P1_U4482
g1772 not P1_U3067 ; P1_U4483
g1773 nand P1_U3033 P1_U3072 ; P1_U4484
g1774 nand P1_R1150_U14 P1_U3994 ; P1_U4485
g1775 nand P1_R1117_U14 P1_U3996 ; P1_U4486
g1776 nand P1_R1138_U111 P1_U3995 ; P1_U4487
g1777 nand P1_R1192_U14 P1_U3992 ; P1_U4488
g1778 nand P1_R1207_U14 P1_U3991 ; P1_U4489
g1779 nand P1_R1171_U111 P1_U4001 ; P1_U4490
g1780 nand P1_R1240_U111 P1_U4000 ; P1_U4491
g1781 not P1_U3390 ; P1_U4492
g1782 nand P1_R1222_U111 P1_U3026 ; P1_U4493
g1783 nand P1_U3025 P1_U3067 ; P1_U4494
g1784 nand P1_R1282_U11 P1_U3023 ; P1_U4495
g1785 nand P1_U3501 P1_U4175 ; P1_U4496
g1786 nand P1_U3698 P1_U4492 ; P1_U4497
g1787 nand P1_U3018 P1_REG2_REG_18__SCAN_IN ; P1_U4498
g1788 nand P1_U3019 P1_REG1_REG_18__SCAN_IN ; P1_U4499
g1789 nand P1_U3020 P1_REG0_REG_18__SCAN_IN ; P1_U4500
g1790 nand P1_ADD_99_U70 P1_U3017 ; P1_U4501
g1791 not P1_U3080 ; P1_U4502
g1792 nand P1_U3033 P1_U3071 ; P1_U4503
g1793 nand P1_R1150_U101 P1_U3994 ; P1_U4504
g1794 nand P1_R1117_U101 P1_U3996 ; P1_U4505
g1795 nand P1_R1138_U13 P1_U3995 ; P1_U4506
g1796 nand P1_R1192_U101 P1_U3992 ; P1_U4507
g1797 nand P1_R1207_U101 P1_U3991 ; P1_U4508
g1798 nand P1_R1171_U13 P1_U4001 ; P1_U4509
g1799 nand P1_R1240_U13 P1_U4000 ; P1_U4510
g1800 not P1_U3391 ; P1_U4511
g1801 nand P1_R1222_U13 P1_U3026 ; P1_U4512
g1802 nand P1_U3025 P1_U3080 ; P1_U4513
g1803 nand P1_R1282_U84 P1_U3023 ; P1_U4514
g1804 nand P1_U3504 P1_U4175 ; P1_U4515
g1805 nand P1_U3702 P1_U4511 ; P1_U4516
g1806 nand P1_U3018 P1_REG2_REG_19__SCAN_IN ; P1_U4517
g1807 nand P1_U3019 P1_REG1_REG_19__SCAN_IN ; P1_U4518
g1808 nand P1_U3020 P1_REG0_REG_19__SCAN_IN ; P1_U4519
g1809 nand P1_ADD_99_U69 P1_U3017 ; P1_U4520
g1810 not P1_U3079 ; P1_U4521
g1811 nand P1_U3033 P1_U3067 ; P1_U4522
g1812 nand P1_R1150_U100 P1_U3994 ; P1_U4523
g1813 nand P1_R1117_U100 P1_U3996 ; P1_U4524
g1814 nand P1_R1138_U110 P1_U3995 ; P1_U4525
g1815 nand P1_R1192_U100 P1_U3992 ; P1_U4526
g1816 nand P1_R1207_U100 P1_U3991 ; P1_U4527
g1817 nand P1_R1171_U110 P1_U4001 ; P1_U4528
g1818 nand P1_R1240_U110 P1_U4000 ; P1_U4529
g1819 not P1_U3392 ; P1_U4530
g1820 nand P1_R1222_U110 P1_U3026 ; P1_U4531
g1821 nand P1_U3025 P1_U3079 ; P1_U4532
g1822 nand P1_R1282_U12 P1_U3023 ; P1_U4533
g1823 nand P1_U3507 P1_U4175 ; P1_U4534
g1824 nand P1_U3706 P1_U4530 ; P1_U4535
g1825 nand P1_U3018 P1_REG2_REG_20__SCAN_IN ; P1_U4536
g1826 nand P1_U3019 P1_REG1_REG_20__SCAN_IN ; P1_U4537
g1827 nand P1_U3020 P1_REG0_REG_20__SCAN_IN ; P1_U4538
g1828 nand P1_ADD_99_U68 P1_U3017 ; P1_U4539
g1829 not P1_U3074 ; P1_U4540
g1830 nand P1_U3033 P1_U3080 ; P1_U4541
g1831 nand P1_R1150_U99 P1_U3994 ; P1_U4542
g1832 nand P1_R1117_U99 P1_U3996 ; P1_U4543
g1833 nand P1_R1138_U109 P1_U3995 ; P1_U4544
g1834 nand P1_R1192_U99 P1_U3992 ; P1_U4545
g1835 nand P1_R1207_U99 P1_U3991 ; P1_U4546
g1836 nand P1_R1171_U109 P1_U4001 ; P1_U4547
g1837 nand P1_R1240_U109 P1_U4000 ; P1_U4548
g1838 not P1_U3393 ; P1_U4549
g1839 nand P1_R1222_U109 P1_U3026 ; P1_U4550
g1840 nand P1_U3025 P1_U3074 ; P1_U4551
g1841 nand P1_R1282_U82 P1_U3023 ; P1_U4552
g1842 nand P1_U3509 P1_U4175 ; P1_U4553
g1843 nand P1_U3710 P1_U4549 ; P1_U4554
g1844 nand P1_U3018 P1_REG2_REG_21__SCAN_IN ; P1_U4555
g1845 nand P1_U3019 P1_REG1_REG_21__SCAN_IN ; P1_U4556
g1846 nand P1_U3020 P1_REG0_REG_21__SCAN_IN ; P1_U4557
g1847 nand P1_ADD_99_U67 P1_U3017 ; P1_U4558
g1848 not P1_U3073 ; P1_U4559
g1849 nand P1_U3033 P1_U3079 ; P1_U4560
g1850 nand P1_R1150_U97 P1_U3994 ; P1_U4561
g1851 nand P1_R1117_U97 P1_U3996 ; P1_U4562
g1852 nand P1_R1138_U14 P1_U3995 ; P1_U4563
g1853 nand P1_R1192_U97 P1_U3992 ; P1_U4564
g1854 nand P1_R1207_U97 P1_U3991 ; P1_U4565
g1855 nand P1_R1171_U14 P1_U4001 ; P1_U4566
g1856 nand P1_R1240_U14 P1_U4000 ; P1_U4567
g1857 not P1_U3395 ; P1_U4568
g1858 nand P1_R1222_U14 P1_U3026 ; P1_U4569
g1859 nand P1_U3025 P1_U3073 ; P1_U4570
g1860 nand P1_R1282_U13 P1_U3023 ; P1_U4571
g1861 nand P1_U4015 P1_U4175 ; P1_U4572
g1862 nand P1_U3714 P1_U4568 ; P1_U4573
g1863 nand P1_U3018 P1_REG2_REG_22__SCAN_IN ; P1_U4574
g1864 nand P1_U3019 P1_REG1_REG_22__SCAN_IN ; P1_U4575
g1865 nand P1_U3020 P1_REG0_REG_22__SCAN_IN ; P1_U4576
g1866 nand P1_ADD_99_U66 P1_U3017 ; P1_U4577
g1867 not P1_U3059 ; P1_U4578
g1868 nand P1_U3033 P1_U3074 ; P1_U4579
g1869 nand P1_R1150_U111 P1_U3994 ; P1_U4580
g1870 nand P1_R1117_U111 P1_U3996 ; P1_U4581
g1871 nand P1_R1138_U15 P1_U3995 ; P1_U4582
g1872 nand P1_R1192_U111 P1_U3992 ; P1_U4583
g1873 nand P1_R1207_U111 P1_U3991 ; P1_U4584
g1874 nand P1_R1171_U15 P1_U4001 ; P1_U4585
g1875 nand P1_R1240_U15 P1_U4000 ; P1_U4586
g1876 not P1_U3397 ; P1_U4587
g1877 nand P1_R1222_U15 P1_U3026 ; P1_U4588
g1878 nand P1_U3025 P1_U3059 ; P1_U4589
g1879 nand P1_R1282_U78 P1_U3023 ; P1_U4590
g1880 nand P1_U4014 P1_U4175 ; P1_U4591
g1881 nand P1_U3718 P1_U4587 ; P1_U4592
g1882 nand P1_U3018 P1_REG2_REG_23__SCAN_IN ; P1_U4593
g1883 nand P1_U3019 P1_REG1_REG_23__SCAN_IN ; P1_U4594
g1884 nand P1_U3020 P1_REG0_REG_23__SCAN_IN ; P1_U4595
g1885 nand P1_ADD_99_U65 P1_U3017 ; P1_U4596
g1886 not P1_U3064 ; P1_U4597
g1887 nand P1_U3033 P1_U3073 ; P1_U4598
g1888 nand P1_R1150_U110 P1_U3994 ; P1_U4599
g1889 nand P1_R1117_U110 P1_U3996 ; P1_U4600
g1890 nand P1_R1138_U108 P1_U3995 ; P1_U4601
g1891 nand P1_R1192_U110 P1_U3992 ; P1_U4602
g1892 nand P1_R1207_U110 P1_U3991 ; P1_U4603
g1893 nand P1_R1171_U108 P1_U4001 ; P1_U4604
g1894 nand P1_R1240_U108 P1_U4000 ; P1_U4605
g1895 not P1_U3399 ; P1_U4606
g1896 nand P1_R1222_U108 P1_U3026 ; P1_U4607
g1897 nand P1_U3025 P1_U3064 ; P1_U4608
g1898 nand P1_R1282_U14 P1_U3023 ; P1_U4609
g1899 nand P1_U4013 P1_U4175 ; P1_U4610
g1900 nand P1_U3722 P1_U4606 ; P1_U4611
g1901 nand P1_U3018 P1_REG2_REG_24__SCAN_IN ; P1_U4612
g1902 nand P1_U3019 P1_REG1_REG_24__SCAN_IN ; P1_U4613
g1903 nand P1_U3020 P1_REG0_REG_24__SCAN_IN ; P1_U4614
g1904 nand P1_ADD_99_U64 P1_U3017 ; P1_U4615
g1905 not P1_U3063 ; P1_U4616
g1906 nand P1_U3033 P1_U3059 ; P1_U4617
g1907 nand P1_R1150_U15 P1_U3994 ; P1_U4618
g1908 nand P1_R1117_U15 P1_U3996 ; P1_U4619
g1909 nand P1_R1138_U107 P1_U3995 ; P1_U4620
g1910 nand P1_R1192_U15 P1_U3992 ; P1_U4621
g1911 nand P1_R1207_U15 P1_U3991 ; P1_U4622
g1912 nand P1_R1171_U107 P1_U4001 ; P1_U4623
g1913 nand P1_R1240_U107 P1_U4000 ; P1_U4624
g1914 not P1_U3401 ; P1_U4625
g1915 nand P1_R1222_U107 P1_U3026 ; P1_U4626
g1916 nand P1_U3025 P1_U3063 ; P1_U4627
g1917 nand P1_R1282_U76 P1_U3023 ; P1_U4628
g1918 nand P1_U4012 P1_U4175 ; P1_U4629
g1919 nand P1_U3726 P1_U4625 ; P1_U4630
g1920 nand P1_U3018 P1_REG2_REG_25__SCAN_IN ; P1_U4631
g1921 nand P1_U3019 P1_REG1_REG_25__SCAN_IN ; P1_U4632
g1922 nand P1_U3020 P1_REG0_REG_25__SCAN_IN ; P1_U4633
g1923 nand P1_ADD_99_U63 P1_U3017 ; P1_U4634
g1924 not P1_U3056 ; P1_U4635
g1925 nand P1_U3033 P1_U3064 ; P1_U4636
g1926 nand P1_R1150_U96 P1_U3994 ; P1_U4637
g1927 nand P1_R1117_U96 P1_U3996 ; P1_U4638
g1928 nand P1_R1138_U106 P1_U3995 ; P1_U4639
g1929 nand P1_R1192_U96 P1_U3992 ; P1_U4640
g1930 nand P1_R1207_U96 P1_U3991 ; P1_U4641
g1931 nand P1_R1171_U106 P1_U4001 ; P1_U4642
g1932 nand P1_R1240_U106 P1_U4000 ; P1_U4643
g1933 not P1_U3403 ; P1_U4644
g1934 nand P1_R1222_U106 P1_U3026 ; P1_U4645
g1935 nand P1_U3025 P1_U3056 ; P1_U4646
g1936 nand P1_R1282_U15 P1_U3023 ; P1_U4647
g1937 nand P1_U4011 P1_U4175 ; P1_U4648
g1938 nand P1_U3730 P1_U4644 ; P1_U4649
g1939 nand P1_U3018 P1_REG2_REG_26__SCAN_IN ; P1_U4650
g1940 nand P1_U3019 P1_REG1_REG_26__SCAN_IN ; P1_U4651
g1941 nand P1_U3020 P1_REG0_REG_26__SCAN_IN ; P1_U4652
g1942 nand P1_ADD_99_U62 P1_U3017 ; P1_U4653
g1943 not P1_U3055 ; P1_U4654
g1944 nand P1_U3033 P1_U3063 ; P1_U4655
g1945 nand P1_R1150_U95 P1_U3994 ; P1_U4656
g1946 nand P1_R1117_U95 P1_U3996 ; P1_U4657
g1947 nand P1_R1138_U105 P1_U3995 ; P1_U4658
g1948 nand P1_R1192_U95 P1_U3992 ; P1_U4659
g1949 nand P1_R1207_U95 P1_U3991 ; P1_U4660
g1950 nand P1_R1171_U105 P1_U4001 ; P1_U4661
g1951 nand P1_R1240_U105 P1_U4000 ; P1_U4662
g1952 not P1_U3405 ; P1_U4663
g1953 nand P1_R1222_U105 P1_U3026 ; P1_U4664
g1954 nand P1_U3025 P1_U3055 ; P1_U4665
g1955 nand P1_R1282_U74 P1_U3023 ; P1_U4666
g1956 nand P1_U4010 P1_U4175 ; P1_U4667
g1957 nand P1_U3734 P1_U4663 ; P1_U4668
g1958 nand P1_U3018 P1_REG2_REG_27__SCAN_IN ; P1_U4669
g1959 nand P1_U3019 P1_REG1_REG_27__SCAN_IN ; P1_U4670
g1960 nand P1_U3020 P1_REG0_REG_27__SCAN_IN ; P1_U4671
g1961 nand P1_ADD_99_U61 P1_U3017 ; P1_U4672
g1962 not P1_U3051 ; P1_U4673
g1963 nand P1_U3033 P1_U3056 ; P1_U4674
g1964 nand P1_R1150_U109 P1_U3994 ; P1_U4675
g1965 nand P1_R1117_U109 P1_U3996 ; P1_U4676
g1966 nand P1_R1138_U16 P1_U3995 ; P1_U4677
g1967 nand P1_R1192_U109 P1_U3992 ; P1_U4678
g1968 nand P1_R1207_U109 P1_U3991 ; P1_U4679
g1969 nand P1_R1171_U16 P1_U4001 ; P1_U4680
g1970 nand P1_R1240_U16 P1_U4000 ; P1_U4681
g1971 not P1_U3407 ; P1_U4682
g1972 nand P1_R1222_U16 P1_U3026 ; P1_U4683
g1973 nand P1_U3025 P1_U3051 ; P1_U4684
g1974 nand P1_R1282_U16 P1_U3023 ; P1_U4685
g1975 nand P1_U4009 P1_U4175 ; P1_U4686
g1976 nand P1_U3738 P1_U4682 ; P1_U4687
g1977 nand P1_U3018 P1_REG2_REG_28__SCAN_IN ; P1_U4688
g1978 nand P1_U3019 P1_REG1_REG_28__SCAN_IN ; P1_U4689
g1979 nand P1_U3020 P1_REG0_REG_28__SCAN_IN ; P1_U4690
g1980 nand P1_ADD_99_U60 P1_U3017 ; P1_U4691
g1981 not P1_U3052 ; P1_U4692
g1982 nand P1_U3033 P1_U3055 ; P1_U4693
g1983 nand P1_R1150_U16 P1_U3994 ; P1_U4694
g1984 nand P1_R1117_U16 P1_U3996 ; P1_U4695
g1985 nand P1_R1138_U104 P1_U3995 ; P1_U4696
g1986 nand P1_R1192_U16 P1_U3992 ; P1_U4697
g1987 nand P1_R1207_U16 P1_U3991 ; P1_U4698
g1988 nand P1_R1171_U104 P1_U4001 ; P1_U4699
g1989 nand P1_R1240_U104 P1_U4000 ; P1_U4700
g1990 not P1_U3409 ; P1_U4701
g1991 nand P1_R1222_U104 P1_U3026 ; P1_U4702
g1992 nand P1_U3025 P1_U3052 ; P1_U4703
g1993 nand P1_R1282_U72 P1_U3023 ; P1_U4704
g1994 nand P1_U4008 P1_U4175 ; P1_U4705
g1995 nand P1_U3742 P1_U4701 ; P1_U4706
g1996 nand P1_ADD_99_U5 P1_U3017 ; P1_U4707
g1997 nand P1_U3018 P1_REG2_REG_29__SCAN_IN ; P1_U4708
g1998 nand P1_U3019 P1_REG1_REG_29__SCAN_IN ; P1_U4709
g1999 nand P1_U3020 P1_REG0_REG_29__SCAN_IN ; P1_U4710
g2000 not P1_U3053 ; P1_U4711
g2001 nand P1_U3033 P1_U3051 ; P1_U4712
g2002 nand P1_R1150_U94 P1_U3994 ; P1_U4713
g2003 nand P1_R1117_U94 P1_U3996 ; P1_U4714
g2004 nand P1_R1138_U103 P1_U3995 ; P1_U4715
g2005 nand P1_R1192_U94 P1_U3992 ; P1_U4716
g2006 nand P1_R1207_U94 P1_U3991 ; P1_U4717
g2007 nand P1_R1171_U103 P1_U4001 ; P1_U4718
g2008 nand P1_R1240_U103 P1_U4000 ; P1_U4719
g2009 not P1_U3411 ; P1_U4720
g2010 nand P1_R1222_U103 P1_U3026 ; P1_U4721
g2011 nand P1_U3025 P1_U3053 ; P1_U4722
g2012 nand P1_R1282_U17 P1_U3023 ; P1_U4723
g2013 nand P1_U4007 P1_U4175 ; P1_U4724
g2014 nand P1_U3746 P1_U4720 ; P1_U4725
g2015 nand P1_U3018 P1_REG2_REG_30__SCAN_IN ; P1_U4726
g2016 nand P1_U3019 P1_REG1_REG_30__SCAN_IN ; P1_U4727
g2017 nand P1_U3020 P1_REG0_REG_30__SCAN_IN ; P1_U4728
g2018 not P1_U3057 ; P1_U4729
g2019 nand P1_U5728 P1_U3358 ; P1_U4730
g2020 nand P1_U3946 P1_U4730 ; P1_U4731
g2021 nand P1_U3747 P1_U3057 ; P1_U4732
g2022 nand P1_U3033 P1_U3052 ; P1_U4733
g2023 nand P1_R1150_U17 P1_U3994 ; P1_U4734
g2024 nand P1_R1117_U17 P1_U3996 ; P1_U4735
g2025 nand P1_R1138_U102 P1_U3995 ; P1_U4736
g2026 nand P1_R1192_U17 P1_U3992 ; P1_U4737
g2027 nand P1_R1207_U17 P1_U3991 ; P1_U4738
g2028 nand P1_R1171_U102 P1_U4001 ; P1_U4739
g2029 nand P1_R1240_U102 P1_U4000 ; P1_U4740
g2030 not P1_U3413 ; P1_U4741
g2031 nand P1_R1222_U102 P1_U3026 ; P1_U4742
g2032 nand P1_R1282_U70 P1_U3023 ; P1_U4743
g2033 nand P1_U4018 P1_U4175 ; P1_U4744
g2034 nand P1_U3751 P1_U4741 ; P1_U4745
g2035 nand P1_U3018 P1_REG2_REG_31__SCAN_IN ; P1_U4746
g2036 nand P1_U3019 P1_REG1_REG_31__SCAN_IN ; P1_U4747
g2037 nand P1_U3020 P1_REG0_REG_31__SCAN_IN ; P1_U4748
g2038 not P1_U3054 ; P1_U4749
g2039 nand P1_R1282_U19 P1_U3023 ; P1_U4750
g2040 nand P1_U4017 P1_U4175 ; P1_U4751
g2041 nand P1_U4751 P1_U3979 P1_U4750 ; P1_U4752
g2042 nand P1_R1282_U68 P1_U3023 ; P1_U4753
g2043 nand P1_U4016 P1_U4175 ; P1_U4754
g2044 nand P1_U4754 P1_U3979 P1_U4753 ; P1_U4755
g2045 nand P1_U3754 P1_U3016 ; P1_U4756
g2046 nand P1_U3418 P1_U4756 ; P1_U4757
g2047 nand P1_U4021 P1_U3442 ; P1_U4758
g2048 not P1_U3422 ; P1_U4759
g2049 nand P1_U3035 P1_U3076 ; P1_U4760
g2050 nand P1_U3032 P1_REG3_REG_0__SCAN_IN ; P1_U4761
g2051 nand P1_U3031 P1_R1222_U96 ; P1_U4762
g2052 nand P1_U3030 P1_U3451 ; P1_U4763
g2053 nand P1_U3029 P1_U3451 ; P1_U4764
g2054 nand P1_U3035 P1_U3066 ; P1_U4765
g2055 nand P1_U3032 P1_REG3_REG_1__SCAN_IN ; P1_U4766
g2056 nand P1_U3031 P1_R1222_U95 ; P1_U4767
g2057 nand P1_U3030 P1_U3456 ; P1_U4768
g2058 nand P1_U3029 P1_R1282_U57 ; P1_U4769
g2059 nand P1_U3035 P1_U3062 ; P1_U4770
g2060 nand P1_U3032 P1_REG3_REG_2__SCAN_IN ; P1_U4771
g2061 nand P1_U3031 P1_R1222_U17 ; P1_U4772
g2062 nand P1_U3030 P1_U3459 ; P1_U4773
g2063 nand P1_U3029 P1_R1282_U18 ; P1_U4774
g2064 nand P1_U3035 P1_U3058 ; P1_U4775
g2065 nand P1_U3032 P1_ADD_99_U4 ; P1_U4776
g2066 nand P1_U3031 P1_R1222_U101 ; P1_U4777
g2067 nand P1_U3030 P1_U3462 ; P1_U4778
g2068 nand P1_U3029 P1_R1282_U20 ; P1_U4779
g2069 nand P1_U3035 P1_U3065 ; P1_U4780
g2070 nand P1_U3032 P1_ADD_99_U59 ; P1_U4781
g2071 nand P1_U3031 P1_R1222_U100 ; P1_U4782
g2072 nand P1_U3030 P1_U3465 ; P1_U4783
g2073 nand P1_U3029 P1_R1282_U21 ; P1_U4784
g2074 nand P1_U3035 P1_U3069 ; P1_U4785
g2075 nand P1_U3032 P1_ADD_99_U58 ; P1_U4786
g2076 nand P1_U3031 P1_R1222_U18 ; P1_U4787
g2077 nand P1_U3030 P1_U3468 ; P1_U4788
g2078 nand P1_U3029 P1_R1282_U65 ; P1_U4789
g2079 nand P1_U3035 P1_U3068 ; P1_U4790
g2080 nand P1_U3032 P1_ADD_99_U57 ; P1_U4791
g2081 nand P1_U3031 P1_R1222_U99 ; P1_U4792
g2082 nand P1_U3030 P1_U3471 ; P1_U4793
g2083 nand P1_U3029 P1_R1282_U22 ; P1_U4794
g2084 nand P1_U3035 P1_U3082 ; P1_U4795
g2085 nand P1_U3032 P1_ADD_99_U56 ; P1_U4796
g2086 nand P1_U3031 P1_R1222_U19 ; P1_U4797
g2087 nand P1_U3030 P1_U3474 ; P1_U4798
g2088 nand P1_U3029 P1_R1282_U23 ; P1_U4799
g2089 nand P1_U3035 P1_U3081 ; P1_U4800
g2090 nand P1_U3032 P1_ADD_99_U55 ; P1_U4801
g2091 nand P1_U3031 P1_R1222_U98 ; P1_U4802
g2092 nand P1_U3030 P1_U3477 ; P1_U4803
g2093 nand P1_U3029 P1_R1282_U24 ; P1_U4804
g2094 nand P1_U3035 P1_U3060 ; P1_U4805
g2095 nand P1_U3032 P1_ADD_99_U54 ; P1_U4806
g2096 nand P1_U3031 P1_R1222_U97 ; P1_U4807
g2097 nand P1_U3030 P1_U3480 ; P1_U4808
g2098 nand P1_U3029 P1_R1282_U63 ; P1_U4809
g2099 nand P1_U3035 P1_U3061 ; P1_U4810
g2100 nand P1_U3032 P1_ADD_99_U78 ; P1_U4811
g2101 nand P1_U3031 P1_R1222_U11 ; P1_U4812
g2102 nand P1_U3030 P1_U3483 ; P1_U4813
g2103 nand P1_U3029 P1_R1282_U6 ; P1_U4814
g2104 nand P1_U3035 P1_U3070 ; P1_U4815
g2105 nand P1_U3032 P1_ADD_99_U77 ; P1_U4816
g2106 nand P1_U3031 P1_R1222_U115 ; P1_U4817
g2107 nand P1_U3030 P1_U3486 ; P1_U4818
g2108 nand P1_U3029 P1_R1282_U7 ; P1_U4819
g2109 nand P1_U3035 P1_U3078 ; P1_U4820
g2110 nand P1_U3032 P1_ADD_99_U76 ; P1_U4821
g2111 nand P1_U3031 P1_R1222_U114 ; P1_U4822
g2112 nand P1_U3030 P1_U3489 ; P1_U4823
g2113 nand P1_U3029 P1_R1282_U8 ; P1_U4824
g2114 nand P1_U3035 P1_U3077 ; P1_U4825
g2115 nand P1_U3032 P1_ADD_99_U75 ; P1_U4826
g2116 nand P1_U3031 P1_R1222_U12 ; P1_U4827
g2117 nand P1_U3030 P1_U3492 ; P1_U4828
g2118 nand P1_U3029 P1_R1282_U86 ; P1_U4829
g2119 nand P1_U3035 P1_U3072 ; P1_U4830
g2120 nand P1_U3032 P1_ADD_99_U74 ; P1_U4831
g2121 nand P1_U3031 P1_R1222_U113 ; P1_U4832
g2122 nand P1_U3030 P1_U3495 ; P1_U4833
g2123 nand P1_U3029 P1_R1282_U9 ; P1_U4834
g2124 nand P1_U3035 P1_U3071 ; P1_U4835
g2125 nand P1_U3032 P1_ADD_99_U73 ; P1_U4836
g2126 nand P1_U3031 P1_R1222_U112 ; P1_U4837
g2127 nand P1_U3030 P1_U3498 ; P1_U4838
g2128 nand P1_U3029 P1_R1282_U10 ; P1_U4839
g2129 nand P1_U3035 P1_U3067 ; P1_U4840
g2130 nand P1_U3032 P1_ADD_99_U72 ; P1_U4841
g2131 nand P1_U3031 P1_R1222_U111 ; P1_U4842
g2132 nand P1_U3030 P1_U3501 ; P1_U4843
g2133 nand P1_U3029 P1_R1282_U11 ; P1_U4844
g2134 nand P1_U3035 P1_U3080 ; P1_U4845
g2135 nand P1_U3032 P1_ADD_99_U71 ; P1_U4846
g2136 nand P1_U3031 P1_R1222_U13 ; P1_U4847
g2137 nand P1_U3030 P1_U3504 ; P1_U4848
g2138 nand P1_U3029 P1_R1282_U84 ; P1_U4849
g2139 nand P1_U3035 P1_U3079 ; P1_U4850
g2140 nand P1_U3032 P1_ADD_99_U70 ; P1_U4851
g2141 nand P1_U3031 P1_R1222_U110 ; P1_U4852
g2142 nand P1_U3030 P1_U3507 ; P1_U4853
g2143 nand P1_U3029 P1_R1282_U12 ; P1_U4854
g2144 nand P1_U3035 P1_U3074 ; P1_U4855
g2145 nand P1_U3032 P1_ADD_99_U69 ; P1_U4856
g2146 nand P1_U3031 P1_R1222_U109 ; P1_U4857
g2147 nand P1_U3030 P1_U3509 ; P1_U4858
g2148 nand P1_U3029 P1_R1282_U82 ; P1_U4859
g2149 nand P1_U3035 P1_U3073 ; P1_U4860
g2150 nand P1_U3032 P1_ADD_99_U68 ; P1_U4861
g2151 nand P1_U3031 P1_R1222_U14 ; P1_U4862
g2152 nand P1_U3030 P1_U4015 ; P1_U4863
g2153 nand P1_U3029 P1_R1282_U13 ; P1_U4864
g2154 nand P1_U3035 P1_U3059 ; P1_U4865
g2155 nand P1_U3032 P1_ADD_99_U67 ; P1_U4866
g2156 nand P1_U3031 P1_R1222_U15 ; P1_U4867
g2157 nand P1_U3030 P1_U4014 ; P1_U4868
g2158 nand P1_U3029 P1_R1282_U78 ; P1_U4869
g2159 nand P1_U3035 P1_U3064 ; P1_U4870
g2160 nand P1_U3032 P1_ADD_99_U66 ; P1_U4871
g2161 nand P1_U3031 P1_R1222_U108 ; P1_U4872
g2162 nand P1_U3030 P1_U4013 ; P1_U4873
g2163 nand P1_U3029 P1_R1282_U14 ; P1_U4874
g2164 nand P1_U3035 P1_U3063 ; P1_U4875
g2165 nand P1_U3032 P1_ADD_99_U65 ; P1_U4876
g2166 nand P1_U3031 P1_R1222_U107 ; P1_U4877
g2167 nand P1_U3030 P1_U4012 ; P1_U4878
g2168 nand P1_U3029 P1_R1282_U76 ; P1_U4879
g2169 nand P1_U3035 P1_U3056 ; P1_U4880
g2170 nand P1_U3032 P1_ADD_99_U64 ; P1_U4881
g2171 nand P1_U3031 P1_R1222_U106 ; P1_U4882
g2172 nand P1_U3030 P1_U4011 ; P1_U4883
g2173 nand P1_U3029 P1_R1282_U15 ; P1_U4884
g2174 nand P1_U3035 P1_U3055 ; P1_U4885
g2175 nand P1_U3032 P1_ADD_99_U63 ; P1_U4886
g2176 nand P1_U3031 P1_R1222_U105 ; P1_U4887
g2177 nand P1_U3030 P1_U4010 ; P1_U4888
g2178 nand P1_U3029 P1_R1282_U74 ; P1_U4889
g2179 nand P1_U3035 P1_U3051 ; P1_U4890
g2180 nand P1_U3032 P1_ADD_99_U62 ; P1_U4891
g2181 nand P1_U3031 P1_R1222_U16 ; P1_U4892
g2182 nand P1_U3030 P1_U4009 ; P1_U4893
g2183 nand P1_U3029 P1_R1282_U16 ; P1_U4894
g2184 nand P1_U3035 P1_U3052 ; P1_U4895
g2185 nand P1_U3032 P1_ADD_99_U61 ; P1_U4896
g2186 nand P1_U3031 P1_R1222_U104 ; P1_U4897
g2187 nand P1_U3030 P1_U4008 ; P1_U4898
g2188 nand P1_U3029 P1_R1282_U72 ; P1_U4899
g2189 nand P1_U3035 P1_U3053 ; P1_U4900
g2190 nand P1_U3032 P1_ADD_99_U60 ; P1_U4901
g2191 nand P1_U3031 P1_R1222_U103 ; P1_U4902
g2192 nand P1_U3030 P1_U4007 ; P1_U4903
g2193 nand P1_U3029 P1_R1282_U17 ; P1_U4904
g2194 nand P1_U3032 P1_ADD_99_U5 ; P1_U4905
g2195 nand P1_U3031 P1_R1222_U102 ; P1_U4906
g2196 nand P1_U3030 P1_U4018 ; P1_U4907
g2197 nand P1_U3029 P1_R1282_U70 ; P1_U4908
g2198 nand P1_U3030 P1_U4017 ; P1_U4909
g2199 nand P1_U3029 P1_R1282_U19 ; P1_U4910
g2200 nand P1_U3030 P1_U4016 ; P1_U4911
g2201 nand P1_U3029 P1_R1282_U68 ; P1_U4912
g2202 nand P1_U3814 P1_U3813 P1_U3816 P1_U4759 P1_U3418 ; P1_U4913
g2203 nand P1_R1105_U13 P1_U3041 ; P1_U4914
g2204 nand P1_U3039 P1_U3443 ; P1_U4915
g2205 nand P1_R1162_U13 P1_U3037 ; P1_U4916
g2206 nand P1_U4915 P1_U4914 P1_U4916 ; P1_U4917
g2207 nand P1_U3046 P1_U3372 ; P1_U4918
g2208 nand P1_U5703 P1_U4918 ; P1_U4919
g2209 nand P1_U4919 P1_U3946 ; P1_U4920
g2210 not P1_U3083 ; P1_U4921
g2211 not P1_U3423 ; P1_U4922
g2212 nand P1_U3043 P1_U4917 ; P1_U4923
g2213 nand P1_U3042 P1_R1105_U13 ; P1_U4924
g2214 nand P1_U3084 P1_REG3_REG_19__SCAN_IN ; P1_U4925
g2215 nand P1_U3040 P1_U3443 ; P1_U4926
g2216 nand P1_U3038 P1_R1162_U13 ; P1_U4927
g2217 nand P1_U4922 P1_ADDR_REG_19__SCAN_IN ; P1_U4928
g2218 nand P1_R1105_U75 P1_U3041 ; P1_U4929
g2219 nand P1_U3039 P1_U3506 ; P1_U4930
g2220 nand P1_R1162_U75 P1_U3037 ; P1_U4931
g2221 nand P1_U4930 P1_U4929 P1_U4931 ; P1_U4932
g2222 nand P1_U3043 P1_U4932 ; P1_U4933
g2223 nand P1_R1105_U75 P1_U3042 ; P1_U4934
g2224 nand P1_U3084 P1_REG3_REG_18__SCAN_IN ; P1_U4935
g2225 nand P1_U3040 P1_U3506 ; P1_U4936
g2226 nand P1_R1162_U75 P1_U3038 ; P1_U4937
g2227 nand P1_U4922 P1_ADDR_REG_18__SCAN_IN ; P1_U4938
g2228 nand P1_R1105_U12 P1_U3041 ; P1_U4939
g2229 nand P1_U3039 P1_U3503 ; P1_U4940
g2230 nand P1_R1162_U12 P1_U3037 ; P1_U4941
g2231 nand P1_U4940 P1_U4939 P1_U4941 ; P1_U4942
g2232 nand P1_U3043 P1_U4942 ; P1_U4943
g2233 nand P1_R1105_U12 P1_U3042 ; P1_U4944
g2234 nand P1_U3084 P1_REG3_REG_17__SCAN_IN ; P1_U4945
g2235 nand P1_U3040 P1_U3503 ; P1_U4946
g2236 nand P1_R1162_U12 P1_U3038 ; P1_U4947
g2237 nand P1_U4922 P1_ADDR_REG_17__SCAN_IN ; P1_U4948
g2238 nand P1_R1105_U76 P1_U3041 ; P1_U4949
g2239 nand P1_U3039 P1_U3500 ; P1_U4950
g2240 nand P1_R1162_U76 P1_U3037 ; P1_U4951
g2241 nand P1_U4950 P1_U4949 P1_U4951 ; P1_U4952
g2242 nand P1_U3043 P1_U4952 ; P1_U4953
g2243 nand P1_R1105_U76 P1_U3042 ; P1_U4954
g2244 nand P1_U3084 P1_REG3_REG_16__SCAN_IN ; P1_U4955
g2245 nand P1_U3040 P1_U3500 ; P1_U4956
g2246 nand P1_R1162_U76 P1_U3038 ; P1_U4957
g2247 nand P1_U4922 P1_ADDR_REG_16__SCAN_IN ; P1_U4958
g2248 nand P1_R1105_U77 P1_U3041 ; P1_U4959
g2249 nand P1_U3039 P1_U3497 ; P1_U4960
g2250 nand P1_R1162_U77 P1_U3037 ; P1_U4961
g2251 nand P1_U4960 P1_U4959 P1_U4961 ; P1_U4962
g2252 nand P1_U3043 P1_U4962 ; P1_U4963
g2253 nand P1_R1105_U77 P1_U3042 ; P1_U4964
g2254 nand P1_U3084 P1_REG3_REG_15__SCAN_IN ; P1_U4965
g2255 nand P1_U3040 P1_U3497 ; P1_U4966
g2256 nand P1_R1162_U77 P1_U3038 ; P1_U4967
g2257 nand P1_U4922 P1_ADDR_REG_15__SCAN_IN ; P1_U4968
g2258 nand P1_R1105_U78 P1_U3041 ; P1_U4969
g2259 nand P1_U3039 P1_U3494 ; P1_U4970
g2260 nand P1_R1162_U78 P1_U3037 ; P1_U4971
g2261 nand P1_U4970 P1_U4969 P1_U4971 ; P1_U4972
g2262 nand P1_U3043 P1_U4972 ; P1_U4973
g2263 nand P1_R1105_U78 P1_U3042 ; P1_U4974
g2264 nand P1_U3084 P1_REG3_REG_14__SCAN_IN ; P1_U4975
g2265 nand P1_U3040 P1_U3494 ; P1_U4976
g2266 nand P1_R1162_U78 P1_U3038 ; P1_U4977
g2267 nand P1_U4922 P1_ADDR_REG_14__SCAN_IN ; P1_U4978
g2268 nand P1_R1105_U11 P1_U3041 ; P1_U4979
g2269 nand P1_U3039 P1_U3491 ; P1_U4980
g2270 nand P1_R1162_U11 P1_U3037 ; P1_U4981
g2271 nand P1_U4980 P1_U4979 P1_U4981 ; P1_U4982
g2272 nand P1_U3043 P1_U4982 ; P1_U4983
g2273 nand P1_R1105_U11 P1_U3042 ; P1_U4984
g2274 nand P1_U3084 P1_REG3_REG_13__SCAN_IN ; P1_U4985
g2275 nand P1_U3040 P1_U3491 ; P1_U4986
g2276 nand P1_R1162_U11 P1_U3038 ; P1_U4987
g2277 nand P1_U4922 P1_ADDR_REG_13__SCAN_IN ; P1_U4988
g2278 nand P1_R1105_U79 P1_U3041 ; P1_U4989
g2279 nand P1_U3039 P1_U3488 ; P1_U4990
g2280 nand P1_R1162_U79 P1_U3037 ; P1_U4991
g2281 nand P1_U4990 P1_U4989 P1_U4991 ; P1_U4992
g2282 nand P1_U3043 P1_U4992 ; P1_U4993
g2283 nand P1_R1105_U79 P1_U3042 ; P1_U4994
g2284 nand P1_U3084 P1_REG3_REG_12__SCAN_IN ; P1_U4995
g2285 nand P1_U3040 P1_U3488 ; P1_U4996
g2286 nand P1_R1162_U79 P1_U3038 ; P1_U4997
g2287 nand P1_U4922 P1_ADDR_REG_12__SCAN_IN ; P1_U4998
g2288 nand P1_R1105_U80 P1_U3041 ; P1_U4999
g2289 nand P1_U3039 P1_U3485 ; P1_U5000
g2290 nand P1_R1162_U80 P1_U3037 ; P1_U5001
g2291 nand P1_U5000 P1_U4999 P1_U5001 ; P1_U5002
g2292 nand P1_U3043 P1_U5002 ; P1_U5003
g2293 nand P1_R1105_U80 P1_U3042 ; P1_U5004
g2294 nand P1_U3084 P1_REG3_REG_11__SCAN_IN ; P1_U5005
g2295 nand P1_U3040 P1_U3485 ; P1_U5006
g2296 nand P1_R1162_U80 P1_U3038 ; P1_U5007
g2297 nand P1_U4922 P1_ADDR_REG_11__SCAN_IN ; P1_U5008
g2298 nand P1_R1105_U10 P1_U3041 ; P1_U5009
g2299 nand P1_U3039 P1_U3482 ; P1_U5010
g2300 nand P1_R1162_U10 P1_U3037 ; P1_U5011
g2301 nand P1_U5010 P1_U5009 P1_U5011 ; P1_U5012
g2302 nand P1_U3043 P1_U5012 ; P1_U5013
g2303 nand P1_R1105_U10 P1_U3042 ; P1_U5014
g2304 nand P1_U3084 P1_REG3_REG_10__SCAN_IN ; P1_U5015
g2305 nand P1_U3040 P1_U3482 ; P1_U5016
g2306 nand P1_R1162_U10 P1_U3038 ; P1_U5017
g2307 nand P1_U4922 P1_ADDR_REG_10__SCAN_IN ; P1_U5018
g2308 nand P1_R1105_U70 P1_U3041 ; P1_U5019
g2309 nand P1_U3039 P1_U3479 ; P1_U5020
g2310 nand P1_R1162_U70 P1_U3037 ; P1_U5021
g2311 nand P1_U5020 P1_U5019 P1_U5021 ; P1_U5022
g2312 nand P1_U3043 P1_U5022 ; P1_U5023
g2313 nand P1_R1105_U70 P1_U3042 ; P1_U5024
g2314 nand P1_U3084 P1_REG3_REG_9__SCAN_IN ; P1_U5025
g2315 nand P1_U3040 P1_U3479 ; P1_U5026
g2316 nand P1_R1162_U70 P1_U3038 ; P1_U5027
g2317 nand P1_U4922 P1_ADDR_REG_9__SCAN_IN ; P1_U5028
g2318 nand P1_R1105_U71 P1_U3041 ; P1_U5029
g2319 nand P1_U3039 P1_U3476 ; P1_U5030
g2320 nand P1_R1162_U71 P1_U3037 ; P1_U5031
g2321 nand P1_U5030 P1_U5029 P1_U5031 ; P1_U5032
g2322 nand P1_U3043 P1_U5032 ; P1_U5033
g2323 nand P1_R1105_U71 P1_U3042 ; P1_U5034
g2324 nand P1_U3084 P1_REG3_REG_8__SCAN_IN ; P1_U5035
g2325 nand P1_U3040 P1_U3476 ; P1_U5036
g2326 nand P1_R1162_U71 P1_U3038 ; P1_U5037
g2327 nand P1_U4922 P1_ADDR_REG_8__SCAN_IN ; P1_U5038
g2328 nand P1_R1105_U16 P1_U3041 ; P1_U5039
g2329 nand P1_U3039 P1_U3473 ; P1_U5040
g2330 nand P1_R1162_U16 P1_U3037 ; P1_U5041
g2331 nand P1_U5040 P1_U5039 P1_U5041 ; P1_U5042
g2332 nand P1_U3043 P1_U5042 ; P1_U5043
g2333 nand P1_R1105_U16 P1_U3042 ; P1_U5044
g2334 nand P1_U3084 P1_REG3_REG_7__SCAN_IN ; P1_U5045
g2335 nand P1_U3040 P1_U3473 ; P1_U5046
g2336 nand P1_R1162_U16 P1_U3038 ; P1_U5047
g2337 nand P1_U4922 P1_ADDR_REG_7__SCAN_IN ; P1_U5048
g2338 nand P1_R1105_U72 P1_U3041 ; P1_U5049
g2339 nand P1_U3039 P1_U3470 ; P1_U5050
g2340 nand P1_R1162_U72 P1_U3037 ; P1_U5051
g2341 nand P1_U5050 P1_U5049 P1_U5051 ; P1_U5052
g2342 nand P1_U3043 P1_U5052 ; P1_U5053
g2343 nand P1_R1105_U72 P1_U3042 ; P1_U5054
g2344 nand P1_U3084 P1_REG3_REG_6__SCAN_IN ; P1_U5055
g2345 nand P1_U3040 P1_U3470 ; P1_U5056
g2346 nand P1_R1162_U72 P1_U3038 ; P1_U5057
g2347 nand P1_U4922 P1_ADDR_REG_6__SCAN_IN ; P1_U5058
g2348 nand P1_R1105_U15 P1_U3041 ; P1_U5059
g2349 nand P1_U3039 P1_U3467 ; P1_U5060
g2350 nand P1_R1162_U15 P1_U3037 ; P1_U5061
g2351 nand P1_U5060 P1_U5059 P1_U5061 ; P1_U5062
g2352 nand P1_U3043 P1_U5062 ; P1_U5063
g2353 nand P1_R1105_U15 P1_U3042 ; P1_U5064
g2354 nand P1_U3084 P1_REG3_REG_5__SCAN_IN ; P1_U5065
g2355 nand P1_U3040 P1_U3467 ; P1_U5066
g2356 nand P1_R1162_U15 P1_U3038 ; P1_U5067
g2357 nand P1_U4922 P1_ADDR_REG_5__SCAN_IN ; P1_U5068
g2358 nand P1_R1105_U73 P1_U3041 ; P1_U5069
g2359 nand P1_U3039 P1_U3464 ; P1_U5070
g2360 nand P1_R1162_U73 P1_U3037 ; P1_U5071
g2361 nand P1_U5070 P1_U5069 P1_U5071 ; P1_U5072
g2362 nand P1_U3043 P1_U5072 ; P1_U5073
g2363 nand P1_R1105_U73 P1_U3042 ; P1_U5074
g2364 nand P1_U3084 P1_REG3_REG_4__SCAN_IN ; P1_U5075
g2365 nand P1_U3040 P1_U3464 ; P1_U5076
g2366 nand P1_R1162_U73 P1_U3038 ; P1_U5077
g2367 nand P1_U4922 P1_ADDR_REG_4__SCAN_IN ; P1_U5078
g2368 nand P1_R1105_U74 P1_U3041 ; P1_U5079
g2369 nand P1_U3039 P1_U3461 ; P1_U5080
g2370 nand P1_R1162_U74 P1_U3037 ; P1_U5081
g2371 nand P1_U5080 P1_U5079 P1_U5081 ; P1_U5082
g2372 nand P1_U3043 P1_U5082 ; P1_U5083
g2373 nand P1_R1105_U74 P1_U3042 ; P1_U5084
g2374 nand P1_U3084 P1_REG3_REG_3__SCAN_IN ; P1_U5085
g2375 nand P1_U3040 P1_U3461 ; P1_U5086
g2376 nand P1_R1162_U74 P1_U3038 ; P1_U5087
g2377 nand P1_U4922 P1_ADDR_REG_3__SCAN_IN ; P1_U5088
g2378 nand P1_R1105_U14 P1_U3041 ; P1_U5089
g2379 nand P1_U3039 P1_U3458 ; P1_U5090
g2380 nand P1_R1162_U14 P1_U3037 ; P1_U5091
g2381 nand P1_U5090 P1_U5089 P1_U5091 ; P1_U5092
g2382 nand P1_U3043 P1_U5092 ; P1_U5093
g2383 nand P1_R1105_U14 P1_U3042 ; P1_U5094
g2384 nand P1_U3084 P1_REG3_REG_2__SCAN_IN ; P1_U5095
g2385 nand P1_U3040 P1_U3458 ; P1_U5096
g2386 nand P1_R1162_U14 P1_U3038 ; P1_U5097
g2387 nand P1_U4922 P1_ADDR_REG_2__SCAN_IN ; P1_U5098
g2388 nand P1_R1105_U68 P1_U3041 ; P1_U5099
g2389 nand P1_U3039 P1_U3455 ; P1_U5100
g2390 nand P1_R1162_U68 P1_U3037 ; P1_U5101
g2391 nand P1_U5100 P1_U5099 P1_U5101 ; P1_U5102
g2392 nand P1_U3043 P1_U5102 ; P1_U5103
g2393 nand P1_R1105_U68 P1_U3042 ; P1_U5104
g2394 nand P1_U3084 P1_REG3_REG_1__SCAN_IN ; P1_U5105
g2395 nand P1_U3040 P1_U3455 ; P1_U5106
g2396 nand P1_R1162_U68 P1_U3038 ; P1_U5107
g2397 nand P1_U4922 P1_ADDR_REG_1__SCAN_IN ; P1_U5108
g2398 nand P1_R1105_U69 P1_U3041 ; P1_U5109
g2399 nand P1_U3039 P1_U3449 ; P1_U5110
g2400 nand P1_R1162_U69 P1_U3037 ; P1_U5111
g2401 nand P1_U5110 P1_U5109 P1_U5111 ; P1_U5112
g2402 nand P1_U3043 P1_U5112 ; P1_U5113
g2403 nand P1_R1105_U69 P1_U3042 ; P1_U5114
g2404 nand P1_U3084 P1_REG3_REG_0__SCAN_IN ; P1_U5115
g2405 nand P1_U3040 P1_U3449 ; P1_U5116
g2406 nand P1_R1162_U69 P1_U3038 ; P1_U5117
g2407 nand P1_U4922 P1_ADDR_REG_0__SCAN_IN ; P1_U5118
g2408 not P1_U3982 ; P1_U5119
g2409 nand P1_U6198 P1_U6197 P1_U3875 ; P1_U5120
g2410 nand P1_U5703 P1_U3427 ; P1_U5121
g2411 nand P1_U3861 P1_U5121 ; P1_U5122
g2412 nand P1_U5122 P1_B_REG_SCAN_IN ; P1_U5123
g2413 nand P1_U3036 P1_U3077 ; P1_U5124
g2414 nand P1_U3034 P1_U3071 ; P1_U5125
g2415 nand P1_ADD_99_U73 P1_U3431 ; P1_U5126
g2416 nand P1_U5126 P1_U5124 P1_U5125 ; P1_U5127
g2417 nand P1_U3363 P1_U3360 P1_U3361 ; P1_U5128
g2418 nand P1_U3365 P1_U3419 P1_U3364 ; P1_U5129
g2419 nand P1_U5710 P1_U5129 ; P1_U5130
g2420 nand P1_U5719 P1_U5128 ; P1_U5131
g2421 nand P1_U5131 P1_U5130 P1_U3877 ; P1_U5132
g2422 nand P1_U5132 P1_U3431 ; P1_U5133
g2423 not P1_U3433 ; P1_U5134
g2424 nand P1_U3498 P1_U5686 ; P1_U5135
g2425 nand P1_ADD_99_U73 P1_U5685 ; P1_U5136
g2426 nand P1_U4027 P1_U5127 ; P1_U5137
g2427 nand P1_R1165_U104 P1_U3027 ; P1_U5138
g2428 nand P1_U3084 P1_REG3_REG_15__SCAN_IN ; P1_U5139
g2429 nand P1_U3036 P1_U3056 ; P1_U5140
g2430 nand P1_U3034 P1_U3051 ; P1_U5141
g2431 nand P1_ADD_99_U62 P1_U3431 ; P1_U5142
g2432 nand P1_U5142 P1_U5140 P1_U5141 ; P1_U5143
g2433 nand P1_U3422 P1_U3431 ; P1_U5144
g2434 nand P1_U5134 P1_U5144 ; P1_U5145
g2435 nand P1_U4005 P1_U3422 ; P1_U5146
g2436 nand P1_U3418 P1_U5146 ; P1_U5147
g2437 nand P1_U3045 P1_U4009 ; P1_U5148
g2438 nand P1_U3044 P1_ADD_99_U62 ; P1_U5149
g2439 nand P1_U4027 P1_U5143 ; P1_U5150
g2440 nand P1_R1165_U13 P1_U3027 ; P1_U5151
g2441 nand P1_U3084 P1_REG3_REG_26__SCAN_IN ; P1_U5152
g2442 nand P1_U3036 P1_U3065 ; P1_U5153
g2443 nand P1_U3034 P1_U3068 ; P1_U5154
g2444 nand P1_ADD_99_U57 P1_U3431 ; P1_U5155
g2445 nand P1_U5154 P1_U5153 P1_U5155 ; P1_U5156
g2446 nand P1_U3471 P1_U5686 ; P1_U5157
g2447 nand P1_ADD_99_U57 P1_U5685 ; P1_U5158
g2448 nand P1_U4027 P1_U5156 ; P1_U5159
g2449 nand P1_R1165_U89 P1_U3027 ; P1_U5160
g2450 nand P1_U3084 P1_REG3_REG_6__SCAN_IN ; P1_U5161
g2451 nand P1_U3036 P1_U3067 ; P1_U5162
g2452 nand P1_U3034 P1_U3079 ; P1_U5163
g2453 nand P1_ADD_99_U70 P1_U3431 ; P1_U5164
g2454 nand P1_U5164 P1_U5162 P1_U5163 ; P1_U5165
g2455 nand P1_U3507 P1_U5686 ; P1_U5166
g2456 nand P1_ADD_99_U70 P1_U5685 ; P1_U5167
g2457 nand P1_U4027 P1_U5165 ; P1_U5168
g2458 nand P1_R1165_U102 P1_U3027 ; P1_U5169
g2459 nand P1_U3084 P1_REG3_REG_18__SCAN_IN ; P1_U5170
g2460 nand P1_U3036 P1_U3076 ; P1_U5171
g2461 nand P1_U3034 P1_U3062 ; P1_U5172
g2462 nand P1_U3431 P1_REG3_REG_2__SCAN_IN ; P1_U5173
g2463 nand P1_U5172 P1_U5171 P1_U5173 ; P1_U5174
g2464 nand P1_U3459 P1_U5686 ; P1_U5175
g2465 nand P1_U5685 P1_REG3_REG_2__SCAN_IN ; P1_U5176
g2466 nand P1_U4027 P1_U5174 ; P1_U5177
g2467 nand P1_R1165_U92 P1_U3027 ; P1_U5178
g2468 nand P1_U3084 P1_REG3_REG_2__SCAN_IN ; P1_U5179
g2469 nand P1_U3036 P1_U3060 ; P1_U5180
g2470 nand P1_U3034 P1_U3070 ; P1_U5181
g2471 nand P1_ADD_99_U77 P1_U3431 ; P1_U5182
g2472 nand P1_U5181 P1_U5180 P1_U5182 ; P1_U5183
g2473 nand P1_U3486 P1_U5686 ; P1_U5184
g2474 nand P1_ADD_99_U77 P1_U5685 ; P1_U5185
g2475 nand P1_U4027 P1_U5183 ; P1_U5186
g2476 nand P1_R1165_U107 P1_U3027 ; P1_U5187
g2477 nand P1_U3084 P1_REG3_REG_11__SCAN_IN ; P1_U5188
g2478 nand P1_U3036 P1_U3073 ; P1_U5189
g2479 nand P1_U3034 P1_U3064 ; P1_U5190
g2480 nand P1_ADD_99_U66 P1_U3431 ; P1_U5191
g2481 nand P1_U5191 P1_U5189 P1_U5190 ; P1_U5192
g2482 nand P1_U3045 P1_U4013 ; P1_U5193
g2483 nand P1_U3044 P1_ADD_99_U66 ; P1_U5194
g2484 nand P1_U4027 P1_U5192 ; P1_U5195
g2485 nand P1_R1165_U98 P1_U3027 ; P1_U5196
g2486 nand P1_U3084 P1_REG3_REG_22__SCAN_IN ; P1_U5197
g2487 nand P1_U3036 P1_U3070 ; P1_U5198
g2488 nand P1_U3034 P1_U3077 ; P1_U5199
g2489 nand P1_ADD_99_U75 P1_U3431 ; P1_U5200
g2490 nand P1_U5200 P1_U5198 P1_U5199 ; P1_U5201
g2491 nand P1_U3492 P1_U5686 ; P1_U5202
g2492 nand P1_ADD_99_U75 P1_U5685 ; P1_U5203
g2493 nand P1_U4027 P1_U5201 ; P1_U5204
g2494 nand P1_R1165_U10 P1_U3027 ; P1_U5205
g2495 nand P1_U3084 P1_REG3_REG_13__SCAN_IN ; P1_U5206
g2496 nand P1_U3036 P1_U3079 ; P1_U5207
g2497 nand P1_U3034 P1_U3073 ; P1_U5208
g2498 nand P1_ADD_99_U68 P1_U3431 ; P1_U5209
g2499 nand P1_U5209 P1_U5207 P1_U5208 ; P1_U5210
g2500 nand P1_U3045 P1_U4015 ; P1_U5211
g2501 nand P1_U3044 P1_ADD_99_U68 ; P1_U5212
g2502 nand P1_U4027 P1_U5210 ; P1_U5213
g2503 nand P1_R1165_U99 P1_U3027 ; P1_U5214
g2504 nand P1_U3084 P1_REG3_REG_20__SCAN_IN ; P1_U5215
g2505 nand P1_U3432 P1_U3430 ; P1_U5216
g2506 nand P1_U5216 P1_U3431 ; P1_U5217
g2507 nand P1_U4028 P1_U5217 ; P1_U5218
g2508 nand P1_U3883 P1_U3034 ; P1_U5219
g2509 nand P1_U3451 P1_U5686 ; P1_U5220
g2510 nand P1_U5218 P1_REG3_REG_0__SCAN_IN ; P1_U5221
g2511 nand P1_R1165_U86 P1_U3027 ; P1_U5222
g2512 nand P1_U3084 P1_REG3_REG_0__SCAN_IN ; P1_U5223
g2513 nand P1_U3036 P1_U3082 ; P1_U5224
g2514 nand P1_U3034 P1_U3060 ; P1_U5225
g2515 nand P1_ADD_99_U54 P1_U3431 ; P1_U5226
g2516 nand P1_U5225 P1_U5224 P1_U5226 ; P1_U5227
g2517 nand P1_U3480 P1_U5686 ; P1_U5228
g2518 nand P1_ADD_99_U54 P1_U5685 ; P1_U5229
g2519 nand P1_U4027 P1_U5227 ; P1_U5230
g2520 nand P1_R1165_U87 P1_U3027 ; P1_U5231
g2521 nand P1_U3084 P1_REG3_REG_9__SCAN_IN ; P1_U5232
g2522 nand P1_U3036 P1_U3062 ; P1_U5233
g2523 nand P1_U3034 P1_U3065 ; P1_U5234
g2524 nand P1_ADD_99_U59 P1_U3431 ; P1_U5235
g2525 nand P1_U5234 P1_U5233 P1_U5235 ; P1_U5236
g2526 nand P1_U3465 P1_U5686 ; P1_U5237
g2527 nand P1_ADD_99_U59 P1_U5685 ; P1_U5238
g2528 nand P1_U4027 P1_U5236 ; P1_U5239
g2529 nand P1_R1165_U91 P1_U3027 ; P1_U5240
g2530 nand P1_U3084 P1_REG3_REG_4__SCAN_IN ; P1_U5241
g2531 nand P1_U3036 P1_U3064 ; P1_U5242
g2532 nand P1_U3034 P1_U3056 ; P1_U5243
g2533 nand P1_ADD_99_U64 P1_U3431 ; P1_U5244
g2534 nand P1_U5244 P1_U5242 P1_U5243 ; P1_U5245
g2535 nand P1_U3045 P1_U4011 ; P1_U5246
g2536 nand P1_U3044 P1_ADD_99_U64 ; P1_U5247
g2537 nand P1_U4027 P1_U5245 ; P1_U5248
g2538 nand P1_R1165_U96 P1_U3027 ; P1_U5249
g2539 nand P1_U3084 P1_REG3_REG_24__SCAN_IN ; P1_U5250
g2540 nand P1_U3036 P1_U3071 ; P1_U5251
g2541 nand P1_U3034 P1_U3080 ; P1_U5252
g2542 nand P1_ADD_99_U71 P1_U3431 ; P1_U5253
g2543 nand P1_U5253 P1_U5251 P1_U5252 ; P1_U5254
g2544 nand P1_U3504 P1_U5686 ; P1_U5255
g2545 nand P1_ADD_99_U71 P1_U5685 ; P1_U5256
g2546 nand P1_U4027 P1_U5254 ; P1_U5257
g2547 nand P1_R1165_U11 P1_U3027 ; P1_U5258
g2548 nand P1_U3084 P1_REG3_REG_17__SCAN_IN ; P1_U5259
g2549 nand P1_U3036 P1_U3058 ; P1_U5260
g2550 nand P1_U3034 P1_U3069 ; P1_U5261
g2551 nand P1_ADD_99_U58 P1_U3431 ; P1_U5262
g2552 nand P1_U5261 P1_U5260 P1_U5262 ; P1_U5263
g2553 nand P1_U3468 P1_U5686 ; P1_U5264
g2554 nand P1_ADD_99_U58 P1_U5685 ; P1_U5265
g2555 nand P1_U4027 P1_U5263 ; P1_U5266
g2556 nand P1_R1165_U90 P1_U3027 ; P1_U5267
g2557 nand P1_U3084 P1_REG3_REG_5__SCAN_IN ; P1_U5268
g2558 nand P1_U3036 P1_U3072 ; P1_U5269
g2559 nand P1_U3034 P1_U3067 ; P1_U5270
g2560 nand P1_ADD_99_U72 P1_U3431 ; P1_U5271
g2561 nand P1_U5271 P1_U5269 P1_U5270 ; P1_U5272
g2562 nand P1_U3501 P1_U5686 ; P1_U5273
g2563 nand P1_ADD_99_U72 P1_U5685 ; P1_U5274
g2564 nand P1_U4027 P1_U5272 ; P1_U5275
g2565 nand P1_R1165_U103 P1_U3027 ; P1_U5276
g2566 nand P1_U3084 P1_REG3_REG_16__SCAN_IN ; P1_U5277
g2567 nand P1_U3036 P1_U3063 ; P1_U5278
g2568 nand P1_U3034 P1_U3055 ; P1_U5279
g2569 nand P1_ADD_99_U63 P1_U3431 ; P1_U5280
g2570 nand P1_U5280 P1_U5278 P1_U5279 ; P1_U5281
g2571 nand P1_U3045 P1_U4010 ; P1_U5282
g2572 nand P1_U3044 P1_ADD_99_U63 ; P1_U5283
g2573 nand P1_U4027 P1_U5281 ; P1_U5284
g2574 nand P1_R1165_U95 P1_U3027 ; P1_U5285
g2575 nand P1_U3084 P1_REG3_REG_25__SCAN_IN ; P1_U5286
g2576 nand P1_U3036 P1_U3061 ; P1_U5287
g2577 nand P1_U3034 P1_U3078 ; P1_U5288
g2578 nand P1_ADD_99_U76 P1_U3431 ; P1_U5289
g2579 nand P1_U5289 P1_U5287 P1_U5288 ; P1_U5290
g2580 nand P1_U3489 P1_U5686 ; P1_U5291
g2581 nand P1_ADD_99_U76 P1_U5685 ; P1_U5292
g2582 nand P1_U4027 P1_U5290 ; P1_U5293
g2583 nand P1_R1165_U106 P1_U3027 ; P1_U5294
g2584 nand P1_U3084 P1_REG3_REG_12__SCAN_IN ; P1_U5295
g2585 nand P1_U3036 P1_U3074 ; P1_U5296
g2586 nand P1_U3034 P1_U3059 ; P1_U5297
g2587 nand P1_ADD_99_U67 P1_U3431 ; P1_U5298
g2588 nand P1_U5298 P1_U5296 P1_U5297 ; P1_U5299
g2589 nand P1_U3045 P1_U4014 ; P1_U5300
g2590 nand P1_U3044 P1_ADD_99_U67 ; P1_U5301
g2591 nand P1_U4027 P1_U5299 ; P1_U5302
g2592 nand P1_R1165_U12 P1_U3027 ; P1_U5303
g2593 nand P1_U3084 P1_REG3_REG_21__SCAN_IN ; P1_U5304
g2594 nand P1_U3036 P1_U3075 ; P1_U5305
g2595 nand P1_U3034 P1_U3066 ; P1_U5306
g2596 nand P1_U3431 P1_REG3_REG_1__SCAN_IN ; P1_U5307
g2597 nand P1_U5306 P1_U5305 P1_U5307 ; P1_U5308
g2598 nand P1_U3456 P1_U5686 ; P1_U5309
g2599 nand P1_U5685 P1_REG3_REG_1__SCAN_IN ; P1_U5310
g2600 nand P1_U4027 P1_U5308 ; P1_U5311
g2601 nand P1_R1165_U100 P1_U3027 ; P1_U5312
g2602 nand P1_U3084 P1_REG3_REG_1__SCAN_IN ; P1_U5313
g2603 nand P1_U3036 P1_U3068 ; P1_U5314
g2604 nand P1_U3034 P1_U3081 ; P1_U5315
g2605 nand P1_ADD_99_U55 P1_U3431 ; P1_U5316
g2606 nand P1_U5315 P1_U5314 P1_U5316 ; P1_U5317
g2607 nand P1_U3477 P1_U5686 ; P1_U5318
g2608 nand P1_ADD_99_U55 P1_U5685 ; P1_U5319
g2609 nand P1_U4027 P1_U5317 ; P1_U5320
g2610 nand P1_R1165_U88 P1_U3027 ; P1_U5321
g2611 nand P1_U3084 P1_REG3_REG_8__SCAN_IN ; P1_U5322
g2612 nand P1_U3036 P1_U3051 ; P1_U5323
g2613 nand P1_U3034 P1_U3053 ; P1_U5324
g2614 nand P1_ADD_99_U60 P1_U3431 ; P1_U5325
g2615 nand P1_U5324 P1_U5323 P1_U5325 ; P1_U5326
g2616 nand P1_U3045 P1_U4007 ; P1_U5327
g2617 nand P1_U3044 P1_ADD_99_U60 ; P1_U5328
g2618 nand P1_U4027 P1_U5326 ; P1_U5329
g2619 nand P1_R1165_U93 P1_U3027 ; P1_U5330
g2620 nand P1_U3084 P1_REG3_REG_28__SCAN_IN ; P1_U5331
g2621 nand P1_U3036 P1_U3080 ; P1_U5332
g2622 nand P1_U3034 P1_U3074 ; P1_U5333
g2623 nand P1_ADD_99_U69 P1_U3431 ; P1_U5334
g2624 nand P1_U5334 P1_U5332 P1_U5333 ; P1_U5335
g2625 nand P1_U3509 P1_U5686 ; P1_U5336
g2626 nand P1_ADD_99_U69 P1_U5685 ; P1_U5337
g2627 nand P1_U4027 P1_U5335 ; P1_U5338
g2628 nand P1_R1165_U101 P1_U3027 ; P1_U5339
g2629 nand P1_U3084 P1_REG3_REG_19__SCAN_IN ; P1_U5340
g2630 nand P1_U3036 P1_U3066 ; P1_U5341
g2631 nand P1_U3034 P1_U3058 ; P1_U5342
g2632 nand P1_ADD_99_U4 P1_U3431 ; P1_U5343
g2633 nand P1_U5342 P1_U5341 P1_U5343 ; P1_U5344
g2634 nand P1_U3462 P1_U5686 ; P1_U5345
g2635 nand P1_ADD_99_U4 P1_U5685 ; P1_U5346
g2636 nand P1_U4027 P1_U5344 ; P1_U5347
g2637 nand P1_R1165_U14 P1_U3027 ; P1_U5348
g2638 nand P1_U3084 P1_REG3_REG_3__SCAN_IN ; P1_U5349
g2639 nand P1_U3036 P1_U3081 ; P1_U5350
g2640 nand P1_U3034 P1_U3061 ; P1_U5351
g2641 nand P1_ADD_99_U78 P1_U3431 ; P1_U5352
g2642 nand P1_U5351 P1_U5350 P1_U5352 ; P1_U5353
g2643 nand P1_U3483 P1_U5686 ; P1_U5354
g2644 nand P1_ADD_99_U78 P1_U5685 ; P1_U5355
g2645 nand P1_U4027 P1_U5353 ; P1_U5356
g2646 nand P1_R1165_U108 P1_U3027 ; P1_U5357
g2647 nand P1_U3084 P1_REG3_REG_10__SCAN_IN ; P1_U5358
g2648 nand P1_U3036 P1_U3059 ; P1_U5359
g2649 nand P1_U3034 P1_U3063 ; P1_U5360
g2650 nand P1_ADD_99_U65 P1_U3431 ; P1_U5361
g2651 nand P1_U5361 P1_U5359 P1_U5360 ; P1_U5362
g2652 nand P1_U3045 P1_U4012 ; P1_U5363
g2653 nand P1_U3044 P1_ADD_99_U65 ; P1_U5364
g2654 nand P1_U4027 P1_U5362 ; P1_U5365
g2655 nand P1_R1165_U97 P1_U3027 ; P1_U5366
g2656 nand P1_U3084 P1_REG3_REG_23__SCAN_IN ; P1_U5367
g2657 nand P1_U3036 P1_U3078 ; P1_U5368
g2658 nand P1_U3034 P1_U3072 ; P1_U5369
g2659 nand P1_ADD_99_U74 P1_U3431 ; P1_U5370
g2660 nand P1_U5370 P1_U5368 P1_U5369 ; P1_U5371
g2661 nand P1_U3495 P1_U5686 ; P1_U5372
g2662 nand P1_ADD_99_U74 P1_U5685 ; P1_U5373
g2663 nand P1_U4027 P1_U5371 ; P1_U5374
g2664 nand P1_R1165_U105 P1_U3027 ; P1_U5375
g2665 nand P1_U3084 P1_REG3_REG_14__SCAN_IN ; P1_U5376
g2666 nand P1_U3036 P1_U3055 ; P1_U5377
g2667 nand P1_U3034 P1_U3052 ; P1_U5378
g2668 nand P1_ADD_99_U61 P1_U3431 ; P1_U5379
g2669 nand P1_U5379 P1_U5377 P1_U5378 ; P1_U5380
g2670 nand P1_U3045 P1_U4008 ; P1_U5381
g2671 nand P1_U3044 P1_ADD_99_U61 ; P1_U5382
g2672 nand P1_U4027 P1_U5380 ; P1_U5383
g2673 nand P1_R1165_U94 P1_U3027 ; P1_U5384
g2674 nand P1_U3084 P1_REG3_REG_27__SCAN_IN ; P1_U5385
g2675 nand P1_U3036 P1_U3069 ; P1_U5386
g2676 nand P1_U3034 P1_U3082 ; P1_U5387
g2677 nand P1_ADD_99_U56 P1_U3431 ; P1_U5388
g2678 nand P1_U5387 P1_U5386 P1_U5388 ; P1_U5389
g2679 nand P1_U3474 P1_U5686 ; P1_U5390
g2680 nand P1_ADD_99_U56 P1_U5685 ; P1_U5391
g2681 nand P1_U4027 P1_U5389 ; P1_U5392
g2682 nand P1_R1165_U15 P1_U3027 ; P1_U5393
g2683 nand P1_U3084 P1_REG3_REG_7__SCAN_IN ; P1_U5394
g2684 nand P1_U3450 P1_U3374 ; P1_U5395
g2685 nand P1_U3447 P1_U5395 ; P1_U5396
g2686 nand P1_U5734 P1_U3447 P1_R1165_U86 ; P1_U5397
g2687 nand P1_U3448 P1_U3442 ; P1_U5398
g2688 nand P1_U3893 P1_U4003 ; P1_U5399
g2689 nand P1_U3369 P1_U3419 ; P1_U5400
g2690 nand P1_U3367 P1_U3362 P1_U3364 ; P1_U5401
g2691 nand P1_U4033 P1_U3421 ; P1_U5402
g2692 nand P1_U5401 P1_U3421 ; P1_U5403
g2693 not P1_U3435 ; P1_U5404
g2694 nand P1_U5404 P1_U4003 ; P1_U5405
g2695 nand P1_U3480 P1_U5405 ; P1_U5406
g2696 nand P1_U3021 P1_U3081 ; P1_U5407
g2697 nand P1_U3477 P1_U5405 ; P1_U5408
g2698 nand P1_U3021 P1_U3082 ; P1_U5409
g2699 nand P1_U3474 P1_U5405 ; P1_U5410
g2700 nand P1_U3021 P1_U3068 ; P1_U5411
g2701 nand P1_U3471 P1_U5405 ; P1_U5412
g2702 nand P1_U3021 P1_U3069 ; P1_U5413
g2703 nand P1_U3468 P1_U5405 ; P1_U5414
g2704 nand P1_U3021 P1_U3065 ; P1_U5415
g2705 nand P1_U3465 P1_U5405 ; P1_U5416
g2706 nand P1_U3021 P1_U3058 ; P1_U5417
g2707 nand P1_U3462 P1_U5405 ; P1_U5418
g2708 nand P1_U3021 P1_U3062 ; P1_U5419
g2709 nand P1_U4007 P1_U5405 ; P1_U5420
g2710 nand P1_U3021 P1_U3052 ; P1_U5421
g2711 nand P1_U4008 P1_U5405 ; P1_U5422
g2712 nand P1_U3021 P1_U3051 ; P1_U5423
g2713 nand P1_U4009 P1_U5405 ; P1_U5424
g2714 nand P1_U3021 P1_U3055 ; P1_U5425
g2715 nand P1_U4010 P1_U5405 ; P1_U5426
g2716 nand P1_U3021 P1_U3056 ; P1_U5427
g2717 nand P1_U4011 P1_U5405 ; P1_U5428
g2718 nand P1_U3021 P1_U3063 ; P1_U5429
g2719 nand P1_U4012 P1_U5405 ; P1_U5430
g2720 nand P1_U3021 P1_U3064 ; P1_U5431
g2721 nand P1_U4013 P1_U5405 ; P1_U5432
g2722 nand P1_U3021 P1_U3059 ; P1_U5433
g2723 nand P1_U4014 P1_U5405 ; P1_U5434
g2724 nand P1_U3021 P1_U3073 ; P1_U5435
g2725 nand P1_U4015 P1_U5405 ; P1_U5436
g2726 nand P1_U3021 P1_U3074 ; P1_U5437
g2727 nand P1_U3459 P1_U5405 ; P1_U5438
g2728 nand P1_U3021 P1_U3066 ; P1_U5439
g2729 nand P1_U3509 P1_U5405 ; P1_U5440
g2730 nand P1_U3021 P1_U3079 ; P1_U5441
g2731 nand P1_U3507 P1_U5405 ; P1_U5442
g2732 nand P1_U3021 P1_U3080 ; P1_U5443
g2733 nand P1_U3504 P1_U5405 ; P1_U5444
g2734 nand P1_U3021 P1_U3067 ; P1_U5445
g2735 nand P1_U3501 P1_U5405 ; P1_U5446
g2736 nand P1_U3021 P1_U3071 ; P1_U5447
g2737 nand P1_U3498 P1_U5405 ; P1_U5448
g2738 nand P1_U3021 P1_U3072 ; P1_U5449
g2739 nand P1_U3495 P1_U5405 ; P1_U5450
g2740 nand P1_U3021 P1_U3077 ; P1_U5451
g2741 nand P1_U3492 P1_U5405 ; P1_U5452
g2742 nand P1_U3021 P1_U3078 ; P1_U5453
g2743 nand P1_U3489 P1_U5405 ; P1_U5454
g2744 nand P1_U3021 P1_U3070 ; P1_U5455
g2745 nand P1_U3486 P1_U5405 ; P1_U5456
g2746 nand P1_U3021 P1_U3061 ; P1_U5457
g2747 nand P1_U3483 P1_U5405 ; P1_U5458
g2748 nand P1_U3021 P1_U3060 ; P1_U5459
g2749 nand P1_U3456 P1_U5405 ; P1_U5460
g2750 nand P1_U3021 P1_U3076 ; P1_U5461
g2751 nand P1_U3451 P1_U5405 ; P1_U5462
g2752 nand P1_U3021 P1_U3075 ; P1_U5463
g2753 nand P1_U4135 P1_REG1_REG_0__SCAN_IN ; P1_U5464
g2754 nand P1_U3021 P1_U3480 ; P1_U5465
g2755 nand P1_U3435 P1_U3081 ; P1_U5466
g2756 nand P1_U3021 P1_U3477 ; P1_U5467
g2757 nand P1_U3435 P1_U3082 ; P1_U5468
g2758 nand P1_U3021 P1_U3474 ; P1_U5469
g2759 nand P1_U3435 P1_U3068 ; P1_U5470
g2760 nand P1_U3021 P1_U3471 ; P1_U5471
g2761 nand P1_U3435 P1_U3069 ; P1_U5472
g2762 nand P1_U3021 P1_U3468 ; P1_U5473
g2763 nand P1_U3435 P1_U3065 ; P1_U5474
g2764 nand P1_U3021 P1_U3465 ; P1_U5475
g2765 nand P1_U3435 P1_U3058 ; P1_U5476
g2766 nand P1_U3021 P1_U3462 ; P1_U5477
g2767 nand P1_U3435 P1_U3062 ; P1_U5478
g2768 nand P1_U3021 P1_U4007 ; P1_U5479
g2769 nand P1_U3435 P1_U3052 ; P1_U5480
g2770 nand P1_U3021 P1_U4008 ; P1_U5481
g2771 nand P1_U3435 P1_U3051 ; P1_U5482
g2772 nand P1_U3021 P1_U4009 ; P1_U5483
g2773 nand P1_U3435 P1_U3055 ; P1_U5484
g2774 nand P1_U3021 P1_U4010 ; P1_U5485
g2775 nand P1_U3435 P1_U3056 ; P1_U5486
g2776 nand P1_U3021 P1_U4011 ; P1_U5487
g2777 nand P1_U3435 P1_U3063 ; P1_U5488
g2778 nand P1_U3021 P1_U4012 ; P1_U5489
g2779 nand P1_U3435 P1_U3064 ; P1_U5490
g2780 nand P1_U3021 P1_U4013 ; P1_U5491
g2781 nand P1_U3435 P1_U3059 ; P1_U5492
g2782 nand P1_U3021 P1_U4014 ; P1_U5493
g2783 nand P1_U3435 P1_U3073 ; P1_U5494
g2784 nand P1_U3021 P1_U4015 ; P1_U5495
g2785 nand P1_U3435 P1_U3074 ; P1_U5496
g2786 nand P1_U3021 P1_U3459 ; P1_U5497
g2787 nand P1_U3435 P1_U3066 ; P1_U5498
g2788 nand P1_U3021 P1_U3509 ; P1_U5499
g2789 nand P1_U3435 P1_U3079 ; P1_U5500
g2790 nand P1_U3021 P1_U3507 ; P1_U5501
g2791 nand P1_U3435 P1_U3080 ; P1_U5502
g2792 nand P1_U3021 P1_U3504 ; P1_U5503
g2793 nand P1_U3435 P1_U3067 ; P1_U5504
g2794 nand P1_U3021 P1_U3501 ; P1_U5505
g2795 nand P1_U3435 P1_U3071 ; P1_U5506
g2796 nand P1_U3021 P1_U3498 ; P1_U5507
g2797 nand P1_U3435 P1_U3072 ; P1_U5508
g2798 nand P1_U3021 P1_U3495 ; P1_U5509
g2799 nand P1_U3435 P1_U3077 ; P1_U5510
g2800 nand P1_U3021 P1_U3492 ; P1_U5511
g2801 nand P1_U3435 P1_U3078 ; P1_U5512
g2802 nand P1_U3021 P1_U3489 ; P1_U5513
g2803 nand P1_U3435 P1_U3070 ; P1_U5514
g2804 nand P1_U3021 P1_U3486 ; P1_U5515
g2805 nand P1_U3435 P1_U3061 ; P1_U5516
g2806 nand P1_U3021 P1_U3483 ; P1_U5517
g2807 nand P1_U3435 P1_U3060 ; P1_U5518
g2808 nand P1_U3021 P1_U3456 ; P1_U5519
g2809 nand P1_U3435 P1_U3076 ; P1_U5520
g2810 nand P1_U3021 P1_U3451 ; P1_U5521
g2811 nand P1_U3435 P1_U3075 ; P1_U5522
g2812 nand P1_U4135 P1_U3449 ; P1_U5523
g2813 nand P1_U3428 P1_U3426 ; P1_U5524
g2814 nand P1_U3986 P1_U3480 ; P1_U5525
g2815 nand P1_U3587 P1_U5524 ; P1_U5526
g2816 nand P1_U3986 P1_U3477 ; P1_U5527
g2817 nand P1_U3588 P1_U5524 ; P1_U5528
g2818 nand P1_U3986 P1_U3474 ; P1_U5529
g2819 nand P1_U3589 P1_U5524 ; P1_U5530
g2820 nand P1_U3986 P1_U3471 ; P1_U5531
g2821 nand P1_U3590 P1_U5524 ; P1_U5532
g2822 nand P1_U3986 P1_U3468 ; P1_U5533
g2823 nand P1_U3591 P1_U5524 ; P1_U5534
g2824 nand P1_U3986 P1_U3465 ; P1_U5535
g2825 nand P1_U3592 P1_U5524 ; P1_U5536
g2826 nand P1_U3594 P1_U5524 ; P1_U5537
g2827 nand P1_U4016 P1_U3986 ; P1_U5538
g2828 nand P1_U3595 P1_U5524 ; P1_U5539
g2829 nand P1_U4017 P1_U3986 ; P1_U5540
g2830 nand P1_U3986 P1_U3462 ; P1_U5541
g2831 nand P1_U3593 P1_U5524 ; P1_U5542
g2832 nand P1_U3597 P1_U5524 ; P1_U5543
g2833 nand P1_U4018 P1_U3986 ; P1_U5544
g2834 nand P1_U3598 P1_U5524 ; P1_U5545
g2835 nand P1_U4007 P1_U3986 ; P1_U5546
g2836 nand P1_U3599 P1_U5524 ; P1_U5547
g2837 nand P1_U4008 P1_U3986 ; P1_U5548
g2838 nand P1_U3600 P1_U5524 ; P1_U5549
g2839 nand P1_U4009 P1_U3986 ; P1_U5550
g2840 nand P1_U3601 P1_U5524 ; P1_U5551
g2841 nand P1_U4010 P1_U3986 ; P1_U5552
g2842 nand P1_U3602 P1_U5524 ; P1_U5553
g2843 nand P1_U4011 P1_U3986 ; P1_U5554
g2844 nand P1_U3603 P1_U5524 ; P1_U5555
g2845 nand P1_U4012 P1_U3986 ; P1_U5556
g2846 nand P1_U3604 P1_U5524 ; P1_U5557
g2847 nand P1_U4013 P1_U3986 ; P1_U5558
g2848 nand P1_U3605 P1_U5524 ; P1_U5559
g2849 nand P1_U4014 P1_U3986 ; P1_U5560
g2850 nand P1_U3606 P1_U5524 ; P1_U5561
g2851 nand P1_U4015 P1_U3986 ; P1_U5562
g2852 nand P1_U3986 P1_U3459 ; P1_U5563
g2853 nand P1_U3596 P1_U5524 ; P1_U5564
g2854 nand P1_U3986 P1_U3509 ; P1_U5565
g2855 nand P1_U3608 P1_U5524 ; P1_U5566
g2856 nand P1_U3986 P1_U3507 ; P1_U5567
g2857 nand P1_U3609 P1_U5524 ; P1_U5568
g2858 nand P1_U3986 P1_U3504 ; P1_U5569
g2859 nand P1_U3610 P1_U5524 ; P1_U5570
g2860 nand P1_U3986 P1_U3501 ; P1_U5571
g2861 nand P1_U3611 P1_U5524 ; P1_U5572
g2862 nand P1_U3986 P1_U3498 ; P1_U5573
g2863 nand P1_U3612 P1_U5524 ; P1_U5574
g2864 nand P1_U3986 P1_U3495 ; P1_U5575
g2865 nand P1_U3613 P1_U5524 ; P1_U5576
g2866 nand P1_U3986 P1_U3492 ; P1_U5577
g2867 nand P1_U3614 P1_U5524 ; P1_U5578
g2868 nand P1_U3986 P1_U3489 ; P1_U5579
g2869 nand P1_U3615 P1_U5524 ; P1_U5580
g2870 nand P1_U3986 P1_U3486 ; P1_U5581
g2871 nand P1_U3616 P1_U5524 ; P1_U5582
g2872 nand P1_U3986 P1_U3483 ; P1_U5583
g2873 nand P1_U3617 P1_U5524 ; P1_U5584
g2874 nand P1_U3986 P1_U3456 ; P1_U5585
g2875 nand P1_U3607 P1_U5524 ; P1_U5586
g2876 nand P1_U3986 P1_U3451 ; P1_U5587
g2877 nand P1_U3618 P1_U5524 ; P1_U5588
g2878 nand P1_U3480 P1_U5524 ; P1_U5589
g2879 nand P1_U3986 P1_U3587 ; P1_U5590
g2880 nand P1_U5703 P1_U3082 ; P1_U5591
g2881 nand P1_U3477 P1_U5524 ; P1_U5592
g2882 nand P1_U3986 P1_U3588 ; P1_U5593
g2883 nand P1_U5703 P1_U3068 ; P1_U5594
g2884 nand P1_U3474 P1_U5524 ; P1_U5595
g2885 nand P1_U3986 P1_U3589 ; P1_U5596
g2886 nand P1_U5703 P1_U3069 ; P1_U5597
g2887 nand P1_U3471 P1_U5524 ; P1_U5598
g2888 nand P1_U3986 P1_U3590 ; P1_U5599
g2889 nand P1_U5703 P1_U3065 ; P1_U5600
g2890 nand P1_U3468 P1_U5524 ; P1_U5601
g2891 nand P1_U3986 P1_U3591 ; P1_U5602
g2892 nand P1_U5703 P1_U3058 ; P1_U5603
g2893 nand P1_U3465 P1_U5524 ; P1_U5604
g2894 nand P1_U3986 P1_U3592 ; P1_U5605
g2895 nand P1_U5703 P1_U3062 ; P1_U5606
g2896 nand P1_U4016 P1_U5524 ; P1_U5607
g2897 nand P1_U3986 P1_U3594 ; P1_U5608
g2898 nand P1_U4017 P1_U5524 ; P1_U5609
g2899 nand P1_U3986 P1_U3595 ; P1_U5610
g2900 nand P1_U3462 P1_U5524 ; P1_U5611
g2901 nand P1_U3986 P1_U3593 ; P1_U5612
g2902 nand P1_U5703 P1_U3066 ; P1_U5613
g2903 nand P1_U4018 P1_U5524 ; P1_U5614
g2904 nand P1_U3986 P1_U3597 ; P1_U5615
g2905 nand P1_U5703 P1_U3052 ; P1_U5616
g2906 nand P1_U4007 P1_U5524 ; P1_U5617
g2907 nand P1_U3986 P1_U3598 ; P1_U5618
g2908 nand P1_U5703 P1_U3051 ; P1_U5619
g2909 nand P1_U4008 P1_U5524 ; P1_U5620
g2910 nand P1_U3986 P1_U3599 ; P1_U5621
g2911 nand P1_U5703 P1_U3055 ; P1_U5622
g2912 nand P1_U4009 P1_U5524 ; P1_U5623
g2913 nand P1_U3986 P1_U3600 ; P1_U5624
g2914 nand P1_U5703 P1_U3056 ; P1_U5625
g2915 nand P1_U4010 P1_U5524 ; P1_U5626
g2916 nand P1_U3986 P1_U3601 ; P1_U5627
g2917 nand P1_U5703 P1_U3063 ; P1_U5628
g2918 nand P1_U4011 P1_U5524 ; P1_U5629
g2919 nand P1_U3986 P1_U3602 ; P1_U5630
g2920 nand P1_U5703 P1_U3064 ; P1_U5631
g2921 nand P1_U4012 P1_U5524 ; P1_U5632
g2922 nand P1_U3986 P1_U3603 ; P1_U5633
g2923 nand P1_U5703 P1_U3059 ; P1_U5634
g2924 nand P1_U4013 P1_U5524 ; P1_U5635
g2925 nand P1_U3986 P1_U3604 ; P1_U5636
g2926 nand P1_U5703 P1_U3073 ; P1_U5637
g2927 nand P1_U4014 P1_U5524 ; P1_U5638
g2928 nand P1_U3986 P1_U3605 ; P1_U5639
g2929 nand P1_U5703 P1_U3074 ; P1_U5640
g2930 nand P1_U4015 P1_U5524 ; P1_U5641
g2931 nand P1_U3986 P1_U3606 ; P1_U5642
g2932 nand P1_U5703 P1_U3079 ; P1_U5643
g2933 nand P1_U3459 P1_U5524 ; P1_U5644
g2934 nand P1_U3986 P1_U3596 ; P1_U5645
g2935 nand P1_U5703 P1_U3076 ; P1_U5646
g2936 nand P1_U3509 P1_U5524 ; P1_U5647
g2937 nand P1_U3986 P1_U3608 ; P1_U5648
g2938 nand P1_U5703 P1_U3080 ; P1_U5649
g2939 nand P1_U3507 P1_U5524 ; P1_U5650
g2940 nand P1_U3986 P1_U3609 ; P1_U5651
g2941 nand P1_U5703 P1_U3067 ; P1_U5652
g2942 nand P1_U3504 P1_U5524 ; P1_U5653
g2943 nand P1_U3986 P1_U3610 ; P1_U5654
g2944 nand P1_U5703 P1_U3071 ; P1_U5655
g2945 nand P1_U3501 P1_U5524 ; P1_U5656
g2946 nand P1_U3986 P1_U3611 ; P1_U5657
g2947 nand P1_U5703 P1_U3072 ; P1_U5658
g2948 nand P1_U3498 P1_U5524 ; P1_U5659
g2949 nand P1_U3986 P1_U3612 ; P1_U5660
g2950 nand P1_U5703 P1_U3077 ; P1_U5661
g2951 nand P1_U3495 P1_U5524 ; P1_U5662
g2952 nand P1_U3986 P1_U3613 ; P1_U5663
g2953 nand P1_U5703 P1_U3078 ; P1_U5664
g2954 nand P1_U3492 P1_U5524 ; P1_U5665
g2955 nand P1_U3986 P1_U3614 ; P1_U5666
g2956 nand P1_U5703 P1_U3070 ; P1_U5667
g2957 nand P1_U3489 P1_U5524 ; P1_U5668
g2958 nand P1_U3986 P1_U3615 ; P1_U5669
g2959 nand P1_U5703 P1_U3061 ; P1_U5670
g2960 nand P1_U3486 P1_U5524 ; P1_U5671
g2961 nand P1_U3986 P1_U3616 ; P1_U5672
g2962 nand P1_U5703 P1_U3060 ; P1_U5673
g2963 nand P1_U3483 P1_U5524 ; P1_U5674
g2964 nand P1_U3986 P1_U3617 ; P1_U5675
g2965 nand P1_U5703 P1_U3081 ; P1_U5676
g2966 nand P1_U3456 P1_U5524 ; P1_U5677
g2967 nand P1_U3986 P1_U3607 ; P1_U5678
g2968 nand P1_U5703 P1_U3075 ; P1_U5679
g2969 nand P1_U3451 P1_U5524 ; P1_U5680
g2970 nand P1_U3986 P1_U3618 ; P1_U5681
g2971 nand P1_U5123 P1_U3084 ; P1_U5682
g2972 nand P1_U4030 P1_U3431 ; P1_U5683
g2973 nand P1_U4005 P1_U4030 ; P1_U5684
g2974 nand P1_U5683 P1_U4028 ; P1_U5685
g2975 nand P1_U5684 P1_U4029 ; P1_U5686
g2976 nand P1_U3439 P1_U3048 P1_U3429 ; P1_U5687
g2977 nand P1_U5692 P1_U5698 ; P1_U5688
g2978 nand P1_U4020 P1_U3442 P1_U3987 P1_LT_201_U14 ; P1_U5689
g2979 nand P1_U3944 P1_IR_REG_24__SCAN_IN ; P1_U5690
g2980 nand P1_SUB_88_U17 P1_IR_REG_31__SCAN_IN ; P1_U5691
g2981 not P1_U3436 ; P1_U5692
g2982 nand P1_U3944 P1_IR_REG_25__SCAN_IN ; P1_U5693
g2983 nand P1_SUB_88_U170 P1_IR_REG_31__SCAN_IN ; P1_U5694
g2984 not P1_U3437 ; P1_U5695
g2985 nand P1_U3944 P1_IR_REG_26__SCAN_IN ; P1_U5696
g2986 nand P1_SUB_88_U18 P1_IR_REG_31__SCAN_IN ; P1_U5697
g2987 not P1_U3438 ; P1_U5698
g2988 nand P1_U3050 P1_U3358 ; P1_U5699
g2989 nand P1_U4036 P1_U5692 P1_B_REG_SCAN_IN ; P1_U5700
g2990 nand P1_U3944 P1_IR_REG_23__SCAN_IN ; P1_U5701
g2991 nand P1_SUB_88_U16 P1_IR_REG_31__SCAN_IN ; P1_U5702
g2992 not P1_U3439 ; P1_U5703
g2993 nand P1_U3945 P1_D_REG_0__SCAN_IN ; P1_U5704
g2994 nand P1_U4025 P1_U4136 ; P1_U5705
g2995 nand P1_U3945 P1_D_REG_1__SCAN_IN ; P1_U5706
g2996 nand P1_U4025 P1_U4137 ; P1_U5707
g2997 nand P1_U3944 P1_IR_REG_22__SCAN_IN ; P1_U5708
g2998 nand P1_SUB_88_U15 P1_IR_REG_31__SCAN_IN ; P1_U5709
g2999 not P1_U3444 ; P1_U5710
g3000 nand P1_U3944 P1_IR_REG_19__SCAN_IN ; P1_U5711
g3001 nand P1_SUB_88_U13 P1_IR_REG_31__SCAN_IN ; P1_U5712
g3002 not P1_U3443 ; P1_U5713
g3003 nand P1_U3944 P1_IR_REG_20__SCAN_IN ; P1_U5714
g3004 nand P1_SUB_88_U14 P1_IR_REG_31__SCAN_IN ; P1_U5715
g3005 not P1_U3442 ; P1_U5716
g3006 nand P1_U3944 P1_IR_REG_21__SCAN_IN ; P1_U5717
g3007 nand P1_SUB_88_U173 P1_IR_REG_31__SCAN_IN ; P1_U5718
g3008 not P1_U3448 ; P1_U5719
g3009 nand P1_U3944 P1_IR_REG_30__SCAN_IN ; P1_U5720
g3010 nand P1_SUB_88_U165 P1_IR_REG_31__SCAN_IN ; P1_U5721
g3011 not P1_U3445 ; P1_U5722
g3012 nand P1_U3944 P1_IR_REG_29__SCAN_IN ; P1_U5723
g3013 nand P1_SUB_88_U20 P1_IR_REG_31__SCAN_IN ; P1_U5724
g3014 not P1_U3446 ; P1_U5725
g3015 nand P1_U3944 P1_IR_REG_28__SCAN_IN ; P1_U5726
g3016 nand P1_SUB_88_U19 P1_IR_REG_31__SCAN_IN ; P1_U5727
g3017 not P1_U3447 ; P1_U5728
g3018 nand P1_U3944 P1_IR_REG_0__SCAN_IN ; P1_U5729
g3019 nand P1_IR_REG_0__SCAN_IN P1_IR_REG_31__SCAN_IN ; P1_U5730
g3020 not P1_U3449 ; P1_U5731
g3021 nand P1_U3944 P1_IR_REG_27__SCAN_IN ; P1_U5732
g3022 nand P1_SUB_88_U42 P1_IR_REG_31__SCAN_IN ; P1_U5733
g3023 not P1_U3450 ; P1_U5734
g3024 nand U88 P1_U3946 ; P1_U5735
g3025 nand P1_U4004 P1_U3449 ; P1_U5736
g3026 not P1_U3451 ; P1_U5737
g3027 nand P1_U3444 P1_U5719 ; P1_U5738
g3028 nand P1_U5710 P1_U4168 ; P1_U5739
g3029 nand P1_U4134 P1_D_REG_1__SCAN_IN ; P1_U5740
g3030 nand P1_U4137 P1_U3359 ; P1_U5741
g3031 not P1_U3453 ; P1_U5742
g3032 nand P1_U5688 P1_U3359 ; P1_U5743
g3033 nand P1_U4134 P1_D_REG_0__SCAN_IN ; P1_U5744
g3034 not P1_U3452 ; P1_U5745
g3035 nand P1_U3947 P1_REG0_REG_0__SCAN_IN ; P1_U5746
g3036 nand P1_U4024 P1_U4188 ; P1_U5747
g3037 nand P1_U3944 P1_IR_REG_1__SCAN_IN ; P1_U5748
g3038 nand P1_SUB_88_U40 P1_IR_REG_31__SCAN_IN ; P1_U5749
g3039 nand U77 P1_U3946 ; P1_U5750
g3040 nand P1_U3455 P1_U4004 ; P1_U5751
g3041 not P1_U3456 ; P1_U5752
g3042 nand P1_U3947 P1_REG0_REG_1__SCAN_IN ; P1_U5753
g3043 nand P1_U4024 P1_U4212 ; P1_U5754
g3044 nand P1_U3944 P1_IR_REG_2__SCAN_IN ; P1_U5755
g3045 nand P1_SUB_88_U21 P1_IR_REG_31__SCAN_IN ; P1_U5756
g3046 nand U66 P1_U3946 ; P1_U5757
g3047 nand P1_U3458 P1_U4004 ; P1_U5758
g3048 not P1_U3459 ; P1_U5759
g3049 nand P1_U3947 P1_REG0_REG_2__SCAN_IN ; P1_U5760
g3050 nand P1_U4024 P1_U4231 ; P1_U5761
g3051 nand P1_U3944 P1_IR_REG_3__SCAN_IN ; P1_U5762
g3052 nand P1_SUB_88_U22 P1_IR_REG_31__SCAN_IN ; P1_U5763
g3053 nand U63 P1_U3946 ; P1_U5764
g3054 nand P1_U3461 P1_U4004 ; P1_U5765
g3055 not P1_U3462 ; P1_U5766
g3056 nand P1_U3947 P1_REG0_REG_3__SCAN_IN ; P1_U5767
g3057 nand P1_U4024 P1_U4250 ; P1_U5768
g3058 nand P1_U3944 P1_IR_REG_4__SCAN_IN ; P1_U5769
g3059 nand P1_SUB_88_U23 P1_IR_REG_31__SCAN_IN ; P1_U5770
g3060 nand U62 P1_U3946 ; P1_U5771
g3061 nand P1_U3464 P1_U4004 ; P1_U5772
g3062 not P1_U3465 ; P1_U5773
g3063 nand P1_U3947 P1_REG0_REG_4__SCAN_IN ; P1_U5774
g3064 nand P1_U4024 P1_U4269 ; P1_U5775
g3065 nand P1_U3944 P1_IR_REG_5__SCAN_IN ; P1_U5776
g3066 nand P1_SUB_88_U162 P1_IR_REG_31__SCAN_IN ; P1_U5777
g3067 nand U61 P1_U3946 ; P1_U5778
g3068 nand P1_U3467 P1_U4004 ; P1_U5779
g3069 not P1_U3468 ; P1_U5780
g3070 nand P1_U3947 P1_REG0_REG_5__SCAN_IN ; P1_U5781
g3071 nand P1_U4024 P1_U4288 ; P1_U5782
g3072 nand P1_U3944 P1_IR_REG_6__SCAN_IN ; P1_U5783
g3073 nand P1_SUB_88_U24 P1_IR_REG_31__SCAN_IN ; P1_U5784
g3074 nand U60 P1_U3946 ; P1_U5785
g3075 nand P1_U3470 P1_U4004 ; P1_U5786
g3076 not P1_U3471 ; P1_U5787
g3077 nand P1_U3947 P1_REG0_REG_6__SCAN_IN ; P1_U5788
g3078 nand P1_U4024 P1_U4307 ; P1_U5789
g3079 nand P1_U3944 P1_IR_REG_7__SCAN_IN ; P1_U5790
g3080 nand P1_SUB_88_U25 P1_IR_REG_31__SCAN_IN ; P1_U5791
g3081 nand U59 P1_U3946 ; P1_U5792
g3082 nand P1_U3473 P1_U4004 ; P1_U5793
g3083 not P1_U3474 ; P1_U5794
g3084 nand P1_U3947 P1_REG0_REG_7__SCAN_IN ; P1_U5795
g3085 nand P1_U4024 P1_U4326 ; P1_U5796
g3086 nand P1_U3944 P1_IR_REG_8__SCAN_IN ; P1_U5797
g3087 nand P1_SUB_88_U26 P1_IR_REG_31__SCAN_IN ; P1_U5798
g3088 nand U58 P1_U3946 ; P1_U5799
g3089 nand P1_U3476 P1_U4004 ; P1_U5800
g3090 not P1_U3477 ; P1_U5801
g3091 nand P1_U3947 P1_REG0_REG_8__SCAN_IN ; P1_U5802
g3092 nand P1_U4024 P1_U4345 ; P1_U5803
g3093 nand P1_U3944 P1_IR_REG_9__SCAN_IN ; P1_U5804
g3094 nand P1_SUB_88_U160 P1_IR_REG_31__SCAN_IN ; P1_U5805
g3095 nand U57 P1_U3946 ; P1_U5806
g3096 nand P1_U3479 P1_U4004 ; P1_U5807
g3097 not P1_U3480 ; P1_U5808
g3098 nand P1_U3947 P1_REG0_REG_9__SCAN_IN ; P1_U5809
g3099 nand P1_U4024 P1_U4364 ; P1_U5810
g3100 nand P1_U3944 P1_IR_REG_10__SCAN_IN ; P1_U5811
g3101 nand P1_SUB_88_U6 P1_IR_REG_31__SCAN_IN ; P1_U5812
g3102 nand U87 P1_U3946 ; P1_U5813
g3103 nand P1_U3482 P1_U4004 ; P1_U5814
g3104 not P1_U3483 ; P1_U5815
g3105 nand P1_U3947 P1_REG0_REG_10__SCAN_IN ; P1_U5816
g3106 nand P1_U4024 P1_U4383 ; P1_U5817
g3107 nand P1_U3944 P1_IR_REG_11__SCAN_IN ; P1_U5818
g3108 nand P1_SUB_88_U7 P1_IR_REG_31__SCAN_IN ; P1_U5819
g3109 nand U86 P1_U3946 ; P1_U5820
g3110 nand P1_U3485 P1_U4004 ; P1_U5821
g3111 not P1_U3486 ; P1_U5822
g3112 nand P1_U3947 P1_REG0_REG_11__SCAN_IN ; P1_U5823
g3113 nand P1_U4024 P1_U4402 ; P1_U5824
g3114 nand P1_U3944 P1_IR_REG_12__SCAN_IN ; P1_U5825
g3115 nand P1_SUB_88_U8 P1_IR_REG_31__SCAN_IN ; P1_U5826
g3116 nand U85 P1_U3946 ; P1_U5827
g3117 nand P1_U3488 P1_U4004 ; P1_U5828
g3118 not P1_U3489 ; P1_U5829
g3119 nand P1_U3947 P1_REG0_REG_12__SCAN_IN ; P1_U5830
g3120 nand P1_U4024 P1_U4421 ; P1_U5831
g3121 nand P1_U3944 P1_IR_REG_13__SCAN_IN ; P1_U5832
g3122 nand P1_SUB_88_U179 P1_IR_REG_31__SCAN_IN ; P1_U5833
g3123 nand U84 P1_U3946 ; P1_U5834
g3124 nand P1_U3491 P1_U4004 ; P1_U5835
g3125 not P1_U3492 ; P1_U5836
g3126 nand P1_U3947 P1_REG0_REG_13__SCAN_IN ; P1_U5837
g3127 nand P1_U4024 P1_U4440 ; P1_U5838
g3128 nand P1_U3944 P1_IR_REG_14__SCAN_IN ; P1_U5839
g3129 nand P1_SUB_88_U9 P1_IR_REG_31__SCAN_IN ; P1_U5840
g3130 nand U83 P1_U3946 ; P1_U5841
g3131 nand P1_U3494 P1_U4004 ; P1_U5842
g3132 not P1_U3495 ; P1_U5843
g3133 nand P1_U3947 P1_REG0_REG_14__SCAN_IN ; P1_U5844
g3134 nand P1_U4024 P1_U4459 ; P1_U5845
g3135 nand P1_U3944 P1_IR_REG_15__SCAN_IN ; P1_U5846
g3136 nand P1_SUB_88_U10 P1_IR_REG_31__SCAN_IN ; P1_U5847
g3137 nand U82 P1_U3946 ; P1_U5848
g3138 nand P1_U3497 P1_U4004 ; P1_U5849
g3139 not P1_U3498 ; P1_U5850
g3140 nand P1_U3947 P1_REG0_REG_15__SCAN_IN ; P1_U5851
g3141 nand P1_U4024 P1_U4478 ; P1_U5852
g3142 nand P1_U3944 P1_IR_REG_16__SCAN_IN ; P1_U5853
g3143 nand P1_SUB_88_U11 P1_IR_REG_31__SCAN_IN ; P1_U5854
g3144 nand U81 P1_U3946 ; P1_U5855
g3145 nand P1_U3500 P1_U4004 ; P1_U5856
g3146 not P1_U3501 ; P1_U5857
g3147 nand P1_U3947 P1_REG0_REG_16__SCAN_IN ; P1_U5858
g3148 nand P1_U4024 P1_U4497 ; P1_U5859
g3149 nand P1_U3944 P1_IR_REG_17__SCAN_IN ; P1_U5860
g3150 nand P1_SUB_88_U177 P1_IR_REG_31__SCAN_IN ; P1_U5861
g3151 nand U80 P1_U3946 ; P1_U5862
g3152 nand P1_U3503 P1_U4004 ; P1_U5863
g3153 not P1_U3504 ; P1_U5864
g3154 nand P1_U3947 P1_REG0_REG_17__SCAN_IN ; P1_U5865
g3155 nand P1_U4024 P1_U4516 ; P1_U5866
g3156 nand P1_U3944 P1_IR_REG_18__SCAN_IN ; P1_U5867
g3157 nand P1_SUB_88_U12 P1_IR_REG_31__SCAN_IN ; P1_U5868
g3158 nand U79 P1_U3946 ; P1_U5869
g3159 nand P1_U3506 P1_U4004 ; P1_U5870
g3160 not P1_U3507 ; P1_U5871
g3161 nand P1_U3947 P1_REG0_REG_18__SCAN_IN ; P1_U5872
g3162 nand P1_U4024 P1_U4535 ; P1_U5873
g3163 nand U78 P1_U3946 ; P1_U5874
g3164 nand P1_U4004 P1_U3443 ; P1_U5875
g3165 not P1_U3509 ; P1_U5876
g3166 nand P1_U3947 P1_REG0_REG_19__SCAN_IN ; P1_U5877
g3167 nand P1_U4024 P1_U4554 ; P1_U5878
g3168 nand P1_U3947 P1_REG0_REG_20__SCAN_IN ; P1_U5879
g3169 nand P1_U4024 P1_U4573 ; P1_U5880
g3170 nand P1_U3947 P1_REG0_REG_21__SCAN_IN ; P1_U5881
g3171 nand P1_U4024 P1_U4592 ; P1_U5882
g3172 nand P1_U3947 P1_REG0_REG_22__SCAN_IN ; P1_U5883
g3173 nand P1_U4024 P1_U4611 ; P1_U5884
g3174 nand P1_U3947 P1_REG0_REG_23__SCAN_IN ; P1_U5885
g3175 nand P1_U4024 P1_U4630 ; P1_U5886
g3176 nand P1_U3947 P1_REG0_REG_24__SCAN_IN ; P1_U5887
g3177 nand P1_U4024 P1_U4649 ; P1_U5888
g3178 nand P1_U3947 P1_REG0_REG_25__SCAN_IN ; P1_U5889
g3179 nand P1_U4024 P1_U4668 ; P1_U5890
g3180 nand P1_U3947 P1_REG0_REG_26__SCAN_IN ; P1_U5891
g3181 nand P1_U4024 P1_U4687 ; P1_U5892
g3182 nand P1_U3947 P1_REG0_REG_27__SCAN_IN ; P1_U5893
g3183 nand P1_U4024 P1_U4706 ; P1_U5894
g3184 nand P1_U3947 P1_REG0_REG_28__SCAN_IN ; P1_U5895
g3185 nand P1_U4024 P1_U4725 ; P1_U5896
g3186 nand P1_U3947 P1_REG0_REG_29__SCAN_IN ; P1_U5897
g3187 nand P1_U4024 P1_U4745 ; P1_U5898
g3188 nand P1_U3947 P1_REG0_REG_30__SCAN_IN ; P1_U5899
g3189 nand P1_U4024 P1_U4752 ; P1_U5900
g3190 nand P1_U3947 P1_REG0_REG_31__SCAN_IN ; P1_U5901
g3191 nand P1_U4024 P1_U4755 ; P1_U5902
g3192 nand P1_U3948 P1_REG1_REG_0__SCAN_IN ; P1_U5903
g3193 nand P1_U4023 P1_U4188 ; P1_U5904
g3194 nand P1_U3948 P1_REG1_REG_1__SCAN_IN ; P1_U5905
g3195 nand P1_U4023 P1_U4212 ; P1_U5906
g3196 nand P1_U3948 P1_REG1_REG_2__SCAN_IN ; P1_U5907
g3197 nand P1_U4023 P1_U4231 ; P1_U5908
g3198 nand P1_U3948 P1_REG1_REG_3__SCAN_IN ; P1_U5909
g3199 nand P1_U4023 P1_U4250 ; P1_U5910
g3200 nand P1_U3948 P1_REG1_REG_4__SCAN_IN ; P1_U5911
g3201 nand P1_U4023 P1_U4269 ; P1_U5912
g3202 nand P1_U3948 P1_REG1_REG_5__SCAN_IN ; P1_U5913
g3203 nand P1_U4023 P1_U4288 ; P1_U5914
g3204 nand P1_U3948 P1_REG1_REG_6__SCAN_IN ; P1_U5915
g3205 nand P1_U4023 P1_U4307 ; P1_U5916
g3206 nand P1_U3948 P1_REG1_REG_7__SCAN_IN ; P1_U5917
g3207 nand P1_U4023 P1_U4326 ; P1_U5918
g3208 nand P1_U3948 P1_REG1_REG_8__SCAN_IN ; P1_U5919
g3209 nand P1_U4023 P1_U4345 ; P1_U5920
g3210 nand P1_U3948 P1_REG1_REG_9__SCAN_IN ; P1_U5921
g3211 nand P1_U4023 P1_U4364 ; P1_U5922
g3212 nand P1_U3948 P1_REG1_REG_10__SCAN_IN ; P1_U5923
g3213 nand P1_U4023 P1_U4383 ; P1_U5924
g3214 nand P1_U3948 P1_REG1_REG_11__SCAN_IN ; P1_U5925
g3215 nand P1_U4023 P1_U4402 ; P1_U5926
g3216 nand P1_U3948 P1_REG1_REG_12__SCAN_IN ; P1_U5927
g3217 nand P1_U4023 P1_U4421 ; P1_U5928
g3218 nand P1_U3948 P1_REG1_REG_13__SCAN_IN ; P1_U5929
g3219 nand P1_U4023 P1_U4440 ; P1_U5930
g3220 nand P1_U3948 P1_REG1_REG_14__SCAN_IN ; P1_U5931
g3221 nand P1_U4023 P1_U4459 ; P1_U5932
g3222 nand P1_U3948 P1_REG1_REG_15__SCAN_IN ; P1_U5933
g3223 nand P1_U4023 P1_U4478 ; P1_U5934
g3224 nand P1_U3948 P1_REG1_REG_16__SCAN_IN ; P1_U5935
g3225 nand P1_U4023 P1_U4497 ; P1_U5936
g3226 nand P1_U3948 P1_REG1_REG_17__SCAN_IN ; P1_U5937
g3227 nand P1_U4023 P1_U4516 ; P1_U5938
g3228 nand P1_U3948 P1_REG1_REG_18__SCAN_IN ; P1_U5939
g3229 nand P1_U4023 P1_U4535 ; P1_U5940
g3230 nand P1_U3948 P1_REG1_REG_19__SCAN_IN ; P1_U5941
g3231 nand P1_U4023 P1_U4554 ; P1_U5942
g3232 nand P1_U3948 P1_REG1_REG_20__SCAN_IN ; P1_U5943
g3233 nand P1_U4023 P1_U4573 ; P1_U5944
g3234 nand P1_U3948 P1_REG1_REG_21__SCAN_IN ; P1_U5945
g3235 nand P1_U4023 P1_U4592 ; P1_U5946
g3236 nand P1_U3948 P1_REG1_REG_22__SCAN_IN ; P1_U5947
g3237 nand P1_U4023 P1_U4611 ; P1_U5948
g3238 nand P1_U3948 P1_REG1_REG_23__SCAN_IN ; P1_U5949
g3239 nand P1_U4023 P1_U4630 ; P1_U5950
g3240 nand P1_U3948 P1_REG1_REG_24__SCAN_IN ; P1_U5951
g3241 nand P1_U4023 P1_U4649 ; P1_U5952
g3242 nand P1_U3948 P1_REG1_REG_25__SCAN_IN ; P1_U5953
g3243 nand P1_U4023 P1_U4668 ; P1_U5954
g3244 nand P1_U3948 P1_REG1_REG_26__SCAN_IN ; P1_U5955
g3245 nand P1_U4023 P1_U4687 ; P1_U5956
g3246 nand P1_U3948 P1_REG1_REG_27__SCAN_IN ; P1_U5957
g3247 nand P1_U4023 P1_U4706 ; P1_U5958
g3248 nand P1_U3948 P1_REG1_REG_28__SCAN_IN ; P1_U5959
g3249 nand P1_U4023 P1_U4725 ; P1_U5960
g3250 nand P1_U3948 P1_REG1_REG_29__SCAN_IN ; P1_U5961
g3251 nand P1_U4023 P1_U4745 ; P1_U5962
g3252 nand P1_U3948 P1_REG1_REG_30__SCAN_IN ; P1_U5963
g3253 nand P1_U4023 P1_U4752 ; P1_U5964
g3254 nand P1_U3948 P1_REG1_REG_31__SCAN_IN ; P1_U5965
g3255 nand P1_U4023 P1_U4755 ; P1_U5966
g3256 nand P1_U3417 P1_REG2_REG_0__SCAN_IN ; P1_U5967
g3257 nand P1_U4022 P1_U3373 ; P1_U5968
g3258 nand P1_U3417 P1_REG2_REG_1__SCAN_IN ; P1_U5969
g3259 nand P1_U4022 P1_U3375 ; P1_U5970
g3260 nand P1_U3417 P1_REG2_REG_2__SCAN_IN ; P1_U5971
g3261 nand P1_U4022 P1_U3376 ; P1_U5972
g3262 nand P1_U3417 P1_REG2_REG_3__SCAN_IN ; P1_U5973
g3263 nand P1_U4022 P1_U3377 ; P1_U5974
g3264 nand P1_U3417 P1_REG2_REG_4__SCAN_IN ; P1_U5975
g3265 nand P1_U4022 P1_U3378 ; P1_U5976
g3266 nand P1_U3417 P1_REG2_REG_5__SCAN_IN ; P1_U5977
g3267 nand P1_U4022 P1_U3379 ; P1_U5978
g3268 nand P1_U3417 P1_REG2_REG_6__SCAN_IN ; P1_U5979
g3269 nand P1_U4022 P1_U3380 ; P1_U5980
g3270 nand P1_U3417 P1_REG2_REG_7__SCAN_IN ; P1_U5981
g3271 nand P1_U4022 P1_U3381 ; P1_U5982
g3272 nand P1_U3417 P1_REG2_REG_8__SCAN_IN ; P1_U5983
g3273 nand P1_U4022 P1_U3382 ; P1_U5984
g3274 nand P1_U3417 P1_REG2_REG_9__SCAN_IN ; P1_U5985
g3275 nand P1_U4022 P1_U3383 ; P1_U5986
g3276 nand P1_U3417 P1_REG2_REG_10__SCAN_IN ; P1_U5987
g3277 nand P1_U4022 P1_U3384 ; P1_U5988
g3278 nand P1_U3417 P1_REG2_REG_11__SCAN_IN ; P1_U5989
g3279 nand P1_U4022 P1_U3385 ; P1_U5990
g3280 nand P1_U3417 P1_REG2_REG_12__SCAN_IN ; P1_U5991
g3281 nand P1_U4022 P1_U3386 ; P1_U5992
g3282 nand P1_U3417 P1_REG2_REG_13__SCAN_IN ; P1_U5993
g3283 nand P1_U4022 P1_U3387 ; P1_U5994
g3284 nand P1_U3417 P1_REG2_REG_14__SCAN_IN ; P1_U5995
g3285 nand P1_U4022 P1_U3388 ; P1_U5996
g3286 nand P1_U3417 P1_REG2_REG_15__SCAN_IN ; P1_U5997
g3287 nand P1_U4022 P1_U3389 ; P1_U5998
g3288 nand P1_U3417 P1_REG2_REG_16__SCAN_IN ; P1_U5999
g3289 nand P1_U4022 P1_U3390 ; P1_U6000
g3290 nand P1_U3417 P1_REG2_REG_17__SCAN_IN ; P1_U6001
g3291 nand P1_U4022 P1_U3391 ; P1_U6002
g3292 nand P1_U3417 P1_REG2_REG_18__SCAN_IN ; P1_U6003
g3293 nand P1_U4022 P1_U3392 ; P1_U6004
g3294 nand P1_U3417 P1_REG2_REG_19__SCAN_IN ; P1_U6005
g3295 nand P1_U4022 P1_U3393 ; P1_U6006
g3296 nand P1_U3417 P1_REG2_REG_20__SCAN_IN ; P1_U6007
g3297 nand P1_U4022 P1_U3395 ; P1_U6008
g3298 nand P1_U3417 P1_REG2_REG_21__SCAN_IN ; P1_U6009
g3299 nand P1_U4022 P1_U3397 ; P1_U6010
g3300 nand P1_U3417 P1_REG2_REG_22__SCAN_IN ; P1_U6011
g3301 nand P1_U4022 P1_U3399 ; P1_U6012
g3302 nand P1_U3417 P1_REG2_REG_23__SCAN_IN ; P1_U6013
g3303 nand P1_U4022 P1_U3401 ; P1_U6014
g3304 nand P1_U3417 P1_REG2_REG_24__SCAN_IN ; P1_U6015
g3305 nand P1_U4022 P1_U3403 ; P1_U6016
g3306 nand P1_U3417 P1_REG2_REG_25__SCAN_IN ; P1_U6017
g3307 nand P1_U4022 P1_U3405 ; P1_U6018
g3308 nand P1_U3417 P1_REG2_REG_26__SCAN_IN ; P1_U6019
g3309 nand P1_U4022 P1_U3407 ; P1_U6020
g3310 nand P1_U3417 P1_REG2_REG_27__SCAN_IN ; P1_U6021
g3311 nand P1_U4022 P1_U3409 ; P1_U6022
g3312 nand P1_U3417 P1_REG2_REG_28__SCAN_IN ; P1_U6023
g3313 nand P1_U4022 P1_U3411 ; P1_U6024
g3314 nand P1_U3417 P1_REG2_REG_29__SCAN_IN ; P1_U6025
g3315 nand P1_U4022 P1_U3413 ; P1_U6026
g3316 nand P1_U3417 P1_REG2_REG_30__SCAN_IN ; P1_U6027
g3317 nand P1_U4026 P1_U4022 ; P1_U6028
g3318 nand P1_U3417 P1_REG2_REG_31__SCAN_IN ; P1_U6029
g3319 nand P1_U4026 P1_U4022 ; P1_U6030
g3320 nand P1_U3425 P1_DATAO_REG_0__SCAN_IN ; P1_U6031
g3321 nand P1_U4006 P1_U3075 ; P1_U6032
g3322 nand P1_U3425 P1_DATAO_REG_1__SCAN_IN ; P1_U6033
g3323 nand P1_U4006 P1_U3076 ; P1_U6034
g3324 nand P1_U3425 P1_DATAO_REG_2__SCAN_IN ; P1_U6035
g3325 nand P1_U4006 P1_U3066 ; P1_U6036
g3326 nand P1_U3425 P1_DATAO_REG_3__SCAN_IN ; P1_U6037
g3327 nand P1_U4006 P1_U3062 ; P1_U6038
g3328 nand P1_U3425 P1_DATAO_REG_4__SCAN_IN ; P1_U6039
g3329 nand P1_U4006 P1_U3058 ; P1_U6040
g3330 nand P1_U3425 P1_DATAO_REG_5__SCAN_IN ; P1_U6041
g3331 nand P1_U4006 P1_U3065 ; P1_U6042
g3332 nand P1_U3425 P1_DATAO_REG_6__SCAN_IN ; P1_U6043
g3333 nand P1_U4006 P1_U3069 ; P1_U6044
g3334 nand P1_U3425 P1_DATAO_REG_7__SCAN_IN ; P1_U6045
g3335 nand P1_U4006 P1_U3068 ; P1_U6046
g3336 nand P1_U3425 P1_DATAO_REG_8__SCAN_IN ; P1_U6047
g3337 nand P1_U4006 P1_U3082 ; P1_U6048
g3338 nand P1_U3425 P1_DATAO_REG_9__SCAN_IN ; P1_U6049
g3339 nand P1_U4006 P1_U3081 ; P1_U6050
g3340 nand P1_U3425 P1_DATAO_REG_10__SCAN_IN ; P1_U6051
g3341 nand P1_U4006 P1_U3060 ; P1_U6052
g3342 nand P1_U3425 P1_DATAO_REG_11__SCAN_IN ; P1_U6053
g3343 nand P1_U4006 P1_U3061 ; P1_U6054
g3344 nand P1_U3425 P1_DATAO_REG_12__SCAN_IN ; P1_U6055
g3345 nand P1_U4006 P1_U3070 ; P1_U6056
g3346 nand P1_U3425 P1_DATAO_REG_13__SCAN_IN ; P1_U6057
g3347 nand P1_U4006 P1_U3078 ; P1_U6058
g3348 nand P1_U3425 P1_DATAO_REG_14__SCAN_IN ; P1_U6059
g3349 nand P1_U4006 P1_U3077 ; P1_U6060
g3350 nand P1_U3425 P1_DATAO_REG_15__SCAN_IN ; P1_U6061
g3351 nand P1_U4006 P1_U3072 ; P1_U6062
g3352 nand P1_U3425 P1_DATAO_REG_16__SCAN_IN ; P1_U6063
g3353 nand P1_U4006 P1_U3071 ; P1_U6064
g3354 nand P1_U3425 P1_DATAO_REG_17__SCAN_IN ; P1_U6065
g3355 nand P1_U4006 P1_U3067 ; P1_U6066
g3356 nand P1_U3425 P1_DATAO_REG_18__SCAN_IN ; P1_U6067
g3357 nand P1_U4006 P1_U3080 ; P1_U6068
g3358 nand P1_U3425 P1_DATAO_REG_19__SCAN_IN ; P1_U6069
g3359 nand P1_U4006 P1_U3079 ; P1_U6070
g3360 nand P1_U3425 P1_DATAO_REG_20__SCAN_IN ; P1_U6071
g3361 nand P1_U4006 P1_U3074 ; P1_U6072
g3362 nand P1_U3425 P1_DATAO_REG_21__SCAN_IN ; P1_U6073
g3363 nand P1_U4006 P1_U3073 ; P1_U6074
g3364 nand P1_U3425 P1_DATAO_REG_22__SCAN_IN ; P1_U6075
g3365 nand P1_U4006 P1_U3059 ; P1_U6076
g3366 nand P1_U3425 P1_DATAO_REG_23__SCAN_IN ; P1_U6077
g3367 nand P1_U4006 P1_U3064 ; P1_U6078
g3368 nand P1_U3425 P1_DATAO_REG_24__SCAN_IN ; P1_U6079
g3369 nand P1_U4006 P1_U3063 ; P1_U6080
g3370 nand P1_U3425 P1_DATAO_REG_25__SCAN_IN ; P1_U6081
g3371 nand P1_U4006 P1_U3056 ; P1_U6082
g3372 nand P1_U3425 P1_DATAO_REG_26__SCAN_IN ; P1_U6083
g3373 nand P1_U4006 P1_U3055 ; P1_U6084
g3374 nand P1_U3425 P1_DATAO_REG_27__SCAN_IN ; P1_U6085
g3375 nand P1_U4006 P1_U3051 ; P1_U6086
g3376 nand P1_U3425 P1_DATAO_REG_28__SCAN_IN ; P1_U6087
g3377 nand P1_U4006 P1_U3052 ; P1_U6088
g3378 nand P1_U3425 P1_DATAO_REG_29__SCAN_IN ; P1_U6089
g3379 nand P1_U4006 P1_U3053 ; P1_U6090
g3380 nand P1_U3425 P1_DATAO_REG_30__SCAN_IN ; P1_U6091
g3381 nand P1_U4006 P1_U3057 ; P1_U6092
g3382 nand P1_U3425 P1_DATAO_REG_31__SCAN_IN ; P1_U6093
g3383 nand P1_U4006 P1_U3054 ; P1_U6094
g3384 nand P1_U4007 P1_U3052 ; P1_U6095
g3385 nand P1_U3410 P1_U4692 ; P1_U6096
g3386 nand P1_U6096 P1_U6095 ; P1_U6097
g3387 nand P1_U4008 P1_U3051 ; P1_U6098
g3388 nand P1_U3408 P1_U4673 ; P1_U6099
g3389 nand P1_U6099 P1_U6098 ; P1_U6100
g3390 nand P1_U4011 P1_U3063 ; P1_U6101
g3391 nand P1_U3402 P1_U4616 ; P1_U6102
g3392 nand P1_U6102 P1_U6101 ; P1_U6103
g3393 nand P1_U4012 P1_U3064 ; P1_U6104
g3394 nand P1_U3400 P1_U4597 ; P1_U6105
g3395 nand P1_U6105 P1_U6104 ; P1_U6106
g3396 nand P1_U4014 P1_U3073 ; P1_U6107
g3397 nand P1_U3396 P1_U4559 ; P1_U6108
g3398 nand P1_U6108 P1_U6107 ; P1_U6109
g3399 nand P1_U4013 P1_U3059 ; P1_U6110
g3400 nand P1_U3398 P1_U4578 ; P1_U6111
g3401 nand P1_U6111 P1_U6110 ; P1_U6112
g3402 nand P1_U4010 P1_U3056 ; P1_U6113
g3403 nand P1_U3404 P1_U4635 ; P1_U6114
g3404 nand P1_U6114 P1_U6113 ; P1_U6115
g3405 nand P1_U4009 P1_U3055 ; P1_U6116
g3406 nand P1_U3406 P1_U4654 ; P1_U6117
g3407 nand P1_U6117 P1_U6116 ; P1_U6118
g3408 nand P1_U5864 P1_U4483 ; P1_U6119
g3409 nand P1_U3504 P1_U3067 ; P1_U6120
g3410 nand P1_U6120 P1_U6119 ; P1_U6121
g3411 nand P1_U5801 P1_U4312 ; P1_U6122
g3412 nand P1_U3477 P1_U3082 ; P1_U6123
g3413 nand P1_U6123 P1_U6122 ; P1_U6124
g3414 nand P1_U5808 P1_U4331 ; P1_U6125
g3415 nand P1_U3480 P1_U3081 ; P1_U6126
g3416 nand P1_U6126 P1_U6125 ; P1_U6127
g3417 nand P1_U5836 P1_U4407 ; P1_U6128
g3418 nand P1_U3492 P1_U3078 ; P1_U6129
g3419 nand P1_U6129 P1_U6128 ; P1_U6130
g3420 nand P1_U5843 P1_U4426 ; P1_U6131
g3421 nand P1_U3495 P1_U3077 ; P1_U6132
g3422 nand P1_U6132 P1_U6131 ; P1_U6133
g3423 nand P1_U5737 P1_U4198 ; P1_U6134
g3424 nand P1_U3451 P1_U3075 ; P1_U6135
g3425 nand P1_U6135 P1_U6134 ; P1_U6136
g3426 nand P1_U5752 P1_U4174 ; P1_U6137
g3427 nand P1_U3456 P1_U3076 ; P1_U6138
g3428 nand P1_U6138 P1_U6137 ; P1_U6139
g3429 nand P1_U5850 P1_U4445 ; P1_U6140
g3430 nand P1_U3498 P1_U3072 ; P1_U6141
g3431 nand P1_U6141 P1_U6140 ; P1_U6142
g3432 nand P1_U5857 P1_U4464 ; P1_U6143
g3433 nand P1_U3501 P1_U3071 ; P1_U6144
g3434 nand P1_U6144 P1_U6143 ; P1_U6145
g3435 nand P1_U5787 P1_U4274 ; P1_U6146
g3436 nand P1_U3471 P1_U3069 ; P1_U6147
g3437 nand P1_U6147 P1_U6146 ; P1_U6148
g3438 nand P1_U5794 P1_U4293 ; P1_U6149
g3439 nand P1_U3474 P1_U3068 ; P1_U6150
g3440 nand P1_U6150 P1_U6149 ; P1_U6151
g3441 nand P1_U5829 P1_U4388 ; P1_U6152
g3442 nand P1_U3489 P1_U3070 ; P1_U6153
g3443 nand P1_U6153 P1_U6152 ; P1_U6154
g3444 nand P1_U5759 P1_U4193 ; P1_U6155
g3445 nand P1_U3459 P1_U3066 ; P1_U6156
g3446 nand P1_U6156 P1_U6155 ; P1_U6157
g3447 nand P1_U5766 P1_U4217 ; P1_U6158
g3448 nand P1_U3462 P1_U3062 ; P1_U6159
g3449 nand P1_U6159 P1_U6158 ; P1_U6160
g3450 nand P1_U5780 P1_U4255 ; P1_U6161
g3451 nand P1_U3468 P1_U3065 ; P1_U6162
g3452 nand P1_U6162 P1_U6161 ; P1_U6163
g3453 nand P1_U5871 P1_U4502 ; P1_U6164
g3454 nand P1_U3507 P1_U3080 ; P1_U6165
g3455 nand P1_U6165 P1_U6164 ; P1_U6166
g3456 nand P1_U4016 P1_U3054 ; P1_U6167
g3457 nand P1_U3415 P1_U4749 ; P1_U6168
g3458 nand P1_U6168 P1_U6167 ; P1_U6169
g3459 nand P1_U5876 P1_U4521 ; P1_U6170
g3460 nand P1_U3509 P1_U3079 ; P1_U6171
g3461 nand P1_U6171 P1_U6170 ; P1_U6172
g3462 nand P1_U5822 P1_U4369 ; P1_U6173
g3463 nand P1_U3486 P1_U3061 ; P1_U6174
g3464 nand P1_U6174 P1_U6173 ; P1_U6175
g3465 nand P1_U5773 P1_U4236 ; P1_U6176
g3466 nand P1_U3465 P1_U3058 ; P1_U6177
g3467 nand P1_U6177 P1_U6176 ; P1_U6178
g3468 nand P1_U5815 P1_U4350 ; P1_U6179
g3469 nand P1_U3483 P1_U3060 ; P1_U6180
g3470 nand P1_U6180 P1_U6179 ; P1_U6181
g3471 nand P1_U4015 P1_U3074 ; P1_U6182
g3472 nand P1_U3394 P1_U4540 ; P1_U6183
g3473 nand P1_U6183 P1_U6182 ; P1_U6184
g3474 nand P1_U4018 P1_U3053 ; P1_U6185
g3475 nand P1_U3412 P1_U4711 ; P1_U6186
g3476 nand P1_U6186 P1_U6185 ; P1_U6187
g3477 nand P1_U4017 P1_U3057 ; P1_U6188
g3478 nand P1_U3414 P1_U4729 ; P1_U6189
g3479 nand P1_U6189 P1_U6188 ; P1_U6190
g3480 nand P1_U5119 P1_U3987 ; P1_U6191
g3481 nand P1_U3354 P1_U3982 ; P1_U6192
g3482 nand P1_U6192 P1_U6191 ; P1_U6193
g3483 nand P1_U3439 P1_U5710 P1_U3983 P1_U3448 ; P1_U6194
g3484 nand P1_U6193 P1_U5719 ; P1_U6195
g3485 nand P1_U6195 P1_U6194 ; P1_U6196
g3486 nand P1_R1375_U14 P1_U3987 P1_U5716 ; P1_U6197
g3487 nand P1_U6196 P1_U3442 ; P1_U6198
g3488 nand P1_U4019 P1_U3022 P1_U3983 ; P1_U6199
g3489 nand P1_U3988 P1_U3992 P1_R1360_U14 ; P1_U6200
g3490 nand P1_U3081 P1_R1352_U6 ; P1_U6201
g3491 nand P1_U3081 P1_U3985 ; P1_U6202
g3492 nand P1_U3082 P1_R1352_U6 ; P1_U6203
g3493 nand P1_U3082 P1_U3985 ; P1_U6204
g3494 nand P1_U3068 P1_R1352_U6 ; P1_U6205
g3495 nand P1_U3068 P1_U3985 ; P1_U6206
g3496 nand P1_U3069 P1_R1352_U6 ; P1_U6207
g3497 nand P1_U3069 P1_U3985 ; P1_U6208
g3498 nand P1_U3065 P1_R1352_U6 ; P1_U6209
g3499 nand P1_U3065 P1_U3985 ; P1_U6210
g3500 nand P1_U3058 P1_R1352_U6 ; P1_U6211
g3501 nand P1_U3058 P1_U3985 ; P1_U6212
g3502 nand P1_U3062 P1_R1352_U6 ; P1_U6213
g3503 nand P1_U3062 P1_U3985 ; P1_U6214
g3504 nand P1_R1309_U8 P1_R1352_U6 ; P1_U6215
g3505 nand P1_U3054 P1_U3985 ; P1_U6216
g3506 nand P1_R1309_U6 P1_R1352_U6 ; P1_U6217
g3507 nand P1_U3057 P1_U3985 ; P1_U6218
g3508 nand P1_U3066 P1_R1352_U6 ; P1_U6219
g3509 nand P1_U3066 P1_U3985 ; P1_U6220
g3510 nand P1_U3053 P1_R1352_U6 ; P1_U6221
g3511 nand P1_U3053 P1_U3985 ; P1_U6222
g3512 nand P1_U3052 P1_R1352_U6 ; P1_U6223
g3513 nand P1_U3052 P1_U3985 ; P1_U6224
g3514 nand P1_U3051 P1_R1352_U6 ; P1_U6225
g3515 nand P1_U3051 P1_U3985 ; P1_U6226
g3516 nand P1_U3055 P1_R1352_U6 ; P1_U6227
g3517 nand P1_U3055 P1_U3985 ; P1_U6228
g3518 nand P1_U3056 P1_R1352_U6 ; P1_U6229
g3519 nand P1_U3056 P1_U3985 ; P1_U6230
g3520 nand P1_U3063 P1_R1352_U6 ; P1_U6231
g3521 nand P1_U3063 P1_U3985 ; P1_U6232
g3522 nand P1_U3064 P1_R1352_U6 ; P1_U6233
g3523 nand P1_U3064 P1_U3985 ; P1_U6234
g3524 nand P1_U3059 P1_R1352_U6 ; P1_U6235
g3525 nand P1_U3059 P1_U3985 ; P1_U6236
g3526 nand P1_U3073 P1_R1352_U6 ; P1_U6237
g3527 nand P1_U3073 P1_U3985 ; P1_U6238
g3528 nand P1_U3074 P1_R1352_U6 ; P1_U6239
g3529 nand P1_U3074 P1_U3985 ; P1_U6240
g3530 nand P1_U3076 P1_R1352_U6 ; P1_U6241
g3531 nand P1_U3076 P1_U3985 ; P1_U6242
g3532 nand P1_U3079 P1_R1352_U6 ; P1_U6243
g3533 nand P1_U3079 P1_U3985 ; P1_U6244
g3534 nand P1_U3080 P1_R1352_U6 ; P1_U6245
g3535 nand P1_U3080 P1_U3985 ; P1_U6246
g3536 nand P1_U3067 P1_R1352_U6 ; P1_U6247
g3537 nand P1_U3067 P1_U3985 ; P1_U6248
g3538 nand P1_U3071 P1_R1352_U6 ; P1_U6249
g3539 nand P1_U3071 P1_U3985 ; P1_U6250
g3540 nand P1_U3072 P1_R1352_U6 ; P1_U6251
g3541 nand P1_U3072 P1_U3985 ; P1_U6252
g3542 nand P1_U3077 P1_R1352_U6 ; P1_U6253
g3543 nand P1_U3077 P1_U3985 ; P1_U6254
g3544 nand P1_U3078 P1_R1352_U6 ; P1_U6255
g3545 nand P1_U3078 P1_U3985 ; P1_U6256
g3546 nand P1_U3070 P1_R1352_U6 ; P1_U6257
g3547 nand P1_U3070 P1_U3985 ; P1_U6258
g3548 nand P1_U3061 P1_R1352_U6 ; P1_U6259
g3549 nand P1_U3061 P1_U3985 ; P1_U6260
g3550 nand P1_U3060 P1_R1352_U6 ; P1_U6261
g3551 nand P1_U3060 P1_U3985 ; P1_U6262
g3552 nand P1_U3075 P1_R1352_U6 ; P1_U6263
g3553 nand P1_U3075 P1_U3985 ; P1_U6264
g3554 nand P1_U3449 P1_U5396 ; P1_U6265
g3555 nand P1_U3015 P1_U5731 P1_REG2_REG_0__SCAN_IN ; P1_U6266
g3556 and P2_U5711 P2_U3441 P2_U3439 ; P2_U3014
g3557 and P2_U3439 P2_U3441 P2_U3445 ; P2_U3015
g3558 and P2_U3954 P2_U5714 ; P2_U3016
g3559 and P2_U3961 P2_U3440 ; P2_U3017
g3560 and P2_U3439 P2_U3445 P2_U3440 ; P2_U3018
g3561 and P2_U5674 P2_U3439 ; P2_U3019
g3562 and P2_U3629 P2_U3624 ; P2_U3020
g3563 and P2_U5733 P2_U3444 ; P2_U3021
g3564 and P2_U3447 P2_U3444 ; P2_U3022
g3565 and P2_U3442 P2_U3443 ; P2_U3023
g3566 and P2_U5723 P2_U3443 ; P2_U3024
g3567 and P2_U5720 P2_U3442 ; P2_U3025
g3568 and P2_U5723 P2_U5720 ; P2_U3026
g3569 and P2_U3048 P2_STATE_REG_SCAN_IN ; P2_U3027
g3570 and P2_U3050 P2_U5708 ; P2_U3028
g3571 and P2_U3811 P2_U3424 ; P2_U3029
g3572 and P2_U3982 P2_U5728 ; P2_U3030
g3573 and P2_U3949 P2_U5714 ; P2_U3031
g3574 and P2_U3890 P2_U3965 ; P2_U3032
g3575 and P2_U3359 P2_STATE_REG_SCAN_IN ; P2_U3033
g3576 and P2_U3956 P2_U3983 ; P2_U3034
g3577 and P2_U3983 P2_U4713 ; P2_U3035
g3578 and P2_U3957 P2_U3983 ; P2_U3036
g3579 and P2_U3751 P2_U3983 ; P2_U3037
g3580 and P2_U3982 P2_U3444 ; P2_U3038
g3581 and P2_U3965 P2_U5728 ; P2_U3039
g3582 and P2_U3983 P2_U3030 ; P2_U3040
g3583 and P2_U3965 P2_U3444 ; P2_U3041
g3584 and P2_U3029 P2_U5733 ; P2_U3042
g3585 and P2_U3029 P2_U5728 ; P2_U3043
g3586 and P2_U3029 P2_U3022 ; P2_U3044
g3587 and P2_U3027 P2_U3424 ; P2_U3045
g3588 and P2_U5196 P2_STATE_REG_SCAN_IN ; P2_U3046
g3589 and P2_U3027 P2_U5198 ; P2_U3047
g3590 and P2_U5701 P2_U3420 ; P2_U3048
g3591 and P2_U3630 P2_U3020 ; P2_U3049
g3592 and P2_U5714 P2_U3445 ; P2_U3050
g3593 and P2_U3950 P2_U4709 ; P2_U3051
g3594 and P2_U3422 P2_STATE_REG_SCAN_IN ; P2_U3052
g3595 nand P2_U4623 P2_U4624 P2_U4622 P2_U4625 ; P2_U3053
g3596 nand P2_U4642 P2_U4643 P2_U4641 P2_U4644 ; P2_U3054
g3597 nand P2_U4663 P2_U4662 P2_U4661 P2_U4660 ; P2_U3055
g3598 nand P2_U4700 P2_U4701 P2_U4699 ; P2_U3056
g3599 nand P2_U4604 P2_U4605 P2_U4603 P2_U4606 ; P2_U3057
g3600 nand P2_U4585 P2_U4586 P2_U4584 P2_U4587 ; P2_U3058
g3601 nand P2_U4680 P2_U4681 P2_U4679 ; P2_U3059
g3602 nand P2_U4188 P2_U4187 P2_U4186 P2_U4185 ; P2_U3060
g3603 nand P2_U4528 P2_U4529 P2_U4527 P2_U4530 ; P2_U3061
g3604 nand P2_U4302 P2_U4301 P2_U4300 P2_U4299 ; P2_U3062
g3605 nand P2_U4321 P2_U4320 P2_U4319 P2_U4318 ; P2_U3063
g3606 nand P2_U4169 P2_U4168 P2_U4167 P2_U4166 ; P2_U3064
g3607 nand P2_U4566 P2_U4567 P2_U4565 P2_U4568 ; P2_U3065
g3608 nand P2_U4547 P2_U4548 P2_U4546 P2_U4549 ; P2_U3066
g3609 nand P2_U4207 P2_U4206 P2_U4205 P2_U4204 ; P2_U3067
g3610 nand P2_U4147 P2_U4146 P2_U5755 P2_U5754 ; P2_U3068
g3611 nand P2_U4433 P2_U4434 P2_U4432 P2_U4435 ; P2_U3069
g3612 nand P2_U4245 P2_U4244 P2_U4243 P2_U4242 ; P2_U3070
g3613 nand P2_U4226 P2_U4225 P2_U4224 P2_U4223 ; P2_U3071
g3614 nand P2_U4340 P2_U4339 P2_U4338 P2_U4337 ; P2_U3072
g3615 nand P2_U4416 P2_U4415 P2_U4414 P2_U4413 ; P2_U3073
g3616 nand P2_U4397 P2_U4396 P2_U4395 P2_U4394 ; P2_U3074
g3617 nand P2_U4509 P2_U4510 P2_U4508 P2_U4511 ; P2_U3075
g3618 nand P2_U4490 P2_U4491 P2_U4489 P2_U4492 ; P2_U3076
g3619 nand P2_U4150 P2_U4149 P2_U5748 P2_U5747 ; P2_U3077
g3620 nand P2_U4129 P2_U4128 P2_U5725 P2_U5724 ; P2_U3078
g3621 nand P2_U4378 P2_U4377 P2_U4376 P2_U4375 ; P2_U3079
g3622 nand P2_U4359 P2_U4358 P2_U4357 P2_U4356 ; P2_U3080
g3623 nand P2_U4471 P2_U4472 P2_U4470 P2_U4473 ; P2_U3081
g3624 nand P2_U4452 P2_U4453 P2_U4451 P2_U4454 ; P2_U3082
g3625 nand P2_U4283 P2_U4282 P2_U4281 P2_U4280 ; P2_U3083
g3626 nand P2_U4264 P2_U4263 P2_U4262 P2_U4261 ; P2_U3084
g3627 nand P2_U5596 P2_U5595 ; P2_U3085
g3628 nand P2_U5598 P2_U5597 ; P2_U3086
g3629 nand P2_U5603 P2_U5604 P2_U5602 ; P2_U3087
g3630 nand P2_U5606 P2_U5607 P2_U5605 ; P2_U3088
g3631 nand P2_U5609 P2_U5610 P2_U5608 ; P2_U3089
g3632 nand P2_U5612 P2_U5613 P2_U5611 ; P2_U3090
g3633 nand P2_U5615 P2_U5616 P2_U5614 ; P2_U3091
g3634 nand P2_U5618 P2_U5619 P2_U5617 ; P2_U3092
g3635 nand P2_U5621 P2_U5622 P2_U5620 ; P2_U3093
g3636 nand P2_U5624 P2_U5625 P2_U5623 ; P2_U3094
g3637 nand P2_U5627 P2_U5628 P2_U5626 ; P2_U3095
g3638 nand P2_U5630 P2_U5631 P2_U5629 ; P2_U3096
g3639 nand P2_U5636 P2_U5637 P2_U5635 ; P2_U3097
g3640 nand P2_U5639 P2_U5640 P2_U5638 ; P2_U3098
g3641 nand P2_U5642 P2_U5643 P2_U5641 ; P2_U3099
g3642 nand P2_U5645 P2_U5646 P2_U5644 ; P2_U3100
g3643 nand P2_U5648 P2_U5649 P2_U5647 ; P2_U3101
g3644 nand P2_U5651 P2_U5652 P2_U5650 ; P2_U3102
g3645 nand P2_U5654 P2_U5655 P2_U5653 ; P2_U3103
g3646 nand P2_U5657 P2_U5658 P2_U5656 ; P2_U3104
g3647 nand P2_U5660 P2_U5659 P2_U5661 ; P2_U3105
g3648 nand P2_U5663 P2_U5662 P2_U5664 ; P2_U3106
g3649 nand P2_U5578 P2_U5577 P2_U5579 ; P2_U3107
g3650 nand P2_U5581 P2_U5580 P2_U5582 ; P2_U3108
g3651 nand P2_U5584 P2_U5583 P2_U5585 ; P2_U3109
g3652 nand P2_U5587 P2_U5586 P2_U5588 ; P2_U3110
g3653 nand P2_U5590 P2_U5589 P2_U5591 ; P2_U3111
g3654 nand P2_U5593 P2_U5592 P2_U5594 ; P2_U3112
g3655 nand P2_U5601 P2_U5599 P2_U5600 ; P2_U3113
g3656 nand P2_U5633 P2_U5632 P2_U5634 ; P2_U3114
g3657 nand P2_U5666 P2_U5665 P2_U5667 ; P2_U3115
g3658 nand P2_U5669 P2_U5668 ; P2_U3116
g3659 nand P2_U5527 P2_U5526 ; P2_U3117
g3660 and P2_U5673 P2_U5672 ; P2_U3118
g3661 nand P2_U3436 P2_U5531 P2_U5532 ; P2_U3119
g3662 nand P2_U3436 P2_U5533 P2_U5534 ; P2_U3120
g3663 nand P2_U3436 P2_U5535 P2_U5536 ; P2_U3121
g3664 nand P2_U3436 P2_U5537 P2_U5538 ; P2_U3122
g3665 nand P2_U3436 P2_U5539 P2_U5540 ; P2_U3123
g3666 nand P2_U3436 P2_U5541 P2_U5542 ; P2_U3124
g3667 nand P2_U3436 P2_U5543 P2_U5544 ; P2_U3125
g3668 nand P2_U3436 P2_U5545 P2_U5546 ; P2_U3126
g3669 nand P2_U3436 P2_U5547 P2_U5548 ; P2_U3127
g3670 nand P2_U3436 P2_U5549 P2_U5550 ; P2_U3128
g3671 nand P2_U5554 P2_U3436 P2_U5553 ; P2_U3129
g3672 nand P2_U5556 P2_U3436 P2_U5555 ; P2_U3130
g3673 nand P2_U5558 P2_U3436 P2_U5557 ; P2_U3131
g3674 nand P2_U5560 P2_U3436 P2_U5559 ; P2_U3132
g3675 nand P2_U5562 P2_U3436 P2_U5561 ; P2_U3133
g3676 nand P2_U5564 P2_U3436 P2_U5563 ; P2_U3134
g3677 nand P2_U5566 P2_U3436 P2_U5565 ; P2_U3135
g3678 nand P2_U5568 P2_U3436 P2_U5567 ; P2_U3136
g3679 nand P2_U3436 P2_U5569 P2_U5570 ; P2_U3137
g3680 nand P2_U3436 P2_U5571 P2_U5572 ; P2_U3138
g3681 nand P2_U3436 P2_U5514 P2_U5515 ; P2_U3139
g3682 nand P2_U3436 P2_U5516 P2_U5517 ; P2_U3140
g3683 nand P2_U3436 P2_U5518 P2_U5519 ; P2_U3141
g3684 nand P2_U3436 P2_U5520 P2_U5521 ; P2_U3142
g3685 nand P2_U3436 P2_U5522 P2_U5523 ; P2_U3143
g3686 nand P2_U3436 P2_U5524 P2_U5525 ; P2_U3144
g3687 nand P2_U3436 P2_U5529 P2_U5530 ; P2_U3145
g3688 nand P2_U3436 P2_U5551 P2_U5552 ; P2_U3146
g3689 nand P2_U3436 P2_U5573 P2_U5574 ; P2_U3147
g3690 nand P2_U3436 P2_U5575 P2_U5576 ; P2_U3148
g3691 nand P2_U3436 P2_U5511 P2_U3440 ; P2_U3149
g3692 nand P2_U3905 P2_U3982 ; P2_U3150
g3693 nand P2_U3903 P2_U5446 ; P2_U3151
g3694 not P2_STATE_REG_SCAN_IN ; P2_U3152
g3695 nand P2_U5463 P2_U5462 ; P2_U3153
g3696 nand P2_U5465 P2_U5464 ; P2_U3154
g3697 nand P2_U5469 P2_U5468 ; P2_U3155
g3698 nand P2_U5471 P2_U5470 ; P2_U3156
g3699 nand P2_U5473 P2_U5472 ; P2_U3157
g3700 nand P2_U5475 P2_U5474 ; P2_U3158
g3701 nand P2_U5477 P2_U5476 ; P2_U3159
g3702 nand P2_U5479 P2_U5478 ; P2_U3160
g3703 nand P2_U5481 P2_U5480 ; P2_U3161
g3704 nand P2_U5483 P2_U5482 ; P2_U3162
g3705 nand P2_U5485 P2_U5484 ; P2_U3163
g3706 nand P2_U5487 P2_U5486 ; P2_U3164
g3707 nand P2_U5490 P2_U5489 ; P2_U3165
g3708 nand P2_U5492 P2_U5491 ; P2_U3166
g3709 nand P2_U5494 P2_U5493 ; P2_U3167
g3710 nand P2_U5496 P2_U5495 ; P2_U3168
g3711 nand P2_U5498 P2_U5497 ; P2_U3169
g3712 nand P2_U5500 P2_U5499 ; P2_U3170
g3713 nand P2_U5502 P2_U5501 ; P2_U3171
g3714 nand P2_U5504 P2_U5503 ; P2_U3172
g3715 nand P2_U5506 P2_U5505 ; P2_U3173
g3716 nand P2_U5508 P2_U5507 ; P2_U3174
g3717 nand P2_U5451 P2_U5450 ; P2_U3175
g3718 nand P2_U5453 P2_U5452 ; P2_U3176
g3719 nand P2_U5455 P2_U5454 ; P2_U3177
g3720 nand P2_U5457 P2_U5456 ; P2_U3178
g3721 nand P2_U5459 P2_U5458 ; P2_U3179
g3722 nand P2_U5461 P2_U5460 ; P2_U3180
g3723 nand P2_U5467 P2_U5466 ; P2_U3181
g3724 and P2_U5683 P2_U5679 ; P2_U3182
g3725 and P2_U5682 P2_U5680 ; P2_U3183
g3726 and P2_U5684 P2_U5681 ; P2_U3184
g3727 and P2_U5448 P2_U3054 ; P2_U3185
g3728 and P2_U5448 P2_U3053 ; P2_U3186
g3729 and P2_U5448 P2_U3057 ; P2_U3187
g3730 and P2_U5448 P2_U3058 ; P2_U3188
g3731 and P2_U5448 P2_U3065 ; P2_U3189
g3732 and P2_U5448 P2_U3066 ; P2_U3190
g3733 and P2_U5448 P2_U3061 ; P2_U3191
g3734 and P2_U5448 P2_U3075 ; P2_U3192
g3735 and P2_U5448 P2_U3076 ; P2_U3193
g3736 and P2_U5448 P2_U3081 ; P2_U3194
g3737 and P2_U5448 P2_U3082 ; P2_U3195
g3738 and P2_U5448 P2_U3069 ; P2_U3196
g3739 and P2_U5448 P2_U3073 ; P2_U3197
g3740 and P2_U5448 P2_U3074 ; P2_U3198
g3741 and P2_U5448 P2_U3079 ; P2_U3199
g3742 and P2_U5448 P2_U3080 ; P2_U3200
g3743 and P2_U5448 P2_U3072 ; P2_U3201
g3744 and P2_U5448 P2_U3063 ; P2_U3202
g3745 and P2_U5448 P2_U3062 ; P2_U3203
g3746 and P2_U5448 P2_U3083 ; P2_U3204
g3747 and P2_U5448 P2_U3084 ; P2_U3205
g3748 and P2_U5448 P2_U3070 ; P2_U3206
g3749 and P2_U5448 P2_U3071 ; P2_U3207
g3750 and P2_U5448 P2_U3067 ; P2_U3208
g3751 and P2_U5448 P2_U3060 ; P2_U3209
g3752 and P2_U5448 P2_U3064 ; P2_U3210
g3753 and P2_U5448 P2_U3068 ; P2_U3211
g3754 and P2_U5448 P2_U3078 ; P2_U3212
g3755 and P2_U5448 P2_U3077 ; P2_U3213
g3756 nand P2_U6270 P2_U6269 P2_U3370 ; P2_U3214
g3757 nand P2_U5442 P2_U5441 P2_U5445 P2_U5443 P2_U5444 ; P2_U3215
g3758 nand P2_U5433 P2_U5434 P2_U5436 P2_U5432 P2_U5435 ; P2_U3216
g3759 nand P2_U5424 P2_U5423 P2_U5427 P2_U5425 P2_U5426 ; P2_U3217
g3760 nand P2_U5415 P2_U5416 P2_U5418 P2_U5414 P2_U5417 ; P2_U3218
g3761 nand P2_U5406 P2_U5405 P2_U5409 P2_U5407 P2_U5408 ; P2_U3219
g3762 nand P2_U3901 P2_U5397 P2_U5398 ; P2_U3220
g3763 nand P2_U5388 P2_U5389 P2_U3900 P2_U5390 ; P2_U3221
g3764 nand P2_U5379 P2_U5380 P2_U5382 P2_U5378 P2_U5381 ; P2_U3222
g3765 nand P2_U5370 P2_U5369 P2_U5373 P2_U5371 P2_U5372 ; P2_U3223
g3766 nand P2_U3898 P2_U5361 P2_U5362 ; P2_U3224
g3767 nand P2_U5352 P2_U5353 P2_U5355 P2_U5351 P2_U5354 ; P2_U3225
g3768 nand P2_U5343 P2_U5342 P2_U5346 P2_U5344 P2_U5345 ; P2_U3226
g3769 nand P2_U5334 P2_U5335 P2_U5337 P2_U5333 P2_U5336 ; P2_U3227
g3770 nand P2_U5325 P2_U5324 P2_U5328 P2_U5326 P2_U5327 ; P2_U3228
g3771 nand P2_U5316 P2_U5315 P2_U5317 P2_U3897 ; P2_U3229
g3772 nand P2_U5307 P2_U5306 P2_U5310 P2_U5308 P2_U5309 ; P2_U3230
g3773 nand P2_U5298 P2_U5299 P2_U5301 P2_U5297 P2_U5300 ; P2_U3231
g3774 nand P2_U5289 P2_U5288 P2_U3896 P2_U5290 ; P2_U3232
g3775 nand P2_U5280 P2_U5279 P2_U5283 P2_U5281 P2_U5282 ; P2_U3233
g3776 nand P2_U3895 P2_U5272 P2_U3894 ; P2_U3234
g3777 nand P2_U5263 P2_U5264 P2_U5266 P2_U5262 P2_U5265 ; P2_U3235
g3778 nand P2_U5254 P2_U5253 P2_U5257 P2_U5255 P2_U5256 ; P2_U3236
g3779 nand P2_U5245 P2_U5246 P2_U5248 P2_U5244 P2_U5247 ; P2_U3237
g3780 nand P2_U5236 P2_U5235 P2_U5239 P2_U5237 P2_U5238 ; P2_U3238
g3781 nand P2_U3891 P2_U5227 P2_U5228 ; P2_U3239
g3782 nand P2_U5218 P2_U5217 P2_U5221 P2_U5219 P2_U5220 ; P2_U3240
g3783 nand P2_U5209 P2_U5208 P2_U5212 P2_U5210 P2_U5211 ; P2_U3241
g3784 nand P2_U5200 P2_U5201 P2_U5203 P2_U5199 P2_U5202 ; P2_U3242
g3785 nand P2_U5187 P2_U5186 P2_U5190 P2_U5188 P2_U5189 ; P2_U3243
g3786 and P2_U5671 P2_U5174 ; P2_U3244
g3787 nand P2_U3872 P2_U3871 ; P2_U3245
g3788 nand P2_U3868 P2_U3867 ; P2_U3246
g3789 nand P2_U3865 P2_U3864 ; P2_U3247
g3790 nand P2_U3862 P2_U3861 ; P2_U3248
g3791 nand P2_U3859 P2_U3858 ; P2_U3249
g3792 nand P2_U3856 P2_U3855 ; P2_U3250
g3793 nand P2_U3853 P2_U3852 ; P2_U3251
g3794 nand P2_U3850 P2_U3849 ; P2_U3252
g3795 nand P2_U3847 P2_U3846 ; P2_U3253
g3796 nand P2_U3843 P2_U3844 P2_U3842 ; P2_U3254
g3797 nand P2_U3840 P2_U3841 P2_U3839 ; P2_U3255
g3798 nand P2_U3837 P2_U3838 P2_U3836 ; P2_U3256
g3799 nand P2_U3834 P2_U3835 P2_U3833 ; P2_U3257
g3800 nand P2_U3831 P2_U3832 P2_U3830 ; P2_U3258
g3801 nand P2_U3828 P2_U3829 P2_U3827 ; P2_U3259
g3802 nand P2_U3825 P2_U3826 P2_U3824 ; P2_U3260
g3803 nand P2_U3822 P2_U3823 P2_U3821 ; P2_U3261
g3804 nand P2_U3819 P2_U3820 P2_U3818 ; P2_U3262
g3805 nand P2_U3816 P2_U3817 P2_U3815 ; P2_U3263
g3806 nand P2_U3813 P2_U3814 P2_U3812 ; P2_U3264
g3807 nand P2_U3944 P2_U4865 P2_U4866 ; P2_U3265
g3808 nand P2_U3943 P2_U4863 P2_U4864 ; P2_U3266
g3809 nand P2_U4860 P2_U4861 P2_U4862 P2_U4859 P2_U3941 ; P2_U3267
g3810 nand P2_U3808 P2_U3809 P2_U4855 P2_U3940 ; P2_U3268
g3811 nand P2_U3806 P2_U3807 P2_U4850 P2_U3939 ; P2_U3269
g3812 nand P2_U3804 P2_U3805 P2_U4845 P2_U3938 ; P2_U3270
g3813 nand P2_U3802 P2_U3803 P2_U4840 P2_U3937 ; P2_U3271
g3814 nand P2_U3800 P2_U3801 P2_U4835 P2_U3936 ; P2_U3272
g3815 nand P2_U3798 P2_U3799 P2_U4830 P2_U3935 ; P2_U3273
g3816 nand P2_U3796 P2_U3797 P2_U4825 P2_U3934 ; P2_U3274
g3817 nand P2_U3794 P2_U3795 P2_U4820 P2_U3933 ; P2_U3275
g3818 nand P2_U3792 P2_U3793 P2_U4815 P2_U3932 ; P2_U3276
g3819 nand P2_U3790 P2_U3791 P2_U4810 P2_U3931 ; P2_U3277
g3820 nand P2_U3788 P2_U3789 P2_U4805 P2_U3930 ; P2_U3278
g3821 nand P2_U3786 P2_U3787 P2_U4800 P2_U3929 ; P2_U3279
g3822 nand P2_U3784 P2_U3785 P2_U4795 P2_U3928 ; P2_U3280
g3823 nand P2_U3782 P2_U3783 P2_U4790 P2_U3927 ; P2_U3281
g3824 nand P2_U3780 P2_U3781 P2_U4785 P2_U3926 ; P2_U3282
g3825 nand P2_U3778 P2_U3779 P2_U4780 P2_U3925 ; P2_U3283
g3826 nand P2_U3776 P2_U3777 P2_U4775 P2_U3924 ; P2_U3284
g3827 nand P2_U3775 P2_U3774 P2_U3923 ; P2_U3285
g3828 nand P2_U3772 P2_U3773 P2_U4765 P2_U3922 ; P2_U3286
g3829 nand P2_U3771 P2_U3770 P2_U3921 ; P2_U3287
g3830 nand P2_U3769 P2_U3768 P2_U3920 ; P2_U3288
g3831 nand P2_U3767 P2_U3766 P2_U3919 ; P2_U3289
g3832 nand P2_U3765 P2_U3764 P2_U3918 ; P2_U3290
g3833 nand P2_U3763 P2_U3762 P2_U3917 ; P2_U3291
g3834 nand P2_U3761 P2_U3760 ; P2_U3292
g3835 nand P2_U3759 P2_U3758 ; P2_U3293
g3836 nand P2_U3757 P2_U3756 ; P2_U3294
g3837 nand P2_U3755 P2_U3754 ; P2_U3295
g3838 nand P2_U3753 P2_U3752 ; P2_U3296
g3839 and P2_U3908 P2_D_REG_31__SCAN_IN ; P2_U3297
g3840 and P2_U3908 P2_D_REG_30__SCAN_IN ; P2_U3298
g3841 and P2_U3908 P2_D_REG_29__SCAN_IN ; P2_U3299
g3842 and P2_U3908 P2_D_REG_28__SCAN_IN ; P2_U3300
g3843 and P2_U3908 P2_D_REG_27__SCAN_IN ; P2_U3301
g3844 and P2_U3908 P2_D_REG_26__SCAN_IN ; P2_U3302
g3845 and P2_U3908 P2_D_REG_25__SCAN_IN ; P2_U3303
g3846 and P2_U3908 P2_D_REG_24__SCAN_IN ; P2_U3304
g3847 and P2_U3908 P2_D_REG_23__SCAN_IN ; P2_U3305
g3848 and P2_U3908 P2_D_REG_22__SCAN_IN ; P2_U3306
g3849 and P2_U3908 P2_D_REG_21__SCAN_IN ; P2_U3307
g3850 and P2_U3908 P2_D_REG_20__SCAN_IN ; P2_U3308
g3851 and P2_U3908 P2_D_REG_19__SCAN_IN ; P2_U3309
g3852 and P2_U3908 P2_D_REG_18__SCAN_IN ; P2_U3310
g3853 and P2_U3908 P2_D_REG_17__SCAN_IN ; P2_U3311
g3854 and P2_U3908 P2_D_REG_16__SCAN_IN ; P2_U3312
g3855 and P2_U3908 P2_D_REG_15__SCAN_IN ; P2_U3313
g3856 and P2_U3908 P2_D_REG_14__SCAN_IN ; P2_U3314
g3857 and P2_U3908 P2_D_REG_13__SCAN_IN ; P2_U3315
g3858 and P2_U3908 P2_D_REG_12__SCAN_IN ; P2_U3316
g3859 and P2_U3908 P2_D_REG_11__SCAN_IN ; P2_U3317
g3860 and P2_U3908 P2_D_REG_10__SCAN_IN ; P2_U3318
g3861 and P2_U3908 P2_D_REG_9__SCAN_IN ; P2_U3319
g3862 and P2_U3908 P2_D_REG_8__SCAN_IN ; P2_U3320
g3863 and P2_U3908 P2_D_REG_7__SCAN_IN ; P2_U3321
g3864 and P2_U3908 P2_D_REG_6__SCAN_IN ; P2_U3322
g3865 and P2_U3908 P2_D_REG_5__SCAN_IN ; P2_U3323
g3866 and P2_U3908 P2_D_REG_4__SCAN_IN ; P2_U3324
g3867 and P2_U3908 P2_D_REG_3__SCAN_IN ; P2_U3325
g3868 and P2_U3908 P2_D_REG_2__SCAN_IN ; P2_U3326
g3869 nand P2_U4091 P2_U4092 P2_U4090 ; P2_U3327
g3870 nand P2_U4088 P2_U4089 P2_U4087 ; P2_U3328
g3871 nand P2_U4085 P2_U4086 P2_U4084 ; P2_U3329
g3872 nand P2_U4082 P2_U4083 P2_U4081 ; P2_U3330
g3873 nand P2_U4079 P2_U4080 P2_U4078 ; P2_U3331
g3874 nand P2_U4076 P2_U4077 P2_U4075 ; P2_U3332
g3875 nand P2_U4073 P2_U4074 P2_U4072 ; P2_U3333
g3876 nand P2_U4070 P2_U4071 P2_U4069 ; P2_U3334
g3877 nand P2_U4067 P2_U4068 P2_U4066 ; P2_U3335
g3878 nand P2_U4064 P2_U4065 P2_U4063 ; P2_U3336
g3879 nand P2_U4061 P2_U4062 P2_U4060 ; P2_U3337
g3880 nand P2_U4058 P2_U4059 P2_U4057 ; P2_U3338
g3881 nand P2_U4055 P2_U4056 P2_U4054 ; P2_U3339
g3882 nand P2_U4052 P2_U4053 P2_U4051 ; P2_U3340
g3883 nand P2_U4049 P2_U4050 P2_U4048 ; P2_U3341
g3884 nand P2_U4046 P2_U4047 P2_U4045 ; P2_U3342
g3885 nand P2_U4043 P2_U4044 P2_U4042 ; P2_U3343
g3886 nand P2_U4040 P2_U4041 P2_U4039 ; P2_U3344
g3887 nand P2_U4037 P2_U4038 P2_U4036 ; P2_U3345
g3888 nand P2_U4034 P2_U4035 P2_U4033 ; P2_U3346
g3889 nand P2_U4031 P2_U4032 P2_U4030 ; P2_U3347
g3890 nand P2_U4028 P2_U4029 P2_U4027 ; P2_U3348
g3891 nand P2_U4025 P2_U4026 P2_U4024 ; P2_U3349
g3892 nand P2_U4022 P2_U4023 P2_U4021 ; P2_U3350
g3893 nand P2_U4019 P2_U4020 P2_U4018 ; P2_U3351
g3894 nand P2_U4016 P2_U4017 P2_U4015 ; P2_U3352
g3895 nand P2_U4013 P2_U4014 P2_U4012 ; P2_U3353
g3896 nand P2_U4010 P2_U4011 P2_U4009 ; P2_U3354
g3897 nand P2_U4007 P2_U4008 P2_U4006 ; P2_U3355
g3898 nand P2_U4004 P2_U4005 P2_U4003 ; P2_U3356
g3899 nand P2_U4001 P2_U4002 P2_U4000 ; P2_U3357
g3900 nand P2_U3998 P2_U3999 P2_U3997 ; P2_U3358
g3901 nand P2_U3907 P2_STATE_REG_SCAN_IN ; P2_U3359
g3902 not P2_B_REG_SCAN_IN ; P2_U3360
g3903 nand P2_U3435 P2_U5692 ; P2_U3361
g3904 nand P2_U3435 P2_U4093 ; P2_U3362
g3905 nand P2_U3050 P2_U3441 ; P2_U3363
g3906 nand P2_U5711 P2_U3439 P2_U3440 ; P2_U3364
g3907 nand P2_U5714 P2_U5711 ; P2_U3365
g3908 nand P2_U3994 P2_U3441 ; P2_U3366
g3909 nand P2_U3961 P2_U5717 ; P2_U3367
g3910 nand P2_U5708 P2_U5711 ; P2_U3368
g3911 nand P2_U3951 P2_U3440 ; P2_U3369
g3912 nand P2_U5708 P2_U5717 ; P2_U3370
g3913 nand P2_U3440 P2_U3441 ; P2_U3371
g3914 nand P2_U5711 P2_U3439 P2_U5717 ; P2_U3372
g3915 nand P2_U4138 P2_U4137 P2_U4139 P2_U3617 P2_U3616 ; P2_U3373
g3916 nand P2_U4153 P2_U4152 P2_U3632 P2_U3634 ; P2_U3374
g3917 nand P2_U4172 P2_U4171 P2_U3636 P2_U3638 ; P2_U3375
g3918 nand P2_U4191 P2_U4190 P2_U3640 P2_U3642 ; P2_U3376
g3919 nand P2_U4210 P2_U4209 P2_U3644 P2_U3646 ; P2_U3377
g3920 nand P2_U4229 P2_U4228 P2_U3648 P2_U3650 ; P2_U3378
g3921 nand P2_U4248 P2_U4247 P2_U3652 P2_U3654 ; P2_U3379
g3922 nand P2_U4267 P2_U4266 P2_U3656 P2_U3658 ; P2_U3380
g3923 nand P2_U4286 P2_U4285 P2_U3660 P2_U3662 ; P2_U3381
g3924 nand P2_U4305 P2_U4304 P2_U3664 P2_U3666 ; P2_U3382
g3925 nand P2_U4324 P2_U4323 P2_U3668 P2_U3670 ; P2_U3383
g3926 nand P2_U4343 P2_U4342 P2_U3672 P2_U3674 ; P2_U3384
g3927 nand P2_U4362 P2_U4361 P2_U3676 P2_U3678 ; P2_U3385
g3928 nand P2_U4381 P2_U4380 P2_U3680 P2_U3682 ; P2_U3386
g3929 nand P2_U4400 P2_U4399 P2_U3684 P2_U3686 ; P2_U3387
g3930 nand P2_U4419 P2_U4418 P2_U3688 P2_U3690 ; P2_U3388
g3931 nand P2_U4438 P2_U4437 P2_U3692 P2_U3694 ; P2_U3389
g3932 nand P2_U4457 P2_U4456 P2_U3696 P2_U3698 ; P2_U3390
g3933 nand P2_U4476 P2_U4475 P2_U3700 P2_U3702 ; P2_U3391
g3934 nand P2_U4495 P2_U4494 P2_U3704 P2_U3706 ; P2_U3392
g3935 nand U44 P2_U3909 ; P2_U3393
g3936 nand P2_U4514 P2_U4513 P2_U3708 P2_U3710 ; P2_U3394
g3937 nand U43 P2_U3909 ; P2_U3395
g3938 nand P2_U4533 P2_U4532 P2_U3712 P2_U3714 ; P2_U3396
g3939 nand U42 P2_U3909 ; P2_U3397
g3940 nand P2_U4552 P2_U4551 P2_U3716 P2_U3718 ; P2_U3398
g3941 nand U41 P2_U3909 ; P2_U3399
g3942 nand P2_U4571 P2_U4570 P2_U3720 P2_U3722 ; P2_U3400
g3943 nand U40 P2_U3909 ; P2_U3401
g3944 nand P2_U4590 P2_U4589 P2_U3724 P2_U3726 ; P2_U3402
g3945 nand U39 P2_U3909 ; P2_U3403
g3946 nand P2_U4609 P2_U4608 P2_U3728 P2_U3730 ; P2_U3404
g3947 nand U38 P2_U3909 ; P2_U3405
g3948 nand P2_U4628 P2_U4627 P2_U3732 P2_U3734 ; P2_U3406
g3949 nand U37 P2_U3909 ; P2_U3407
g3950 nand P2_U4647 P2_U4646 P2_U3736 P2_U3738 ; P2_U3408
g3951 nand U36 P2_U3909 ; P2_U3409
g3952 nand P2_U4666 P2_U4665 P2_U4667 P2_U4668 P2_U3741 ; P2_U3410
g3953 nand U35 P2_U3909 ; P2_U3411
g3954 nand P2_U4686 P2_U4685 P2_U4687 P2_U3744 P2_U3746 ; P2_U3412
g3955 nand U33 P2_U3909 ; P2_U3413
g3956 nand U32 P2_U3909 ; P2_U3414
g3957 nand P2_U3445 P2_U5717 ; P2_U3415
g3958 nand P2_U5674 P2_U5714 ; P2_U3416
g3959 nand P2_U3027 P2_U4711 ; P2_U3417
g3960 nand P2_U3960 P2_U5708 ; P2_U3418
g3961 nand P2_U3031 P2_U5711 ; P2_U3419
g3962 nand P2_U3434 P2_U3435 P2_U3433 ; P2_U3420
g3963 nand P2_U3371 P2_U3909 ; P2_U3421
g3964 nand P2_U3981 P2_U5701 ; P2_U3422
g3965 nand P2_U3995 P2_STATE_REG_SCAN_IN ; P2_U3423
g3966 nand P2_U3810 P2_U3052 ; P2_U3424
g3967 nand P2_U3017 P2_U3022 ; P2_U3425
g3968 nand P2_U3027 P2_U4713 ; P2_U3426
g3969 nand P2_U3887 P2_U3020 ; P2_U3427
g3970 nand P2_U5708 P2_U3440 ; P2_U3428
g3971 nand P2_U3017 P2_U3027 ; P2_U3429
g3972 nand P2_U5184 P2_U3889 ; P2_U3430
g3973 nand P2_U3951 P2_U3369 ; P2_U3431
g3974 nand P2_U3993 P2_U3445 ; P2_U3432
g3975 nand P2_U5688 P2_U5687 ; P2_U3433
g3976 nand P2_U5691 P2_U5690 ; P2_U3434
g3977 nand P2_U5694 P2_U5693 ; P2_U3435
g3978 nand P2_U5700 P2_U5699 ; P2_U3436
g3979 nand P2_U5703 P2_U5702 ; P2_U3437
g3980 nand P2_U5705 P2_U5704 ; P2_U3438
g3981 nand P2_U5713 P2_U5712 ; P2_U3439
g3982 nand P2_U5716 P2_U5715 ; P2_U3440
g3983 nand P2_U5707 P2_U5706 ; P2_U3441
g3984 nand P2_U5722 P2_U5721 ; P2_U3442
g3985 nand P2_U5719 P2_U5718 ; P2_U3443
g3986 nand P2_U5727 P2_U5726 ; P2_U3444
g3987 nand P2_U5710 P2_U5709 ; P2_U3445
g3988 nand P2_U5730 P2_U5729 ; P2_U3446
g3989 nand P2_U5732 P2_U5731 ; P2_U3447
g3990 nand P2_U5735 P2_U5734 ; P2_U3448
g3991 nand P2_U5743 P2_U5742 ; P2_U3449
g3992 nand P2_U5740 P2_U5739 ; P2_U3450
g3993 nand P2_U5746 P2_U5745 ; P2_U3451
g3994 nand P2_U5750 P2_U5749 ; P2_U3452
g3995 nand P2_U5752 P2_U5751 ; P2_U3453
g3996 nand P2_U5757 P2_U5756 ; P2_U3454
g3997 nand P2_U5759 P2_U5758 ; P2_U3455
g3998 nand P2_U5761 P2_U5760 ; P2_U3456
g3999 nand P2_U5764 P2_U5763 ; P2_U3457
g4000 nand P2_U5766 P2_U5765 ; P2_U3458
g4001 nand P2_U5768 P2_U5767 ; P2_U3459
g4002 nand P2_U5771 P2_U5770 ; P2_U3460
g4003 nand P2_U5773 P2_U5772 ; P2_U3461
g4004 nand P2_U5775 P2_U5774 ; P2_U3462
g4005 nand P2_U5778 P2_U5777 ; P2_U3463
g4006 nand P2_U5780 P2_U5779 ; P2_U3464
g4007 nand P2_U5782 P2_U5781 ; P2_U3465
g4008 nand P2_U5785 P2_U5784 ; P2_U3466
g4009 nand P2_U5787 P2_U5786 ; P2_U3467
g4010 nand P2_U5789 P2_U5788 ; P2_U3468
g4011 nand P2_U5792 P2_U5791 ; P2_U3469
g4012 nand P2_U5794 P2_U5793 ; P2_U3470
g4013 nand P2_U5796 P2_U5795 ; P2_U3471
g4014 nand P2_U5799 P2_U5798 ; P2_U3472
g4015 nand P2_U5801 P2_U5800 ; P2_U3473
g4016 nand P2_U5803 P2_U5802 ; P2_U3474
g4017 nand P2_U5806 P2_U5805 ; P2_U3475
g4018 nand P2_U5808 P2_U5807 ; P2_U3476
g4019 nand P2_U5810 P2_U5809 ; P2_U3477
g4020 nand P2_U5813 P2_U5812 ; P2_U3478
g4021 nand P2_U5815 P2_U5814 ; P2_U3479
g4022 nand P2_U5817 P2_U5816 ; P2_U3480
g4023 nand P2_U5820 P2_U5819 ; P2_U3481
g4024 nand P2_U5822 P2_U5821 ; P2_U3482
g4025 nand P2_U5824 P2_U5823 ; P2_U3483
g4026 nand P2_U5827 P2_U5826 ; P2_U3484
g4027 nand P2_U5829 P2_U5828 ; P2_U3485
g4028 nand P2_U5831 P2_U5830 ; P2_U3486
g4029 nand P2_U5834 P2_U5833 ; P2_U3487
g4030 nand P2_U5836 P2_U5835 ; P2_U3488
g4031 nand P2_U5838 P2_U5837 ; P2_U3489
g4032 nand P2_U5841 P2_U5840 ; P2_U3490
g4033 nand P2_U5843 P2_U5842 ; P2_U3491
g4034 nand P2_U5845 P2_U5844 ; P2_U3492
g4035 nand P2_U5848 P2_U5847 ; P2_U3493
g4036 nand P2_U5850 P2_U5849 ; P2_U3494
g4037 nand P2_U5852 P2_U5851 ; P2_U3495
g4038 nand P2_U5855 P2_U5854 ; P2_U3496
g4039 nand P2_U5857 P2_U5856 ; P2_U3497
g4040 nand P2_U5859 P2_U5858 ; P2_U3498
g4041 nand P2_U5862 P2_U5861 ; P2_U3499
g4042 nand P2_U5864 P2_U5863 ; P2_U3500
g4043 nand P2_U5866 P2_U5865 ; P2_U3501
g4044 nand P2_U5869 P2_U5868 ; P2_U3502
g4045 nand P2_U5871 P2_U5870 ; P2_U3503
g4046 nand P2_U5873 P2_U5872 ; P2_U3504
g4047 nand P2_U5876 P2_U5875 ; P2_U3505
g4048 nand P2_U5878 P2_U5877 ; P2_U3506
g4049 nand P2_U5881 P2_U5880 ; P2_U3507
g4050 nand P2_U5883 P2_U5882 ; P2_U3508
g4051 nand P2_U5885 P2_U5884 ; P2_U3509
g4052 nand P2_U5887 P2_U5886 ; P2_U3510
g4053 nand P2_U5889 P2_U5888 ; P2_U3511
g4054 nand P2_U5891 P2_U5890 ; P2_U3512
g4055 nand P2_U5893 P2_U5892 ; P2_U3513
g4056 nand P2_U5895 P2_U5894 ; P2_U3514
g4057 nand P2_U5897 P2_U5896 ; P2_U3515
g4058 nand P2_U5899 P2_U5898 ; P2_U3516
g4059 nand P2_U5901 P2_U5900 ; P2_U3517
g4060 nand P2_U5903 P2_U5902 ; P2_U3518
g4061 nand P2_U5905 P2_U5904 ; P2_U3519
g4062 nand P2_U5907 P2_U5906 ; P2_U3520
g4063 nand P2_U5909 P2_U5908 ; P2_U3521
g4064 nand P2_U5911 P2_U5910 ; P2_U3522
g4065 nand P2_U5913 P2_U5912 ; P2_U3523
g4066 nand P2_U5915 P2_U5914 ; P2_U3524
g4067 nand P2_U5917 P2_U5916 ; P2_U3525
g4068 nand P2_U5919 P2_U5918 ; P2_U3526
g4069 nand P2_U5921 P2_U5920 ; P2_U3527
g4070 nand P2_U5923 P2_U5922 ; P2_U3528
g4071 nand P2_U5925 P2_U5924 ; P2_U3529
g4072 nand P2_U5927 P2_U5926 ; P2_U3530
g4073 nand P2_U5929 P2_U5928 ; P2_U3531
g4074 nand P2_U5931 P2_U5930 ; P2_U3532
g4075 nand P2_U5933 P2_U5932 ; P2_U3533
g4076 nand P2_U5935 P2_U5934 ; P2_U3534
g4077 nand P2_U5937 P2_U5936 ; P2_U3535
g4078 nand P2_U5939 P2_U5938 ; P2_U3536
g4079 nand P2_U5941 P2_U5940 ; P2_U3537
g4080 nand P2_U5943 P2_U5942 ; P2_U3538
g4081 nand P2_U5945 P2_U5944 ; P2_U3539
g4082 nand P2_U5947 P2_U5946 ; P2_U3540
g4083 nand P2_U5949 P2_U5948 ; P2_U3541
g4084 nand P2_U5951 P2_U5950 ; P2_U3542
g4085 nand P2_U5953 P2_U5952 ; P2_U3543
g4086 nand P2_U5955 P2_U5954 ; P2_U3544
g4087 nand P2_U5957 P2_U5956 ; P2_U3545
g4088 nand P2_U5959 P2_U5958 ; P2_U3546
g4089 nand P2_U5961 P2_U5960 ; P2_U3547
g4090 nand P2_U5963 P2_U5962 ; P2_U3548
g4091 nand P2_U5965 P2_U5964 ; P2_U3549
g4092 nand P2_U5967 P2_U5966 ; P2_U3550
g4093 nand P2_U5969 P2_U5968 ; P2_U3551
g4094 nand P2_U6035 P2_U6034 ; P2_U3552
g4095 nand P2_U6037 P2_U6036 ; P2_U3553
g4096 nand P2_U6039 P2_U6038 ; P2_U3554
g4097 nand P2_U6041 P2_U6040 ; P2_U3555
g4098 nand P2_U6043 P2_U6042 ; P2_U3556
g4099 nand P2_U6045 P2_U6044 ; P2_U3557
g4100 nand P2_U6047 P2_U6046 ; P2_U3558
g4101 nand P2_U6049 P2_U6048 ; P2_U3559
g4102 nand P2_U6051 P2_U6050 ; P2_U3560
g4103 nand P2_U6053 P2_U6052 ; P2_U3561
g4104 nand P2_U6055 P2_U6054 ; P2_U3562
g4105 nand P2_U6057 P2_U6056 ; P2_U3563
g4106 nand P2_U6059 P2_U6058 ; P2_U3564
g4107 nand P2_U6061 P2_U6060 ; P2_U3565
g4108 nand P2_U6063 P2_U6062 ; P2_U3566
g4109 nand P2_U6065 P2_U6064 ; P2_U3567
g4110 nand P2_U6067 P2_U6066 ; P2_U3568
g4111 nand P2_U6069 P2_U6068 ; P2_U3569
g4112 nand P2_U6071 P2_U6070 ; P2_U3570
g4113 nand P2_U6073 P2_U6072 ; P2_U3571
g4114 nand P2_U6075 P2_U6074 ; P2_U3572
g4115 nand P2_U6077 P2_U6076 ; P2_U3573
g4116 nand P2_U6079 P2_U6078 ; P2_U3574
g4117 nand P2_U6081 P2_U6080 ; P2_U3575
g4118 nand P2_U6083 P2_U6082 ; P2_U3576
g4119 nand P2_U6085 P2_U6084 ; P2_U3577
g4120 nand P2_U6087 P2_U6086 ; P2_U3578
g4121 nand P2_U6089 P2_U6088 ; P2_U3579
g4122 nand P2_U6091 P2_U6090 ; P2_U3580
g4123 nand P2_U6093 P2_U6092 ; P2_U3581
g4124 nand P2_U6095 P2_U6094 ; P2_U3582
g4125 nand P2_U6097 P2_U6096 ; P2_U3583
g4126 nand P2_U6203 P2_U6202 ; P2_U3584
g4127 nand P2_U6205 P2_U6204 ; P2_U3585
g4128 nand P2_U6207 P2_U6206 ; P2_U3586
g4129 nand P2_U6209 P2_U6208 ; P2_U3587
g4130 nand P2_U6211 P2_U6210 ; P2_U3588
g4131 nand P2_U6213 P2_U6212 ; P2_U3589
g4132 nand P2_U6215 P2_U6214 ; P2_U3590
g4133 nand P2_U6217 P2_U6216 ; P2_U3591
g4134 nand P2_U6219 P2_U6218 ; P2_U3592
g4135 nand P2_U6221 P2_U6220 ; P2_U3593
g4136 nand P2_U6224 P2_U6223 ; P2_U3594
g4137 nand P2_U6226 P2_U6225 ; P2_U3595
g4138 nand P2_U6228 P2_U6227 ; P2_U3596
g4139 nand P2_U6230 P2_U6229 ; P2_U3597
g4140 nand P2_U6232 P2_U6231 ; P2_U3598
g4141 nand P2_U6234 P2_U6233 ; P2_U3599
g4142 nand P2_U6236 P2_U6235 ; P2_U3600
g4143 nand P2_U6238 P2_U6237 ; P2_U3601
g4144 nand P2_U6240 P2_U6239 ; P2_U3602
g4145 nand P2_U6242 P2_U6241 ; P2_U3603
g4146 nand P2_U6244 P2_U6243 ; P2_U3604
g4147 nand P2_U6247 P2_U6246 ; P2_U3605
g4148 nand P2_U6249 P2_U6248 ; P2_U3606
g4149 nand P2_U6251 P2_U6250 ; P2_U3607
g4150 nand P2_U6253 P2_U6252 ; P2_U3608
g4151 nand P2_U6255 P2_U6254 ; P2_U3609
g4152 nand P2_U6257 P2_U6256 ; P2_U3610
g4153 nand P2_U6259 P2_U6258 ; P2_U3611
g4154 nand P2_U6261 P2_U6260 ; P2_U3612
g4155 nand P2_U6263 P2_U6262 ; P2_U3613
g4156 nand P2_U6265 P2_U6264 ; P2_U3614
g4157 nand P2_U6267 P2_U6266 ; P2_U3615
g4158 and P2_U4134 P2_U4133 ; P2_U3616
g4159 and P2_U4136 P2_U4135 ; P2_U3617
g4160 and P2_U4143 P2_U4141 ; P2_U3618
g4161 and P2_U4144 P2_U4142 P2_U3618 ; P2_U3619
g4162 and P2_U4100 P2_U4099 P2_U4098 P2_U4097 ; P2_U3620
g4163 and P2_U4104 P2_U4103 P2_U4102 P2_U4101 ; P2_U3621
g4164 and P2_U4108 P2_U4107 P2_U4106 P2_U4105 ; P2_U3622
g4165 and P2_U4110 P2_U4109 P2_U4111 ; P2_U3623
g4166 and P2_U3623 P2_U3622 P2_U3621 P2_U3620 ; P2_U3624
g4167 and P2_U4115 P2_U4114 P2_U4113 P2_U4112 ; P2_U3625
g4168 and P2_U4119 P2_U4118 P2_U4117 P2_U4116 ; P2_U3626
g4169 and P2_U4123 P2_U4122 P2_U4121 P2_U4120 ; P2_U3627
g4170 and P2_U4125 P2_U4124 P2_U4126 ; P2_U3628
g4171 and P2_U3628 P2_U3627 P2_U3626 P2_U3625 ; P2_U3629
g4172 and P2_U5741 P2_U4127 ; P2_U3630
g4173 and P2_U5744 P2_U3027 ; P2_U3631
g4174 and P2_U4155 P2_U4154 ; P2_U3632
g4175 and P2_U4157 P2_U4156 ; P2_U3633
g4176 and P2_U4159 P2_U4158 P2_U3633 ; P2_U3634
g4177 and P2_U4162 P2_U4161 P2_U4164 P2_U4163 ; P2_U3635
g4178 and P2_U4174 P2_U4173 ; P2_U3636
g4179 and P2_U4176 P2_U4175 ; P2_U3637
g4180 and P2_U4178 P2_U4177 P2_U3637 ; P2_U3638
g4181 and P2_U4181 P2_U4180 P2_U4183 P2_U4182 ; P2_U3639
g4182 and P2_U4193 P2_U4192 ; P2_U3640
g4183 and P2_U4195 P2_U4194 ; P2_U3641
g4184 and P2_U4197 P2_U4196 P2_U3641 ; P2_U3642
g4185 and P2_U4200 P2_U4199 P2_U4202 P2_U4201 ; P2_U3643
g4186 and P2_U4212 P2_U4211 ; P2_U3644
g4187 and P2_U4214 P2_U4213 ; P2_U3645
g4188 and P2_U4216 P2_U4215 P2_U3645 ; P2_U3646
g4189 and P2_U4219 P2_U4218 P2_U4221 P2_U4220 ; P2_U3647
g4190 and P2_U4231 P2_U4230 ; P2_U3648
g4191 and P2_U4233 P2_U4232 ; P2_U3649
g4192 and P2_U4235 P2_U4234 P2_U3649 ; P2_U3650
g4193 and P2_U4238 P2_U4237 P2_U4240 P2_U4239 ; P2_U3651
g4194 and P2_U4250 P2_U4249 ; P2_U3652
g4195 and P2_U4252 P2_U4251 ; P2_U3653
g4196 and P2_U4254 P2_U4253 P2_U3653 ; P2_U3654
g4197 and P2_U4257 P2_U4256 P2_U4259 P2_U4258 ; P2_U3655
g4198 and P2_U4269 P2_U4268 ; P2_U3656
g4199 and P2_U4271 P2_U4270 ; P2_U3657
g4200 and P2_U4273 P2_U4272 P2_U3657 ; P2_U3658
g4201 and P2_U4276 P2_U4275 P2_U4278 P2_U4277 ; P2_U3659
g4202 and P2_U4288 P2_U4287 ; P2_U3660
g4203 and P2_U4290 P2_U4289 ; P2_U3661
g4204 and P2_U4292 P2_U4291 P2_U3661 ; P2_U3662
g4205 and P2_U4295 P2_U4294 P2_U4297 P2_U4296 ; P2_U3663
g4206 and P2_U4307 P2_U4306 ; P2_U3664
g4207 and P2_U4309 P2_U4308 ; P2_U3665
g4208 and P2_U4311 P2_U4310 P2_U3665 ; P2_U3666
g4209 and P2_U4314 P2_U4313 P2_U4316 P2_U4315 ; P2_U3667
g4210 and P2_U4326 P2_U4325 ; P2_U3668
g4211 and P2_U4328 P2_U4327 ; P2_U3669
g4212 and P2_U4330 P2_U4329 P2_U3669 ; P2_U3670
g4213 and P2_U4333 P2_U4332 P2_U4335 P2_U4334 ; P2_U3671
g4214 and P2_U4345 P2_U4344 ; P2_U3672
g4215 and P2_U4347 P2_U4346 ; P2_U3673
g4216 and P2_U4349 P2_U4348 P2_U3673 ; P2_U3674
g4217 and P2_U4352 P2_U4351 P2_U4354 P2_U4353 ; P2_U3675
g4218 and P2_U4364 P2_U4363 ; P2_U3676
g4219 and P2_U4366 P2_U4365 ; P2_U3677
g4220 and P2_U4368 P2_U4367 P2_U3677 ; P2_U3678
g4221 and P2_U4371 P2_U4370 P2_U4373 P2_U4372 ; P2_U3679
g4222 and P2_U4383 P2_U4382 ; P2_U3680
g4223 and P2_U4385 P2_U4384 ; P2_U3681
g4224 and P2_U4387 P2_U4386 P2_U3681 ; P2_U3682
g4225 and P2_U4390 P2_U4389 P2_U4392 P2_U4391 ; P2_U3683
g4226 and P2_U4402 P2_U4401 ; P2_U3684
g4227 and P2_U4404 P2_U4403 ; P2_U3685
g4228 and P2_U4406 P2_U4405 P2_U3685 ; P2_U3686
g4229 and P2_U4409 P2_U4408 P2_U4411 P2_U4410 ; P2_U3687
g4230 and P2_U4421 P2_U4420 ; P2_U3688
g4231 and P2_U4423 P2_U4422 ; P2_U3689
g4232 and P2_U4425 P2_U4424 P2_U3689 ; P2_U3690
g4233 and P2_U4428 P2_U4427 P2_U4430 P2_U4429 ; P2_U3691
g4234 and P2_U4440 P2_U4439 ; P2_U3692
g4235 and P2_U4442 P2_U4441 ; P2_U3693
g4236 and P2_U4444 P2_U4443 P2_U3693 ; P2_U3694
g4237 and P2_U4447 P2_U4446 P2_U4449 P2_U4448 ; P2_U3695
g4238 and P2_U4459 P2_U4458 ; P2_U3696
g4239 and P2_U4461 P2_U4460 ; P2_U3697
g4240 and P2_U4463 P2_U4462 P2_U3697 ; P2_U3698
g4241 and P2_U4466 P2_U4465 P2_U4468 P2_U4467 ; P2_U3699
g4242 and P2_U4478 P2_U4477 ; P2_U3700
g4243 and P2_U4480 P2_U4479 ; P2_U3701
g4244 and P2_U4482 P2_U4481 P2_U3701 ; P2_U3702
g4245 and P2_U4485 P2_U4484 P2_U4487 P2_U4486 ; P2_U3703
g4246 and P2_U4497 P2_U4496 ; P2_U3704
g4247 and P2_U4499 P2_U4498 ; P2_U3705
g4248 and P2_U4501 P2_U4500 P2_U3705 ; P2_U3706
g4249 and P2_U4504 P2_U4503 P2_U4506 P2_U4505 ; P2_U3707
g4250 and P2_U4516 P2_U4515 ; P2_U3708
g4251 and P2_U4518 P2_U4517 ; P2_U3709
g4252 and P2_U4520 P2_U4519 P2_U3709 ; P2_U3710
g4253 and P2_U4523 P2_U4522 P2_U4525 P2_U4524 ; P2_U3711
g4254 and P2_U4535 P2_U4534 ; P2_U3712
g4255 and P2_U4537 P2_U4536 ; P2_U3713
g4256 and P2_U4539 P2_U4538 P2_U3713 ; P2_U3714
g4257 and P2_U4542 P2_U4541 P2_U4544 P2_U4543 ; P2_U3715
g4258 and P2_U4554 P2_U4553 ; P2_U3716
g4259 and P2_U4556 P2_U4555 ; P2_U3717
g4260 and P2_U4558 P2_U4557 P2_U3717 ; P2_U3718
g4261 and P2_U4561 P2_U4560 P2_U4563 P2_U4562 ; P2_U3719
g4262 and P2_U4573 P2_U4572 ; P2_U3720
g4263 and P2_U4575 P2_U4574 ; P2_U3721
g4264 and P2_U4577 P2_U4576 P2_U3721 ; P2_U3722
g4265 and P2_U4580 P2_U4579 P2_U4582 P2_U4581 ; P2_U3723
g4266 and P2_U4592 P2_U4591 ; P2_U3724
g4267 and P2_U4594 P2_U4593 ; P2_U3725
g4268 and P2_U4596 P2_U4595 P2_U3725 ; P2_U3726
g4269 and P2_U4599 P2_U4598 P2_U4601 P2_U4600 ; P2_U3727
g4270 and P2_U4611 P2_U4610 ; P2_U3728
g4271 and P2_U4613 P2_U4612 ; P2_U3729
g4272 and P2_U4615 P2_U4614 P2_U3729 ; P2_U3730
g4273 and P2_U4618 P2_U4617 P2_U4620 P2_U4619 ; P2_U3731
g4274 and P2_U4630 P2_U4629 ; P2_U3732
g4275 and P2_U4632 P2_U4631 ; P2_U3733
g4276 and P2_U4634 P2_U4633 P2_U3733 ; P2_U3734
g4277 and P2_U4637 P2_U4636 P2_U4639 P2_U4638 ; P2_U3735
g4278 and P2_U4649 P2_U4648 ; P2_U3736
g4279 and P2_U4651 P2_U4650 ; P2_U3737
g4280 and P2_U4653 P2_U4652 P2_U3737 ; P2_U3738
g4281 and P2_U4656 P2_U4655 P2_U4658 P2_U4657 ; P2_U3739
g4282 and P2_U4670 P2_U4669 ; P2_U3740
g4283 and P2_U4672 P2_U4671 P2_U3740 ; P2_U3741
g4284 and P2_U4675 P2_U4674 P2_U4677 P2_U4676 ; P2_U3742
g4285 and P2_U4684 P2_U3982 ; P2_U3743
g4286 and P2_U4689 P2_U4688 ; P2_U3744
g4287 and P2_U4691 P2_U4690 ; P2_U3745
g4288 and P2_U4693 P2_U4692 P2_U3745 ; P2_U3746
g4289 and P2_U4697 P2_U4695 P2_U4696 ; P2_U3747
g4290 and P2_U3982 P2_U4684 ; P2_U3748
g4291 and P2_U3027 P2_U3449 ; P2_U3749
g4292 and P2_U5744 P2_U3051 P2_U3450 ; P2_U3750
g4293 and P2_U3445 P2_U5714 P2_U3440 ; P2_U3751
g4294 and P2_U4715 P2_U4714 P2_U4716 ; P2_U3752
g4295 and P2_U4718 P2_U4717 P2_U3912 ; P2_U3753
g4296 and P2_U4720 P2_U4719 P2_U4721 ; P2_U3754
g4297 and P2_U4723 P2_U4722 P2_U3913 ; P2_U3755
g4298 and P2_U4725 P2_U4724 P2_U4726 ; P2_U3756
g4299 and P2_U4728 P2_U4727 P2_U3914 ; P2_U3757
g4300 and P2_U4730 P2_U4729 P2_U4731 ; P2_U3758
g4301 and P2_U4733 P2_U4732 P2_U3915 ; P2_U3759
g4302 and P2_U4735 P2_U4734 P2_U4736 ; P2_U3760
g4303 and P2_U4738 P2_U4737 P2_U3916 ; P2_U3761
g4304 and P2_U4740 P2_U4739 P2_U4741 ; P2_U3762
g4305 and P2_U4743 P2_U4742 ; P2_U3763
g4306 and P2_U4745 P2_U4744 P2_U4746 ; P2_U3764
g4307 and P2_U4748 P2_U4747 ; P2_U3765
g4308 and P2_U4750 P2_U4749 P2_U4751 ; P2_U3766
g4309 and P2_U4753 P2_U4752 ; P2_U3767
g4310 and P2_U4755 P2_U4754 P2_U4756 ; P2_U3768
g4311 and P2_U4758 P2_U4757 ; P2_U3769
g4312 and P2_U4760 P2_U4759 P2_U4761 ; P2_U3770
g4313 and P2_U4763 P2_U4762 ; P2_U3771
g4314 and P2_U4766 P2_U4764 ; P2_U3772
g4315 and P2_U4768 P2_U4767 ; P2_U3773
g4316 and P2_U4770 P2_U4769 P2_U4771 ; P2_U3774
g4317 and P2_U4773 P2_U4772 ; P2_U3775
g4318 and P2_U4776 P2_U4774 ; P2_U3776
g4319 and P2_U4778 P2_U4777 ; P2_U3777
g4320 and P2_U4781 P2_U4779 ; P2_U3778
g4321 and P2_U4783 P2_U4782 ; P2_U3779
g4322 and P2_U4786 P2_U4784 ; P2_U3780
g4323 and P2_U4788 P2_U4787 ; P2_U3781
g4324 and P2_U4791 P2_U4789 ; P2_U3782
g4325 and P2_U4793 P2_U4792 ; P2_U3783
g4326 and P2_U4796 P2_U4794 ; P2_U3784
g4327 and P2_U4798 P2_U4797 ; P2_U3785
g4328 and P2_U4801 P2_U4799 ; P2_U3786
g4329 and P2_U4803 P2_U4802 ; P2_U3787
g4330 and P2_U4806 P2_U4804 ; P2_U3788
g4331 and P2_U4808 P2_U4807 ; P2_U3789
g4332 and P2_U4811 P2_U4809 ; P2_U3790
g4333 and P2_U4813 P2_U4812 ; P2_U3791
g4334 and P2_U4816 P2_U4814 ; P2_U3792
g4335 and P2_U4818 P2_U4817 ; P2_U3793
g4336 and P2_U4821 P2_U4819 ; P2_U3794
g4337 and P2_U4823 P2_U4822 ; P2_U3795
g4338 and P2_U4826 P2_U4824 ; P2_U3796
g4339 and P2_U4828 P2_U4827 ; P2_U3797
g4340 and P2_U4831 P2_U4829 ; P2_U3798
g4341 and P2_U4833 P2_U4832 ; P2_U3799
g4342 and P2_U4836 P2_U4834 ; P2_U3800
g4343 and P2_U4838 P2_U4837 ; P2_U3801
g4344 and P2_U4841 P2_U4839 ; P2_U3802
g4345 and P2_U4843 P2_U4842 ; P2_U3803
g4346 and P2_U4846 P2_U4844 ; P2_U3804
g4347 and P2_U4848 P2_U4847 ; P2_U3805
g4348 and P2_U4851 P2_U4849 ; P2_U3806
g4349 and P2_U4853 P2_U4852 ; P2_U3807
g4350 and P2_U4856 P2_U4854 ; P2_U3808
g4351 and P2_U4858 P2_U4857 ; P2_U3809
g4352 and P2_U5686 P2_U3421 ; P2_U3810
g4353 and P2_U3436 P2_STATE_REG_SCAN_IN ; P2_U3811
g4354 and P2_U4877 P2_U4876 ; P2_U3812
g4355 and P2_U4879 P2_U4878 ; P2_U3813
g4356 and P2_U4882 P2_U4880 P2_U4881 ; P2_U3814
g4357 and P2_U4892 P2_U4891 ; P2_U3815
g4358 and P2_U4894 P2_U4893 ; P2_U3816
g4359 and P2_U4897 P2_U4895 P2_U4896 ; P2_U3817
g4360 and P2_U4907 P2_U4906 ; P2_U3818
g4361 and P2_U4909 P2_U4908 ; P2_U3819
g4362 and P2_U4912 P2_U4910 P2_U4911 ; P2_U3820
g4363 and P2_U4922 P2_U4921 ; P2_U3821
g4364 and P2_U4924 P2_U4923 ; P2_U3822
g4365 and P2_U4927 P2_U4925 P2_U4926 ; P2_U3823
g4366 and P2_U4937 P2_U4936 ; P2_U3824
g4367 and P2_U4939 P2_U4938 ; P2_U3825
g4368 and P2_U4942 P2_U4940 P2_U4941 ; P2_U3826
g4369 and P2_U4952 P2_U4951 ; P2_U3827
g4370 and P2_U4954 P2_U4953 ; P2_U3828
g4371 and P2_U4957 P2_U4955 P2_U4956 ; P2_U3829
g4372 and P2_U4967 P2_U4966 ; P2_U3830
g4373 and P2_U4969 P2_U4968 ; P2_U3831
g4374 and P2_U4972 P2_U4970 P2_U4971 ; P2_U3832
g4375 and P2_U4982 P2_U4981 ; P2_U3833
g4376 and P2_U4984 P2_U4983 ; P2_U3834
g4377 and P2_U4987 P2_U4985 P2_U4986 ; P2_U3835
g4378 and P2_U4997 P2_U4996 ; P2_U3836
g4379 and P2_U4999 P2_U4998 ; P2_U3837
g4380 and P2_U5002 P2_U5000 P2_U5001 ; P2_U3838
g4381 and P2_U5012 P2_U5011 ; P2_U3839
g4382 and P2_U5014 P2_U5013 ; P2_U3840
g4383 and P2_U5017 P2_U5015 P2_U5016 ; P2_U3841
g4384 and P2_U5027 P2_U5026 ; P2_U3842
g4385 and P2_U5029 P2_U5028 ; P2_U3843
g4386 and P2_U5032 P2_U5030 P2_U5031 ; P2_U3844
g4387 and P2_U5042 P2_U5041 ; P2_U3845
g4388 and P2_U5044 P2_U5043 P2_U3845 ; P2_U3846
g4389 and P2_U5046 P2_U5045 P2_U5047 ; P2_U3847
g4390 and P2_U5057 P2_U5056 ; P2_U3848
g4391 and P2_U5059 P2_U5058 P2_U3848 ; P2_U3849
g4392 and P2_U5061 P2_U5060 P2_U5062 ; P2_U3850
g4393 and P2_U5072 P2_U5071 ; P2_U3851
g4394 and P2_U5074 P2_U5073 P2_U3851 ; P2_U3852
g4395 and P2_U5076 P2_U5075 P2_U5077 ; P2_U3853
g4396 and P2_U5087 P2_U5086 ; P2_U3854
g4397 and P2_U5089 P2_U5088 P2_U3854 ; P2_U3855
g4398 and P2_U5091 P2_U5090 P2_U5092 ; P2_U3856
g4399 and P2_U5102 P2_U5101 ; P2_U3857
g4400 and P2_U5104 P2_U5103 P2_U3857 ; P2_U3858
g4401 and P2_U5106 P2_U5105 P2_U5107 ; P2_U3859
g4402 and P2_U5117 P2_U5116 ; P2_U3860
g4403 and P2_U5119 P2_U5118 P2_U3860 ; P2_U3861
g4404 and P2_U5121 P2_U5120 P2_U5122 ; P2_U3862
g4405 and P2_U5132 P2_U5131 ; P2_U3863
g4406 and P2_U5134 P2_U5133 P2_U3863 ; P2_U3864
g4407 and P2_U5136 P2_U5135 P2_U5137 ; P2_U3865
g4408 and P2_U5147 P2_U5146 ; P2_U3866
g4409 and P2_U5149 P2_U5148 P2_U3866 ; P2_U3867
g4410 and P2_U5151 P2_U5150 P2_U5152 ; P2_U3868
g4411 and P2_U5154 P2_U5155 ; P2_U3869
g4412 and P2_U5162 P2_U5161 ; P2_U3870
g4413 and P2_U5164 P2_U5163 P2_U3870 ; P2_U3871
g4414 and P2_U5166 P2_U5165 P2_U5167 ; P2_U3872
g4415 and P2_U6157 P2_U6154 P2_U6160 ; P2_U3873
g4416 and P2_U3873 P2_U3875 ; P2_U3874
g4417 and P2_U6151 P2_U6148 P2_U6145 P2_U6142 ; P2_U3875
g4418 and P2_U6169 P2_U6166 P2_U6172 ; P2_U3876
g4419 and P2_U6178 P2_U6175 P2_U6181 ; P2_U3877
g4420 and P2_U3877 P2_U3876 P2_U6163 ; P2_U3878
g4421 and P2_U3884 P2_U3883 P2_U6112 P2_U6109 P2_U6106 ; P2_U3879
g4422 and P2_U6196 P2_U6193 P2_U6190 P2_U6187 P2_U6199 ; P2_U3880
g4423 and P2_U3878 P2_U3874 P2_U6139 P2_U6184 P2_U3880 ; P2_U3881
g4424 and P2_U6133 P2_U3879 ; P2_U3882
g4425 and P2_U6124 P2_U6121 P2_U6118 P2_U6115 ; P2_U3883
g4426 and P2_U6130 P2_U6127 ; P2_U3884
g4427 and P2_U5173 P2_U5177 P2_U5172 ; P2_U3885
g4428 and P2_U5670 P2_U5176 ; P2_U3886
g4429 and P2_U3449 P2_U3450 ; P2_U3887
g4430 and P2_U3432 P2_U3952 ; P2_U3888
g4431 and P2_U5701 P2_U3051 P2_U3422 ; P2_U3889
g4432 and P2_U3027 P2_U5183 ; P2_U3890
g4433 and P2_U3892 P2_U5226 ; P2_U3891
g4434 and P2_U5230 P2_U5229 ; P2_U3892
g4435 and P2_U3988 P2_U3078 ; P2_U3893
g4436 and P2_U5271 P2_U5270 ; P2_U3894
g4437 and P2_U5274 P2_U5273 ; P2_U3895
g4438 and P2_U5292 P2_U5291 ; P2_U3896
g4439 and P2_U5319 P2_U5318 ; P2_U3897
g4440 and P2_U3899 P2_U5360 ; P2_U3898
g4441 and P2_U5364 P2_U5363 ; P2_U3899
g4442 and P2_U5391 P2_U5387 ; P2_U3900
g4443 and P2_U3902 P2_U5396 ; P2_U3901
g4444 and P2_U5400 P2_U5399 ; P2_U3902
g4445 and P2_U5447 P2_STATE_REG_SCAN_IN ; P2_U3903
g4446 and P2_U5717 P2_U3415 ; P2_U3904
g4447 and P2_U5711 P2_U5701 ; P2_U3905
g4448 and P2_U3440 P2_U5512 ; P2_U3906
g4449 not P2_IR_REG_31__SCAN_IN ; P2_U3907
g4450 nand P2_U3027 P2_U3362 ; P2_U3908
g4451 nand P2_U5733 P2_U5728 ; P2_U3909
g4452 nand P2_U3631 P2_U3049 ; P2_U3910
g4453 nand P2_U3749 P2_U3049 ; P2_U3911
g4454 and P2_U5971 P2_U5970 ; P2_U3912
g4455 and P2_U5973 P2_U5972 ; P2_U3913
g4456 and P2_U5975 P2_U5974 ; P2_U3914
g4457 and P2_U5977 P2_U5976 ; P2_U3915
g4458 and P2_U5979 P2_U5978 ; P2_U3916
g4459 and P2_U5981 P2_U5980 ; P2_U3917
g4460 and P2_U5983 P2_U5982 ; P2_U3918
g4461 and P2_U5985 P2_U5984 ; P2_U3919
g4462 and P2_U5987 P2_U5986 ; P2_U3920
g4463 and P2_U5989 P2_U5988 ; P2_U3921
g4464 and P2_U5991 P2_U5990 ; P2_U3922
g4465 and P2_U5993 P2_U5992 ; P2_U3923
g4466 and P2_U5995 P2_U5994 ; P2_U3924
g4467 and P2_U5997 P2_U5996 ; P2_U3925
g4468 and P2_U5999 P2_U5998 ; P2_U3926
g4469 and P2_U6001 P2_U6000 ; P2_U3927
g4470 and P2_U6003 P2_U6002 ; P2_U3928
g4471 and P2_U6005 P2_U6004 ; P2_U3929
g4472 and P2_U6007 P2_U6006 ; P2_U3930
g4473 and P2_U6009 P2_U6008 ; P2_U3931
g4474 and P2_U6011 P2_U6010 ; P2_U3932
g4475 and P2_U6013 P2_U6012 ; P2_U3933
g4476 and P2_U6015 P2_U6014 ; P2_U3934
g4477 and P2_U6017 P2_U6016 ; P2_U3935
g4478 and P2_U6019 P2_U6018 ; P2_U3936
g4479 and P2_U6021 P2_U6020 ; P2_U3937
g4480 and P2_U6023 P2_U6022 ; P2_U3938
g4481 and P2_U6025 P2_U6024 ; P2_U3939
g4482 and P2_U6027 P2_U6026 ; P2_U3940
g4483 and P2_U6029 P2_U6028 ; P2_U3941
g4484 nand P2_U3748 P2_U3056 ; P2_U3942
g4485 and P2_U6031 P2_U6030 ; P2_U3943
g4486 and P2_U6033 P2_U6032 ; P2_U3944
g4487 not P2_R1312_U21 ; P2_U3945
g4488 and P2_U6103 P2_U6102 ; P2_U3946
g4489 nand P2_U3881 P2_U6136 P2_U3882 ; P2_U3947
g4490 not P2_R1299_U6 ; P2_U3948
g4491 not P2_U3370 ; P2_U3949
g4492 nand P2_U3982 P2_U3445 ; P2_U3950
g4493 not P2_U3368 ; P2_U3951
g4494 nand P2_U5674 P2_U3441 ; P2_U3952
g4495 not P2_U3432 ; P2_U3953
g4496 not P2_U3369 ; P2_U3954
g4497 not P2_U3363 ; P2_U3955
g4498 not P2_U3419 ; P2_U3956
g4499 not P2_U3418 ; P2_U3957
g4500 nand P2_U3962 P2_U5708 ; P2_U3958
g4501 not P2_U3367 ; P2_U3959
g4502 not P2_U3416 ; P2_U3960
g4503 not P2_U3366 ; P2_U3961
g4504 not P2_U3372 ; P2_U3962
g4505 not P2_U3364 ; P2_U3963
g4506 not P2_U3909 ; P2_U3964
g4507 not P2_U3427 ; P2_U3965
g4508 not P2_U3423 ; P2_U3966
g4509 not P2_U3421 ; P2_U3967
g4510 not P2_U3409 ; P2_U3968
g4511 not P2_U3407 ; P2_U3969
g4512 not P2_U3405 ; P2_U3970
g4513 not P2_U3403 ; P2_U3971
g4514 not P2_U3401 ; P2_U3972
g4515 not P2_U3399 ; P2_U3973
g4516 not P2_U3397 ; P2_U3974
g4517 not P2_U3395 ; P2_U3975
g4518 not P2_U3393 ; P2_U3976
g4519 not P2_U3414 ; P2_U3977
g4520 not P2_U3413 ; P2_U3978
g4521 not P2_U3411 ; P2_U3979
g4522 not P2_U3425 ; P2_U3980
g4523 not P2_U3420 ; P2_U3981
g4524 not P2_U3371 ; P2_U3982
g4525 not P2_U3417 ; P2_U3983
g4526 not P2_U3911 ; P2_U3984
g4527 not P2_U3910 ; P2_U3985
g4528 not P2_U3908 ; P2_U3986
g4529 not P2_U3942 ; P2_U3987
g4530 not P2_U3429 ; P2_U3988
g4531 nand P2_U3430 P2_STATE_REG_SCAN_IN ; P2_U3989
g4532 nand P2_U3957 P2_U3027 ; P2_U3990
g4533 not P2_U3426 ; P2_U3991
g4534 not P2_U3361 ; P2_U3992
g4535 not P2_U3428 ; P2_U3993
g4536 not P2_U3365 ; P2_U3994
g4537 not P2_U3422 ; P2_U3995
g4538 not P2_U3359 ; P2_U3996
g4539 nand U56 P2_U3152 ; P2_U3997
g4540 nand P2_U3033 P2_IR_REG_0__SCAN_IN ; P2_U3998
g4541 nand P2_U3996 P2_IR_REG_0__SCAN_IN ; P2_U3999
g4542 nand U45 P2_U3152 ; P2_U4000
g4543 nand P2_SUB_598_U49 P2_U3033 ; P2_U4001
g4544 nand P2_U3996 P2_IR_REG_1__SCAN_IN ; P2_U4002
g4545 nand U34 P2_U3152 ; P2_U4003
g4546 nand P2_SUB_598_U24 P2_U3033 ; P2_U4004
g4547 nand P2_U3996 P2_IR_REG_2__SCAN_IN ; P2_U4005
g4548 nand U31 P2_U3152 ; P2_U4006
g4549 nand P2_SUB_598_U25 P2_U3033 ; P2_U4007
g4550 nand P2_U3996 P2_IR_REG_3__SCAN_IN ; P2_U4008
g4551 nand U30 P2_U3152 ; P2_U4009
g4552 nand P2_SUB_598_U26 P2_U3033 ; P2_U4010
g4553 nand P2_U3996 P2_IR_REG_4__SCAN_IN ; P2_U4011
g4554 nand U29 P2_U3152 ; P2_U4012
g4555 nand P2_SUB_598_U74 P2_U3033 ; P2_U4013
g4556 nand P2_U3996 P2_IR_REG_5__SCAN_IN ; P2_U4014
g4557 nand U28 P2_U3152 ; P2_U4015
g4558 nand P2_SUB_598_U27 P2_U3033 ; P2_U4016
g4559 nand P2_U3996 P2_IR_REG_6__SCAN_IN ; P2_U4017
g4560 nand U27 P2_U3152 ; P2_U4018
g4561 nand P2_SUB_598_U28 P2_U3033 ; P2_U4019
g4562 nand P2_U3996 P2_IR_REG_7__SCAN_IN ; P2_U4020
g4563 nand U26 P2_U3152 ; P2_U4021
g4564 nand P2_SUB_598_U29 P2_U3033 ; P2_U4022
g4565 nand P2_U3996 P2_IR_REG_8__SCAN_IN ; P2_U4023
g4566 nand U25 P2_U3152 ; P2_U4024
g4567 nand P2_SUB_598_U72 P2_U3033 ; P2_U4025
g4568 nand P2_U3996 P2_IR_REG_9__SCAN_IN ; P2_U4026
g4569 nand U55 P2_U3152 ; P2_U4027
g4570 nand P2_SUB_598_U11 P2_U3033 ; P2_U4028
g4571 nand P2_U3996 P2_IR_REG_10__SCAN_IN ; P2_U4029
g4572 nand U54 P2_U3152 ; P2_U4030
g4573 nand P2_SUB_598_U12 P2_U3033 ; P2_U4031
g4574 nand P2_U3996 P2_IR_REG_11__SCAN_IN ; P2_U4032
g4575 nand U53 P2_U3152 ; P2_U4033
g4576 nand P2_SUB_598_U13 P2_U3033 ; P2_U4034
g4577 nand P2_U3996 P2_IR_REG_12__SCAN_IN ; P2_U4035
g4578 nand U52 P2_U3152 ; P2_U4036
g4579 nand P2_SUB_598_U99 P2_U3033 ; P2_U4037
g4580 nand P2_U3996 P2_IR_REG_13__SCAN_IN ; P2_U4038
g4581 nand U51 P2_U3152 ; P2_U4039
g4582 nand P2_SUB_598_U14 P2_U3033 ; P2_U4040
g4583 nand P2_U3996 P2_IR_REG_14__SCAN_IN ; P2_U4041
g4584 nand U50 P2_U3152 ; P2_U4042
g4585 nand P2_SUB_598_U15 P2_U3033 ; P2_U4043
g4586 nand P2_U3996 P2_IR_REG_15__SCAN_IN ; P2_U4044
g4587 nand U49 P2_U3152 ; P2_U4045
g4588 nand P2_SUB_598_U16 P2_U3033 ; P2_U4046
g4589 nand P2_U3996 P2_IR_REG_16__SCAN_IN ; P2_U4047
g4590 nand U48 P2_U3152 ; P2_U4048
g4591 nand P2_SUB_598_U97 P2_U3033 ; P2_U4049
g4592 nand P2_U3996 P2_IR_REG_17__SCAN_IN ; P2_U4050
g4593 nand U47 P2_U3152 ; P2_U4051
g4594 nand P2_SUB_598_U17 P2_U3033 ; P2_U4052
g4595 nand P2_U3996 P2_IR_REG_18__SCAN_IN ; P2_U4053
g4596 nand U46 P2_U3152 ; P2_U4054
g4597 nand P2_SUB_598_U18 P2_U3033 ; P2_U4055
g4598 nand P2_U3996 P2_IR_REG_19__SCAN_IN ; P2_U4056
g4599 nand U44 P2_U3152 ; P2_U4057
g4600 nand P2_SUB_598_U19 P2_U3033 ; P2_U4058
g4601 nand P2_U3996 P2_IR_REG_20__SCAN_IN ; P2_U4059
g4602 nand U43 P2_U3152 ; P2_U4060
g4603 nand P2_SUB_598_U92 P2_U3033 ; P2_U4061
g4604 nand P2_U3996 P2_IR_REG_21__SCAN_IN ; P2_U4062
g4605 nand U42 P2_U3152 ; P2_U4063
g4606 nand P2_SUB_598_U20 P2_U3033 ; P2_U4064
g4607 nand P2_U3996 P2_IR_REG_22__SCAN_IN ; P2_U4065
g4608 nand U41 P2_U3152 ; P2_U4066
g4609 nand P2_SUB_598_U21 P2_U3033 ; P2_U4067
g4610 nand P2_U3996 P2_IR_REG_23__SCAN_IN ; P2_U4068
g4611 nand U40 P2_U3152 ; P2_U4069
g4612 nand P2_SUB_598_U90 P2_U3033 ; P2_U4070
g4613 nand P2_U3996 P2_IR_REG_24__SCAN_IN ; P2_U4071
g4614 nand U39 P2_U3152 ; P2_U4072
g4615 nand P2_SUB_598_U22 P2_U3033 ; P2_U4073
g4616 nand P2_U3996 P2_IR_REG_25__SCAN_IN ; P2_U4074
g4617 nand U38 P2_U3152 ; P2_U4075
g4618 nand P2_SUB_598_U23 P2_U3033 ; P2_U4076
g4619 nand P2_U3996 P2_IR_REG_26__SCAN_IN ; P2_U4077
g4620 nand U37 P2_U3152 ; P2_U4078
g4621 nand P2_SUB_598_U87 P2_U3033 ; P2_U4079
g4622 nand P2_U3996 P2_IR_REG_27__SCAN_IN ; P2_U4080
g4623 nand U36 P2_U3152 ; P2_U4081
g4624 nand P2_SUB_598_U84 P2_U3033 ; P2_U4082
g4625 nand P2_U3996 P2_IR_REG_28__SCAN_IN ; P2_U4083
g4626 nand U35 P2_U3152 ; P2_U4084
g4627 nand P2_SUB_598_U81 P2_U3033 ; P2_U4085
g4628 nand P2_U3996 P2_IR_REG_29__SCAN_IN ; P2_U4086
g4629 nand U33 P2_U3152 ; P2_U4087
g4630 nand P2_SUB_598_U79 P2_U3033 ; P2_U4088
g4631 nand P2_U3996 P2_IR_REG_30__SCAN_IN ; P2_U4089
g4632 nand U32 P2_U3152 ; P2_U4090
g4633 nand P2_SUB_598_U77 P2_U3033 ; P2_U4091
g4634 nand P2_U3996 P2_IR_REG_31__SCAN_IN ; P2_U4092
g4635 nand P2_U3992 P2_U5698 ; P2_U4093
g4636 not P2_U3362 ; P2_U4094
g4637 nand P2_U3361 P2_U5689 ; P2_U4095
g4638 nand P2_U3361 P2_U5692 ; P2_U4096
g4639 nand P2_U4094 P2_D_REG_10__SCAN_IN ; P2_U4097
g4640 nand P2_U4094 P2_D_REG_11__SCAN_IN ; P2_U4098
g4641 nand P2_U4094 P2_D_REG_12__SCAN_IN ; P2_U4099
g4642 nand P2_U4094 P2_D_REG_13__SCAN_IN ; P2_U4100
g4643 nand P2_U4094 P2_D_REG_14__SCAN_IN ; P2_U4101
g4644 nand P2_U4094 P2_D_REG_15__SCAN_IN ; P2_U4102
g4645 nand P2_U4094 P2_D_REG_16__SCAN_IN ; P2_U4103
g4646 nand P2_U4094 P2_D_REG_17__SCAN_IN ; P2_U4104
g4647 nand P2_U4094 P2_D_REG_18__SCAN_IN ; P2_U4105
g4648 nand P2_U4094 P2_D_REG_19__SCAN_IN ; P2_U4106
g4649 nand P2_U4094 P2_D_REG_20__SCAN_IN ; P2_U4107
g4650 nand P2_U4094 P2_D_REG_21__SCAN_IN ; P2_U4108
g4651 nand P2_U4094 P2_D_REG_22__SCAN_IN ; P2_U4109
g4652 nand P2_U4094 P2_D_REG_23__SCAN_IN ; P2_U4110
g4653 nand P2_U4094 P2_D_REG_24__SCAN_IN ; P2_U4111
g4654 nand P2_U4094 P2_D_REG_25__SCAN_IN ; P2_U4112
g4655 nand P2_U4094 P2_D_REG_26__SCAN_IN ; P2_U4113
g4656 nand P2_U4094 P2_D_REG_27__SCAN_IN ; P2_U4114
g4657 nand P2_U4094 P2_D_REG_28__SCAN_IN ; P2_U4115
g4658 nand P2_U4094 P2_D_REG_29__SCAN_IN ; P2_U4116
g4659 nand P2_U4094 P2_D_REG_2__SCAN_IN ; P2_U4117
g4660 nand P2_U4094 P2_D_REG_30__SCAN_IN ; P2_U4118
g4661 nand P2_U4094 P2_D_REG_31__SCAN_IN ; P2_U4119
g4662 nand P2_U4094 P2_D_REG_3__SCAN_IN ; P2_U4120
g4663 nand P2_U4094 P2_D_REG_4__SCAN_IN ; P2_U4121
g4664 nand P2_U4094 P2_D_REG_5__SCAN_IN ; P2_U4122
g4665 nand P2_U4094 P2_D_REG_6__SCAN_IN ; P2_U4123
g4666 nand P2_U4094 P2_D_REG_7__SCAN_IN ; P2_U4124
g4667 nand P2_U4094 P2_D_REG_8__SCAN_IN ; P2_U4125
g4668 nand P2_U4094 P2_D_REG_9__SCAN_IN ; P2_U4126
g4669 nand P2_U3365 P2_U3428 P2_U5738 P2_U5737 ; P2_U4127
g4670 nand P2_U3025 P2_REG1_REG_1__SCAN_IN ; P2_U4128
g4671 nand P2_U3026 P2_REG0_REG_1__SCAN_IN ; P2_U4129
g4672 not P2_U3078 ; P2_U4130
g4673 nand P2_U3949 P2_U3445 ; P2_U4131
g4674 nand P2_U3958 P2_U4131 ; P2_U4132
g4675 nand P2_U3955 P2_R1146_U19 ; P2_U4133
g4676 nand P2_U3015 P2_R1113_U19 ; P2_U4134
g4677 nand P2_U3014 P2_R1131_U95 ; P2_U4135
g4678 nand P2_U3018 P2_R1179_U19 ; P2_U4136
g4679 nand P2_U3963 P2_R1203_U19 ; P2_U4137
g4680 nand P2_U3959 P2_R1164_U95 ; P2_U4138
g4681 nand P2_U3016 P2_R1233_U95 ; P2_U4139
g4682 not P2_U3373 ; P2_U4140
g4683 nand P2_U3448 P2_U3031 ; P2_U4141
g4684 nand P2_U3030 P2_U3078 ; P2_U4142
g4685 nand P2_R1215_U95 P2_U3028 ; P2_U4143
g4686 nand P2_U3448 P2_U4132 ; P2_U4144
g4687 nand P2_U3619 P2_U4140 ; P2_U4145
g4688 nand P2_U3025 P2_REG1_REG_2__SCAN_IN ; P2_U4146
g4689 nand P2_U3026 P2_REG0_REG_2__SCAN_IN ; P2_U4147
g4690 not P2_U3068 ; P2_U4148
g4691 nand P2_U3025 P2_REG1_REG_0__SCAN_IN ; P2_U4149
g4692 nand P2_U3026 P2_REG0_REG_0__SCAN_IN ; P2_U4150
g4693 not P2_U3077 ; P2_U4151
g4694 nand P2_U3038 P2_U3077 ; P2_U4152
g4695 nand P2_R1146_U94 P2_U3955 ; P2_U4153
g4696 nand P2_R1113_U94 P2_U3015 ; P2_U4154
g4697 nand P2_R1131_U94 P2_U3014 ; P2_U4155
g4698 nand P2_R1179_U94 P2_U3018 ; P2_U4156
g4699 nand P2_R1203_U94 P2_U3963 ; P2_U4157
g4700 nand P2_R1164_U94 P2_U3959 ; P2_U4158
g4701 nand P2_R1233_U94 P2_U3016 ; P2_U4159
g4702 not P2_U3374 ; P2_U4160
g4703 nand P2_R1275_U55 P2_U3031 ; P2_U4161
g4704 nand P2_U3030 P2_U3068 ; P2_U4162
g4705 nand P2_R1215_U94 P2_U3028 ; P2_U4163
g4706 nand P2_U3453 P2_U4132 ; P2_U4164
g4707 nand P2_U3635 P2_U4160 ; P2_U4165
g4708 nand P2_U3024 P2_REG2_REG_3__SCAN_IN ; P2_U4166
g4709 nand P2_U3025 P2_REG1_REG_3__SCAN_IN ; P2_U4167
g4710 nand P2_U3026 P2_REG0_REG_3__SCAN_IN ; P2_U4168
g4711 nand P2_ADD_609_U4 P2_U3023 ; P2_U4169
g4712 not P2_U3064 ; P2_U4170
g4713 nand P2_U3038 P2_U3078 ; P2_U4171
g4714 nand P2_R1146_U104 P2_U3955 ; P2_U4172
g4715 nand P2_R1113_U104 P2_U3015 ; P2_U4173
g4716 nand P2_R1131_U16 P2_U3014 ; P2_U4174
g4717 nand P2_R1179_U104 P2_U3018 ; P2_U4175
g4718 nand P2_R1203_U104 P2_U3963 ; P2_U4176
g4719 nand P2_R1164_U16 P2_U3959 ; P2_U4177
g4720 nand P2_R1233_U16 P2_U3016 ; P2_U4178
g4721 not P2_U3375 ; P2_U4179
g4722 nand P2_R1275_U18 P2_U3031 ; P2_U4180
g4723 nand P2_U3030 P2_U3064 ; P2_U4181
g4724 nand P2_R1215_U16 P2_U3028 ; P2_U4182
g4725 nand P2_U3456 P2_U4132 ; P2_U4183
g4726 nand P2_U3639 P2_U4179 ; P2_U4184
g4727 nand P2_U3024 P2_REG2_REG_4__SCAN_IN ; P2_U4185
g4728 nand P2_U3025 P2_REG1_REG_4__SCAN_IN ; P2_U4186
g4729 nand P2_U3026 P2_REG0_REG_4__SCAN_IN ; P2_U4187
g4730 nand P2_ADD_609_U54 P2_U3023 ; P2_U4188
g4731 not P2_U3060 ; P2_U4189
g4732 nand P2_U3038 P2_U3068 ; P2_U4190
g4733 nand P2_R1146_U16 P2_U3955 ; P2_U4191
g4734 nand P2_R1113_U16 P2_U3015 ; P2_U4192
g4735 nand P2_R1131_U100 P2_U3014 ; P2_U4193
g4736 nand P2_R1179_U16 P2_U3018 ; P2_U4194
g4737 nand P2_R1203_U16 P2_U3963 ; P2_U4195
g4738 nand P2_R1164_U100 P2_U3959 ; P2_U4196
g4739 nand P2_R1233_U100 P2_U3016 ; P2_U4197
g4740 not P2_U3376 ; P2_U4198
g4741 nand P2_R1275_U20 P2_U3031 ; P2_U4199
g4742 nand P2_U3030 P2_U3060 ; P2_U4200
g4743 nand P2_R1215_U100 P2_U3028 ; P2_U4201
g4744 nand P2_U3459 P2_U4132 ; P2_U4202
g4745 nand P2_U3643 P2_U4198 ; P2_U4203
g4746 nand P2_U3024 P2_REG2_REG_5__SCAN_IN ; P2_U4204
g4747 nand P2_U3025 P2_REG1_REG_5__SCAN_IN ; P2_U4205
g4748 nand P2_U3026 P2_REG0_REG_5__SCAN_IN ; P2_U4206
g4749 nand P2_ADD_609_U53 P2_U3023 ; P2_U4207
g4750 not P2_U3067 ; P2_U4208
g4751 nand P2_U3038 P2_U3064 ; P2_U4209
g4752 nand P2_R1146_U103 P2_U3955 ; P2_U4210
g4753 nand P2_R1113_U103 P2_U3015 ; P2_U4211
g4754 nand P2_R1131_U99 P2_U3014 ; P2_U4212
g4755 nand P2_R1179_U103 P2_U3018 ; P2_U4213
g4756 nand P2_R1203_U103 P2_U3963 ; P2_U4214
g4757 nand P2_R1164_U99 P2_U3959 ; P2_U4215
g4758 nand P2_R1233_U99 P2_U3016 ; P2_U4216
g4759 not P2_U3377 ; P2_U4217
g4760 nand P2_R1275_U21 P2_U3031 ; P2_U4218
g4761 nand P2_U3030 P2_U3067 ; P2_U4219
g4762 nand P2_R1215_U99 P2_U3028 ; P2_U4220
g4763 nand P2_U3462 P2_U4132 ; P2_U4221
g4764 nand P2_U3647 P2_U4217 ; P2_U4222
g4765 nand P2_U3024 P2_REG2_REG_6__SCAN_IN ; P2_U4223
g4766 nand P2_U3025 P2_REG1_REG_6__SCAN_IN ; P2_U4224
g4767 nand P2_U3026 P2_REG0_REG_6__SCAN_IN ; P2_U4225
g4768 nand P2_ADD_609_U52 P2_U3023 ; P2_U4226
g4769 not P2_U3071 ; P2_U4227
g4770 nand P2_U3038 P2_U3060 ; P2_U4228
g4771 nand P2_R1146_U102 P2_U3955 ; P2_U4229
g4772 nand P2_R1113_U102 P2_U3015 ; P2_U4230
g4773 nand P2_R1131_U17 P2_U3014 ; P2_U4231
g4774 nand P2_R1179_U102 P2_U3018 ; P2_U4232
g4775 nand P2_R1203_U102 P2_U3963 ; P2_U4233
g4776 nand P2_R1164_U17 P2_U3959 ; P2_U4234
g4777 nand P2_R1233_U17 P2_U3016 ; P2_U4235
g4778 not P2_U3378 ; P2_U4236
g4779 nand P2_R1275_U65 P2_U3031 ; P2_U4237
g4780 nand P2_U3030 P2_U3071 ; P2_U4238
g4781 nand P2_R1215_U17 P2_U3028 ; P2_U4239
g4782 nand P2_U3465 P2_U4132 ; P2_U4240
g4783 nand P2_U3651 P2_U4236 ; P2_U4241
g4784 nand P2_U3024 P2_REG2_REG_7__SCAN_IN ; P2_U4242
g4785 nand P2_U3025 P2_REG1_REG_7__SCAN_IN ; P2_U4243
g4786 nand P2_U3026 P2_REG0_REG_7__SCAN_IN ; P2_U4244
g4787 nand P2_ADD_609_U51 P2_U3023 ; P2_U4245
g4788 not P2_U3070 ; P2_U4246
g4789 nand P2_U3038 P2_U3067 ; P2_U4247
g4790 nand P2_R1146_U17 P2_U3955 ; P2_U4248
g4791 nand P2_R1113_U17 P2_U3015 ; P2_U4249
g4792 nand P2_R1131_U98 P2_U3014 ; P2_U4250
g4793 nand P2_R1179_U17 P2_U3018 ; P2_U4251
g4794 nand P2_R1203_U17 P2_U3963 ; P2_U4252
g4795 nand P2_R1164_U98 P2_U3959 ; P2_U4253
g4796 nand P2_R1233_U98 P2_U3016 ; P2_U4254
g4797 not P2_U3379 ; P2_U4255
g4798 nand P2_R1275_U22 P2_U3031 ; P2_U4256
g4799 nand P2_U3030 P2_U3070 ; P2_U4257
g4800 nand P2_R1215_U98 P2_U3028 ; P2_U4258
g4801 nand P2_U3468 P2_U4132 ; P2_U4259
g4802 nand P2_U3655 P2_U4255 ; P2_U4260
g4803 nand P2_U3024 P2_REG2_REG_8__SCAN_IN ; P2_U4261
g4804 nand P2_U3025 P2_REG1_REG_8__SCAN_IN ; P2_U4262
g4805 nand P2_U3026 P2_REG0_REG_8__SCAN_IN ; P2_U4263
g4806 nand P2_ADD_609_U50 P2_U3023 ; P2_U4264
g4807 not P2_U3084 ; P2_U4265
g4808 nand P2_U3038 P2_U3071 ; P2_U4266
g4809 nand P2_R1146_U101 P2_U3955 ; P2_U4267
g4810 nand P2_R1113_U101 P2_U3015 ; P2_U4268
g4811 nand P2_R1131_U18 P2_U3014 ; P2_U4269
g4812 nand P2_R1179_U101 P2_U3018 ; P2_U4270
g4813 nand P2_R1203_U101 P2_U3963 ; P2_U4271
g4814 nand P2_R1164_U18 P2_U3959 ; P2_U4272
g4815 nand P2_R1233_U18 P2_U3016 ; P2_U4273
g4816 not P2_U3380 ; P2_U4274
g4817 nand P2_R1275_U23 P2_U3031 ; P2_U4275
g4818 nand P2_U3030 P2_U3084 ; P2_U4276
g4819 nand P2_R1215_U18 P2_U3028 ; P2_U4277
g4820 nand P2_U3471 P2_U4132 ; P2_U4278
g4821 nand P2_U3659 P2_U4274 ; P2_U4279
g4822 nand P2_U3024 P2_REG2_REG_9__SCAN_IN ; P2_U4280
g4823 nand P2_U3025 P2_REG1_REG_9__SCAN_IN ; P2_U4281
g4824 nand P2_U3026 P2_REG0_REG_9__SCAN_IN ; P2_U4282
g4825 nand P2_ADD_609_U49 P2_U3023 ; P2_U4283
g4826 not P2_U3083 ; P2_U4284
g4827 nand P2_U3038 P2_U3070 ; P2_U4285
g4828 nand P2_R1146_U18 P2_U3955 ; P2_U4286
g4829 nand P2_R1113_U18 P2_U3015 ; P2_U4287
g4830 nand P2_R1131_U97 P2_U3014 ; P2_U4288
g4831 nand P2_R1179_U18 P2_U3018 ; P2_U4289
g4832 nand P2_R1203_U18 P2_U3963 ; P2_U4290
g4833 nand P2_R1164_U97 P2_U3959 ; P2_U4291
g4834 nand P2_R1233_U97 P2_U3016 ; P2_U4292
g4835 not P2_U3381 ; P2_U4293
g4836 nand P2_R1275_U24 P2_U3031 ; P2_U4294
g4837 nand P2_U3030 P2_U3083 ; P2_U4295
g4838 nand P2_R1215_U97 P2_U3028 ; P2_U4296
g4839 nand P2_U3474 P2_U4132 ; P2_U4297
g4840 nand P2_U3663 P2_U4293 ; P2_U4298
g4841 nand P2_U3024 P2_REG2_REG_10__SCAN_IN ; P2_U4299
g4842 nand P2_U3025 P2_REG1_REG_10__SCAN_IN ; P2_U4300
g4843 nand P2_U3026 P2_REG0_REG_10__SCAN_IN ; P2_U4301
g4844 nand P2_ADD_609_U73 P2_U3023 ; P2_U4302
g4845 not P2_U3062 ; P2_U4303
g4846 nand P2_U3038 P2_U3084 ; P2_U4304
g4847 nand P2_R1146_U100 P2_U3955 ; P2_U4305
g4848 nand P2_R1113_U100 P2_U3015 ; P2_U4306
g4849 nand P2_R1131_U96 P2_U3014 ; P2_U4307
g4850 nand P2_R1179_U100 P2_U3018 ; P2_U4308
g4851 nand P2_R1203_U100 P2_U3963 ; P2_U4309
g4852 nand P2_R1164_U96 P2_U3959 ; P2_U4310
g4853 nand P2_R1233_U96 P2_U3016 ; P2_U4311
g4854 not P2_U3382 ; P2_U4312
g4855 nand P2_R1275_U63 P2_U3031 ; P2_U4313
g4856 nand P2_U3030 P2_U3062 ; P2_U4314
g4857 nand P2_R1215_U96 P2_U3028 ; P2_U4315
g4858 nand P2_U3477 P2_U4132 ; P2_U4316
g4859 nand P2_U3667 P2_U4312 ; P2_U4317
g4860 nand P2_U3024 P2_REG2_REG_11__SCAN_IN ; P2_U4318
g4861 nand P2_U3025 P2_REG1_REG_11__SCAN_IN ; P2_U4319
g4862 nand P2_U3026 P2_REG0_REG_11__SCAN_IN ; P2_U4320
g4863 nand P2_ADD_609_U72 P2_U3023 ; P2_U4321
g4864 not P2_U3063 ; P2_U4322
g4865 nand P2_U3038 P2_U3083 ; P2_U4323
g4866 nand P2_R1146_U110 P2_U3955 ; P2_U4324
g4867 nand P2_R1113_U110 P2_U3015 ; P2_U4325
g4868 nand P2_R1131_U10 P2_U3014 ; P2_U4326
g4869 nand P2_R1179_U110 P2_U3018 ; P2_U4327
g4870 nand P2_R1203_U110 P2_U3963 ; P2_U4328
g4871 nand P2_R1164_U10 P2_U3959 ; P2_U4329
g4872 nand P2_R1233_U10 P2_U3016 ; P2_U4330
g4873 not P2_U3383 ; P2_U4331
g4874 nand P2_R1275_U6 P2_U3031 ; P2_U4332
g4875 nand P2_U3030 P2_U3063 ; P2_U4333
g4876 nand P2_R1215_U10 P2_U3028 ; P2_U4334
g4877 nand P2_U3480 P2_U4132 ; P2_U4335
g4878 nand P2_U3671 P2_U4331 ; P2_U4336
g4879 nand P2_U3024 P2_REG2_REG_12__SCAN_IN ; P2_U4337
g4880 nand P2_U3025 P2_REG1_REG_12__SCAN_IN ; P2_U4338
g4881 nand P2_U3026 P2_REG0_REG_12__SCAN_IN ; P2_U4339
g4882 nand P2_ADD_609_U71 P2_U3023 ; P2_U4340
g4883 not P2_U3072 ; P2_U4341
g4884 nand P2_U3038 P2_U3062 ; P2_U4342
g4885 nand P2_R1146_U11 P2_U3955 ; P2_U4343
g4886 nand P2_R1113_U11 P2_U3015 ; P2_U4344
g4887 nand P2_R1131_U114 P2_U3014 ; P2_U4345
g4888 nand P2_R1179_U11 P2_U3018 ; P2_U4346
g4889 nand P2_R1203_U11 P2_U3963 ; P2_U4347
g4890 nand P2_R1164_U114 P2_U3959 ; P2_U4348
g4891 nand P2_R1233_U114 P2_U3016 ; P2_U4349
g4892 not P2_U3384 ; P2_U4350
g4893 nand P2_R1275_U7 P2_U3031 ; P2_U4351
g4894 nand P2_U3030 P2_U3072 ; P2_U4352
g4895 nand P2_R1215_U114 P2_U3028 ; P2_U4353
g4896 nand P2_U3483 P2_U4132 ; P2_U4354
g4897 nand P2_U3675 P2_U4350 ; P2_U4355
g4898 nand P2_U3024 P2_REG2_REG_13__SCAN_IN ; P2_U4356
g4899 nand P2_U3025 P2_REG1_REG_13__SCAN_IN ; P2_U4357
g4900 nand P2_U3026 P2_REG0_REG_13__SCAN_IN ; P2_U4358
g4901 nand P2_ADD_609_U70 P2_U3023 ; P2_U4359
g4902 not P2_U3080 ; P2_U4360
g4903 nand P2_U3038 P2_U3063 ; P2_U4361
g4904 nand P2_R1146_U99 P2_U3955 ; P2_U4362
g4905 nand P2_R1113_U99 P2_U3015 ; P2_U4363
g4906 nand P2_R1131_U113 P2_U3014 ; P2_U4364
g4907 nand P2_R1179_U99 P2_U3018 ; P2_U4365
g4908 nand P2_R1203_U99 P2_U3963 ; P2_U4366
g4909 nand P2_R1164_U113 P2_U3959 ; P2_U4367
g4910 nand P2_R1233_U113 P2_U3016 ; P2_U4368
g4911 not P2_U3385 ; P2_U4369
g4912 nand P2_R1275_U8 P2_U3031 ; P2_U4370
g4913 nand P2_U3030 P2_U3080 ; P2_U4371
g4914 nand P2_R1215_U113 P2_U3028 ; P2_U4372
g4915 nand P2_U3486 P2_U4132 ; P2_U4373
g4916 nand P2_U3679 P2_U4369 ; P2_U4374
g4917 nand P2_U3024 P2_REG2_REG_14__SCAN_IN ; P2_U4375
g4918 nand P2_U3025 P2_REG1_REG_14__SCAN_IN ; P2_U4376
g4919 nand P2_U3026 P2_REG0_REG_14__SCAN_IN ; P2_U4377
g4920 nand P2_ADD_609_U69 P2_U3023 ; P2_U4378
g4921 not P2_U3079 ; P2_U4379
g4922 nand P2_U3038 P2_U3072 ; P2_U4380
g4923 nand P2_R1146_U98 P2_U3955 ; P2_U4381
g4924 nand P2_R1113_U98 P2_U3015 ; P2_U4382
g4925 nand P2_R1131_U11 P2_U3014 ; P2_U4383
g4926 nand P2_R1179_U98 P2_U3018 ; P2_U4384
g4927 nand P2_R1203_U98 P2_U3963 ; P2_U4385
g4928 nand P2_R1164_U11 P2_U3959 ; P2_U4386
g4929 nand P2_R1233_U11 P2_U3016 ; P2_U4387
g4930 not P2_U3386 ; P2_U4388
g4931 nand P2_R1275_U86 P2_U3031 ; P2_U4389
g4932 nand P2_U3030 P2_U3079 ; P2_U4390
g4933 nand P2_R1215_U11 P2_U3028 ; P2_U4391
g4934 nand P2_U3489 P2_U4132 ; P2_U4392
g4935 nand P2_U3683 P2_U4388 ; P2_U4393
g4936 nand P2_U3024 P2_REG2_REG_15__SCAN_IN ; P2_U4394
g4937 nand P2_U3025 P2_REG1_REG_15__SCAN_IN ; P2_U4395
g4938 nand P2_U3026 P2_REG0_REG_15__SCAN_IN ; P2_U4396
g4939 nand P2_ADD_609_U68 P2_U3023 ; P2_U4397
g4940 not P2_U3074 ; P2_U4398
g4941 nand P2_U3038 P2_U3080 ; P2_U4399
g4942 nand P2_R1146_U109 P2_U3955 ; P2_U4400
g4943 nand P2_R1113_U109 P2_U3015 ; P2_U4401
g4944 nand P2_R1131_U112 P2_U3014 ; P2_U4402
g4945 nand P2_R1179_U109 P2_U3018 ; P2_U4403
g4946 nand P2_R1203_U109 P2_U3963 ; P2_U4404
g4947 nand P2_R1164_U112 P2_U3959 ; P2_U4405
g4948 nand P2_R1233_U112 P2_U3016 ; P2_U4406
g4949 not P2_U3387 ; P2_U4407
g4950 nand P2_R1275_U9 P2_U3031 ; P2_U4408
g4951 nand P2_U3030 P2_U3074 ; P2_U4409
g4952 nand P2_R1215_U112 P2_U3028 ; P2_U4410
g4953 nand P2_U3492 P2_U4132 ; P2_U4411
g4954 nand P2_U3687 P2_U4407 ; P2_U4412
g4955 nand P2_U3024 P2_REG2_REG_16__SCAN_IN ; P2_U4413
g4956 nand P2_U3025 P2_REG1_REG_16__SCAN_IN ; P2_U4414
g4957 nand P2_U3026 P2_REG0_REG_16__SCAN_IN ; P2_U4415
g4958 nand P2_ADD_609_U67 P2_U3023 ; P2_U4416
g4959 not P2_U3073 ; P2_U4417
g4960 nand P2_U3038 P2_U3079 ; P2_U4418
g4961 nand P2_R1146_U108 P2_U3955 ; P2_U4419
g4962 nand P2_R1113_U108 P2_U3015 ; P2_U4420
g4963 nand P2_R1131_U111 P2_U3014 ; P2_U4421
g4964 nand P2_R1179_U108 P2_U3018 ; P2_U4422
g4965 nand P2_R1203_U108 P2_U3963 ; P2_U4423
g4966 nand P2_R1164_U111 P2_U3959 ; P2_U4424
g4967 nand P2_R1233_U111 P2_U3016 ; P2_U4425
g4968 not P2_U3388 ; P2_U4426
g4969 nand P2_R1275_U10 P2_U3031 ; P2_U4427
g4970 nand P2_U3030 P2_U3073 ; P2_U4428
g4971 nand P2_R1215_U111 P2_U3028 ; P2_U4429
g4972 nand P2_U3495 P2_U4132 ; P2_U4430
g4973 nand P2_U3691 P2_U4426 ; P2_U4431
g4974 nand P2_U3024 P2_REG2_REG_17__SCAN_IN ; P2_U4432
g4975 nand P2_U3025 P2_REG1_REG_17__SCAN_IN ; P2_U4433
g4976 nand P2_U3026 P2_REG0_REG_17__SCAN_IN ; P2_U4434
g4977 nand P2_ADD_609_U66 P2_U3023 ; P2_U4435
g4978 not P2_U3069 ; P2_U4436
g4979 nand P2_U3038 P2_U3074 ; P2_U4437
g4980 nand P2_R1146_U12 P2_U3955 ; P2_U4438
g4981 nand P2_R1113_U12 P2_U3015 ; P2_U4439
g4982 nand P2_R1131_U110 P2_U3014 ; P2_U4440
g4983 nand P2_R1179_U12 P2_U3018 ; P2_U4441
g4984 nand P2_R1203_U12 P2_U3963 ; P2_U4442
g4985 nand P2_R1164_U110 P2_U3959 ; P2_U4443
g4986 nand P2_R1233_U110 P2_U3016 ; P2_U4444
g4987 not P2_U3389 ; P2_U4445
g4988 nand P2_R1275_U11 P2_U3031 ; P2_U4446
g4989 nand P2_U3030 P2_U3069 ; P2_U4447
g4990 nand P2_R1215_U110 P2_U3028 ; P2_U4448
g4991 nand P2_U3498 P2_U4132 ; P2_U4449
g4992 nand P2_U3695 P2_U4445 ; P2_U4450
g4993 nand P2_U3024 P2_REG2_REG_18__SCAN_IN ; P2_U4451
g4994 nand P2_U3025 P2_REG1_REG_18__SCAN_IN ; P2_U4452
g4995 nand P2_U3026 P2_REG0_REG_18__SCAN_IN ; P2_U4453
g4996 nand P2_ADD_609_U65 P2_U3023 ; P2_U4454
g4997 not P2_U3082 ; P2_U4455
g4998 nand P2_U3038 P2_U3073 ; P2_U4456
g4999 nand P2_R1146_U97 P2_U3955 ; P2_U4457
g5000 nand P2_R1113_U97 P2_U3015 ; P2_U4458
g5001 nand P2_R1131_U12 P2_U3014 ; P2_U4459
g5002 nand P2_R1179_U97 P2_U3018 ; P2_U4460
g5003 nand P2_R1203_U97 P2_U3963 ; P2_U4461
g5004 nand P2_R1164_U12 P2_U3959 ; P2_U4462
g5005 nand P2_R1233_U12 P2_U3016 ; P2_U4463
g5006 not P2_U3390 ; P2_U4464
g5007 nand P2_R1275_U84 P2_U3031 ; P2_U4465
g5008 nand P2_U3030 P2_U3082 ; P2_U4466
g5009 nand P2_R1215_U12 P2_U3028 ; P2_U4467
g5010 nand P2_U3501 P2_U4132 ; P2_U4468
g5011 nand P2_U3699 P2_U4464 ; P2_U4469
g5012 nand P2_U3024 P2_REG2_REG_19__SCAN_IN ; P2_U4470
g5013 nand P2_U3025 P2_REG1_REG_19__SCAN_IN ; P2_U4471
g5014 nand P2_U3026 P2_REG0_REG_19__SCAN_IN ; P2_U4472
g5015 nand P2_ADD_609_U64 P2_U3023 ; P2_U4473
g5016 not P2_U3081 ; P2_U4474
g5017 nand P2_U3038 P2_U3069 ; P2_U4475
g5018 nand P2_R1146_U96 P2_U3955 ; P2_U4476
g5019 nand P2_R1113_U96 P2_U3015 ; P2_U4477
g5020 nand P2_R1131_U109 P2_U3014 ; P2_U4478
g5021 nand P2_R1179_U96 P2_U3018 ; P2_U4479
g5022 nand P2_R1203_U96 P2_U3963 ; P2_U4480
g5023 nand P2_R1164_U109 P2_U3959 ; P2_U4481
g5024 nand P2_R1233_U109 P2_U3016 ; P2_U4482
g5025 not P2_U3391 ; P2_U4483
g5026 nand P2_R1275_U12 P2_U3031 ; P2_U4484
g5027 nand P2_U3030 P2_U3081 ; P2_U4485
g5028 nand P2_R1215_U109 P2_U3028 ; P2_U4486
g5029 nand P2_U3504 P2_U4132 ; P2_U4487
g5030 nand P2_U3703 P2_U4483 ; P2_U4488
g5031 nand P2_U3024 P2_REG2_REG_20__SCAN_IN ; P2_U4489
g5032 nand P2_U3025 P2_REG1_REG_20__SCAN_IN ; P2_U4490
g5033 nand P2_U3026 P2_REG0_REG_20__SCAN_IN ; P2_U4491
g5034 nand P2_ADD_609_U63 P2_U3023 ; P2_U4492
g5035 not P2_U3076 ; P2_U4493
g5036 nand P2_U3038 P2_U3082 ; P2_U4494
g5037 nand P2_R1146_U95 P2_U3955 ; P2_U4495
g5038 nand P2_R1113_U95 P2_U3015 ; P2_U4496
g5039 nand P2_R1131_U108 P2_U3014 ; P2_U4497
g5040 nand P2_R1179_U95 P2_U3018 ; P2_U4498
g5041 nand P2_R1203_U95 P2_U3963 ; P2_U4499
g5042 nand P2_R1164_U108 P2_U3959 ; P2_U4500
g5043 nand P2_R1233_U108 P2_U3016 ; P2_U4501
g5044 not P2_U3392 ; P2_U4502
g5045 nand P2_R1275_U82 P2_U3031 ; P2_U4503
g5046 nand P2_U3030 P2_U3076 ; P2_U4504
g5047 nand P2_R1215_U108 P2_U3028 ; P2_U4505
g5048 nand P2_U3506 P2_U4132 ; P2_U4506
g5049 nand P2_U3707 P2_U4502 ; P2_U4507
g5050 nand P2_U3024 P2_REG2_REG_21__SCAN_IN ; P2_U4508
g5051 nand P2_U3025 P2_REG1_REG_21__SCAN_IN ; P2_U4509
g5052 nand P2_U3026 P2_REG0_REG_21__SCAN_IN ; P2_U4510
g5053 nand P2_ADD_609_U62 P2_U3023 ; P2_U4511
g5054 not P2_U3075 ; P2_U4512
g5055 nand P2_U3038 P2_U3081 ; P2_U4513
g5056 nand P2_R1146_U93 P2_U3955 ; P2_U4514
g5057 nand P2_R1113_U93 P2_U3015 ; P2_U4515
g5058 nand P2_R1131_U13 P2_U3014 ; P2_U4516
g5059 nand P2_R1179_U93 P2_U3018 ; P2_U4517
g5060 nand P2_R1203_U93 P2_U3963 ; P2_U4518
g5061 nand P2_R1164_U13 P2_U3959 ; P2_U4519
g5062 nand P2_R1233_U13 P2_U3016 ; P2_U4520
g5063 not P2_U3394 ; P2_U4521
g5064 nand P2_R1275_U13 P2_U3031 ; P2_U4522
g5065 nand P2_U3030 P2_U3075 ; P2_U4523
g5066 nand P2_R1215_U13 P2_U3028 ; P2_U4524
g5067 nand P2_U3976 P2_U4132 ; P2_U4525
g5068 nand P2_U3711 P2_U4521 ; P2_U4526
g5069 nand P2_U3024 P2_REG2_REG_22__SCAN_IN ; P2_U4527
g5070 nand P2_U3025 P2_REG1_REG_22__SCAN_IN ; P2_U4528
g5071 nand P2_U3026 P2_REG0_REG_22__SCAN_IN ; P2_U4529
g5072 nand P2_ADD_609_U61 P2_U3023 ; P2_U4530
g5073 not P2_U3061 ; P2_U4531
g5074 nand P2_U3038 P2_U3076 ; P2_U4532
g5075 nand P2_R1146_U107 P2_U3955 ; P2_U4533
g5076 nand P2_R1113_U107 P2_U3015 ; P2_U4534
g5077 nand P2_R1131_U14 P2_U3014 ; P2_U4535
g5078 nand P2_R1179_U107 P2_U3018 ; P2_U4536
g5079 nand P2_R1203_U107 P2_U3963 ; P2_U4537
g5080 nand P2_R1164_U14 P2_U3959 ; P2_U4538
g5081 nand P2_R1233_U14 P2_U3016 ; P2_U4539
g5082 not P2_U3396 ; P2_U4540
g5083 nand P2_R1275_U78 P2_U3031 ; P2_U4541
g5084 nand P2_U3030 P2_U3061 ; P2_U4542
g5085 nand P2_R1215_U14 P2_U3028 ; P2_U4543
g5086 nand P2_U3975 P2_U4132 ; P2_U4544
g5087 nand P2_U3715 P2_U4540 ; P2_U4545
g5088 nand P2_U3024 P2_REG2_REG_23__SCAN_IN ; P2_U4546
g5089 nand P2_U3025 P2_REG1_REG_23__SCAN_IN ; P2_U4547
g5090 nand P2_U3026 P2_REG0_REG_23__SCAN_IN ; P2_U4548
g5091 nand P2_ADD_609_U60 P2_U3023 ; P2_U4549
g5092 not P2_U3066 ; P2_U4550
g5093 nand P2_U3038 P2_U3075 ; P2_U4551
g5094 nand P2_R1146_U106 P2_U3955 ; P2_U4552
g5095 nand P2_R1113_U106 P2_U3015 ; P2_U4553
g5096 nand P2_R1131_U107 P2_U3014 ; P2_U4554
g5097 nand P2_R1179_U106 P2_U3018 ; P2_U4555
g5098 nand P2_R1203_U106 P2_U3963 ; P2_U4556
g5099 nand P2_R1164_U107 P2_U3959 ; P2_U4557
g5100 nand P2_R1233_U107 P2_U3016 ; P2_U4558
g5101 not P2_U3398 ; P2_U4559
g5102 nand P2_R1275_U14 P2_U3031 ; P2_U4560
g5103 nand P2_U3030 P2_U3066 ; P2_U4561
g5104 nand P2_R1215_U107 P2_U3028 ; P2_U4562
g5105 nand P2_U3974 P2_U4132 ; P2_U4563
g5106 nand P2_U3719 P2_U4559 ; P2_U4564
g5107 nand P2_U3024 P2_REG2_REG_24__SCAN_IN ; P2_U4565
g5108 nand P2_U3025 P2_REG1_REG_24__SCAN_IN ; P2_U4566
g5109 nand P2_U3026 P2_REG0_REG_24__SCAN_IN ; P2_U4567
g5110 nand P2_ADD_609_U59 P2_U3023 ; P2_U4568
g5111 not P2_U3065 ; P2_U4569
g5112 nand P2_U3038 P2_U3061 ; P2_U4570
g5113 nand P2_R1146_U13 P2_U3955 ; P2_U4571
g5114 nand P2_R1113_U13 P2_U3015 ; P2_U4572
g5115 nand P2_R1131_U106 P2_U3014 ; P2_U4573
g5116 nand P2_R1179_U13 P2_U3018 ; P2_U4574
g5117 nand P2_R1203_U13 P2_U3963 ; P2_U4575
g5118 nand P2_R1164_U106 P2_U3959 ; P2_U4576
g5119 nand P2_R1233_U106 P2_U3016 ; P2_U4577
g5120 not P2_U3400 ; P2_U4578
g5121 nand P2_R1275_U76 P2_U3031 ; P2_U4579
g5122 nand P2_U3030 P2_U3065 ; P2_U4580
g5123 nand P2_R1215_U106 P2_U3028 ; P2_U4581
g5124 nand P2_U3973 P2_U4132 ; P2_U4582
g5125 nand P2_U3723 P2_U4578 ; P2_U4583
g5126 nand P2_U3024 P2_REG2_REG_25__SCAN_IN ; P2_U4584
g5127 nand P2_U3025 P2_REG1_REG_25__SCAN_IN ; P2_U4585
g5128 nand P2_U3026 P2_REG0_REG_25__SCAN_IN ; P2_U4586
g5129 nand P2_ADD_609_U58 P2_U3023 ; P2_U4587
g5130 not P2_U3058 ; P2_U4588
g5131 nand P2_U3038 P2_U3066 ; P2_U4589
g5132 nand P2_R1146_U92 P2_U3955 ; P2_U4590
g5133 nand P2_R1113_U92 P2_U3015 ; P2_U4591
g5134 nand P2_R1131_U105 P2_U3014 ; P2_U4592
g5135 nand P2_R1179_U92 P2_U3018 ; P2_U4593
g5136 nand P2_R1203_U92 P2_U3963 ; P2_U4594
g5137 nand P2_R1164_U105 P2_U3959 ; P2_U4595
g5138 nand P2_R1233_U105 P2_U3016 ; P2_U4596
g5139 not P2_U3402 ; P2_U4597
g5140 nand P2_R1275_U15 P2_U3031 ; P2_U4598
g5141 nand P2_U3030 P2_U3058 ; P2_U4599
g5142 nand P2_R1215_U105 P2_U3028 ; P2_U4600
g5143 nand P2_U3972 P2_U4132 ; P2_U4601
g5144 nand P2_U3727 P2_U4597 ; P2_U4602
g5145 nand P2_U3024 P2_REG2_REG_26__SCAN_IN ; P2_U4603
g5146 nand P2_U3025 P2_REG1_REG_26__SCAN_IN ; P2_U4604
g5147 nand P2_U3026 P2_REG0_REG_26__SCAN_IN ; P2_U4605
g5148 nand P2_ADD_609_U57 P2_U3023 ; P2_U4606
g5149 not P2_U3057 ; P2_U4607
g5150 nand P2_U3038 P2_U3065 ; P2_U4608
g5151 nand P2_R1146_U91 P2_U3955 ; P2_U4609
g5152 nand P2_R1113_U91 P2_U3015 ; P2_U4610
g5153 nand P2_R1131_U104 P2_U3014 ; P2_U4611
g5154 nand P2_R1179_U91 P2_U3018 ; P2_U4612
g5155 nand P2_R1203_U91 P2_U3963 ; P2_U4613
g5156 nand P2_R1164_U104 P2_U3959 ; P2_U4614
g5157 nand P2_R1233_U104 P2_U3016 ; P2_U4615
g5158 not P2_U3404 ; P2_U4616
g5159 nand P2_R1275_U74 P2_U3031 ; P2_U4617
g5160 nand P2_U3030 P2_U3057 ; P2_U4618
g5161 nand P2_R1215_U104 P2_U3028 ; P2_U4619
g5162 nand P2_U3971 P2_U4132 ; P2_U4620
g5163 nand P2_U3731 P2_U4616 ; P2_U4621
g5164 nand P2_U3024 P2_REG2_REG_27__SCAN_IN ; P2_U4622
g5165 nand P2_U3025 P2_REG1_REG_27__SCAN_IN ; P2_U4623
g5166 nand P2_U3026 P2_REG0_REG_27__SCAN_IN ; P2_U4624
g5167 nand P2_ADD_609_U56 P2_U3023 ; P2_U4625
g5168 not P2_U3053 ; P2_U4626
g5169 nand P2_U3038 P2_U3058 ; P2_U4627
g5170 nand P2_R1146_U105 P2_U3955 ; P2_U4628
g5171 nand P2_R1113_U105 P2_U3015 ; P2_U4629
g5172 nand P2_R1131_U15 P2_U3014 ; P2_U4630
g5173 nand P2_R1179_U105 P2_U3018 ; P2_U4631
g5174 nand P2_R1203_U105 P2_U3963 ; P2_U4632
g5175 nand P2_R1164_U15 P2_U3959 ; P2_U4633
g5176 nand P2_R1233_U15 P2_U3016 ; P2_U4634
g5177 not P2_U3406 ; P2_U4635
g5178 nand P2_R1275_U16 P2_U3031 ; P2_U4636
g5179 nand P2_U3030 P2_U3053 ; P2_U4637
g5180 nand P2_R1215_U15 P2_U3028 ; P2_U4638
g5181 nand P2_U3970 P2_U4132 ; P2_U4639
g5182 nand P2_U3735 P2_U4635 ; P2_U4640
g5183 nand P2_U3024 P2_REG2_REG_28__SCAN_IN ; P2_U4641
g5184 nand P2_U3025 P2_REG1_REG_28__SCAN_IN ; P2_U4642
g5185 nand P2_U3026 P2_REG0_REG_28__SCAN_IN ; P2_U4643
g5186 nand P2_ADD_609_U55 P2_U3023 ; P2_U4644
g5187 not P2_U3054 ; P2_U4645
g5188 nand P2_U3038 P2_U3057 ; P2_U4646
g5189 nand P2_R1146_U14 P2_U3955 ; P2_U4647
g5190 nand P2_R1113_U14 P2_U3015 ; P2_U4648
g5191 nand P2_R1131_U103 P2_U3014 ; P2_U4649
g5192 nand P2_R1179_U14 P2_U3018 ; P2_U4650
g5193 nand P2_R1203_U14 P2_U3963 ; P2_U4651
g5194 nand P2_R1164_U103 P2_U3959 ; P2_U4652
g5195 nand P2_R1233_U103 P2_U3016 ; P2_U4653
g5196 not P2_U3408 ; P2_U4654
g5197 nand P2_R1275_U72 P2_U3031 ; P2_U4655
g5198 nand P2_U3030 P2_U3054 ; P2_U4656
g5199 nand P2_R1215_U103 P2_U3028 ; P2_U4657
g5200 nand P2_U3969 P2_U4132 ; P2_U4658
g5201 nand P2_U3739 P2_U4654 ; P2_U4659
g5202 nand P2_ADD_609_U5 P2_U3023 ; P2_U4660
g5203 nand P2_U3024 P2_REG2_REG_29__SCAN_IN ; P2_U4661
g5204 nand P2_U3025 P2_REG1_REG_29__SCAN_IN ; P2_U4662
g5205 nand P2_U3026 P2_REG0_REG_29__SCAN_IN ; P2_U4663
g5206 not P2_U3055 ; P2_U4664
g5207 nand P2_U3038 P2_U3053 ; P2_U4665
g5208 nand P2_R1146_U90 P2_U3955 ; P2_U4666
g5209 nand P2_R1113_U90 P2_U3015 ; P2_U4667
g5210 nand P2_R1131_U102 P2_U3014 ; P2_U4668
g5211 nand P2_R1179_U90 P2_U3018 ; P2_U4669
g5212 nand P2_R1203_U90 P2_U3963 ; P2_U4670
g5213 nand P2_R1164_U102 P2_U3959 ; P2_U4671
g5214 nand P2_R1233_U102 P2_U3016 ; P2_U4672
g5215 not P2_U3410 ; P2_U4673
g5216 nand P2_R1275_U17 P2_U3031 ; P2_U4674
g5217 nand P2_U3030 P2_U3055 ; P2_U4675
g5218 nand P2_R1215_U102 P2_U3028 ; P2_U4676
g5219 nand P2_U3968 P2_U4132 ; P2_U4677
g5220 nand P2_U3742 P2_U4673 ; P2_U4678
g5221 nand P2_U3024 P2_REG2_REG_30__SCAN_IN ; P2_U4679
g5222 nand P2_U3025 P2_REG1_REG_30__SCAN_IN ; P2_U4680
g5223 nand P2_U3026 P2_REG0_REG_30__SCAN_IN ; P2_U4681
g5224 not P2_U3059 ; P2_U4682
g5225 nand P2_U5728 P2_U3360 ; P2_U4683
g5226 nand P2_U3909 P2_U4683 ; P2_U4684
g5227 nand P2_U3743 P2_U3059 ; P2_U4685
g5228 nand P2_U3038 P2_U3054 ; P2_U4686
g5229 nand P2_R1146_U15 P2_U3955 ; P2_U4687
g5230 nand P2_R1113_U15 P2_U3015 ; P2_U4688
g5231 nand P2_R1131_U101 P2_U3014 ; P2_U4689
g5232 nand P2_R1179_U15 P2_U3018 ; P2_U4690
g5233 nand P2_R1203_U15 P2_U3963 ; P2_U4691
g5234 nand P2_R1164_U101 P2_U3959 ; P2_U4692
g5235 nand P2_R1233_U101 P2_U3016 ; P2_U4693
g5236 not P2_U3412 ; P2_U4694
g5237 nand P2_R1275_U70 P2_U3031 ; P2_U4695
g5238 nand P2_R1215_U101 P2_U3028 ; P2_U4696
g5239 nand P2_U3979 P2_U4132 ; P2_U4697
g5240 nand P2_U3747 P2_U4694 ; P2_U4698
g5241 nand P2_U3024 P2_REG2_REG_31__SCAN_IN ; P2_U4699
g5242 nand P2_U3025 P2_REG1_REG_31__SCAN_IN ; P2_U4700
g5243 nand P2_U3026 P2_REG0_REG_31__SCAN_IN ; P2_U4701
g5244 not P2_U3056 ; P2_U4702
g5245 nand P2_R1275_U19 P2_U3031 ; P2_U4703
g5246 nand P2_U3978 P2_U4132 ; P2_U4704
g5247 nand P2_U4704 P2_U3942 P2_U4703 ; P2_U4705
g5248 nand P2_R1275_U68 P2_U3031 ; P2_U4706
g5249 nand P2_U3977 P2_U4132 ; P2_U4707
g5250 nand P2_U4707 P2_U3942 P2_U4706 ; P2_U4708
g5251 nand P2_U3982 P2_U3439 ; P2_U4709
g5252 nand P2_U3020 P2_U3750 ; P2_U4710
g5253 nand P2_U3418 P2_U4710 ; P2_U4711
g5254 nand P2_U3019 P2_U5708 ; P2_U4712
g5255 nand P2_U3958 P2_U4712 ; P2_U4713
g5256 nand P2_U3040 P2_U3078 ; P2_U4714
g5257 nand P2_U3037 P2_R1215_U95 ; P2_U4715
g5258 nand P2_U3036 P2_REG3_REG_0__SCAN_IN ; P2_U4716
g5259 nand P2_U3035 P2_U3448 ; P2_U4717
g5260 nand P2_U3034 P2_U3448 ; P2_U4718
g5261 nand P2_U3040 P2_U3068 ; P2_U4719
g5262 nand P2_U3037 P2_R1215_U94 ; P2_U4720
g5263 nand P2_U3036 P2_REG3_REG_1__SCAN_IN ; P2_U4721
g5264 nand P2_U3035 P2_U3453 ; P2_U4722
g5265 nand P2_U3034 P2_R1275_U55 ; P2_U4723
g5266 nand P2_U3040 P2_U3064 ; P2_U4724
g5267 nand P2_U3037 P2_R1215_U16 ; P2_U4725
g5268 nand P2_U3036 P2_REG3_REG_2__SCAN_IN ; P2_U4726
g5269 nand P2_U3035 P2_U3456 ; P2_U4727
g5270 nand P2_U3034 P2_R1275_U18 ; P2_U4728
g5271 nand P2_U3040 P2_U3060 ; P2_U4729
g5272 nand P2_U3037 P2_R1215_U100 ; P2_U4730
g5273 nand P2_U3036 P2_ADD_609_U4 ; P2_U4731
g5274 nand P2_U3035 P2_U3459 ; P2_U4732
g5275 nand P2_U3034 P2_R1275_U20 ; P2_U4733
g5276 nand P2_U3040 P2_U3067 ; P2_U4734
g5277 nand P2_U3037 P2_R1215_U99 ; P2_U4735
g5278 nand P2_U3036 P2_ADD_609_U54 ; P2_U4736
g5279 nand P2_U3035 P2_U3462 ; P2_U4737
g5280 nand P2_U3034 P2_R1275_U21 ; P2_U4738
g5281 nand P2_U3040 P2_U3071 ; P2_U4739
g5282 nand P2_U3037 P2_R1215_U17 ; P2_U4740
g5283 nand P2_U3036 P2_ADD_609_U53 ; P2_U4741
g5284 nand P2_U3035 P2_U3465 ; P2_U4742
g5285 nand P2_U3034 P2_R1275_U65 ; P2_U4743
g5286 nand P2_U3040 P2_U3070 ; P2_U4744
g5287 nand P2_U3037 P2_R1215_U98 ; P2_U4745
g5288 nand P2_U3036 P2_ADD_609_U52 ; P2_U4746
g5289 nand P2_U3035 P2_U3468 ; P2_U4747
g5290 nand P2_U3034 P2_R1275_U22 ; P2_U4748
g5291 nand P2_U3040 P2_U3084 ; P2_U4749
g5292 nand P2_U3037 P2_R1215_U18 ; P2_U4750
g5293 nand P2_U3036 P2_ADD_609_U51 ; P2_U4751
g5294 nand P2_U3035 P2_U3471 ; P2_U4752
g5295 nand P2_U3034 P2_R1275_U23 ; P2_U4753
g5296 nand P2_U3040 P2_U3083 ; P2_U4754
g5297 nand P2_U3037 P2_R1215_U97 ; P2_U4755
g5298 nand P2_U3036 P2_ADD_609_U50 ; P2_U4756
g5299 nand P2_U3035 P2_U3474 ; P2_U4757
g5300 nand P2_U3034 P2_R1275_U24 ; P2_U4758
g5301 nand P2_U3040 P2_U3062 ; P2_U4759
g5302 nand P2_U3037 P2_R1215_U96 ; P2_U4760
g5303 nand P2_U3036 P2_ADD_609_U49 ; P2_U4761
g5304 nand P2_U3035 P2_U3477 ; P2_U4762
g5305 nand P2_U3034 P2_R1275_U63 ; P2_U4763
g5306 nand P2_U3040 P2_U3063 ; P2_U4764
g5307 nand P2_U3037 P2_R1215_U10 ; P2_U4765
g5308 nand P2_U3036 P2_ADD_609_U73 ; P2_U4766
g5309 nand P2_U3035 P2_U3480 ; P2_U4767
g5310 nand P2_U3034 P2_R1275_U6 ; P2_U4768
g5311 nand P2_U3040 P2_U3072 ; P2_U4769
g5312 nand P2_U3037 P2_R1215_U114 ; P2_U4770
g5313 nand P2_U3036 P2_ADD_609_U72 ; P2_U4771
g5314 nand P2_U3035 P2_U3483 ; P2_U4772
g5315 nand P2_U3034 P2_R1275_U7 ; P2_U4773
g5316 nand P2_U3040 P2_U3080 ; P2_U4774
g5317 nand P2_U3037 P2_R1215_U113 ; P2_U4775
g5318 nand P2_U3036 P2_ADD_609_U71 ; P2_U4776
g5319 nand P2_U3035 P2_U3486 ; P2_U4777
g5320 nand P2_U3034 P2_R1275_U8 ; P2_U4778
g5321 nand P2_U3040 P2_U3079 ; P2_U4779
g5322 nand P2_U3037 P2_R1215_U11 ; P2_U4780
g5323 nand P2_U3036 P2_ADD_609_U70 ; P2_U4781
g5324 nand P2_U3035 P2_U3489 ; P2_U4782
g5325 nand P2_U3034 P2_R1275_U86 ; P2_U4783
g5326 nand P2_U3040 P2_U3074 ; P2_U4784
g5327 nand P2_U3037 P2_R1215_U112 ; P2_U4785
g5328 nand P2_U3036 P2_ADD_609_U69 ; P2_U4786
g5329 nand P2_U3035 P2_U3492 ; P2_U4787
g5330 nand P2_U3034 P2_R1275_U9 ; P2_U4788
g5331 nand P2_U3040 P2_U3073 ; P2_U4789
g5332 nand P2_U3037 P2_R1215_U111 ; P2_U4790
g5333 nand P2_U3036 P2_ADD_609_U68 ; P2_U4791
g5334 nand P2_U3035 P2_U3495 ; P2_U4792
g5335 nand P2_U3034 P2_R1275_U10 ; P2_U4793
g5336 nand P2_U3040 P2_U3069 ; P2_U4794
g5337 nand P2_U3037 P2_R1215_U110 ; P2_U4795
g5338 nand P2_U3036 P2_ADD_609_U67 ; P2_U4796
g5339 nand P2_U3035 P2_U3498 ; P2_U4797
g5340 nand P2_U3034 P2_R1275_U11 ; P2_U4798
g5341 nand P2_U3040 P2_U3082 ; P2_U4799
g5342 nand P2_U3037 P2_R1215_U12 ; P2_U4800
g5343 nand P2_U3036 P2_ADD_609_U66 ; P2_U4801
g5344 nand P2_U3035 P2_U3501 ; P2_U4802
g5345 nand P2_U3034 P2_R1275_U84 ; P2_U4803
g5346 nand P2_U3040 P2_U3081 ; P2_U4804
g5347 nand P2_U3037 P2_R1215_U109 ; P2_U4805
g5348 nand P2_U3036 P2_ADD_609_U65 ; P2_U4806
g5349 nand P2_U3035 P2_U3504 ; P2_U4807
g5350 nand P2_U3034 P2_R1275_U12 ; P2_U4808
g5351 nand P2_U3040 P2_U3076 ; P2_U4809
g5352 nand P2_U3037 P2_R1215_U108 ; P2_U4810
g5353 nand P2_U3036 P2_ADD_609_U64 ; P2_U4811
g5354 nand P2_U3035 P2_U3506 ; P2_U4812
g5355 nand P2_U3034 P2_R1275_U82 ; P2_U4813
g5356 nand P2_U3040 P2_U3075 ; P2_U4814
g5357 nand P2_U3037 P2_R1215_U13 ; P2_U4815
g5358 nand P2_U3036 P2_ADD_609_U63 ; P2_U4816
g5359 nand P2_U3035 P2_U3976 ; P2_U4817
g5360 nand P2_U3034 P2_R1275_U13 ; P2_U4818
g5361 nand P2_U3040 P2_U3061 ; P2_U4819
g5362 nand P2_U3037 P2_R1215_U14 ; P2_U4820
g5363 nand P2_U3036 P2_ADD_609_U62 ; P2_U4821
g5364 nand P2_U3035 P2_U3975 ; P2_U4822
g5365 nand P2_U3034 P2_R1275_U78 ; P2_U4823
g5366 nand P2_U3040 P2_U3066 ; P2_U4824
g5367 nand P2_U3037 P2_R1215_U107 ; P2_U4825
g5368 nand P2_U3036 P2_ADD_609_U61 ; P2_U4826
g5369 nand P2_U3035 P2_U3974 ; P2_U4827
g5370 nand P2_U3034 P2_R1275_U14 ; P2_U4828
g5371 nand P2_U3040 P2_U3065 ; P2_U4829
g5372 nand P2_U3037 P2_R1215_U106 ; P2_U4830
g5373 nand P2_U3036 P2_ADD_609_U60 ; P2_U4831
g5374 nand P2_U3035 P2_U3973 ; P2_U4832
g5375 nand P2_U3034 P2_R1275_U76 ; P2_U4833
g5376 nand P2_U3040 P2_U3058 ; P2_U4834
g5377 nand P2_U3037 P2_R1215_U105 ; P2_U4835
g5378 nand P2_U3036 P2_ADD_609_U59 ; P2_U4836
g5379 nand P2_U3035 P2_U3972 ; P2_U4837
g5380 nand P2_U3034 P2_R1275_U15 ; P2_U4838
g5381 nand P2_U3040 P2_U3057 ; P2_U4839
g5382 nand P2_U3037 P2_R1215_U104 ; P2_U4840
g5383 nand P2_U3036 P2_ADD_609_U58 ; P2_U4841
g5384 nand P2_U3035 P2_U3971 ; P2_U4842
g5385 nand P2_U3034 P2_R1275_U74 ; P2_U4843
g5386 nand P2_U3040 P2_U3053 ; P2_U4844
g5387 nand P2_U3037 P2_R1215_U15 ; P2_U4845
g5388 nand P2_U3036 P2_ADD_609_U57 ; P2_U4846
g5389 nand P2_U3035 P2_U3970 ; P2_U4847
g5390 nand P2_U3034 P2_R1275_U16 ; P2_U4848
g5391 nand P2_U3040 P2_U3054 ; P2_U4849
g5392 nand P2_U3037 P2_R1215_U103 ; P2_U4850
g5393 nand P2_U3036 P2_ADD_609_U56 ; P2_U4851
g5394 nand P2_U3035 P2_U3969 ; P2_U4852
g5395 nand P2_U3034 P2_R1275_U72 ; P2_U4853
g5396 nand P2_U3040 P2_U3055 ; P2_U4854
g5397 nand P2_U3037 P2_R1215_U102 ; P2_U4855
g5398 nand P2_U3036 P2_ADD_609_U55 ; P2_U4856
g5399 nand P2_U3035 P2_U3968 ; P2_U4857
g5400 nand P2_U3034 P2_R1275_U17 ; P2_U4858
g5401 nand P2_U3037 P2_R1215_U101 ; P2_U4859
g5402 nand P2_U3036 P2_ADD_609_U5 ; P2_U4860
g5403 nand P2_U3035 P2_U3979 ; P2_U4861
g5404 nand P2_U3034 P2_R1275_U70 ; P2_U4862
g5405 nand P2_U3035 P2_U3978 ; P2_U4863
g5406 nand P2_U3034 P2_R1275_U19 ; P2_U4864
g5407 nand P2_U3035 P2_U3977 ; P2_U4865
g5408 nand P2_U3034 P2_R1275_U68 ; P2_U4866
g5409 nand P2_R1170_U13 P2_U3022 ; P2_U4867
g5410 nand P2_U5728 P2_U3445 ; P2_U4868
g5411 nand P2_R1209_U13 P2_U5733 ; P2_U4869
g5412 nand P2_U4868 P2_U4867 P2_U4869 ; P2_U4870
g5413 nand P2_R1170_U13 P2_U3022 ; P2_U4871
g5414 nand P2_U3021 P2_R1209_U13 ; P2_U4872
g5415 nand P2_U5728 P2_U3445 ; P2_U4873
g5416 nand P2_U4872 P2_U4871 P2_U4873 ; P2_U4874
g5417 not P2_U3424 ; P2_U4875
g5418 nand P2_U3045 P2_U4870 ; P2_U4876
g5419 nand P2_U3966 P2_U4874 ; P2_U4877
g5420 nand P2_U3044 P2_R1170_U13 ; P2_U4878
g5421 nand P2_U3152 P2_REG3_REG_19__SCAN_IN ; P2_U4879
g5422 nand P2_U3043 P2_U3445 ; P2_U4880
g5423 nand P2_U3042 P2_R1209_U13 ; P2_U4881
g5424 nand P2_U4875 P2_ADDR_REG_19__SCAN_IN ; P2_U4882
g5425 nand P2_R1170_U75 P2_U3022 ; P2_U4883
g5426 nand P2_U5728 P2_U3503 ; P2_U4884
g5427 nand P2_R1209_U75 P2_U5733 ; P2_U4885
g5428 nand P2_U4884 P2_U4883 P2_U4885 ; P2_U4886
g5429 nand P2_R1170_U75 P2_U3022 ; P2_U4887
g5430 nand P2_R1209_U75 P2_U3021 ; P2_U4888
g5431 nand P2_U5728 P2_U3503 ; P2_U4889
g5432 nand P2_U4888 P2_U4887 P2_U4889 ; P2_U4890
g5433 nand P2_U3045 P2_U4886 ; P2_U4891
g5434 nand P2_U3966 P2_U4890 ; P2_U4892
g5435 nand P2_R1170_U75 P2_U3044 ; P2_U4893
g5436 nand P2_U3152 P2_REG3_REG_18__SCAN_IN ; P2_U4894
g5437 nand P2_U3043 P2_U3503 ; P2_U4895
g5438 nand P2_R1209_U75 P2_U3042 ; P2_U4896
g5439 nand P2_U4875 P2_ADDR_REG_18__SCAN_IN ; P2_U4897
g5440 nand P2_R1170_U12 P2_U3022 ; P2_U4898
g5441 nand P2_U5728 P2_U3500 ; P2_U4899
g5442 nand P2_R1209_U12 P2_U5733 ; P2_U4900
g5443 nand P2_U4899 P2_U4898 P2_U4900 ; P2_U4901
g5444 nand P2_R1170_U12 P2_U3022 ; P2_U4902
g5445 nand P2_R1209_U12 P2_U3021 ; P2_U4903
g5446 nand P2_U5728 P2_U3500 ; P2_U4904
g5447 nand P2_U4903 P2_U4902 P2_U4904 ; P2_U4905
g5448 nand P2_U3045 P2_U4901 ; P2_U4906
g5449 nand P2_U3966 P2_U4905 ; P2_U4907
g5450 nand P2_R1170_U12 P2_U3044 ; P2_U4908
g5451 nand P2_U3152 P2_REG3_REG_17__SCAN_IN ; P2_U4909
g5452 nand P2_U3043 P2_U3500 ; P2_U4910
g5453 nand P2_R1209_U12 P2_U3042 ; P2_U4911
g5454 nand P2_U4875 P2_ADDR_REG_17__SCAN_IN ; P2_U4912
g5455 nand P2_R1170_U76 P2_U3022 ; P2_U4913
g5456 nand P2_U5728 P2_U3497 ; P2_U4914
g5457 nand P2_R1209_U76 P2_U5733 ; P2_U4915
g5458 nand P2_U4914 P2_U4913 P2_U4915 ; P2_U4916
g5459 nand P2_R1170_U76 P2_U3022 ; P2_U4917
g5460 nand P2_R1209_U76 P2_U3021 ; P2_U4918
g5461 nand P2_U5728 P2_U3497 ; P2_U4919
g5462 nand P2_U4918 P2_U4917 P2_U4919 ; P2_U4920
g5463 nand P2_U3045 P2_U4916 ; P2_U4921
g5464 nand P2_U3966 P2_U4920 ; P2_U4922
g5465 nand P2_R1170_U76 P2_U3044 ; P2_U4923
g5466 nand P2_U3152 P2_REG3_REG_16__SCAN_IN ; P2_U4924
g5467 nand P2_U3043 P2_U3497 ; P2_U4925
g5468 nand P2_R1209_U76 P2_U3042 ; P2_U4926
g5469 nand P2_U4875 P2_ADDR_REG_16__SCAN_IN ; P2_U4927
g5470 nand P2_R1170_U77 P2_U3022 ; P2_U4928
g5471 nand P2_U5728 P2_U3494 ; P2_U4929
g5472 nand P2_R1209_U77 P2_U5733 ; P2_U4930
g5473 nand P2_U4929 P2_U4928 P2_U4930 ; P2_U4931
g5474 nand P2_R1170_U77 P2_U3022 ; P2_U4932
g5475 nand P2_R1209_U77 P2_U3021 ; P2_U4933
g5476 nand P2_U5728 P2_U3494 ; P2_U4934
g5477 nand P2_U4933 P2_U4932 P2_U4934 ; P2_U4935
g5478 nand P2_U3045 P2_U4931 ; P2_U4936
g5479 nand P2_U3966 P2_U4935 ; P2_U4937
g5480 nand P2_R1170_U77 P2_U3044 ; P2_U4938
g5481 nand P2_U3152 P2_REG3_REG_15__SCAN_IN ; P2_U4939
g5482 nand P2_U3043 P2_U3494 ; P2_U4940
g5483 nand P2_R1209_U77 P2_U3042 ; P2_U4941
g5484 nand P2_U4875 P2_ADDR_REG_15__SCAN_IN ; P2_U4942
g5485 nand P2_R1170_U78 P2_U3022 ; P2_U4943
g5486 nand P2_U5728 P2_U3491 ; P2_U4944
g5487 nand P2_R1209_U78 P2_U5733 ; P2_U4945
g5488 nand P2_U4944 P2_U4943 P2_U4945 ; P2_U4946
g5489 nand P2_R1170_U78 P2_U3022 ; P2_U4947
g5490 nand P2_R1209_U78 P2_U3021 ; P2_U4948
g5491 nand P2_U5728 P2_U3491 ; P2_U4949
g5492 nand P2_U4948 P2_U4947 P2_U4949 ; P2_U4950
g5493 nand P2_U3045 P2_U4946 ; P2_U4951
g5494 nand P2_U3966 P2_U4950 ; P2_U4952
g5495 nand P2_R1170_U78 P2_U3044 ; P2_U4953
g5496 nand P2_U3152 P2_REG3_REG_14__SCAN_IN ; P2_U4954
g5497 nand P2_U3043 P2_U3491 ; P2_U4955
g5498 nand P2_R1209_U78 P2_U3042 ; P2_U4956
g5499 nand P2_U4875 P2_ADDR_REG_14__SCAN_IN ; P2_U4957
g5500 nand P2_R1170_U11 P2_U3022 ; P2_U4958
g5501 nand P2_U5728 P2_U3488 ; P2_U4959
g5502 nand P2_R1209_U11 P2_U5733 ; P2_U4960
g5503 nand P2_U4959 P2_U4958 P2_U4960 ; P2_U4961
g5504 nand P2_R1170_U11 P2_U3022 ; P2_U4962
g5505 nand P2_R1209_U11 P2_U3021 ; P2_U4963
g5506 nand P2_U5728 P2_U3488 ; P2_U4964
g5507 nand P2_U4963 P2_U4962 P2_U4964 ; P2_U4965
g5508 nand P2_U3045 P2_U4961 ; P2_U4966
g5509 nand P2_U3966 P2_U4965 ; P2_U4967
g5510 nand P2_R1170_U11 P2_U3044 ; P2_U4968
g5511 nand P2_U3152 P2_REG3_REG_13__SCAN_IN ; P2_U4969
g5512 nand P2_U3043 P2_U3488 ; P2_U4970
g5513 nand P2_R1209_U11 P2_U3042 ; P2_U4971
g5514 nand P2_U4875 P2_ADDR_REG_13__SCAN_IN ; P2_U4972
g5515 nand P2_R1170_U79 P2_U3022 ; P2_U4973
g5516 nand P2_U5728 P2_U3485 ; P2_U4974
g5517 nand P2_R1209_U79 P2_U5733 ; P2_U4975
g5518 nand P2_U4974 P2_U4973 P2_U4975 ; P2_U4976
g5519 nand P2_R1170_U79 P2_U3022 ; P2_U4977
g5520 nand P2_R1209_U79 P2_U3021 ; P2_U4978
g5521 nand P2_U5728 P2_U3485 ; P2_U4979
g5522 nand P2_U4978 P2_U4977 P2_U4979 ; P2_U4980
g5523 nand P2_U3045 P2_U4976 ; P2_U4981
g5524 nand P2_U3966 P2_U4980 ; P2_U4982
g5525 nand P2_R1170_U79 P2_U3044 ; P2_U4983
g5526 nand P2_U3152 P2_REG3_REG_12__SCAN_IN ; P2_U4984
g5527 nand P2_U3043 P2_U3485 ; P2_U4985
g5528 nand P2_R1209_U79 P2_U3042 ; P2_U4986
g5529 nand P2_U4875 P2_ADDR_REG_12__SCAN_IN ; P2_U4987
g5530 nand P2_R1170_U80 P2_U3022 ; P2_U4988
g5531 nand P2_U5728 P2_U3482 ; P2_U4989
g5532 nand P2_R1209_U80 P2_U5733 ; P2_U4990
g5533 nand P2_U4989 P2_U4988 P2_U4990 ; P2_U4991
g5534 nand P2_R1170_U80 P2_U3022 ; P2_U4992
g5535 nand P2_R1209_U80 P2_U3021 ; P2_U4993
g5536 nand P2_U5728 P2_U3482 ; P2_U4994
g5537 nand P2_U4993 P2_U4992 P2_U4994 ; P2_U4995
g5538 nand P2_U3045 P2_U4991 ; P2_U4996
g5539 nand P2_U3966 P2_U4995 ; P2_U4997
g5540 nand P2_R1170_U80 P2_U3044 ; P2_U4998
g5541 nand P2_U3152 P2_REG3_REG_11__SCAN_IN ; P2_U4999
g5542 nand P2_U3043 P2_U3482 ; P2_U5000
g5543 nand P2_R1209_U80 P2_U3042 ; P2_U5001
g5544 nand P2_U4875 P2_ADDR_REG_11__SCAN_IN ; P2_U5002
g5545 nand P2_R1170_U10 P2_U3022 ; P2_U5003
g5546 nand P2_U5728 P2_U3479 ; P2_U5004
g5547 nand P2_R1209_U10 P2_U5733 ; P2_U5005
g5548 nand P2_U5004 P2_U5003 P2_U5005 ; P2_U5006
g5549 nand P2_R1170_U10 P2_U3022 ; P2_U5007
g5550 nand P2_R1209_U10 P2_U3021 ; P2_U5008
g5551 nand P2_U5728 P2_U3479 ; P2_U5009
g5552 nand P2_U5008 P2_U5007 P2_U5009 ; P2_U5010
g5553 nand P2_U3045 P2_U5006 ; P2_U5011
g5554 nand P2_U3966 P2_U5010 ; P2_U5012
g5555 nand P2_R1170_U10 P2_U3044 ; P2_U5013
g5556 nand P2_U3152 P2_REG3_REG_10__SCAN_IN ; P2_U5014
g5557 nand P2_U3043 P2_U3479 ; P2_U5015
g5558 nand P2_R1209_U10 P2_U3042 ; P2_U5016
g5559 nand P2_U4875 P2_ADDR_REG_10__SCAN_IN ; P2_U5017
g5560 nand P2_R1170_U70 P2_U3022 ; P2_U5018
g5561 nand P2_U5728 P2_U3476 ; P2_U5019
g5562 nand P2_R1209_U70 P2_U5733 ; P2_U5020
g5563 nand P2_U5019 P2_U5018 P2_U5020 ; P2_U5021
g5564 nand P2_R1170_U70 P2_U3022 ; P2_U5022
g5565 nand P2_R1209_U70 P2_U3021 ; P2_U5023
g5566 nand P2_U5728 P2_U3476 ; P2_U5024
g5567 nand P2_U5023 P2_U5022 P2_U5024 ; P2_U5025
g5568 nand P2_U3045 P2_U5021 ; P2_U5026
g5569 nand P2_U3966 P2_U5025 ; P2_U5027
g5570 nand P2_R1170_U70 P2_U3044 ; P2_U5028
g5571 nand P2_U3152 P2_REG3_REG_9__SCAN_IN ; P2_U5029
g5572 nand P2_U3043 P2_U3476 ; P2_U5030
g5573 nand P2_R1209_U70 P2_U3042 ; P2_U5031
g5574 nand P2_U4875 P2_ADDR_REG_9__SCAN_IN ; P2_U5032
g5575 nand P2_R1170_U71 P2_U3022 ; P2_U5033
g5576 nand P2_U5728 P2_U3473 ; P2_U5034
g5577 nand P2_R1209_U71 P2_U5733 ; P2_U5035
g5578 nand P2_U5034 P2_U5033 P2_U5035 ; P2_U5036
g5579 nand P2_R1170_U71 P2_U3022 ; P2_U5037
g5580 nand P2_R1209_U71 P2_U3021 ; P2_U5038
g5581 nand P2_U5728 P2_U3473 ; P2_U5039
g5582 nand P2_U5038 P2_U5037 P2_U5039 ; P2_U5040
g5583 nand P2_U3045 P2_U5036 ; P2_U5041
g5584 nand P2_U3966 P2_U5040 ; P2_U5042
g5585 nand P2_R1170_U71 P2_U3044 ; P2_U5043
g5586 nand P2_U3152 P2_REG3_REG_8__SCAN_IN ; P2_U5044
g5587 nand P2_U3043 P2_U3473 ; P2_U5045
g5588 nand P2_R1209_U71 P2_U3042 ; P2_U5046
g5589 nand P2_U4875 P2_ADDR_REG_8__SCAN_IN ; P2_U5047
g5590 nand P2_R1170_U16 P2_U3022 ; P2_U5048
g5591 nand P2_U5728 P2_U3470 ; P2_U5049
g5592 nand P2_R1209_U16 P2_U5733 ; P2_U5050
g5593 nand P2_U5049 P2_U5048 P2_U5050 ; P2_U5051
g5594 nand P2_R1170_U16 P2_U3022 ; P2_U5052
g5595 nand P2_R1209_U16 P2_U3021 ; P2_U5053
g5596 nand P2_U5728 P2_U3470 ; P2_U5054
g5597 nand P2_U5053 P2_U5052 P2_U5054 ; P2_U5055
g5598 nand P2_U3045 P2_U5051 ; P2_U5056
g5599 nand P2_U3966 P2_U5055 ; P2_U5057
g5600 nand P2_R1170_U16 P2_U3044 ; P2_U5058
g5601 nand P2_U3152 P2_REG3_REG_7__SCAN_IN ; P2_U5059
g5602 nand P2_U3043 P2_U3470 ; P2_U5060
g5603 nand P2_R1209_U16 P2_U3042 ; P2_U5061
g5604 nand P2_U4875 P2_ADDR_REG_7__SCAN_IN ; P2_U5062
g5605 nand P2_R1170_U72 P2_U3022 ; P2_U5063
g5606 nand P2_U5728 P2_U3467 ; P2_U5064
g5607 nand P2_R1209_U72 P2_U5733 ; P2_U5065
g5608 nand P2_U5064 P2_U5063 P2_U5065 ; P2_U5066
g5609 nand P2_R1170_U72 P2_U3022 ; P2_U5067
g5610 nand P2_R1209_U72 P2_U3021 ; P2_U5068
g5611 nand P2_U5728 P2_U3467 ; P2_U5069
g5612 nand P2_U5068 P2_U5067 P2_U5069 ; P2_U5070
g5613 nand P2_U3045 P2_U5066 ; P2_U5071
g5614 nand P2_U3966 P2_U5070 ; P2_U5072
g5615 nand P2_R1170_U72 P2_U3044 ; P2_U5073
g5616 nand P2_U3152 P2_REG3_REG_6__SCAN_IN ; P2_U5074
g5617 nand P2_U3043 P2_U3467 ; P2_U5075
g5618 nand P2_R1209_U72 P2_U3042 ; P2_U5076
g5619 nand P2_U4875 P2_ADDR_REG_6__SCAN_IN ; P2_U5077
g5620 nand P2_R1170_U15 P2_U3022 ; P2_U5078
g5621 nand P2_U5728 P2_U3464 ; P2_U5079
g5622 nand P2_R1209_U15 P2_U5733 ; P2_U5080
g5623 nand P2_U5079 P2_U5078 P2_U5080 ; P2_U5081
g5624 nand P2_R1170_U15 P2_U3022 ; P2_U5082
g5625 nand P2_R1209_U15 P2_U3021 ; P2_U5083
g5626 nand P2_U5728 P2_U3464 ; P2_U5084
g5627 nand P2_U5083 P2_U5082 P2_U5084 ; P2_U5085
g5628 nand P2_U3045 P2_U5081 ; P2_U5086
g5629 nand P2_U3966 P2_U5085 ; P2_U5087
g5630 nand P2_R1170_U15 P2_U3044 ; P2_U5088
g5631 nand P2_U3152 P2_REG3_REG_5__SCAN_IN ; P2_U5089
g5632 nand P2_U3043 P2_U3464 ; P2_U5090
g5633 nand P2_R1209_U15 P2_U3042 ; P2_U5091
g5634 nand P2_U4875 P2_ADDR_REG_5__SCAN_IN ; P2_U5092
g5635 nand P2_R1170_U73 P2_U3022 ; P2_U5093
g5636 nand P2_U5728 P2_U3461 ; P2_U5094
g5637 nand P2_R1209_U73 P2_U5733 ; P2_U5095
g5638 nand P2_U5094 P2_U5093 P2_U5095 ; P2_U5096
g5639 nand P2_R1170_U73 P2_U3022 ; P2_U5097
g5640 nand P2_R1209_U73 P2_U3021 ; P2_U5098
g5641 nand P2_U5728 P2_U3461 ; P2_U5099
g5642 nand P2_U5098 P2_U5097 P2_U5099 ; P2_U5100
g5643 nand P2_U3045 P2_U5096 ; P2_U5101
g5644 nand P2_U3966 P2_U5100 ; P2_U5102
g5645 nand P2_R1170_U73 P2_U3044 ; P2_U5103
g5646 nand P2_U3152 P2_REG3_REG_4__SCAN_IN ; P2_U5104
g5647 nand P2_U3043 P2_U3461 ; P2_U5105
g5648 nand P2_R1209_U73 P2_U3042 ; P2_U5106
g5649 nand P2_U4875 P2_ADDR_REG_4__SCAN_IN ; P2_U5107
g5650 nand P2_R1170_U74 P2_U3022 ; P2_U5108
g5651 nand P2_U5728 P2_U3458 ; P2_U5109
g5652 nand P2_R1209_U74 P2_U5733 ; P2_U5110
g5653 nand P2_U5109 P2_U5108 P2_U5110 ; P2_U5111
g5654 nand P2_R1170_U74 P2_U3022 ; P2_U5112
g5655 nand P2_R1209_U74 P2_U3021 ; P2_U5113
g5656 nand P2_U5728 P2_U3458 ; P2_U5114
g5657 nand P2_U5113 P2_U5112 P2_U5114 ; P2_U5115
g5658 nand P2_U3045 P2_U5111 ; P2_U5116
g5659 nand P2_U3966 P2_U5115 ; P2_U5117
g5660 nand P2_R1170_U74 P2_U3044 ; P2_U5118
g5661 nand P2_U3152 P2_REG3_REG_3__SCAN_IN ; P2_U5119
g5662 nand P2_U3043 P2_U3458 ; P2_U5120
g5663 nand P2_R1209_U74 P2_U3042 ; P2_U5121
g5664 nand P2_U4875 P2_ADDR_REG_3__SCAN_IN ; P2_U5122
g5665 nand P2_R1170_U14 P2_U3022 ; P2_U5123
g5666 nand P2_U5728 P2_U3455 ; P2_U5124
g5667 nand P2_R1209_U14 P2_U5733 ; P2_U5125
g5668 nand P2_U5124 P2_U5123 P2_U5125 ; P2_U5126
g5669 nand P2_R1170_U14 P2_U3022 ; P2_U5127
g5670 nand P2_R1209_U14 P2_U3021 ; P2_U5128
g5671 nand P2_U5728 P2_U3455 ; P2_U5129
g5672 nand P2_U5128 P2_U5127 P2_U5129 ; P2_U5130
g5673 nand P2_U3045 P2_U5126 ; P2_U5131
g5674 nand P2_U3966 P2_U5130 ; P2_U5132
g5675 nand P2_R1170_U14 P2_U3044 ; P2_U5133
g5676 nand P2_U3152 P2_REG3_REG_2__SCAN_IN ; P2_U5134
g5677 nand P2_U3043 P2_U3455 ; P2_U5135
g5678 nand P2_R1209_U14 P2_U3042 ; P2_U5136
g5679 nand P2_U4875 P2_ADDR_REG_2__SCAN_IN ; P2_U5137
g5680 nand P2_R1170_U68 P2_U3022 ; P2_U5138
g5681 nand P2_U5728 P2_U3452 ; P2_U5139
g5682 nand P2_R1209_U68 P2_U5733 ; P2_U5140
g5683 nand P2_U5139 P2_U5138 P2_U5140 ; P2_U5141
g5684 nand P2_R1170_U68 P2_U3022 ; P2_U5142
g5685 nand P2_R1209_U68 P2_U3021 ; P2_U5143
g5686 nand P2_U5728 P2_U3452 ; P2_U5144
g5687 nand P2_U5143 P2_U5142 P2_U5144 ; P2_U5145
g5688 nand P2_U3045 P2_U5141 ; P2_U5146
g5689 nand P2_U3966 P2_U5145 ; P2_U5147
g5690 nand P2_R1170_U68 P2_U3044 ; P2_U5148
g5691 nand P2_U3152 P2_REG3_REG_1__SCAN_IN ; P2_U5149
g5692 nand P2_U3043 P2_U3452 ; P2_U5150
g5693 nand P2_R1209_U68 P2_U3042 ; P2_U5151
g5694 nand P2_U4875 P2_ADDR_REG_1__SCAN_IN ; P2_U5152
g5695 nand P2_R1170_U69 P2_U3022 ; P2_U5153
g5696 nand P2_U5728 P2_U3446 ; P2_U5154
g5697 nand P2_R1209_U69 P2_U5733 ; P2_U5155
g5698 nand P2_U3869 P2_U5153 ; P2_U5156
g5699 nand P2_R1170_U69 P2_U3022 ; P2_U5157
g5700 nand P2_R1209_U69 P2_U3021 ; P2_U5158
g5701 nand P2_U5728 P2_U3446 ; P2_U5159
g5702 nand P2_U5158 P2_U5157 P2_U5159 ; P2_U5160
g5703 nand P2_U3045 P2_U5156 ; P2_U5161
g5704 nand P2_U3966 P2_U5160 ; P2_U5162
g5705 nand P2_R1170_U69 P2_U3044 ; P2_U5163
g5706 nand P2_U3152 P2_REG3_REG_0__SCAN_IN ; P2_U5164
g5707 nand P2_U3043 P2_U3446 ; P2_U5165
g5708 nand P2_R1209_U69 P2_U3042 ; P2_U5166
g5709 nand P2_U4875 P2_ADDR_REG_0__SCAN_IN ; P2_U5167
g5710 not P2_U3947 ; P2_U5168
g5711 nand P2_U3363 P2_U3416 ; P2_U5169
g5712 nand P2_U3366 P2_U3428 ; P2_U5170
g5713 nand P2_U3419 P2_U3364 ; P2_U5171
g5714 nand P2_U6099 P2_U6098 P2_U3018 ; P2_U5172
g5715 nand P2_R1340_U6 P2_U5171 ; P2_U5173
g5716 nand P2_U6201 P2_U6200 P2_U3946 P2_U3885 ; P2_U5174
g5717 nand P2_U6101 P2_U6100 P2_U3052 ; P2_U5175
g5718 nand P2_U3980 P2_U3027 ; P2_U5176
g5719 nand P2_U5175 P2_B_REG_SCAN_IN ; P2_U5177
g5720 nand P2_U3041 P2_U3079 ; P2_U5178
g5721 nand P2_U3039 P2_U3073 ; P2_U5179
g5722 nand P2_ADD_609_U68 P2_U3427 ; P2_U5180
g5723 nand P2_U5179 P2_U5178 P2_U5180 ; P2_U5181
g5724 nand P2_U3014 P2_U5717 ; P2_U5182
g5725 nand P2_U3369 P2_U3367 P2_U5182 P2_U3888 P2_U3419 ; P2_U5183
g5726 nand P2_U5183 P2_U3427 ; P2_U5184
g5727 not P2_U3430 ; P2_U5185
g5728 nand P2_U3495 P2_U5678 ; P2_U5186
g5729 nand P2_ADD_609_U68 P2_U5677 ; P2_U5187
g5730 nand P2_U3988 P2_U5181 ; P2_U5188
g5731 nand P2_R1176_U102 P2_U3032 ; P2_U5189
g5732 nand P2_U3152 P2_REG3_REG_15__SCAN_IN ; P2_U5190
g5733 nand P2_U3041 P2_U3058 ; P2_U5191
g5734 nand P2_U3039 P2_U3053 ; P2_U5192
g5735 nand P2_ADD_609_U57 P2_U3427 ; P2_U5193
g5736 nand P2_U5193 P2_U5191 P2_U5192 ; P2_U5194
g5737 nand P2_U4713 P2_U3427 ; P2_U5195
g5738 nand P2_U5185 P2_U5195 ; P2_U5196
g5739 nand P2_U3965 P2_U4713 ; P2_U5197
g5740 nand P2_U3418 P2_U5197 ; P2_U5198
g5741 nand P2_U3047 P2_U3970 ; P2_U5199
g5742 nand P2_U3046 P2_ADD_609_U57 ; P2_U5200
g5743 nand P2_U3988 P2_U5194 ; P2_U5201
g5744 nand P2_R1176_U12 P2_U3032 ; P2_U5202
g5745 nand P2_U3152 P2_REG3_REG_26__SCAN_IN ; P2_U5203
g5746 nand P2_U3041 P2_U3067 ; P2_U5204
g5747 nand P2_U3039 P2_U3070 ; P2_U5205
g5748 nand P2_ADD_609_U52 P2_U3427 ; P2_U5206
g5749 nand P2_U5205 P2_U5204 P2_U5206 ; P2_U5207
g5750 nand P2_U3468 P2_U5678 ; P2_U5208
g5751 nand P2_ADD_609_U52 P2_U5677 ; P2_U5209
g5752 nand P2_U3988 P2_U5207 ; P2_U5210
g5753 nand P2_R1176_U87 P2_U3032 ; P2_U5211
g5754 nand P2_U3152 P2_REG3_REG_6__SCAN_IN ; P2_U5212
g5755 nand P2_U3041 P2_U3069 ; P2_U5213
g5756 nand P2_U3039 P2_U3081 ; P2_U5214
g5757 nand P2_ADD_609_U65 P2_U3427 ; P2_U5215
g5758 nand P2_U5214 P2_U5213 P2_U5215 ; P2_U5216
g5759 nand P2_U3504 P2_U5678 ; P2_U5217
g5760 nand P2_ADD_609_U65 P2_U5677 ; P2_U5218
g5761 nand P2_U3988 P2_U5216 ; P2_U5219
g5762 nand P2_R1176_U100 P2_U3032 ; P2_U5220
g5763 nand P2_U3152 P2_REG3_REG_18__SCAN_IN ; P2_U5221
g5764 nand P2_U3041 P2_U3078 ; P2_U5222
g5765 nand P2_U3039 P2_U3064 ; P2_U5223
g5766 nand P2_U3427 P2_REG3_REG_2__SCAN_IN ; P2_U5224
g5767 nand P2_U5223 P2_U5222 P2_U5224 ; P2_U5225
g5768 nand P2_U3456 P2_U5678 ; P2_U5226
g5769 nand P2_U5677 P2_REG3_REG_2__SCAN_IN ; P2_U5227
g5770 nand P2_U3988 P2_U5225 ; P2_U5228
g5771 nand P2_R1176_U90 P2_U3032 ; P2_U5229
g5772 nand P2_U3152 P2_REG3_REG_2__SCAN_IN ; P2_U5230
g5773 nand P2_U3041 P2_U3062 ; P2_U5231
g5774 nand P2_U3039 P2_U3072 ; P2_U5232
g5775 nand P2_ADD_609_U72 P2_U3427 ; P2_U5233
g5776 nand P2_U5232 P2_U5231 P2_U5233 ; P2_U5234
g5777 nand P2_U3483 P2_U5678 ; P2_U5235
g5778 nand P2_ADD_609_U72 P2_U5677 ; P2_U5236
g5779 nand P2_U3988 P2_U5234 ; P2_U5237
g5780 nand P2_R1176_U105 P2_U3032 ; P2_U5238
g5781 nand P2_U3152 P2_REG3_REG_11__SCAN_IN ; P2_U5239
g5782 nand P2_U3041 P2_U3075 ; P2_U5240
g5783 nand P2_U3039 P2_U3066 ; P2_U5241
g5784 nand P2_ADD_609_U61 P2_U3427 ; P2_U5242
g5785 nand P2_U5242 P2_U5240 P2_U5241 ; P2_U5243
g5786 nand P2_U3047 P2_U3974 ; P2_U5244
g5787 nand P2_U3046 P2_ADD_609_U61 ; P2_U5245
g5788 nand P2_U3988 P2_U5243 ; P2_U5246
g5789 nand P2_R1176_U96 P2_U3032 ; P2_U5247
g5790 nand P2_U3152 P2_REG3_REG_22__SCAN_IN ; P2_U5248
g5791 nand P2_U3041 P2_U3072 ; P2_U5249
g5792 nand P2_U3039 P2_U3079 ; P2_U5250
g5793 nand P2_ADD_609_U70 P2_U3427 ; P2_U5251
g5794 nand P2_U5250 P2_U5249 P2_U5251 ; P2_U5252
g5795 nand P2_U3489 P2_U5678 ; P2_U5253
g5796 nand P2_ADD_609_U70 P2_U5677 ; P2_U5254
g5797 nand P2_U3988 P2_U5252 ; P2_U5255
g5798 nand P2_R1176_U9 P2_U3032 ; P2_U5256
g5799 nand P2_U3152 P2_REG3_REG_13__SCAN_IN ; P2_U5257
g5800 nand P2_U3041 P2_U3081 ; P2_U5258
g5801 nand P2_U3039 P2_U3075 ; P2_U5259
g5802 nand P2_ADD_609_U63 P2_U3427 ; P2_U5260
g5803 nand P2_U5259 P2_U5258 P2_U5260 ; P2_U5261
g5804 nand P2_U3047 P2_U3976 ; P2_U5262
g5805 nand P2_U3046 P2_ADD_609_U63 ; P2_U5263
g5806 nand P2_U3988 P2_U5261 ; P2_U5264
g5807 nand P2_R1176_U97 P2_U3032 ; P2_U5265
g5808 nand P2_U3152 P2_REG3_REG_20__SCAN_IN ; P2_U5266
g5809 nand P2_U3429 P2_U3426 ; P2_U5267
g5810 nand P2_U5267 P2_U3427 ; P2_U5268
g5811 nand P2_U3989 P2_U5268 ; P2_U5269
g5812 nand P2_U3893 P2_U3039 ; P2_U5270
g5813 nand P2_U3448 P2_U5678 ; P2_U5271
g5814 nand P2_U5269 P2_REG3_REG_0__SCAN_IN ; P2_U5272
g5815 nand P2_R1176_U84 P2_U3032 ; P2_U5273
g5816 nand P2_U3152 P2_REG3_REG_0__SCAN_IN ; P2_U5274
g5817 nand P2_U3041 P2_U3084 ; P2_U5275
g5818 nand P2_U3039 P2_U3062 ; P2_U5276
g5819 nand P2_ADD_609_U49 P2_U3427 ; P2_U5277
g5820 nand P2_U5276 P2_U5275 P2_U5277 ; P2_U5278
g5821 nand P2_U3477 P2_U5678 ; P2_U5279
g5822 nand P2_ADD_609_U49 P2_U5677 ; P2_U5280
g5823 nand P2_U3988 P2_U5278 ; P2_U5281
g5824 nand P2_R1176_U85 P2_U3032 ; P2_U5282
g5825 nand P2_U3152 P2_REG3_REG_9__SCAN_IN ; P2_U5283
g5826 nand P2_U3041 P2_U3064 ; P2_U5284
g5827 nand P2_U3039 P2_U3067 ; P2_U5285
g5828 nand P2_ADD_609_U54 P2_U3427 ; P2_U5286
g5829 nand P2_U5285 P2_U5284 P2_U5286 ; P2_U5287
g5830 nand P2_U3462 P2_U5678 ; P2_U5288
g5831 nand P2_ADD_609_U54 P2_U5677 ; P2_U5289
g5832 nand P2_U3988 P2_U5287 ; P2_U5290
g5833 nand P2_R1176_U89 P2_U3032 ; P2_U5291
g5834 nand P2_U3152 P2_REG3_REG_4__SCAN_IN ; P2_U5292
g5835 nand P2_U3041 P2_U3066 ; P2_U5293
g5836 nand P2_U3039 P2_U3058 ; P2_U5294
g5837 nand P2_ADD_609_U59 P2_U3427 ; P2_U5295
g5838 nand P2_U5295 P2_U5293 P2_U5294 ; P2_U5296
g5839 nand P2_U3047 P2_U3972 ; P2_U5297
g5840 nand P2_U3046 P2_ADD_609_U59 ; P2_U5298
g5841 nand P2_U3988 P2_U5296 ; P2_U5299
g5842 nand P2_R1176_U94 P2_U3032 ; P2_U5300
g5843 nand P2_U3152 P2_REG3_REG_24__SCAN_IN ; P2_U5301
g5844 nand P2_U3041 P2_U3073 ; P2_U5302
g5845 nand P2_U3039 P2_U3082 ; P2_U5303
g5846 nand P2_ADD_609_U66 P2_U3427 ; P2_U5304
g5847 nand P2_U5303 P2_U5302 P2_U5304 ; P2_U5305
g5848 nand P2_U3501 P2_U5678 ; P2_U5306
g5849 nand P2_ADD_609_U66 P2_U5677 ; P2_U5307
g5850 nand P2_U3988 P2_U5305 ; P2_U5308
g5851 nand P2_R1176_U10 P2_U3032 ; P2_U5309
g5852 nand P2_U3152 P2_REG3_REG_17__SCAN_IN ; P2_U5310
g5853 nand P2_U3041 P2_U3060 ; P2_U5311
g5854 nand P2_U3039 P2_U3071 ; P2_U5312
g5855 nand P2_ADD_609_U53 P2_U3427 ; P2_U5313
g5856 nand P2_U5312 P2_U5311 P2_U5313 ; P2_U5314
g5857 nand P2_U3465 P2_U5678 ; P2_U5315
g5858 nand P2_ADD_609_U53 P2_U5677 ; P2_U5316
g5859 nand P2_U3988 P2_U5314 ; P2_U5317
g5860 nand P2_R1176_U88 P2_U3032 ; P2_U5318
g5861 nand P2_U3152 P2_REG3_REG_5__SCAN_IN ; P2_U5319
g5862 nand P2_U3041 P2_U3074 ; P2_U5320
g5863 nand P2_U3039 P2_U3069 ; P2_U5321
g5864 nand P2_ADD_609_U67 P2_U3427 ; P2_U5322
g5865 nand P2_U5321 P2_U5320 P2_U5322 ; P2_U5323
g5866 nand P2_U3498 P2_U5678 ; P2_U5324
g5867 nand P2_ADD_609_U67 P2_U5677 ; P2_U5325
g5868 nand P2_U3988 P2_U5323 ; P2_U5326
g5869 nand P2_R1176_U101 P2_U3032 ; P2_U5327
g5870 nand P2_U3152 P2_REG3_REG_16__SCAN_IN ; P2_U5328
g5871 nand P2_U3041 P2_U3065 ; P2_U5329
g5872 nand P2_U3039 P2_U3057 ; P2_U5330
g5873 nand P2_ADD_609_U58 P2_U3427 ; P2_U5331
g5874 nand P2_U5331 P2_U5329 P2_U5330 ; P2_U5332
g5875 nand P2_U3047 P2_U3971 ; P2_U5333
g5876 nand P2_U3046 P2_ADD_609_U58 ; P2_U5334
g5877 nand P2_U3988 P2_U5332 ; P2_U5335
g5878 nand P2_R1176_U93 P2_U3032 ; P2_U5336
g5879 nand P2_U3152 P2_REG3_REG_25__SCAN_IN ; P2_U5337
g5880 nand P2_U3041 P2_U3063 ; P2_U5338
g5881 nand P2_U3039 P2_U3080 ; P2_U5339
g5882 nand P2_ADD_609_U71 P2_U3427 ; P2_U5340
g5883 nand P2_U5339 P2_U5338 P2_U5340 ; P2_U5341
g5884 nand P2_U3486 P2_U5678 ; P2_U5342
g5885 nand P2_ADD_609_U71 P2_U5677 ; P2_U5343
g5886 nand P2_U3988 P2_U5341 ; P2_U5344
g5887 nand P2_R1176_U104 P2_U3032 ; P2_U5345
g5888 nand P2_U3152 P2_REG3_REG_12__SCAN_IN ; P2_U5346
g5889 nand P2_U3041 P2_U3076 ; P2_U5347
g5890 nand P2_U3039 P2_U3061 ; P2_U5348
g5891 nand P2_ADD_609_U62 P2_U3427 ; P2_U5349
g5892 nand P2_U5348 P2_U5347 P2_U5349 ; P2_U5350
g5893 nand P2_U3047 P2_U3975 ; P2_U5351
g5894 nand P2_U3046 P2_ADD_609_U62 ; P2_U5352
g5895 nand P2_U3988 P2_U5350 ; P2_U5353
g5896 nand P2_R1176_U11 P2_U3032 ; P2_U5354
g5897 nand P2_U3152 P2_REG3_REG_21__SCAN_IN ; P2_U5355
g5898 nand P2_U3041 P2_U3077 ; P2_U5356
g5899 nand P2_U3039 P2_U3068 ; P2_U5357
g5900 nand P2_U3427 P2_REG3_REG_1__SCAN_IN ; P2_U5358
g5901 nand P2_U5357 P2_U5356 P2_U5358 ; P2_U5359
g5902 nand P2_U3453 P2_U5678 ; P2_U5360
g5903 nand P2_U5677 P2_REG3_REG_1__SCAN_IN ; P2_U5361
g5904 nand P2_U3988 P2_U5359 ; P2_U5362
g5905 nand P2_R1176_U98 P2_U3032 ; P2_U5363
g5906 nand P2_U3152 P2_REG3_REG_1__SCAN_IN ; P2_U5364
g5907 nand P2_U3041 P2_U3070 ; P2_U5365
g5908 nand P2_U3039 P2_U3083 ; P2_U5366
g5909 nand P2_ADD_609_U50 P2_U3427 ; P2_U5367
g5910 nand P2_U5366 P2_U5365 P2_U5367 ; P2_U5368
g5911 nand P2_U3474 P2_U5678 ; P2_U5369
g5912 nand P2_ADD_609_U50 P2_U5677 ; P2_U5370
g5913 nand P2_U3988 P2_U5368 ; P2_U5371
g5914 nand P2_R1176_U86 P2_U3032 ; P2_U5372
g5915 nand P2_U3152 P2_REG3_REG_8__SCAN_IN ; P2_U5373
g5916 nand P2_U3041 P2_U3053 ; P2_U5374
g5917 nand P2_U3039 P2_U3055 ; P2_U5375
g5918 nand P2_ADD_609_U55 P2_U3427 ; P2_U5376
g5919 nand P2_U5375 P2_U5376 P2_U5374 ; P2_U5377
g5920 nand P2_U3047 P2_U3968 ; P2_U5378
g5921 nand P2_U3046 P2_ADD_609_U55 ; P2_U5379
g5922 nand P2_U3988 P2_U5377 ; P2_U5380
g5923 nand P2_R1176_U91 P2_U3032 ; P2_U5381
g5924 nand P2_U3152 P2_REG3_REG_28__SCAN_IN ; P2_U5382
g5925 nand P2_U3041 P2_U3082 ; P2_U5383
g5926 nand P2_U3039 P2_U3076 ; P2_U5384
g5927 nand P2_ADD_609_U64 P2_U3427 ; P2_U5385
g5928 nand P2_U5384 P2_U5383 P2_U5385 ; P2_U5386
g5929 nand P2_U3506 P2_U5678 ; P2_U5387
g5930 nand P2_ADD_609_U64 P2_U5677 ; P2_U5388
g5931 nand P2_U3988 P2_U5386 ; P2_U5389
g5932 nand P2_R1176_U99 P2_U3032 ; P2_U5390
g5933 nand P2_U3152 P2_REG3_REG_19__SCAN_IN ; P2_U5391
g5934 nand P2_U3041 P2_U3068 ; P2_U5392
g5935 nand P2_U3039 P2_U3060 ; P2_U5393
g5936 nand P2_ADD_609_U4 P2_U3427 ; P2_U5394
g5937 nand P2_U5393 P2_U5392 P2_U5394 ; P2_U5395
g5938 nand P2_U3459 P2_U5678 ; P2_U5396
g5939 nand P2_ADD_609_U4 P2_U5677 ; P2_U5397
g5940 nand P2_U3988 P2_U5395 ; P2_U5398
g5941 nand P2_R1176_U13 P2_U3032 ; P2_U5399
g5942 nand P2_U3152 P2_REG3_REG_3__SCAN_IN ; P2_U5400
g5943 nand P2_U3041 P2_U3083 ; P2_U5401
g5944 nand P2_U3039 P2_U3063 ; P2_U5402
g5945 nand P2_ADD_609_U73 P2_U3427 ; P2_U5403
g5946 nand P2_U5402 P2_U5401 P2_U5403 ; P2_U5404
g5947 nand P2_U3480 P2_U5678 ; P2_U5405
g5948 nand P2_ADD_609_U73 P2_U5677 ; P2_U5406
g5949 nand P2_U3988 P2_U5404 ; P2_U5407
g5950 nand P2_R1176_U106 P2_U3032 ; P2_U5408
g5951 nand P2_U3152 P2_REG3_REG_10__SCAN_IN ; P2_U5409
g5952 nand P2_U3041 P2_U3061 ; P2_U5410
g5953 nand P2_U3039 P2_U3065 ; P2_U5411
g5954 nand P2_ADD_609_U60 P2_U3427 ; P2_U5412
g5955 nand P2_U5412 P2_U5410 P2_U5411 ; P2_U5413
g5956 nand P2_U3047 P2_U3973 ; P2_U5414
g5957 nand P2_U3046 P2_ADD_609_U60 ; P2_U5415
g5958 nand P2_U3988 P2_U5413 ; P2_U5416
g5959 nand P2_R1176_U95 P2_U3032 ; P2_U5417
g5960 nand P2_U3152 P2_REG3_REG_23__SCAN_IN ; P2_U5418
g5961 nand P2_U3041 P2_U3080 ; P2_U5419
g5962 nand P2_U3039 P2_U3074 ; P2_U5420
g5963 nand P2_ADD_609_U69 P2_U3427 ; P2_U5421
g5964 nand P2_U5420 P2_U5419 P2_U5421 ; P2_U5422
g5965 nand P2_U3492 P2_U5678 ; P2_U5423
g5966 nand P2_ADD_609_U69 P2_U5677 ; P2_U5424
g5967 nand P2_U3988 P2_U5422 ; P2_U5425
g5968 nand P2_R1176_U103 P2_U3032 ; P2_U5426
g5969 nand P2_U3152 P2_REG3_REG_14__SCAN_IN ; P2_U5427
g5970 nand P2_U3041 P2_U3057 ; P2_U5428
g5971 nand P2_U3039 P2_U3054 ; P2_U5429
g5972 nand P2_ADD_609_U56 P2_U3427 ; P2_U5430
g5973 nand P2_U5430 P2_U5428 P2_U5429 ; P2_U5431
g5974 nand P2_U3047 P2_U3969 ; P2_U5432
g5975 nand P2_U3046 P2_ADD_609_U56 ; P2_U5433
g5976 nand P2_U3988 P2_U5431 ; P2_U5434
g5977 nand P2_R1176_U92 P2_U3032 ; P2_U5435
g5978 nand P2_U3152 P2_REG3_REG_27__SCAN_IN ; P2_U5436
g5979 nand P2_U3041 P2_U3071 ; P2_U5437
g5980 nand P2_U3039 P2_U3084 ; P2_U5438
g5981 nand P2_ADD_609_U51 P2_U3427 ; P2_U5439
g5982 nand P2_U5438 P2_U5437 P2_U5439 ; P2_U5440
g5983 nand P2_U3471 P2_U5678 ; P2_U5441
g5984 nand P2_ADD_609_U51 P2_U5677 ; P2_U5442
g5985 nand P2_U3988 P2_U5440 ; P2_U5443
g5986 nand P2_R1176_U14 P2_U3032 ; P2_U5444
g5987 nand P2_U3152 P2_REG3_REG_7__SCAN_IN ; P2_U5445
g5988 nand P2_U3967 P2_U3048 ; P2_U5446
g5989 nand P2_U3436 P2_U3909 ; P2_U5447
g5990 nand P2_U3372 P2_U3366 P2_U3904 ; P2_U5448
g5991 not P2_U3431 ; P2_U5449
g5992 nand P2_U3584 P2_U3431 ; P2_U5450
g5993 nand P2_U5717 P2_U3083 ; P2_U5451
g5994 nand P2_U3585 P2_U3431 ; P2_U5452
g5995 nand P2_U5717 P2_U3084 ; P2_U5453
g5996 nand P2_U3586 P2_U3431 ; P2_U5454
g5997 nand P2_U5717 P2_U3070 ; P2_U5455
g5998 nand P2_U3587 P2_U3431 ; P2_U5456
g5999 nand P2_U5717 P2_U3071 ; P2_U5457
g6000 nand P2_U3588 P2_U3431 ; P2_U5458
g6001 nand P2_U5717 P2_U3067 ; P2_U5459
g6002 nand P2_U3589 P2_U3431 ; P2_U5460
g6003 nand P2_U5717 P2_U3060 ; P2_U5461
g6004 nand P2_U3591 P2_U3431 ; P2_U5462
g6005 nand P2_U5717 P2_U3056 ; P2_U5463
g6006 nand P2_U3592 P2_U3431 ; P2_U5464
g6007 nand P2_U5717 P2_U3059 ; P2_U5465
g6008 nand P2_U3590 P2_U3431 ; P2_U5466
g6009 nand P2_U5717 P2_U3064 ; P2_U5467
g6010 nand P2_U3594 P2_U3431 ; P2_U5468
g6011 nand P2_U5717 P2_U3055 ; P2_U5469
g6012 nand P2_U3595 P2_U3431 ; P2_U5470
g6013 nand P2_U5717 P2_U3054 ; P2_U5471
g6014 nand P2_U3596 P2_U3431 ; P2_U5472
g6015 nand P2_U5717 P2_U3053 ; P2_U5473
g6016 nand P2_U3597 P2_U3431 ; P2_U5474
g6017 nand P2_U5717 P2_U3057 ; P2_U5475
g6018 nand P2_U3598 P2_U3431 ; P2_U5476
g6019 nand P2_U5717 P2_U3058 ; P2_U5477
g6020 nand P2_U3599 P2_U3431 ; P2_U5478
g6021 nand P2_U5717 P2_U3065 ; P2_U5479
g6022 nand P2_U3600 P2_U3431 ; P2_U5480
g6023 nand P2_U5717 P2_U3066 ; P2_U5481
g6024 nand P2_U3601 P2_U3431 ; P2_U5482
g6025 nand P2_U5717 P2_U3061 ; P2_U5483
g6026 nand P2_U3602 P2_U3431 ; P2_U5484
g6027 nand P2_U5717 P2_U3075 ; P2_U5485
g6028 nand P2_U3603 P2_U3431 ; P2_U5486
g6029 nand P2_U5717 P2_U3076 ; P2_U5487
g6030 nand P2_U5717 P2_U3068 ; P2_U5488
g6031 nand P2_U3605 P2_U3431 ; P2_U5489
g6032 nand P2_U5717 P2_U3081 ; P2_U5490
g6033 nand P2_U3606 P2_U3431 ; P2_U5491
g6034 nand P2_U5717 P2_U3082 ; P2_U5492
g6035 nand P2_U3607 P2_U3431 ; P2_U5493
g6036 nand P2_U5717 P2_U3069 ; P2_U5494
g6037 nand P2_U3608 P2_U3431 ; P2_U5495
g6038 nand P2_U5717 P2_U3073 ; P2_U5496
g6039 nand P2_U3609 P2_U3431 ; P2_U5497
g6040 nand P2_U5717 P2_U3074 ; P2_U5498
g6041 nand P2_U3610 P2_U3431 ; P2_U5499
g6042 nand P2_U5717 P2_U3079 ; P2_U5500
g6043 nand P2_U3611 P2_U3431 ; P2_U5501
g6044 nand P2_U5717 P2_U3080 ; P2_U5502
g6045 nand P2_U3612 P2_U3431 ; P2_U5503
g6046 nand P2_U5717 P2_U3072 ; P2_U5504
g6047 nand P2_U3613 P2_U3431 ; P2_U5505
g6048 nand P2_U5717 P2_U3063 ; P2_U5506
g6049 nand P2_U3614 P2_U3431 ; P2_U5507
g6050 nand P2_U5717 P2_U3062 ; P2_U5508
g6051 nand P2_U5717 P2_U3078 ; P2_U5509
g6052 nand P2_U5717 P2_U3077 ; P2_U5510
g6053 nand P2_U5708 P2_U3445 ; P2_U5511
g6054 nand P2_U3436 P2_U5711 ; P2_U5512
g6055 nand P2_U3368 P2_U3950 P2_U3906 ; P2_U5513
g6056 nand P2_U3953 P2_U3477 ; P2_U5514
g6057 nand P2_U5513 P2_U3083 ; P2_U5515
g6058 nand P2_U3953 P2_U3474 ; P2_U5516
g6059 nand P2_U5513 P2_U3084 ; P2_U5517
g6060 nand P2_U3953 P2_U3471 ; P2_U5518
g6061 nand P2_U5513 P2_U3070 ; P2_U5519
g6062 nand P2_U3953 P2_U3468 ; P2_U5520
g6063 nand P2_U5513 P2_U3071 ; P2_U5521
g6064 nand P2_U3953 P2_U3465 ; P2_U5522
g6065 nand P2_U5513 P2_U3067 ; P2_U5523
g6066 nand P2_U3953 P2_U3462 ; P2_U5524
g6067 nand P2_U5513 P2_U3060 ; P2_U5525
g6068 nand P2_U5513 P2_U3056 ; P2_U5526
g6069 nand P2_U3953 P2_U3977 ; P2_U5527
g6070 nand P2_U5513 P2_U3059 ; P2_U5528
g6071 nand P2_U3953 P2_U3459 ; P2_U5529
g6072 nand P2_U5513 P2_U3064 ; P2_U5530
g6073 nand P2_U5513 P2_U3055 ; P2_U5531
g6074 nand P2_U3953 P2_U3979 ; P2_U5532
g6075 nand P2_U5513 P2_U3054 ; P2_U5533
g6076 nand P2_U3953 P2_U3968 ; P2_U5534
g6077 nand P2_U5513 P2_U3053 ; P2_U5535
g6078 nand P2_U3953 P2_U3969 ; P2_U5536
g6079 nand P2_U5513 P2_U3057 ; P2_U5537
g6080 nand P2_U3953 P2_U3970 ; P2_U5538
g6081 nand P2_U5513 P2_U3058 ; P2_U5539
g6082 nand P2_U3953 P2_U3971 ; P2_U5540
g6083 nand P2_U5513 P2_U3065 ; P2_U5541
g6084 nand P2_U3953 P2_U3972 ; P2_U5542
g6085 nand P2_U5513 P2_U3066 ; P2_U5543
g6086 nand P2_U3953 P2_U3973 ; P2_U5544
g6087 nand P2_U5513 P2_U3061 ; P2_U5545
g6088 nand P2_U3953 P2_U3974 ; P2_U5546
g6089 nand P2_U5513 P2_U3075 ; P2_U5547
g6090 nand P2_U3953 P2_U3975 ; P2_U5548
g6091 nand P2_U5513 P2_U3076 ; P2_U5549
g6092 nand P2_U3953 P2_U3976 ; P2_U5550
g6093 nand P2_U3953 P2_U3456 ; P2_U5551
g6094 nand P2_U5513 P2_U3068 ; P2_U5552
g6095 nand P2_U3953 P2_U3506 ; P2_U5553
g6096 nand P2_U5513 P2_U3081 ; P2_U5554
g6097 nand P2_U3953 P2_U3504 ; P2_U5555
g6098 nand P2_U5513 P2_U3082 ; P2_U5556
g6099 nand P2_U3953 P2_U3501 ; P2_U5557
g6100 nand P2_U5513 P2_U3069 ; P2_U5558
g6101 nand P2_U3953 P2_U3498 ; P2_U5559
g6102 nand P2_U5513 P2_U3073 ; P2_U5560
g6103 nand P2_U3953 P2_U3495 ; P2_U5561
g6104 nand P2_U5513 P2_U3074 ; P2_U5562
g6105 nand P2_U3953 P2_U3492 ; P2_U5563
g6106 nand P2_U5513 P2_U3079 ; P2_U5564
g6107 nand P2_U3953 P2_U3489 ; P2_U5565
g6108 nand P2_U5513 P2_U3080 ; P2_U5566
g6109 nand P2_U3953 P2_U3486 ; P2_U5567
g6110 nand P2_U5513 P2_U3072 ; P2_U5568
g6111 nand P2_U3953 P2_U3483 ; P2_U5569
g6112 nand P2_U5513 P2_U3063 ; P2_U5570
g6113 nand P2_U3953 P2_U3480 ; P2_U5571
g6114 nand P2_U5513 P2_U3062 ; P2_U5572
g6115 nand P2_U3953 P2_U3453 ; P2_U5573
g6116 nand P2_U5513 P2_U3078 ; P2_U5574
g6117 nand P2_U3953 P2_U3448 ; P2_U5575
g6118 nand P2_U5513 P2_U3077 ; P2_U5576
g6119 nand P2_U3477 P2_U5513 ; P2_U5577
g6120 nand P2_U3953 P2_U3083 ; P2_U5578
g6121 nand P2_U5701 P2_U3084 ; P2_U5579
g6122 nand P2_U3474 P2_U5513 ; P2_U5580
g6123 nand P2_U3953 P2_U3084 ; P2_U5581
g6124 nand P2_U5701 P2_U3070 ; P2_U5582
g6125 nand P2_U3471 P2_U5513 ; P2_U5583
g6126 nand P2_U3953 P2_U3070 ; P2_U5584
g6127 nand P2_U5701 P2_U3071 ; P2_U5585
g6128 nand P2_U3468 P2_U5513 ; P2_U5586
g6129 nand P2_U3953 P2_U3071 ; P2_U5587
g6130 nand P2_U5701 P2_U3067 ; P2_U5588
g6131 nand P2_U3465 P2_U5513 ; P2_U5589
g6132 nand P2_U3953 P2_U3067 ; P2_U5590
g6133 nand P2_U5701 P2_U3060 ; P2_U5591
g6134 nand P2_U3462 P2_U5513 ; P2_U5592
g6135 nand P2_U3953 P2_U3060 ; P2_U5593
g6136 nand P2_U5701 P2_U3064 ; P2_U5594
g6137 nand P2_U3977 P2_U5513 ; P2_U5595
g6138 nand P2_U3953 P2_U3056 ; P2_U5596
g6139 nand P2_U3978 P2_U5513 ; P2_U5597
g6140 nand P2_U3953 P2_U3059 ; P2_U5598
g6141 nand P2_U3459 P2_U5513 ; P2_U5599
g6142 nand P2_U3953 P2_U3064 ; P2_U5600
g6143 nand P2_U5701 P2_U3068 ; P2_U5601
g6144 nand P2_U3979 P2_U5513 ; P2_U5602
g6145 nand P2_U3953 P2_U3055 ; P2_U5603
g6146 nand P2_U5701 P2_U3054 ; P2_U5604
g6147 nand P2_U3968 P2_U5513 ; P2_U5605
g6148 nand P2_U3953 P2_U3054 ; P2_U5606
g6149 nand P2_U5701 P2_U3053 ; P2_U5607
g6150 nand P2_U3969 P2_U5513 ; P2_U5608
g6151 nand P2_U3953 P2_U3053 ; P2_U5609
g6152 nand P2_U5701 P2_U3057 ; P2_U5610
g6153 nand P2_U3970 P2_U5513 ; P2_U5611
g6154 nand P2_U3953 P2_U3057 ; P2_U5612
g6155 nand P2_U5701 P2_U3058 ; P2_U5613
g6156 nand P2_U3971 P2_U5513 ; P2_U5614
g6157 nand P2_U3953 P2_U3058 ; P2_U5615
g6158 nand P2_U5701 P2_U3065 ; P2_U5616
g6159 nand P2_U3972 P2_U5513 ; P2_U5617
g6160 nand P2_U3953 P2_U3065 ; P2_U5618
g6161 nand P2_U5701 P2_U3066 ; P2_U5619
g6162 nand P2_U3973 P2_U5513 ; P2_U5620
g6163 nand P2_U3953 P2_U3066 ; P2_U5621
g6164 nand P2_U5701 P2_U3061 ; P2_U5622
g6165 nand P2_U3974 P2_U5513 ; P2_U5623
g6166 nand P2_U3953 P2_U3061 ; P2_U5624
g6167 nand P2_U5701 P2_U3075 ; P2_U5625
g6168 nand P2_U3975 P2_U5513 ; P2_U5626
g6169 nand P2_U3953 P2_U3075 ; P2_U5627
g6170 nand P2_U5701 P2_U3076 ; P2_U5628
g6171 nand P2_U3976 P2_U5513 ; P2_U5629
g6172 nand P2_U3953 P2_U3076 ; P2_U5630
g6173 nand P2_U5701 P2_U3081 ; P2_U5631
g6174 nand P2_U3456 P2_U5513 ; P2_U5632
g6175 nand P2_U3953 P2_U3068 ; P2_U5633
g6176 nand P2_U5701 P2_U3078 ; P2_U5634
g6177 nand P2_U3506 P2_U5513 ; P2_U5635
g6178 nand P2_U3953 P2_U3081 ; P2_U5636
g6179 nand P2_U5701 P2_U3082 ; P2_U5637
g6180 nand P2_U3504 P2_U5513 ; P2_U5638
g6181 nand P2_U3953 P2_U3082 ; P2_U5639
g6182 nand P2_U5701 P2_U3069 ; P2_U5640
g6183 nand P2_U3501 P2_U5513 ; P2_U5641
g6184 nand P2_U3953 P2_U3069 ; P2_U5642
g6185 nand P2_U5701 P2_U3073 ; P2_U5643
g6186 nand P2_U3498 P2_U5513 ; P2_U5644
g6187 nand P2_U3953 P2_U3073 ; P2_U5645
g6188 nand P2_U5701 P2_U3074 ; P2_U5646
g6189 nand P2_U3495 P2_U5513 ; P2_U5647
g6190 nand P2_U3953 P2_U3074 ; P2_U5648
g6191 nand P2_U5701 P2_U3079 ; P2_U5649
g6192 nand P2_U3492 P2_U5513 ; P2_U5650
g6193 nand P2_U3953 P2_U3079 ; P2_U5651
g6194 nand P2_U5701 P2_U3080 ; P2_U5652
g6195 nand P2_U3489 P2_U5513 ; P2_U5653
g6196 nand P2_U3953 P2_U3080 ; P2_U5654
g6197 nand P2_U5701 P2_U3072 ; P2_U5655
g6198 nand P2_U3486 P2_U5513 ; P2_U5656
g6199 nand P2_U3953 P2_U3072 ; P2_U5657
g6200 nand P2_U5701 P2_U3063 ; P2_U5658
g6201 nand P2_U3483 P2_U5513 ; P2_U5659
g6202 nand P2_U3953 P2_U3063 ; P2_U5660
g6203 nand P2_U5701 P2_U3062 ; P2_U5661
g6204 nand P2_U3480 P2_U5513 ; P2_U5662
g6205 nand P2_U3953 P2_U3062 ; P2_U5663
g6206 nand P2_U5701 P2_U3083 ; P2_U5664
g6207 nand P2_U3453 P2_U5513 ; P2_U5665
g6208 nand P2_U3953 P2_U3078 ; P2_U5666
g6209 nand P2_U5701 P2_U3077 ; P2_U5667
g6210 nand P2_U3448 P2_U5513 ; P2_U5668
g6211 nand P2_U3953 P2_U3077 ; P2_U5669
g6212 nand P2_U3436 P2_STATE_REG_SCAN_IN ; P2_U5670
g6213 nand P2_U3886 P2_U5177 ; P2_U5671
g6214 nand P2_U5528 P2_U3413 ; P2_U5672
g6215 nand P2_U3432 P2_U5528 ; P2_U5673
g6216 not P2_U3415 ; P2_U5674
g6217 nand P2_U3991 P2_U3427 ; P2_U5675
g6218 nand P2_U3965 P2_U3991 ; P2_U5676
g6219 nand P2_U5675 P2_U3989 ; P2_U5677
g6220 nand P2_U5676 P2_U3990 ; P2_U5678
g6221 nand P2_U6222 P2_U5488 ; P2_U5679
g6222 nand P2_U6245 P2_U5509 ; P2_U5680
g6223 nand P2_U6268 P2_U5510 ; P2_U5681
g6224 nand P2_U5449 P2_U5509 ; P2_U5682
g6225 nand P2_U5449 P2_U5488 ; P2_U5683
g6226 nand P2_U5449 P2_U5510 ; P2_U5684
g6227 nand P2_U5695 P2_U5689 ; P2_U5685
g6228 nand P2_U3436 P2_U3909 ; P2_U5686
g6229 nand P2_U3907 P2_IR_REG_24__SCAN_IN ; P2_U5687
g6230 nand P2_SUB_598_U90 P2_IR_REG_31__SCAN_IN ; P2_U5688
g6231 not P2_U3433 ; P2_U5689
g6232 nand P2_U3907 P2_IR_REG_25__SCAN_IN ; P2_U5690
g6233 nand P2_SUB_598_U22 P2_IR_REG_31__SCAN_IN ; P2_U5691
g6234 not P2_U3434 ; P2_U5692
g6235 nand P2_U3907 P2_IR_REG_26__SCAN_IN ; P2_U5693
g6236 nand P2_SUB_598_U23 P2_IR_REG_31__SCAN_IN ; P2_U5694
g6237 not P2_U3435 ; P2_U5695
g6238 nand P2_U5689 P2_B_REG_SCAN_IN ; P2_U5696
g6239 nand P2_U3433 P2_U3360 ; P2_U5697
g6240 nand P2_U5697 P2_U5696 ; P2_U5698
g6241 nand P2_U3907 P2_IR_REG_23__SCAN_IN ; P2_U5699
g6242 nand P2_SUB_598_U21 P2_IR_REG_31__SCAN_IN ; P2_U5700
g6243 not P2_U3436 ; P2_U5701
g6244 nand P2_U3908 P2_D_REG_0__SCAN_IN ; P2_U5702
g6245 nand P2_U3986 P2_U4095 ; P2_U5703
g6246 nand P2_U3908 P2_D_REG_1__SCAN_IN ; P2_U5704
g6247 nand P2_U3986 P2_U4096 ; P2_U5705
g6248 nand P2_U3907 P2_IR_REG_22__SCAN_IN ; P2_U5706
g6249 nand P2_SUB_598_U20 P2_IR_REG_31__SCAN_IN ; P2_U5707
g6250 not P2_U3441 ; P2_U5708
g6251 nand P2_U3907 P2_IR_REG_19__SCAN_IN ; P2_U5709
g6252 nand P2_SUB_598_U18 P2_IR_REG_31__SCAN_IN ; P2_U5710
g6253 not P2_U3445 ; P2_U5711
g6254 nand P2_U3907 P2_IR_REG_20__SCAN_IN ; P2_U5712
g6255 nand P2_SUB_598_U19 P2_IR_REG_31__SCAN_IN ; P2_U5713
g6256 not P2_U3439 ; P2_U5714
g6257 nand P2_U3907 P2_IR_REG_21__SCAN_IN ; P2_U5715
g6258 nand P2_SUB_598_U92 P2_IR_REG_31__SCAN_IN ; P2_U5716
g6259 not P2_U3440 ; P2_U5717
g6260 nand P2_U3907 P2_IR_REG_30__SCAN_IN ; P2_U5718
g6261 nand P2_SUB_598_U79 P2_IR_REG_31__SCAN_IN ; P2_U5719
g6262 not P2_U3443 ; P2_U5720
g6263 nand P2_U3907 P2_IR_REG_29__SCAN_IN ; P2_U5721
g6264 nand P2_SUB_598_U81 P2_IR_REG_31__SCAN_IN ; P2_U5722
g6265 not P2_U3442 ; P2_U5723
g6266 nand P2_U3443 P2_U5723 P2_REG2_REG_1__SCAN_IN ; P2_U5724
g6267 nand P2_U3443 P2_U3442 P2_REG3_REG_1__SCAN_IN ; P2_U5725
g6268 nand P2_U3907 P2_IR_REG_28__SCAN_IN ; P2_U5726
g6269 nand P2_SUB_598_U84 P2_IR_REG_31__SCAN_IN ; P2_U5727
g6270 not P2_U3444 ; P2_U5728
g6271 nand P2_U3907 P2_IR_REG_0__SCAN_IN ; P2_U5729
g6272 nand P2_IR_REG_0__SCAN_IN P2_IR_REG_31__SCAN_IN ; P2_U5730
g6273 nand P2_U3907 P2_IR_REG_27__SCAN_IN ; P2_U5731
g6274 nand P2_SUB_598_U87 P2_IR_REG_31__SCAN_IN ; P2_U5732
g6275 not P2_U3447 ; P2_U5733
g6276 nand U56 P2_U3909 ; P2_U5734
g6277 nand P2_U3964 P2_U3446 ; P2_U5735
g6278 not P2_U3448 ; P2_U5736
g6279 nand P2_U3441 P2_U5717 ; P2_U5737
g6280 nand P2_U3439 P2_U5708 ; P2_U5738
g6281 nand P2_U4094 P2_D_REG_1__SCAN_IN ; P2_U5739
g6282 nand P2_U4096 P2_U3362 ; P2_U5740
g6283 not P2_U3450 ; P2_U5741
g6284 nand P2_U5685 P2_U3362 ; P2_U5742
g6285 nand P2_U4094 P2_D_REG_0__SCAN_IN ; P2_U5743
g6286 not P2_U3449 ; P2_U5744
g6287 nand P2_U3910 P2_REG0_REG_0__SCAN_IN ; P2_U5745
g6288 nand P2_U3985 P2_U4145 ; P2_U5746
g6289 nand P2_U3443 P2_U5723 P2_REG2_REG_0__SCAN_IN ; P2_U5747
g6290 nand P2_U3443 P2_U3442 P2_REG3_REG_0__SCAN_IN ; P2_U5748
g6291 nand P2_U3907 P2_IR_REG_1__SCAN_IN ; P2_U5749
g6292 nand P2_SUB_598_U49 P2_IR_REG_31__SCAN_IN ; P2_U5750
g6293 nand U45 P2_U3909 ; P2_U5751
g6294 nand P2_U3452 P2_U3964 ; P2_U5752
g6295 not P2_U3453 ; P2_U5753
g6296 nand P2_U3443 P2_U5723 P2_REG2_REG_2__SCAN_IN ; P2_U5754
g6297 nand P2_U3443 P2_U3442 P2_REG3_REG_2__SCAN_IN ; P2_U5755
g6298 nand P2_U3910 P2_REG0_REG_1__SCAN_IN ; P2_U5756
g6299 nand P2_U3985 P2_U4165 ; P2_U5757
g6300 nand P2_U3907 P2_IR_REG_2__SCAN_IN ; P2_U5758
g6301 nand P2_SUB_598_U24 P2_IR_REG_31__SCAN_IN ; P2_U5759
g6302 nand U34 P2_U3909 ; P2_U5760
g6303 nand P2_U3455 P2_U3964 ; P2_U5761
g6304 not P2_U3456 ; P2_U5762
g6305 nand P2_U3910 P2_REG0_REG_2__SCAN_IN ; P2_U5763
g6306 nand P2_U3985 P2_U4184 ; P2_U5764
g6307 nand P2_U3907 P2_IR_REG_3__SCAN_IN ; P2_U5765
g6308 nand P2_SUB_598_U25 P2_IR_REG_31__SCAN_IN ; P2_U5766
g6309 nand U31 P2_U3909 ; P2_U5767
g6310 nand P2_U3458 P2_U3964 ; P2_U5768
g6311 not P2_U3459 ; P2_U5769
g6312 nand P2_U3910 P2_REG0_REG_3__SCAN_IN ; P2_U5770
g6313 nand P2_U3985 P2_U4203 ; P2_U5771
g6314 nand P2_U3907 P2_IR_REG_4__SCAN_IN ; P2_U5772
g6315 nand P2_SUB_598_U26 P2_IR_REG_31__SCAN_IN ; P2_U5773
g6316 nand U30 P2_U3909 ; P2_U5774
g6317 nand P2_U3461 P2_U3964 ; P2_U5775
g6318 not P2_U3462 ; P2_U5776
g6319 nand P2_U3910 P2_REG0_REG_4__SCAN_IN ; P2_U5777
g6320 nand P2_U3985 P2_U4222 ; P2_U5778
g6321 nand P2_U3907 P2_IR_REG_5__SCAN_IN ; P2_U5779
g6322 nand P2_SUB_598_U74 P2_IR_REG_31__SCAN_IN ; P2_U5780
g6323 nand U29 P2_U3909 ; P2_U5781
g6324 nand P2_U3464 P2_U3964 ; P2_U5782
g6325 not P2_U3465 ; P2_U5783
g6326 nand P2_U3910 P2_REG0_REG_5__SCAN_IN ; P2_U5784
g6327 nand P2_U3985 P2_U4241 ; P2_U5785
g6328 nand P2_U3907 P2_IR_REG_6__SCAN_IN ; P2_U5786
g6329 nand P2_SUB_598_U27 P2_IR_REG_31__SCAN_IN ; P2_U5787
g6330 nand U28 P2_U3909 ; P2_U5788
g6331 nand P2_U3467 P2_U3964 ; P2_U5789
g6332 not P2_U3468 ; P2_U5790
g6333 nand P2_U3910 P2_REG0_REG_6__SCAN_IN ; P2_U5791
g6334 nand P2_U3985 P2_U4260 ; P2_U5792
g6335 nand P2_U3907 P2_IR_REG_7__SCAN_IN ; P2_U5793
g6336 nand P2_SUB_598_U28 P2_IR_REG_31__SCAN_IN ; P2_U5794
g6337 nand U27 P2_U3909 ; P2_U5795
g6338 nand P2_U3470 P2_U3964 ; P2_U5796
g6339 not P2_U3471 ; P2_U5797
g6340 nand P2_U3910 P2_REG0_REG_7__SCAN_IN ; P2_U5798
g6341 nand P2_U3985 P2_U4279 ; P2_U5799
g6342 nand P2_U3907 P2_IR_REG_8__SCAN_IN ; P2_U5800
g6343 nand P2_SUB_598_U29 P2_IR_REG_31__SCAN_IN ; P2_U5801
g6344 nand U26 P2_U3909 ; P2_U5802
g6345 nand P2_U3473 P2_U3964 ; P2_U5803
g6346 not P2_U3474 ; P2_U5804
g6347 nand P2_U3910 P2_REG0_REG_8__SCAN_IN ; P2_U5805
g6348 nand P2_U3985 P2_U4298 ; P2_U5806
g6349 nand P2_U3907 P2_IR_REG_9__SCAN_IN ; P2_U5807
g6350 nand P2_SUB_598_U72 P2_IR_REG_31__SCAN_IN ; P2_U5808
g6351 nand U25 P2_U3909 ; P2_U5809
g6352 nand P2_U3476 P2_U3964 ; P2_U5810
g6353 not P2_U3477 ; P2_U5811
g6354 nand P2_U3910 P2_REG0_REG_9__SCAN_IN ; P2_U5812
g6355 nand P2_U3985 P2_U4317 ; P2_U5813
g6356 nand P2_U3907 P2_IR_REG_10__SCAN_IN ; P2_U5814
g6357 nand P2_SUB_598_U11 P2_IR_REG_31__SCAN_IN ; P2_U5815
g6358 nand U55 P2_U3909 ; P2_U5816
g6359 nand P2_U3479 P2_U3964 ; P2_U5817
g6360 not P2_U3480 ; P2_U5818
g6361 nand P2_U3910 P2_REG0_REG_10__SCAN_IN ; P2_U5819
g6362 nand P2_U3985 P2_U4336 ; P2_U5820
g6363 nand P2_U3907 P2_IR_REG_11__SCAN_IN ; P2_U5821
g6364 nand P2_SUB_598_U12 P2_IR_REG_31__SCAN_IN ; P2_U5822
g6365 nand U54 P2_U3909 ; P2_U5823
g6366 nand P2_U3482 P2_U3964 ; P2_U5824
g6367 not P2_U3483 ; P2_U5825
g6368 nand P2_U3910 P2_REG0_REG_11__SCAN_IN ; P2_U5826
g6369 nand P2_U3985 P2_U4355 ; P2_U5827
g6370 nand P2_U3907 P2_IR_REG_12__SCAN_IN ; P2_U5828
g6371 nand P2_SUB_598_U13 P2_IR_REG_31__SCAN_IN ; P2_U5829
g6372 nand U53 P2_U3909 ; P2_U5830
g6373 nand P2_U3485 P2_U3964 ; P2_U5831
g6374 not P2_U3486 ; P2_U5832
g6375 nand P2_U3910 P2_REG0_REG_12__SCAN_IN ; P2_U5833
g6376 nand P2_U3985 P2_U4374 ; P2_U5834
g6377 nand P2_U3907 P2_IR_REG_13__SCAN_IN ; P2_U5835
g6378 nand P2_SUB_598_U99 P2_IR_REG_31__SCAN_IN ; P2_U5836
g6379 nand U52 P2_U3909 ; P2_U5837
g6380 nand P2_U3488 P2_U3964 ; P2_U5838
g6381 not P2_U3489 ; P2_U5839
g6382 nand P2_U3910 P2_REG0_REG_13__SCAN_IN ; P2_U5840
g6383 nand P2_U3985 P2_U4393 ; P2_U5841
g6384 nand P2_U3907 P2_IR_REG_14__SCAN_IN ; P2_U5842
g6385 nand P2_SUB_598_U14 P2_IR_REG_31__SCAN_IN ; P2_U5843
g6386 nand U51 P2_U3909 ; P2_U5844
g6387 nand P2_U3491 P2_U3964 ; P2_U5845
g6388 not P2_U3492 ; P2_U5846
g6389 nand P2_U3910 P2_REG0_REG_14__SCAN_IN ; P2_U5847
g6390 nand P2_U3985 P2_U4412 ; P2_U5848
g6391 nand P2_U3907 P2_IR_REG_15__SCAN_IN ; P2_U5849
g6392 nand P2_SUB_598_U15 P2_IR_REG_31__SCAN_IN ; P2_U5850
g6393 nand U50 P2_U3909 ; P2_U5851
g6394 nand P2_U3494 P2_U3964 ; P2_U5852
g6395 not P2_U3495 ; P2_U5853
g6396 nand P2_U3910 P2_REG0_REG_15__SCAN_IN ; P2_U5854
g6397 nand P2_U3985 P2_U4431 ; P2_U5855
g6398 nand P2_U3907 P2_IR_REG_16__SCAN_IN ; P2_U5856
g6399 nand P2_SUB_598_U16 P2_IR_REG_31__SCAN_IN ; P2_U5857
g6400 nand U49 P2_U3909 ; P2_U5858
g6401 nand P2_U3497 P2_U3964 ; P2_U5859
g6402 not P2_U3498 ; P2_U5860
g6403 nand P2_U3910 P2_REG0_REG_16__SCAN_IN ; P2_U5861
g6404 nand P2_U3985 P2_U4450 ; P2_U5862
g6405 nand P2_U3907 P2_IR_REG_17__SCAN_IN ; P2_U5863
g6406 nand P2_SUB_598_U97 P2_IR_REG_31__SCAN_IN ; P2_U5864
g6407 nand U48 P2_U3909 ; P2_U5865
g6408 nand P2_U3500 P2_U3964 ; P2_U5866
g6409 not P2_U3501 ; P2_U5867
g6410 nand P2_U3910 P2_REG0_REG_17__SCAN_IN ; P2_U5868
g6411 nand P2_U3985 P2_U4469 ; P2_U5869
g6412 nand P2_U3907 P2_IR_REG_18__SCAN_IN ; P2_U5870
g6413 nand P2_SUB_598_U17 P2_IR_REG_31__SCAN_IN ; P2_U5871
g6414 nand U47 P2_U3909 ; P2_U5872
g6415 nand P2_U3503 P2_U3964 ; P2_U5873
g6416 not P2_U3504 ; P2_U5874
g6417 nand P2_U3910 P2_REG0_REG_18__SCAN_IN ; P2_U5875
g6418 nand P2_U3985 P2_U4488 ; P2_U5876
g6419 nand U46 P2_U3909 ; P2_U5877
g6420 nand P2_U3964 P2_U3445 ; P2_U5878
g6421 not P2_U3506 ; P2_U5879
g6422 nand P2_U3910 P2_REG0_REG_19__SCAN_IN ; P2_U5880
g6423 nand P2_U3985 P2_U4507 ; P2_U5881
g6424 nand P2_U3910 P2_REG0_REG_20__SCAN_IN ; P2_U5882
g6425 nand P2_U3985 P2_U4526 ; P2_U5883
g6426 nand P2_U3910 P2_REG0_REG_21__SCAN_IN ; P2_U5884
g6427 nand P2_U3985 P2_U4545 ; P2_U5885
g6428 nand P2_U3910 P2_REG0_REG_22__SCAN_IN ; P2_U5886
g6429 nand P2_U3985 P2_U4564 ; P2_U5887
g6430 nand P2_U3910 P2_REG0_REG_23__SCAN_IN ; P2_U5888
g6431 nand P2_U3985 P2_U4583 ; P2_U5889
g6432 nand P2_U3910 P2_REG0_REG_24__SCAN_IN ; P2_U5890
g6433 nand P2_U3985 P2_U4602 ; P2_U5891
g6434 nand P2_U3910 P2_REG0_REG_25__SCAN_IN ; P2_U5892
g6435 nand P2_U3985 P2_U4621 ; P2_U5893
g6436 nand P2_U3910 P2_REG0_REG_26__SCAN_IN ; P2_U5894
g6437 nand P2_U3985 P2_U4640 ; P2_U5895
g6438 nand P2_U3910 P2_REG0_REG_27__SCAN_IN ; P2_U5896
g6439 nand P2_U3985 P2_U4659 ; P2_U5897
g6440 nand P2_U3910 P2_REG0_REG_28__SCAN_IN ; P2_U5898
g6441 nand P2_U3985 P2_U4678 ; P2_U5899
g6442 nand P2_U3910 P2_REG0_REG_29__SCAN_IN ; P2_U5900
g6443 nand P2_U3985 P2_U4698 ; P2_U5901
g6444 nand P2_U3910 P2_REG0_REG_30__SCAN_IN ; P2_U5902
g6445 nand P2_U3985 P2_U4705 ; P2_U5903
g6446 nand P2_U3910 P2_REG0_REG_31__SCAN_IN ; P2_U5904
g6447 nand P2_U3985 P2_U4708 ; P2_U5905
g6448 nand P2_U3911 P2_REG1_REG_0__SCAN_IN ; P2_U5906
g6449 nand P2_U3984 P2_U4145 ; P2_U5907
g6450 nand P2_U3911 P2_REG1_REG_1__SCAN_IN ; P2_U5908
g6451 nand P2_U3984 P2_U4165 ; P2_U5909
g6452 nand P2_U3911 P2_REG1_REG_2__SCAN_IN ; P2_U5910
g6453 nand P2_U3984 P2_U4184 ; P2_U5911
g6454 nand P2_U3911 P2_REG1_REG_3__SCAN_IN ; P2_U5912
g6455 nand P2_U3984 P2_U4203 ; P2_U5913
g6456 nand P2_U3911 P2_REG1_REG_4__SCAN_IN ; P2_U5914
g6457 nand P2_U3984 P2_U4222 ; P2_U5915
g6458 nand P2_U3911 P2_REG1_REG_5__SCAN_IN ; P2_U5916
g6459 nand P2_U3984 P2_U4241 ; P2_U5917
g6460 nand P2_U3911 P2_REG1_REG_6__SCAN_IN ; P2_U5918
g6461 nand P2_U3984 P2_U4260 ; P2_U5919
g6462 nand P2_U3911 P2_REG1_REG_7__SCAN_IN ; P2_U5920
g6463 nand P2_U3984 P2_U4279 ; P2_U5921
g6464 nand P2_U3911 P2_REG1_REG_8__SCAN_IN ; P2_U5922
g6465 nand P2_U3984 P2_U4298 ; P2_U5923
g6466 nand P2_U3911 P2_REG1_REG_9__SCAN_IN ; P2_U5924
g6467 nand P2_U3984 P2_U4317 ; P2_U5925
g6468 nand P2_U3911 P2_REG1_REG_10__SCAN_IN ; P2_U5926
g6469 nand P2_U3984 P2_U4336 ; P2_U5927
g6470 nand P2_U3911 P2_REG1_REG_11__SCAN_IN ; P2_U5928
g6471 nand P2_U3984 P2_U4355 ; P2_U5929
g6472 nand P2_U3911 P2_REG1_REG_12__SCAN_IN ; P2_U5930
g6473 nand P2_U3984 P2_U4374 ; P2_U5931
g6474 nand P2_U3911 P2_REG1_REG_13__SCAN_IN ; P2_U5932
g6475 nand P2_U3984 P2_U4393 ; P2_U5933
g6476 nand P2_U3911 P2_REG1_REG_14__SCAN_IN ; P2_U5934
g6477 nand P2_U3984 P2_U4412 ; P2_U5935
g6478 nand P2_U3911 P2_REG1_REG_15__SCAN_IN ; P2_U5936
g6479 nand P2_U3984 P2_U4431 ; P2_U5937
g6480 nand P2_U3911 P2_REG1_REG_16__SCAN_IN ; P2_U5938
g6481 nand P2_U3984 P2_U4450 ; P2_U5939
g6482 nand P2_U3911 P2_REG1_REG_17__SCAN_IN ; P2_U5940
g6483 nand P2_U3984 P2_U4469 ; P2_U5941
g6484 nand P2_U3911 P2_REG1_REG_18__SCAN_IN ; P2_U5942
g6485 nand P2_U3984 P2_U4488 ; P2_U5943
g6486 nand P2_U3911 P2_REG1_REG_19__SCAN_IN ; P2_U5944
g6487 nand P2_U3984 P2_U4507 ; P2_U5945
g6488 nand P2_U3911 P2_REG1_REG_20__SCAN_IN ; P2_U5946
g6489 nand P2_U3984 P2_U4526 ; P2_U5947
g6490 nand P2_U3911 P2_REG1_REG_21__SCAN_IN ; P2_U5948
g6491 nand P2_U3984 P2_U4545 ; P2_U5949
g6492 nand P2_U3911 P2_REG1_REG_22__SCAN_IN ; P2_U5950
g6493 nand P2_U3984 P2_U4564 ; P2_U5951
g6494 nand P2_U3911 P2_REG1_REG_23__SCAN_IN ; P2_U5952
g6495 nand P2_U3984 P2_U4583 ; P2_U5953
g6496 nand P2_U3911 P2_REG1_REG_24__SCAN_IN ; P2_U5954
g6497 nand P2_U3984 P2_U4602 ; P2_U5955
g6498 nand P2_U3911 P2_REG1_REG_25__SCAN_IN ; P2_U5956
g6499 nand P2_U3984 P2_U4621 ; P2_U5957
g6500 nand P2_U3911 P2_REG1_REG_26__SCAN_IN ; P2_U5958
g6501 nand P2_U3984 P2_U4640 ; P2_U5959
g6502 nand P2_U3911 P2_REG1_REG_27__SCAN_IN ; P2_U5960
g6503 nand P2_U3984 P2_U4659 ; P2_U5961
g6504 nand P2_U3911 P2_REG1_REG_28__SCAN_IN ; P2_U5962
g6505 nand P2_U3984 P2_U4678 ; P2_U5963
g6506 nand P2_U3911 P2_REG1_REG_29__SCAN_IN ; P2_U5964
g6507 nand P2_U3984 P2_U4698 ; P2_U5965
g6508 nand P2_U3911 P2_REG1_REG_30__SCAN_IN ; P2_U5966
g6509 nand P2_U3984 P2_U4705 ; P2_U5967
g6510 nand P2_U3911 P2_REG1_REG_31__SCAN_IN ; P2_U5968
g6511 nand P2_U3984 P2_U4708 ; P2_U5969
g6512 nand P2_U3417 P2_REG2_REG_0__SCAN_IN ; P2_U5970
g6513 nand P2_U3983 P2_U3373 ; P2_U5971
g6514 nand P2_U3417 P2_REG2_REG_1__SCAN_IN ; P2_U5972
g6515 nand P2_U3983 P2_U3374 ; P2_U5973
g6516 nand P2_U3417 P2_REG2_REG_2__SCAN_IN ; P2_U5974
g6517 nand P2_U3983 P2_U3375 ; P2_U5975
g6518 nand P2_U3417 P2_REG2_REG_3__SCAN_IN ; P2_U5976
g6519 nand P2_U3983 P2_U3376 ; P2_U5977
g6520 nand P2_U3417 P2_REG2_REG_4__SCAN_IN ; P2_U5978
g6521 nand P2_U3983 P2_U3377 ; P2_U5979
g6522 nand P2_U3417 P2_REG2_REG_5__SCAN_IN ; P2_U5980
g6523 nand P2_U3983 P2_U3378 ; P2_U5981
g6524 nand P2_U3417 P2_REG2_REG_6__SCAN_IN ; P2_U5982
g6525 nand P2_U3983 P2_U3379 ; P2_U5983
g6526 nand P2_U3417 P2_REG2_REG_7__SCAN_IN ; P2_U5984
g6527 nand P2_U3983 P2_U3380 ; P2_U5985
g6528 nand P2_U3417 P2_REG2_REG_8__SCAN_IN ; P2_U5986
g6529 nand P2_U3983 P2_U3381 ; P2_U5987
g6530 nand P2_U3417 P2_REG2_REG_9__SCAN_IN ; P2_U5988
g6531 nand P2_U3983 P2_U3382 ; P2_U5989
g6532 nand P2_U3417 P2_REG2_REG_10__SCAN_IN ; P2_U5990
g6533 nand P2_U3983 P2_U3383 ; P2_U5991
g6534 nand P2_U3417 P2_REG2_REG_11__SCAN_IN ; P2_U5992
g6535 nand P2_U3983 P2_U3384 ; P2_U5993
g6536 nand P2_U3417 P2_REG2_REG_12__SCAN_IN ; P2_U5994
g6537 nand P2_U3983 P2_U3385 ; P2_U5995
g6538 nand P2_U3417 P2_REG2_REG_13__SCAN_IN ; P2_U5996
g6539 nand P2_U3983 P2_U3386 ; P2_U5997
g6540 nand P2_U3417 P2_REG2_REG_14__SCAN_IN ; P2_U5998
g6541 nand P2_U3983 P2_U3387 ; P2_U5999
g6542 nand P2_U3417 P2_REG2_REG_15__SCAN_IN ; P2_U6000
g6543 nand P2_U3983 P2_U3388 ; P2_U6001
g6544 nand P2_U3417 P2_REG2_REG_16__SCAN_IN ; P2_U6002
g6545 nand P2_U3983 P2_U3389 ; P2_U6003
g6546 nand P2_U3417 P2_REG2_REG_17__SCAN_IN ; P2_U6004
g6547 nand P2_U3983 P2_U3390 ; P2_U6005
g6548 nand P2_U3417 P2_REG2_REG_18__SCAN_IN ; P2_U6006
g6549 nand P2_U3983 P2_U3391 ; P2_U6007
g6550 nand P2_U3417 P2_REG2_REG_19__SCAN_IN ; P2_U6008
g6551 nand P2_U3983 P2_U3392 ; P2_U6009
g6552 nand P2_U3417 P2_REG2_REG_20__SCAN_IN ; P2_U6010
g6553 nand P2_U3983 P2_U3394 ; P2_U6011
g6554 nand P2_U3417 P2_REG2_REG_21__SCAN_IN ; P2_U6012
g6555 nand P2_U3983 P2_U3396 ; P2_U6013
g6556 nand P2_U3417 P2_REG2_REG_22__SCAN_IN ; P2_U6014
g6557 nand P2_U3983 P2_U3398 ; P2_U6015
g6558 nand P2_U3417 P2_REG2_REG_23__SCAN_IN ; P2_U6016
g6559 nand P2_U3983 P2_U3400 ; P2_U6017
g6560 nand P2_U3417 P2_REG2_REG_24__SCAN_IN ; P2_U6018
g6561 nand P2_U3983 P2_U3402 ; P2_U6019
g6562 nand P2_U3417 P2_REG2_REG_25__SCAN_IN ; P2_U6020
g6563 nand P2_U3983 P2_U3404 ; P2_U6021
g6564 nand P2_U3417 P2_REG2_REG_26__SCAN_IN ; P2_U6022
g6565 nand P2_U3983 P2_U3406 ; P2_U6023
g6566 nand P2_U3417 P2_REG2_REG_27__SCAN_IN ; P2_U6024
g6567 nand P2_U3983 P2_U3408 ; P2_U6025
g6568 nand P2_U3417 P2_REG2_REG_28__SCAN_IN ; P2_U6026
g6569 nand P2_U3983 P2_U3410 ; P2_U6027
g6570 nand P2_U3417 P2_REG2_REG_29__SCAN_IN ; P2_U6028
g6571 nand P2_U3983 P2_U3412 ; P2_U6029
g6572 nand P2_U3417 P2_REG2_REG_30__SCAN_IN ; P2_U6030
g6573 nand P2_U3987 P2_U3983 ; P2_U6031
g6574 nand P2_U3417 P2_REG2_REG_31__SCAN_IN ; P2_U6032
g6575 nand P2_U3987 P2_U3983 ; P2_U6033
g6576 nand P2_U3423 P2_DATAO_REG_0__SCAN_IN ; P2_U6034
g6577 nand P2_U3966 P2_U3077 ; P2_U6035
g6578 nand P2_U3423 P2_DATAO_REG_1__SCAN_IN ; P2_U6036
g6579 nand P2_U3966 P2_U3078 ; P2_U6037
g6580 nand P2_U3423 P2_DATAO_REG_2__SCAN_IN ; P2_U6038
g6581 nand P2_U3966 P2_U3068 ; P2_U6039
g6582 nand P2_U3423 P2_DATAO_REG_3__SCAN_IN ; P2_U6040
g6583 nand P2_U3966 P2_U3064 ; P2_U6041
g6584 nand P2_U3423 P2_DATAO_REG_4__SCAN_IN ; P2_U6042
g6585 nand P2_U3966 P2_U3060 ; P2_U6043
g6586 nand P2_U3423 P2_DATAO_REG_5__SCAN_IN ; P2_U6044
g6587 nand P2_U3966 P2_U3067 ; P2_U6045
g6588 nand P2_U3423 P2_DATAO_REG_6__SCAN_IN ; P2_U6046
g6589 nand P2_U3966 P2_U3071 ; P2_U6047
g6590 nand P2_U3423 P2_DATAO_REG_7__SCAN_IN ; P2_U6048
g6591 nand P2_U3966 P2_U3070 ; P2_U6049
g6592 nand P2_U3423 P2_DATAO_REG_8__SCAN_IN ; P2_U6050
g6593 nand P2_U3966 P2_U3084 ; P2_U6051
g6594 nand P2_U3423 P2_DATAO_REG_9__SCAN_IN ; P2_U6052
g6595 nand P2_U3966 P2_U3083 ; P2_U6053
g6596 nand P2_U3423 P2_DATAO_REG_10__SCAN_IN ; P2_U6054
g6597 nand P2_U3966 P2_U3062 ; P2_U6055
g6598 nand P2_U3423 P2_DATAO_REG_11__SCAN_IN ; P2_U6056
g6599 nand P2_U3966 P2_U3063 ; P2_U6057
g6600 nand P2_U3423 P2_DATAO_REG_12__SCAN_IN ; P2_U6058
g6601 nand P2_U3966 P2_U3072 ; P2_U6059
g6602 nand P2_U3423 P2_DATAO_REG_13__SCAN_IN ; P2_U6060
g6603 nand P2_U3966 P2_U3080 ; P2_U6061
g6604 nand P2_U3423 P2_DATAO_REG_14__SCAN_IN ; P2_U6062
g6605 nand P2_U3966 P2_U3079 ; P2_U6063
g6606 nand P2_U3423 P2_DATAO_REG_15__SCAN_IN ; P2_U6064
g6607 nand P2_U3966 P2_U3074 ; P2_U6065
g6608 nand P2_U3423 P2_DATAO_REG_16__SCAN_IN ; P2_U6066
g6609 nand P2_U3966 P2_U3073 ; P2_U6067
g6610 nand P2_U3423 P2_DATAO_REG_17__SCAN_IN ; P2_U6068
g6611 nand P2_U3966 P2_U3069 ; P2_U6069
g6612 nand P2_U3423 P2_DATAO_REG_18__SCAN_IN ; P2_U6070
g6613 nand P2_U3966 P2_U3082 ; P2_U6071
g6614 nand P2_U3423 P2_DATAO_REG_19__SCAN_IN ; P2_U6072
g6615 nand P2_U3966 P2_U3081 ; P2_U6073
g6616 nand P2_U3423 P2_DATAO_REG_20__SCAN_IN ; P2_U6074
g6617 nand P2_U3966 P2_U3076 ; P2_U6075
g6618 nand P2_U3423 P2_DATAO_REG_21__SCAN_IN ; P2_U6076
g6619 nand P2_U3966 P2_U3075 ; P2_U6077
g6620 nand P2_U3423 P2_DATAO_REG_22__SCAN_IN ; P2_U6078
g6621 nand P2_U3966 P2_U3061 ; P2_U6079
g6622 nand P2_U3423 P2_DATAO_REG_23__SCAN_IN ; P2_U6080
g6623 nand P2_U3966 P2_U3066 ; P2_U6081
g6624 nand P2_U3423 P2_DATAO_REG_24__SCAN_IN ; P2_U6082
g6625 nand P2_U3966 P2_U3065 ; P2_U6083
g6626 nand P2_U3423 P2_DATAO_REG_25__SCAN_IN ; P2_U6084
g6627 nand P2_U3966 P2_U3058 ; P2_U6085
g6628 nand P2_U3423 P2_DATAO_REG_26__SCAN_IN ; P2_U6086
g6629 nand P2_U3966 P2_U3057 ; P2_U6087
g6630 nand P2_U3423 P2_DATAO_REG_27__SCAN_IN ; P2_U6088
g6631 nand P2_U3966 P2_U3053 ; P2_U6089
g6632 nand P2_U3423 P2_DATAO_REG_28__SCAN_IN ; P2_U6090
g6633 nand P2_U3966 P2_U3054 ; P2_U6091
g6634 nand P2_U3423 P2_DATAO_REG_29__SCAN_IN ; P2_U6092
g6635 nand P2_U3966 P2_U3055 ; P2_U6093
g6636 nand P2_U3423 P2_DATAO_REG_30__SCAN_IN ; P2_U6094
g6637 nand P2_U3966 P2_U3059 ; P2_U6095
g6638 nand P2_U3423 P2_DATAO_REG_31__SCAN_IN ; P2_U6096
g6639 nand P2_U3966 P2_U3056 ; P2_U6097
g6640 nand P2_U5708 P2_R1340_U6 ; P2_U6098
g6641 nand P2_LT_719_U11 P2_U3441 ; P2_U6099
g6642 nand P2_U5701 P2_U3425 ; P2_U6100
g6643 nand P2_U3441 P2_U3436 ; P2_U6101
g6644 nand P2_R1312_U21 P2_U5169 ; P2_U6102
g6645 nand P2_U5714 P2_U5170 P2_U3945 ; P2_U6103
g6646 nand P2_U3979 P2_U3055 ; P2_U6104
g6647 nand P2_U3411 P2_U4664 ; P2_U6105
g6648 nand P2_U6105 P2_U6104 ; P2_U6106
g6649 nand P2_U3968 P2_U3054 ; P2_U6107
g6650 nand P2_U3409 P2_U4645 ; P2_U6108
g6651 nand P2_U6108 P2_U6107 ; P2_U6109
g6652 nand P2_U3969 P2_U3053 ; P2_U6110
g6653 nand P2_U3407 P2_U4626 ; P2_U6111
g6654 nand P2_U6111 P2_U6110 ; P2_U6112
g6655 nand P2_U3972 P2_U3065 ; P2_U6113
g6656 nand P2_U3401 P2_U4569 ; P2_U6114
g6657 nand P2_U6114 P2_U6113 ; P2_U6115
g6658 nand P2_U3973 P2_U3066 ; P2_U6116
g6659 nand P2_U3399 P2_U4550 ; P2_U6117
g6660 nand P2_U6117 P2_U6116 ; P2_U6118
g6661 nand P2_U3975 P2_U3075 ; P2_U6119
g6662 nand P2_U3395 P2_U4512 ; P2_U6120
g6663 nand P2_U6120 P2_U6119 ; P2_U6121
g6664 nand P2_U3974 P2_U3061 ; P2_U6122
g6665 nand P2_U3397 P2_U4531 ; P2_U6123
g6666 nand P2_U6123 P2_U6122 ; P2_U6124
g6667 nand P2_U3971 P2_U3058 ; P2_U6125
g6668 nand P2_U3403 P2_U4588 ; P2_U6126
g6669 nand P2_U6126 P2_U6125 ; P2_U6127
g6670 nand P2_U3970 P2_U3057 ; P2_U6128
g6671 nand P2_U3405 P2_U4607 ; P2_U6129
g6672 nand P2_U6129 P2_U6128 ; P2_U6130
g6673 nand P2_U3978 P2_U3059 ; P2_U6131
g6674 nand P2_U3413 P2_U4682 ; P2_U6132
g6675 nand P2_U6132 P2_U6131 ; P2_U6133
g6676 nand P2_U3977 P2_U3056 ; P2_U6134
g6677 nand P2_U3414 P2_U4702 ; P2_U6135
g6678 nand P2_U6135 P2_U6134 ; P2_U6136
g6679 nand P2_U5867 P2_U4436 ; P2_U6137
g6680 nand P2_U3501 P2_U3069 ; P2_U6138
g6681 nand P2_U6138 P2_U6137 ; P2_U6139
g6682 nand P2_U5846 P2_U4379 ; P2_U6140
g6683 nand P2_U3492 P2_U3079 ; P2_U6141
g6684 nand P2_U6141 P2_U6140 ; P2_U6142
g6685 nand P2_U5753 P2_U4130 ; P2_U6143
g6686 nand P2_U3453 P2_U3078 ; P2_U6144
g6687 nand P2_U6144 P2_U6143 ; P2_U6145
g6688 nand P2_U5736 P2_U4151 ; P2_U6146
g6689 nand P2_U3448 P2_U3077 ; P2_U6147
g6690 nand P2_U6147 P2_U6146 ; P2_U6148
g6691 nand P2_U5853 P2_U4398 ; P2_U6149
g6692 nand P2_U3495 P2_U3074 ; P2_U6150
g6693 nand P2_U6150 P2_U6149 ; P2_U6151
g6694 nand P2_U5804 P2_U4265 ; P2_U6152
g6695 nand P2_U3474 P2_U3084 ; P2_U6153
g6696 nand P2_U6153 P2_U6152 ; P2_U6154
g6697 nand P2_U5811 P2_U4284 ; P2_U6155
g6698 nand P2_U3477 P2_U3083 ; P2_U6156
g6699 nand P2_U6156 P2_U6155 ; P2_U6157
g6700 nand P2_U5839 P2_U4360 ; P2_U6158
g6701 nand P2_U3489 P2_U3080 ; P2_U6159
g6702 nand P2_U6159 P2_U6158 ; P2_U6160
g6703 nand P2_U5860 P2_U4417 ; P2_U6161
g6704 nand P2_U3498 P2_U3073 ; P2_U6162
g6705 nand P2_U6162 P2_U6161 ; P2_U6163
g6706 nand P2_U5790 P2_U4227 ; P2_U6164
g6707 nand P2_U3468 P2_U3071 ; P2_U6165
g6708 nand P2_U6165 P2_U6164 ; P2_U6166
g6709 nand P2_U5797 P2_U4246 ; P2_U6167
g6710 nand P2_U3471 P2_U3070 ; P2_U6168
g6711 nand P2_U6168 P2_U6167 ; P2_U6169
g6712 nand P2_U5832 P2_U4341 ; P2_U6170
g6713 nand P2_U3486 P2_U3072 ; P2_U6171
g6714 nand P2_U6171 P2_U6170 ; P2_U6172
g6715 nand P2_U5783 P2_U4208 ; P2_U6173
g6716 nand P2_U3465 P2_U3067 ; P2_U6174
g6717 nand P2_U6174 P2_U6173 ; P2_U6175
g6718 nand P2_U5769 P2_U4170 ; P2_U6176
g6719 nand P2_U3459 P2_U3064 ; P2_U6177
g6720 nand P2_U6177 P2_U6176 ; P2_U6178
g6721 nand P2_U5762 P2_U4148 ; P2_U6179
g6722 nand P2_U3456 P2_U3068 ; P2_U6180
g6723 nand P2_U6180 P2_U6179 ; P2_U6181
g6724 nand P2_U5874 P2_U4455 ; P2_U6182
g6725 nand P2_U3504 P2_U3082 ; P2_U6183
g6726 nand P2_U6183 P2_U6182 ; P2_U6184
g6727 nand P2_U5879 P2_U4474 ; P2_U6185
g6728 nand P2_U3506 P2_U3081 ; P2_U6186
g6729 nand P2_U6186 P2_U6185 ; P2_U6187
g6730 nand P2_U5776 P2_U4189 ; P2_U6188
g6731 nand P2_U3462 P2_U3060 ; P2_U6189
g6732 nand P2_U6189 P2_U6188 ; P2_U6190
g6733 nand P2_U5825 P2_U4322 ; P2_U6191
g6734 nand P2_U3483 P2_U3063 ; P2_U6192
g6735 nand P2_U6192 P2_U6191 ; P2_U6193
g6736 nand P2_U5818 P2_U4303 ; P2_U6194
g6737 nand P2_U3480 P2_U3062 ; P2_U6195
g6738 nand P2_U6195 P2_U6194 ; P2_U6196
g6739 nand P2_U3976 P2_U3076 ; P2_U6197
g6740 nand P2_U3393 P2_U4493 ; P2_U6198
g6741 nand P2_U6198 P2_U6197 ; P2_U6199
g6742 nand P2_U3019 P2_U3947 ; P2_U6200
g6743 nand P2_U5168 P2_U3962 ; P2_U6201
g6744 nand P2_U3083 P2_R1299_U6 ; P2_U6202
g6745 nand P2_U3083 P2_U3948 ; P2_U6203
g6746 nand P2_U3084 P2_R1299_U6 ; P2_U6204
g6747 nand P2_U3084 P2_U3948 ; P2_U6205
g6748 nand P2_U3070 P2_R1299_U6 ; P2_U6206
g6749 nand P2_U3070 P2_U3948 ; P2_U6207
g6750 nand P2_U3071 P2_R1299_U6 ; P2_U6208
g6751 nand P2_U3071 P2_U3948 ; P2_U6209
g6752 nand P2_U3067 P2_R1299_U6 ; P2_U6210
g6753 nand P2_U3067 P2_U3948 ; P2_U6211
g6754 nand P2_U3060 P2_R1299_U6 ; P2_U6212
g6755 nand P2_U3060 P2_U3948 ; P2_U6213
g6756 nand P2_U3064 P2_R1299_U6 ; P2_U6214
g6757 nand P2_U3064 P2_U3948 ; P2_U6215
g6758 nand P2_R1335_U8 P2_R1299_U6 ; P2_U6216
g6759 nand P2_U3056 P2_U3948 ; P2_U6217
g6760 nand P2_R1335_U6 P2_R1299_U6 ; P2_U6218
g6761 nand P2_U3059 P2_U3948 ; P2_U6219
g6762 nand P2_U3068 P2_R1299_U6 ; P2_U6220
g6763 nand P2_U3068 P2_U3948 ; P2_U6221
g6764 not P2_U3593 ; P2_U6222
g6765 nand P2_U3055 P2_R1299_U6 ; P2_U6223
g6766 nand P2_U3055 P2_U3948 ; P2_U6224
g6767 nand P2_U3054 P2_R1299_U6 ; P2_U6225
g6768 nand P2_U3054 P2_U3948 ; P2_U6226
g6769 nand P2_U3053 P2_R1299_U6 ; P2_U6227
g6770 nand P2_U3053 P2_U3948 ; P2_U6228
g6771 nand P2_U3057 P2_R1299_U6 ; P2_U6229
g6772 nand P2_U3057 P2_U3948 ; P2_U6230
g6773 nand P2_U3058 P2_R1299_U6 ; P2_U6231
g6774 nand P2_U3058 P2_U3948 ; P2_U6232
g6775 nand P2_U3065 P2_R1299_U6 ; P2_U6233
g6776 nand P2_U3065 P2_U3948 ; P2_U6234
g6777 nand P2_U3066 P2_R1299_U6 ; P2_U6235
g6778 nand P2_U3066 P2_U3948 ; P2_U6236
g6779 nand P2_U3061 P2_R1299_U6 ; P2_U6237
g6780 nand P2_U3061 P2_U3948 ; P2_U6238
g6781 nand P2_U3075 P2_R1299_U6 ; P2_U6239
g6782 nand P2_U3075 P2_U3948 ; P2_U6240
g6783 nand P2_U3076 P2_R1299_U6 ; P2_U6241
g6784 nand P2_U3076 P2_U3948 ; P2_U6242
g6785 nand P2_U3078 P2_R1299_U6 ; P2_U6243
g6786 nand P2_U3078 P2_U3948 ; P2_U6244
g6787 not P2_U3604 ; P2_U6245
g6788 nand P2_U3081 P2_R1299_U6 ; P2_U6246
g6789 nand P2_U3081 P2_U3948 ; P2_U6247
g6790 nand P2_U3082 P2_R1299_U6 ; P2_U6248
g6791 nand P2_U3082 P2_U3948 ; P2_U6249
g6792 nand P2_U3069 P2_R1299_U6 ; P2_U6250
g6793 nand P2_U3069 P2_U3948 ; P2_U6251
g6794 nand P2_U3073 P2_R1299_U6 ; P2_U6252
g6795 nand P2_U3073 P2_U3948 ; P2_U6253
g6796 nand P2_U3074 P2_R1299_U6 ; P2_U6254
g6797 nand P2_U3074 P2_U3948 ; P2_U6255
g6798 nand P2_U3079 P2_R1299_U6 ; P2_U6256
g6799 nand P2_U3079 P2_U3948 ; P2_U6257
g6800 nand P2_U3080 P2_R1299_U6 ; P2_U6258
g6801 nand P2_U3080 P2_U3948 ; P2_U6259
g6802 nand P2_U3072 P2_R1299_U6 ; P2_U6260
g6803 nand P2_U3072 P2_U3948 ; P2_U6261
g6804 nand P2_U3063 P2_R1299_U6 ; P2_U6262
g6805 nand P2_U3063 P2_U3948 ; P2_U6263
g6806 nand P2_U3062 P2_R1299_U6 ; P2_U6264
g6807 nand P2_U3062 P2_U3948 ; P2_U6265
g6808 nand P2_U3077 P2_R1299_U6 ; P2_U6266
g6809 nand P2_U3077 P2_U3948 ; P2_U6267
g6810 not P2_U3615 ; P2_U6268
g6811 nand P2_U3445 P2_U5717 ; P2_U6269
g6812 nand P2_U3440 P2_U3439 ; P2_U6270
g6813 not P1_ADDR_REG_19__SCAN_IN ; LT_1079_U6
g6814 and ADD_1071_U159 ADD_1071_U155 ; ADD_1071_U4
g6815 nand ADD_1071_U221 ADD_1071_U220 ADD_1071_U160 ; ADD_1071_U5
g6816 not P1_ADDR_REG_0__SCAN_IN ; ADD_1071_U6
g6817 not P2_ADDR_REG_0__SCAN_IN ; ADD_1071_U7
g6818 not P2_ADDR_REG_1__SCAN_IN ; ADD_1071_U8
g6819 nand P1_ADDR_REG_0__SCAN_IN P2_ADDR_REG_0__SCAN_IN ; ADD_1071_U9
g6820 not P1_ADDR_REG_1__SCAN_IN ; ADD_1071_U10
g6821 not P1_ADDR_REG_2__SCAN_IN ; ADD_1071_U11
g6822 not P2_ADDR_REG_2__SCAN_IN ; ADD_1071_U12
g6823 not P1_ADDR_REG_3__SCAN_IN ; ADD_1071_U13
g6824 not P2_ADDR_REG_3__SCAN_IN ; ADD_1071_U14
g6825 not P1_ADDR_REG_4__SCAN_IN ; ADD_1071_U15
g6826 not P2_ADDR_REG_4__SCAN_IN ; ADD_1071_U16
g6827 not P1_ADDR_REG_5__SCAN_IN ; ADD_1071_U17
g6828 not P2_ADDR_REG_5__SCAN_IN ; ADD_1071_U18
g6829 not P1_ADDR_REG_6__SCAN_IN ; ADD_1071_U19
g6830 not P2_ADDR_REG_6__SCAN_IN ; ADD_1071_U20
g6831 not P1_ADDR_REG_7__SCAN_IN ; ADD_1071_U21
g6832 not P2_ADDR_REG_7__SCAN_IN ; ADD_1071_U22
g6833 not P1_ADDR_REG_8__SCAN_IN ; ADD_1071_U23
g6834 not P2_ADDR_REG_8__SCAN_IN ; ADD_1071_U24
g6835 not P2_ADDR_REG_9__SCAN_IN ; ADD_1071_U25
g6836 not P1_ADDR_REG_9__SCAN_IN ; ADD_1071_U26
g6837 not P1_ADDR_REG_10__SCAN_IN ; ADD_1071_U27
g6838 not P2_ADDR_REG_10__SCAN_IN ; ADD_1071_U28
g6839 not P1_ADDR_REG_11__SCAN_IN ; ADD_1071_U29
g6840 not P2_ADDR_REG_11__SCAN_IN ; ADD_1071_U30
g6841 not P1_ADDR_REG_12__SCAN_IN ; ADD_1071_U31
g6842 not P2_ADDR_REG_12__SCAN_IN ; ADD_1071_U32
g6843 not P1_ADDR_REG_13__SCAN_IN ; ADD_1071_U33
g6844 not P2_ADDR_REG_13__SCAN_IN ; ADD_1071_U34
g6845 not P1_ADDR_REG_14__SCAN_IN ; ADD_1071_U35
g6846 not P2_ADDR_REG_14__SCAN_IN ; ADD_1071_U36
g6847 not P1_ADDR_REG_15__SCAN_IN ; ADD_1071_U37
g6848 not P2_ADDR_REG_15__SCAN_IN ; ADD_1071_U38
g6849 not P1_ADDR_REG_16__SCAN_IN ; ADD_1071_U39
g6850 not P2_ADDR_REG_16__SCAN_IN ; ADD_1071_U40
g6851 not P1_ADDR_REG_17__SCAN_IN ; ADD_1071_U41
g6852 not P2_ADDR_REG_17__SCAN_IN ; ADD_1071_U42
g6853 not P1_ADDR_REG_18__SCAN_IN ; ADD_1071_U43
g6854 not P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U44
g6855 nand ADD_1071_U150 ADD_1071_U149 ; ADD_1071_U45
g6856 nand ADD_1071_U291 ADD_1071_U290 ; ADD_1071_U46
g6857 nand ADD_1071_U167 ADD_1071_U166 ; ADD_1071_U47
g6858 nand ADD_1071_U174 ADD_1071_U173 ; ADD_1071_U48
g6859 nand ADD_1071_U181 ADD_1071_U180 ; ADD_1071_U49
g6860 nand ADD_1071_U188 ADD_1071_U187 ; ADD_1071_U50
g6861 nand ADD_1071_U195 ADD_1071_U194 ; ADD_1071_U51
g6862 nand ADD_1071_U202 ADD_1071_U201 ; ADD_1071_U52
g6863 nand ADD_1071_U209 ADD_1071_U208 ; ADD_1071_U53
g6864 nand ADD_1071_U216 ADD_1071_U215 ; ADD_1071_U54
g6865 nand ADD_1071_U233 ADD_1071_U232 ; ADD_1071_U55
g6866 nand ADD_1071_U240 ADD_1071_U239 ; ADD_1071_U56
g6867 nand ADD_1071_U247 ADD_1071_U246 ; ADD_1071_U57
g6868 nand ADD_1071_U254 ADD_1071_U253 ; ADD_1071_U58
g6869 nand ADD_1071_U261 ADD_1071_U260 ; ADD_1071_U59
g6870 nand ADD_1071_U268 ADD_1071_U267 ; ADD_1071_U60
g6871 nand ADD_1071_U275 ADD_1071_U274 ; ADD_1071_U61
g6872 nand ADD_1071_U282 ADD_1071_U281 ; ADD_1071_U62
g6873 nand ADD_1071_U289 ADD_1071_U288 ; ADD_1071_U63
g6874 nand ADD_1071_U114 ADD_1071_U113 ; ADD_1071_U64
g6875 nand ADD_1071_U110 ADD_1071_U109 ; ADD_1071_U65
g6876 nand ADD_1071_U106 ADD_1071_U105 ; ADD_1071_U66
g6877 nand ADD_1071_U102 ADD_1071_U101 ; ADD_1071_U67
g6878 nand ADD_1071_U98 ADD_1071_U97 ; ADD_1071_U68
g6879 nand ADD_1071_U94 ADD_1071_U93 ; ADD_1071_U69
g6880 nand ADD_1071_U90 ADD_1071_U89 ; ADD_1071_U70
g6881 nand ADD_1071_U72 ADD_1071_U86 ; ADD_1071_U71
g6882 nand ADD_1071_U84 P1_ADDR_REG_1__SCAN_IN ; ADD_1071_U72
g6883 not P2_ADDR_REG_19__SCAN_IN ; ADD_1071_U73
g6884 not P1_ADDR_REG_19__SCAN_IN ; ADD_1071_U74
g6885 nand ADD_1071_U146 ADD_1071_U145 ; ADD_1071_U75
g6886 nand ADD_1071_U142 ADD_1071_U141 ; ADD_1071_U76
g6887 nand ADD_1071_U138 ADD_1071_U137 ; ADD_1071_U77
g6888 nand ADD_1071_U134 ADD_1071_U133 ; ADD_1071_U78
g6889 nand ADD_1071_U130 ADD_1071_U129 ; ADD_1071_U79
g6890 nand ADD_1071_U126 ADD_1071_U125 ; ADD_1071_U80
g6891 nand ADD_1071_U122 ADD_1071_U121 ; ADD_1071_U81
g6892 nand ADD_1071_U118 ADD_1071_U117 ; ADD_1071_U82
g6893 not ADD_1071_U72 ; ADD_1071_U83
g6894 not ADD_1071_U9 ; ADD_1071_U84
g6895 nand ADD_1071_U10 ADD_1071_U9 ; ADD_1071_U85
g6896 nand ADD_1071_U85 P2_ADDR_REG_1__SCAN_IN ; ADD_1071_U86
g6897 not ADD_1071_U71 ; ADD_1071_U87
g6898 or P1_ADDR_REG_2__SCAN_IN P2_ADDR_REG_2__SCAN_IN ; ADD_1071_U88
g6899 nand ADD_1071_U88 ADD_1071_U71 ; ADD_1071_U89
g6900 nand P1_ADDR_REG_2__SCAN_IN P2_ADDR_REG_2__SCAN_IN ; ADD_1071_U90
g6901 not ADD_1071_U70 ; ADD_1071_U91
g6902 or P1_ADDR_REG_3__SCAN_IN P2_ADDR_REG_3__SCAN_IN ; ADD_1071_U92
g6903 nand ADD_1071_U92 ADD_1071_U70 ; ADD_1071_U93
g6904 nand P1_ADDR_REG_3__SCAN_IN P2_ADDR_REG_3__SCAN_IN ; ADD_1071_U94
g6905 not ADD_1071_U69 ; ADD_1071_U95
g6906 or P1_ADDR_REG_4__SCAN_IN P2_ADDR_REG_4__SCAN_IN ; ADD_1071_U96
g6907 nand ADD_1071_U96 ADD_1071_U69 ; ADD_1071_U97
g6908 nand P1_ADDR_REG_4__SCAN_IN P2_ADDR_REG_4__SCAN_IN ; ADD_1071_U98
g6909 not ADD_1071_U68 ; ADD_1071_U99
g6910 or P1_ADDR_REG_5__SCAN_IN P2_ADDR_REG_5__SCAN_IN ; ADD_1071_U100
g6911 nand ADD_1071_U100 ADD_1071_U68 ; ADD_1071_U101
g6912 nand P1_ADDR_REG_5__SCAN_IN P2_ADDR_REG_5__SCAN_IN ; ADD_1071_U102
g6913 not ADD_1071_U67 ; ADD_1071_U103
g6914 or P1_ADDR_REG_6__SCAN_IN P2_ADDR_REG_6__SCAN_IN ; ADD_1071_U104
g6915 nand ADD_1071_U104 ADD_1071_U67 ; ADD_1071_U105
g6916 nand P1_ADDR_REG_6__SCAN_IN P2_ADDR_REG_6__SCAN_IN ; ADD_1071_U106
g6917 not ADD_1071_U66 ; ADD_1071_U107
g6918 or P1_ADDR_REG_7__SCAN_IN P2_ADDR_REG_7__SCAN_IN ; ADD_1071_U108
g6919 nand ADD_1071_U108 ADD_1071_U66 ; ADD_1071_U109
g6920 nand P1_ADDR_REG_7__SCAN_IN P2_ADDR_REG_7__SCAN_IN ; ADD_1071_U110
g6921 not ADD_1071_U65 ; ADD_1071_U111
g6922 or P1_ADDR_REG_8__SCAN_IN P2_ADDR_REG_8__SCAN_IN ; ADD_1071_U112
g6923 nand ADD_1071_U112 ADD_1071_U65 ; ADD_1071_U113
g6924 nand P1_ADDR_REG_8__SCAN_IN P2_ADDR_REG_8__SCAN_IN ; ADD_1071_U114
g6925 not ADD_1071_U64 ; ADD_1071_U115
g6926 or P1_ADDR_REG_9__SCAN_IN P2_ADDR_REG_9__SCAN_IN ; ADD_1071_U116
g6927 nand ADD_1071_U116 ADD_1071_U64 ; ADD_1071_U117
g6928 nand P1_ADDR_REG_9__SCAN_IN P2_ADDR_REG_9__SCAN_IN ; ADD_1071_U118
g6929 not ADD_1071_U82 ; ADD_1071_U119
g6930 or P1_ADDR_REG_10__SCAN_IN P2_ADDR_REG_10__SCAN_IN ; ADD_1071_U120
g6931 nand ADD_1071_U120 ADD_1071_U82 ; ADD_1071_U121
g6932 nand P1_ADDR_REG_10__SCAN_IN P2_ADDR_REG_10__SCAN_IN ; ADD_1071_U122
g6933 not ADD_1071_U81 ; ADD_1071_U123
g6934 or P1_ADDR_REG_11__SCAN_IN P2_ADDR_REG_11__SCAN_IN ; ADD_1071_U124
g6935 nand ADD_1071_U124 ADD_1071_U81 ; ADD_1071_U125
g6936 nand P1_ADDR_REG_11__SCAN_IN P2_ADDR_REG_11__SCAN_IN ; ADD_1071_U126
g6937 not ADD_1071_U80 ; ADD_1071_U127
g6938 or P1_ADDR_REG_12__SCAN_IN P2_ADDR_REG_12__SCAN_IN ; ADD_1071_U128
g6939 nand ADD_1071_U128 ADD_1071_U80 ; ADD_1071_U129
g6940 nand P1_ADDR_REG_12__SCAN_IN P2_ADDR_REG_12__SCAN_IN ; ADD_1071_U130
g6941 not ADD_1071_U79 ; ADD_1071_U131
g6942 or P1_ADDR_REG_13__SCAN_IN P2_ADDR_REG_13__SCAN_IN ; ADD_1071_U132
g6943 nand ADD_1071_U132 ADD_1071_U79 ; ADD_1071_U133
g6944 nand P1_ADDR_REG_13__SCAN_IN P2_ADDR_REG_13__SCAN_IN ; ADD_1071_U134
g6945 not ADD_1071_U78 ; ADD_1071_U135
g6946 or P1_ADDR_REG_14__SCAN_IN P2_ADDR_REG_14__SCAN_IN ; ADD_1071_U136
g6947 nand ADD_1071_U136 ADD_1071_U78 ; ADD_1071_U137
g6948 nand P1_ADDR_REG_14__SCAN_IN P2_ADDR_REG_14__SCAN_IN ; ADD_1071_U138
g6949 not ADD_1071_U77 ; ADD_1071_U139
g6950 or P1_ADDR_REG_15__SCAN_IN P2_ADDR_REG_15__SCAN_IN ; ADD_1071_U140
g6951 nand ADD_1071_U140 ADD_1071_U77 ; ADD_1071_U141
g6952 nand P1_ADDR_REG_15__SCAN_IN P2_ADDR_REG_15__SCAN_IN ; ADD_1071_U142
g6953 not ADD_1071_U76 ; ADD_1071_U143
g6954 or P1_ADDR_REG_16__SCAN_IN P2_ADDR_REG_16__SCAN_IN ; ADD_1071_U144
g6955 nand ADD_1071_U144 ADD_1071_U76 ; ADD_1071_U145
g6956 nand P1_ADDR_REG_16__SCAN_IN P2_ADDR_REG_16__SCAN_IN ; ADD_1071_U146
g6957 not ADD_1071_U75 ; ADD_1071_U147
g6958 or P1_ADDR_REG_17__SCAN_IN P2_ADDR_REG_17__SCAN_IN ; ADD_1071_U148
g6959 nand ADD_1071_U148 ADD_1071_U75 ; ADD_1071_U149
g6960 nand P1_ADDR_REG_17__SCAN_IN P2_ADDR_REG_17__SCAN_IN ; ADD_1071_U150
g6961 not ADD_1071_U45 ; ADD_1071_U151
g6962 or P1_ADDR_REG_18__SCAN_IN P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U152
g6963 nand ADD_1071_U152 ADD_1071_U45 ; ADD_1071_U153
g6964 nand P1_ADDR_REG_18__SCAN_IN P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U154
g6965 nand ADD_1071_U223 ADD_1071_U222 ADD_1071_U154 ADD_1071_U153 ; ADD_1071_U155
g6966 nand P1_ADDR_REG_18__SCAN_IN P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U156
g6967 nand ADD_1071_U151 ADD_1071_U156 ; ADD_1071_U157
g6968 or P1_ADDR_REG_18__SCAN_IN P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U158
g6969 nand ADD_1071_U158 ADD_1071_U226 ADD_1071_U157 ; ADD_1071_U159
g6970 nand ADD_1071_U219 ADD_1071_U10 ; ADD_1071_U160
g6971 nand ADD_1071_U26 P2_ADDR_REG_9__SCAN_IN ; ADD_1071_U161
g6972 nand ADD_1071_U25 P1_ADDR_REG_9__SCAN_IN ; ADD_1071_U162
g6973 nand ADD_1071_U26 P2_ADDR_REG_9__SCAN_IN ; ADD_1071_U163
g6974 nand ADD_1071_U25 P1_ADDR_REG_9__SCAN_IN ; ADD_1071_U164
g6975 nand ADD_1071_U164 ADD_1071_U163 ; ADD_1071_U165
g6976 nand ADD_1071_U162 ADD_1071_U161 ADD_1071_U64 ; ADD_1071_U166
g6977 nand ADD_1071_U115 ADD_1071_U165 ; ADD_1071_U167
g6978 nand ADD_1071_U23 P2_ADDR_REG_8__SCAN_IN ; ADD_1071_U168
g6979 nand ADD_1071_U24 P1_ADDR_REG_8__SCAN_IN ; ADD_1071_U169
g6980 nand ADD_1071_U23 P2_ADDR_REG_8__SCAN_IN ; ADD_1071_U170
g6981 nand ADD_1071_U24 P1_ADDR_REG_8__SCAN_IN ; ADD_1071_U171
g6982 nand ADD_1071_U171 ADD_1071_U170 ; ADD_1071_U172
g6983 nand ADD_1071_U169 ADD_1071_U168 ADD_1071_U65 ; ADD_1071_U173
g6984 nand ADD_1071_U111 ADD_1071_U172 ; ADD_1071_U174
g6985 nand ADD_1071_U21 P2_ADDR_REG_7__SCAN_IN ; ADD_1071_U175
g6986 nand ADD_1071_U22 P1_ADDR_REG_7__SCAN_IN ; ADD_1071_U176
g6987 nand ADD_1071_U21 P2_ADDR_REG_7__SCAN_IN ; ADD_1071_U177
g6988 nand ADD_1071_U22 P1_ADDR_REG_7__SCAN_IN ; ADD_1071_U178
g6989 nand ADD_1071_U178 ADD_1071_U177 ; ADD_1071_U179
g6990 nand ADD_1071_U176 ADD_1071_U175 ADD_1071_U66 ; ADD_1071_U180
g6991 nand ADD_1071_U107 ADD_1071_U179 ; ADD_1071_U181
g6992 nand ADD_1071_U19 P2_ADDR_REG_6__SCAN_IN ; ADD_1071_U182
g6993 nand ADD_1071_U20 P1_ADDR_REG_6__SCAN_IN ; ADD_1071_U183
g6994 nand ADD_1071_U19 P2_ADDR_REG_6__SCAN_IN ; ADD_1071_U184
g6995 nand ADD_1071_U20 P1_ADDR_REG_6__SCAN_IN ; ADD_1071_U185
g6996 nand ADD_1071_U185 ADD_1071_U184 ; ADD_1071_U186
g6997 nand ADD_1071_U183 ADD_1071_U182 ADD_1071_U67 ; ADD_1071_U187
g6998 nand ADD_1071_U103 ADD_1071_U186 ; ADD_1071_U188
g6999 nand ADD_1071_U17 P2_ADDR_REG_5__SCAN_IN ; ADD_1071_U189
g7000 nand ADD_1071_U18 P1_ADDR_REG_5__SCAN_IN ; ADD_1071_U190
g7001 nand ADD_1071_U17 P2_ADDR_REG_5__SCAN_IN ; ADD_1071_U191
g7002 nand ADD_1071_U18 P1_ADDR_REG_5__SCAN_IN ; ADD_1071_U192
g7003 nand ADD_1071_U192 ADD_1071_U191 ; ADD_1071_U193
g7004 nand ADD_1071_U190 ADD_1071_U189 ADD_1071_U68 ; ADD_1071_U194
g7005 nand ADD_1071_U99 ADD_1071_U193 ; ADD_1071_U195
g7006 nand ADD_1071_U15 P2_ADDR_REG_4__SCAN_IN ; ADD_1071_U196
g7007 nand ADD_1071_U16 P1_ADDR_REG_4__SCAN_IN ; ADD_1071_U197
g7008 nand ADD_1071_U15 P2_ADDR_REG_4__SCAN_IN ; ADD_1071_U198
g7009 nand ADD_1071_U16 P1_ADDR_REG_4__SCAN_IN ; ADD_1071_U199
g7010 nand ADD_1071_U199 ADD_1071_U198 ; ADD_1071_U200
g7011 nand ADD_1071_U197 ADD_1071_U196 ADD_1071_U69 ; ADD_1071_U201
g7012 nand ADD_1071_U95 ADD_1071_U200 ; ADD_1071_U202
g7013 nand ADD_1071_U13 P2_ADDR_REG_3__SCAN_IN ; ADD_1071_U203
g7014 nand ADD_1071_U14 P1_ADDR_REG_3__SCAN_IN ; ADD_1071_U204
g7015 nand ADD_1071_U13 P2_ADDR_REG_3__SCAN_IN ; ADD_1071_U205
g7016 nand ADD_1071_U14 P1_ADDR_REG_3__SCAN_IN ; ADD_1071_U206
g7017 nand ADD_1071_U206 ADD_1071_U205 ; ADD_1071_U207
g7018 nand ADD_1071_U204 ADD_1071_U203 ADD_1071_U70 ; ADD_1071_U208
g7019 nand ADD_1071_U91 ADD_1071_U207 ; ADD_1071_U209
g7020 nand ADD_1071_U11 P2_ADDR_REG_2__SCAN_IN ; ADD_1071_U210
g7021 nand ADD_1071_U12 P1_ADDR_REG_2__SCAN_IN ; ADD_1071_U211
g7022 nand ADD_1071_U11 P2_ADDR_REG_2__SCAN_IN ; ADD_1071_U212
g7023 nand ADD_1071_U12 P1_ADDR_REG_2__SCAN_IN ; ADD_1071_U213
g7024 nand ADD_1071_U213 ADD_1071_U212 ; ADD_1071_U214
g7025 nand ADD_1071_U211 ADD_1071_U210 ADD_1071_U71 ; ADD_1071_U215
g7026 nand ADD_1071_U87 ADD_1071_U214 ; ADD_1071_U216
g7027 nand ADD_1071_U9 P2_ADDR_REG_1__SCAN_IN ; ADD_1071_U217
g7028 nand ADD_1071_U84 ADD_1071_U8 ; ADD_1071_U218
g7029 nand ADD_1071_U218 ADD_1071_U217 ; ADD_1071_U219
g7030 nand ADD_1071_U9 ADD_1071_U8 P1_ADDR_REG_1__SCAN_IN ; ADD_1071_U220
g7031 nand ADD_1071_U83 P2_ADDR_REG_1__SCAN_IN ; ADD_1071_U221
g7032 nand ADD_1071_U74 P2_ADDR_REG_19__SCAN_IN ; ADD_1071_U222
g7033 nand ADD_1071_U73 P1_ADDR_REG_19__SCAN_IN ; ADD_1071_U223
g7034 nand ADD_1071_U74 P2_ADDR_REG_19__SCAN_IN ; ADD_1071_U224
g7035 nand ADD_1071_U73 P1_ADDR_REG_19__SCAN_IN ; ADD_1071_U225
g7036 nand ADD_1071_U225 ADD_1071_U224 ; ADD_1071_U226
g7037 nand ADD_1071_U43 P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U227
g7038 nand ADD_1071_U44 P1_ADDR_REG_18__SCAN_IN ; ADD_1071_U228
g7039 nand ADD_1071_U43 P2_ADDR_REG_18__SCAN_IN ; ADD_1071_U229
g7040 nand ADD_1071_U44 P1_ADDR_REG_18__SCAN_IN ; ADD_1071_U230
g7041 nand ADD_1071_U230 ADD_1071_U229 ; ADD_1071_U231
g7042 nand ADD_1071_U228 ADD_1071_U227 ADD_1071_U45 ; ADD_1071_U232
g7043 nand ADD_1071_U231 ADD_1071_U151 ; ADD_1071_U233
g7044 nand ADD_1071_U41 P2_ADDR_REG_17__SCAN_IN ; ADD_1071_U234
g7045 nand ADD_1071_U42 P1_ADDR_REG_17__SCAN_IN ; ADD_1071_U235
g7046 nand ADD_1071_U41 P2_ADDR_REG_17__SCAN_IN ; ADD_1071_U236
g7047 nand ADD_1071_U42 P1_ADDR_REG_17__SCAN_IN ; ADD_1071_U237
g7048 nand ADD_1071_U237 ADD_1071_U236 ; ADD_1071_U238
g7049 nand ADD_1071_U235 ADD_1071_U234 ADD_1071_U75 ; ADD_1071_U239
g7050 nand ADD_1071_U147 ADD_1071_U238 ; ADD_1071_U240
g7051 nand ADD_1071_U39 P2_ADDR_REG_16__SCAN_IN ; ADD_1071_U241
g7052 nand ADD_1071_U40 P1_ADDR_REG_16__SCAN_IN ; ADD_1071_U242
g7053 nand ADD_1071_U39 P2_ADDR_REG_16__SCAN_IN ; ADD_1071_U243
g7054 nand ADD_1071_U40 P1_ADDR_REG_16__SCAN_IN ; ADD_1071_U244
g7055 nand ADD_1071_U244 ADD_1071_U243 ; ADD_1071_U245
g7056 nand ADD_1071_U242 ADD_1071_U241 ADD_1071_U76 ; ADD_1071_U246
g7057 nand ADD_1071_U143 ADD_1071_U245 ; ADD_1071_U247
g7058 nand ADD_1071_U37 P2_ADDR_REG_15__SCAN_IN ; ADD_1071_U248
g7059 nand ADD_1071_U38 P1_ADDR_REG_15__SCAN_IN ; ADD_1071_U249
g7060 nand ADD_1071_U37 P2_ADDR_REG_15__SCAN_IN ; ADD_1071_U250
g7061 nand ADD_1071_U38 P1_ADDR_REG_15__SCAN_IN ; ADD_1071_U251
g7062 nand ADD_1071_U251 ADD_1071_U250 ; ADD_1071_U252
g7063 nand ADD_1071_U249 ADD_1071_U248 ADD_1071_U77 ; ADD_1071_U253
g7064 nand ADD_1071_U139 ADD_1071_U252 ; ADD_1071_U254
g7065 nand ADD_1071_U35 P2_ADDR_REG_14__SCAN_IN ; ADD_1071_U255
g7066 nand ADD_1071_U36 P1_ADDR_REG_14__SCAN_IN ; ADD_1071_U256
g7067 nand ADD_1071_U35 P2_ADDR_REG_14__SCAN_IN ; ADD_1071_U257
g7068 nand ADD_1071_U36 P1_ADDR_REG_14__SCAN_IN ; ADD_1071_U258
g7069 nand ADD_1071_U258 ADD_1071_U257 ; ADD_1071_U259
g7070 nand ADD_1071_U256 ADD_1071_U255 ADD_1071_U78 ; ADD_1071_U260
g7071 nand ADD_1071_U135 ADD_1071_U259 ; ADD_1071_U261
g7072 nand ADD_1071_U33 P2_ADDR_REG_13__SCAN_IN ; ADD_1071_U262
g7073 nand ADD_1071_U34 P1_ADDR_REG_13__SCAN_IN ; ADD_1071_U263
g7074 nand ADD_1071_U33 P2_ADDR_REG_13__SCAN_IN ; ADD_1071_U264
g7075 nand ADD_1071_U34 P1_ADDR_REG_13__SCAN_IN ; ADD_1071_U265
g7076 nand ADD_1071_U265 ADD_1071_U264 ; ADD_1071_U266
g7077 nand ADD_1071_U263 ADD_1071_U262 ADD_1071_U79 ; ADD_1071_U267
g7078 nand ADD_1071_U131 ADD_1071_U266 ; ADD_1071_U268
g7079 nand ADD_1071_U31 P2_ADDR_REG_12__SCAN_IN ; ADD_1071_U269
g7080 nand ADD_1071_U32 P1_ADDR_REG_12__SCAN_IN ; ADD_1071_U270
g7081 nand ADD_1071_U31 P2_ADDR_REG_12__SCAN_IN ; ADD_1071_U271
g7082 nand ADD_1071_U32 P1_ADDR_REG_12__SCAN_IN ; ADD_1071_U272
g7083 nand ADD_1071_U272 ADD_1071_U271 ; ADD_1071_U273
g7084 nand ADD_1071_U270 ADD_1071_U269 ADD_1071_U80 ; ADD_1071_U274
g7085 nand ADD_1071_U127 ADD_1071_U273 ; ADD_1071_U275
g7086 nand ADD_1071_U29 P2_ADDR_REG_11__SCAN_IN ; ADD_1071_U276
g7087 nand ADD_1071_U30 P1_ADDR_REG_11__SCAN_IN ; ADD_1071_U277
g7088 nand ADD_1071_U29 P2_ADDR_REG_11__SCAN_IN ; ADD_1071_U278
g7089 nand ADD_1071_U30 P1_ADDR_REG_11__SCAN_IN ; ADD_1071_U279
g7090 nand ADD_1071_U279 ADD_1071_U278 ; ADD_1071_U280
g7091 nand ADD_1071_U277 ADD_1071_U276 ADD_1071_U81 ; ADD_1071_U281
g7092 nand ADD_1071_U123 ADD_1071_U280 ; ADD_1071_U282
g7093 nand ADD_1071_U27 P2_ADDR_REG_10__SCAN_IN ; ADD_1071_U283
g7094 nand ADD_1071_U28 P1_ADDR_REG_10__SCAN_IN ; ADD_1071_U284
g7095 nand ADD_1071_U27 P2_ADDR_REG_10__SCAN_IN ; ADD_1071_U285
g7096 nand ADD_1071_U28 P1_ADDR_REG_10__SCAN_IN ; ADD_1071_U286
g7097 nand ADD_1071_U286 ADD_1071_U285 ; ADD_1071_U287
g7098 nand ADD_1071_U284 ADD_1071_U283 ADD_1071_U82 ; ADD_1071_U288
g7099 nand ADD_1071_U119 ADD_1071_U287 ; ADD_1071_U289
g7100 nand ADD_1071_U6 P2_ADDR_REG_0__SCAN_IN ; ADD_1071_U290
g7101 nand ADD_1071_U7 P1_ADDR_REG_0__SCAN_IN ; ADD_1071_U291
g7102 and R140_U197 R140_U195 ; R140_U4
g7103 and R140_U203 R140_U201 ; R140_U5
g7104 and R140_U5 R140_U205 ; R140_U6
g7105 and R140_U213 R140_U209 ; R140_U7
g7106 and R140_U7 R140_U216 ; R140_U8
g7107 and R140_U378 R140_U377 ; R140_U9
g7108 nand R140_U469 R140_U468 R140_U324 ; R140_U10
g7109 and R140_U124 R140_U323 ; R140_U11
g7110 not SI_8_ ; R140_U12
g7111 not U90 ; R140_U13
g7112 not SI_7_ ; R140_U14
g7113 not U91 ; R140_U15
g7114 nand U91 SI_7_ ; R140_U16
g7115 not SI_6_ ; R140_U17
g7116 not U92 ; R140_U18
g7117 not SI_5_ ; R140_U19
g7118 not U93 ; R140_U20
g7119 not SI_4_ ; R140_U21
g7120 not U94 ; R140_U22
g7121 nand U94 SI_4_ ; R140_U23
g7122 not SI_3_ ; R140_U24
g7123 not U97 ; R140_U25
g7124 not SI_2_ ; R140_U26
g7125 not U108 ; R140_U27
g7126 nand U108 SI_2_ ; R140_U28
g7127 not SI_1_ ; R140_U29
g7128 not SI_0_ ; R140_U30
g7129 not U120 ; R140_U31
g7130 not U119 ; R140_U32
g7131 not U89 ; R140_U33
g7132 not SI_9_ ; R140_U34
g7133 nand R140_U288 R140_U198 ; R140_U35
g7134 not SI_14_ ; R140_U36
g7135 not U114 ; R140_U37
g7136 not SI_10_ ; R140_U38
g7137 not U118 ; R140_U39
g7138 not SI_13_ ; R140_U40
g7139 not U115 ; R140_U41
g7140 not SI_12_ ; R140_U42
g7141 not U116 ; R140_U43
g7142 not SI_11_ ; R140_U44
g7143 not U117 ; R140_U45
g7144 nand U117 SI_11_ ; R140_U46
g7145 not SI_15_ ; R140_U47
g7146 not U113 ; R140_U48
g7147 not SI_16_ ; R140_U49
g7148 not U112 ; R140_U50
g7149 not SI_17_ ; R140_U51
g7150 not U111 ; R140_U52
g7151 not SI_18_ ; R140_U53
g7152 not U110 ; R140_U54
g7153 not SI_19_ ; R140_U55
g7154 not U109 ; R140_U56
g7155 not SI_20_ ; R140_U57
g7156 not U107 ; R140_U58
g7157 not SI_21_ ; R140_U59
g7158 not U106 ; R140_U60
g7159 not SI_22_ ; R140_U61
g7160 not U105 ; R140_U62
g7161 not SI_23_ ; R140_U63
g7162 not U104 ; R140_U64
g7163 not SI_24_ ; R140_U65
g7164 not U103 ; R140_U66
g7165 not SI_25_ ; R140_U67
g7166 not U102 ; R140_U68
g7167 not SI_26_ ; R140_U69
g7168 not U101 ; R140_U70
g7169 not SI_27_ ; R140_U71
g7170 not U100 ; R140_U72
g7171 not SI_28_ ; R140_U73
g7172 not U99 ; R140_U74
g7173 not SI_29_ ; R140_U75
g7174 not U98 ; R140_U76
g7175 not SI_30_ ; R140_U77
g7176 not U96 ; R140_U78
g7177 nand SI_0_ SI_1_ U120 ; R140_U79
g7178 nand R140_U300 R140_U217 ; R140_U80
g7179 nand R140_U297 R140_U214 ; R140_U81
g7180 nand R140_U293 R140_U206 ; R140_U82
g7181 nand R140_U541 R140_U540 ; R140_U83
g7182 nand R140_U331 R140_U330 ; R140_U84
g7183 nand R140_U338 R140_U337 ; R140_U85
g7184 nand R140_U345 R140_U344 ; R140_U86
g7185 nand R140_U352 R140_U351 ; R140_U87
g7186 nand R140_U359 R140_U358 ; R140_U88
g7187 nand R140_U366 R140_U365 ; R140_U89
g7188 nand R140_U373 R140_U372 ; R140_U90
g7189 nand R140_U387 R140_U386 ; R140_U91
g7190 nand R140_U394 R140_U393 ; R140_U92
g7191 nand R140_U401 R140_U400 ; R140_U93
g7192 nand R140_U408 R140_U407 ; R140_U94
g7193 nand R140_U415 R140_U414 ; R140_U95
g7194 nand R140_U422 R140_U421 ; R140_U96
g7195 nand R140_U429 R140_U428 ; R140_U97
g7196 nand R140_U436 R140_U435 ; R140_U98
g7197 nand R140_U443 R140_U442 ; R140_U99
g7198 nand R140_U450 R140_U449 ; R140_U100
g7199 nand R140_U457 R140_U456 ; R140_U101
g7200 nand R140_U464 R140_U463 ; R140_U102
g7201 nand R140_U476 R140_U475 ; R140_U103
g7202 nand R140_U483 R140_U482 ; R140_U104
g7203 nand R140_U490 R140_U489 ; R140_U105
g7204 nand R140_U497 R140_U496 ; R140_U106
g7205 nand R140_U504 R140_U503 ; R140_U107
g7206 nand R140_U511 R140_U510 ; R140_U108
g7207 nand R140_U518 R140_U517 ; R140_U109
g7208 nand R140_U525 R140_U524 ; R140_U110
g7209 nand R140_U532 R140_U531 ; R140_U111
g7210 nand R140_U539 R140_U538 ; R140_U112
g7211 and R140_U189 R140_U193 ; R140_U113
g7212 and R140_U287 R140_U194 ; R140_U114
g7213 and R140_U4 R140_U199 ; R140_U115
g7214 and R140_U290 R140_U200 ; R140_U116
g7215 and R140_U291 R140_U204 ; R140_U117
g7216 and R140_U6 R140_U207 ; R140_U118
g7217 and R140_U295 R140_U208 ; R140_U119
g7218 and R140_U8 R140_U219 ; R140_U120
g7219 and R140_U303 R140_U220 ; R140_U121
g7220 and R140_U9 R140_U282 R140_U280 ; R140_U122
g7221 and R140_U283 R140_U376 ; R140_U123
g7222 and R140_U141 R140_U284 ; R140_U124
g7223 and R140_U326 R140_U325 ; R140_U125
g7224 nand R140_U117 R140_U309 ; R140_U126
g7225 and R140_U333 R140_U332 ; R140_U127
g7226 nand R140_U307 R140_U16 ; R140_U128
g7227 and R140_U340 R140_U339 ; R140_U129
g7228 nand R140_U116 R140_U319 ; R140_U130
g7229 and R140_U347 R140_U346 ; R140_U131
g7230 nand R140_U289 R140_U317 ; R140_U132
g7231 and R140_U354 R140_U353 ; R140_U133
g7232 nand R140_U315 R140_U23 ; R140_U134
g7233 and R140_U361 R140_U360 ; R140_U135
g7234 nand R140_U114 R140_U321 ; R140_U136
g7235 and R140_U368 R140_U367 ; R140_U137
g7236 nand R140_U28 R140_U190 ; R140_U138
g7237 not U95 ; R140_U139
g7238 not SI_31_ ; R140_U140
g7239 and R140_U380 R140_U379 ; R140_U141
g7240 and R140_U382 R140_U381 ; R140_U142
g7241 nand R140_U280 R140_U279 ; R140_U143
g7242 nand R140_U286 R140_U79 R140_U285 ; R140_U144
g7243 and R140_U396 R140_U395 ; R140_U145
g7244 nand R140_U276 R140_U275 ; R140_U146
g7245 and R140_U403 R140_U402 ; R140_U147
g7246 nand R140_U272 R140_U271 ; R140_U148
g7247 and R140_U410 R140_U409 ; R140_U149
g7248 nand R140_U268 R140_U267 ; R140_U150
g7249 and R140_U417 R140_U416 ; R140_U151
g7250 nand R140_U264 R140_U263 ; R140_U152
g7251 and R140_U424 R140_U423 ; R140_U153
g7252 nand R140_U260 R140_U259 ; R140_U154
g7253 and R140_U431 R140_U430 ; R140_U155
g7254 nand R140_U256 R140_U255 ; R140_U156
g7255 and R140_U438 R140_U437 ; R140_U157
g7256 nand R140_U252 R140_U251 ; R140_U158
g7257 and R140_U445 R140_U444 ; R140_U159
g7258 nand R140_U248 R140_U247 ; R140_U160
g7259 and R140_U452 R140_U451 ; R140_U161
g7260 nand R140_U244 R140_U243 ; R140_U162
g7261 and R140_U459 R140_U458 ; R140_U163
g7262 nand R140_U240 R140_U239 ; R140_U164
g7263 nand U120 SI_0_ ; R140_U165
g7264 and R140_U471 R140_U470 ; R140_U166
g7265 nand R140_U236 R140_U235 ; R140_U167
g7266 and R140_U478 R140_U477 ; R140_U168
g7267 nand R140_U232 R140_U231 ; R140_U169
g7268 and R140_U485 R140_U484 ; R140_U170
g7269 nand R140_U228 R140_U227 ; R140_U171
g7270 and R140_U492 R140_U491 ; R140_U172
g7271 nand R140_U224 R140_U223 ; R140_U173
g7272 and R140_U499 R140_U498 ; R140_U174
g7273 nand R140_U121 R140_U302 ; R140_U175
g7274 and R140_U506 R140_U505 ; R140_U176
g7275 nand R140_U301 R140_U299 ; R140_U177
g7276 and R140_U513 R140_U512 ; R140_U178
g7277 nand R140_U298 R140_U296 ; R140_U179
g7278 and R140_U520 R140_U519 ; R140_U180
g7279 nand R140_U46 R140_U210 ; R140_U181
g7280 and R140_U527 R140_U526 ; R140_U182
g7281 nand R140_U119 R140_U313 ; R140_U183
g7282 and R140_U534 R140_U533 ; R140_U184
g7283 nand R140_U294 R140_U311 ; R140_U185
g7284 not R140_U79 ; R140_U186
g7285 not R140_U165 ; R140_U187
g7286 not R140_U144 ; R140_U188
g7287 or SI_2_ U108 ; R140_U189
g7288 nand R140_U304 R140_U189 ; R140_U190
g7289 not R140_U28 ; R140_U191
g7290 not R140_U138 ; R140_U192
g7291 or SI_3_ U97 ; R140_U193
g7292 nand U97 SI_3_ ; R140_U194
g7293 or SI_4_ U94 ; R140_U195
g7294 not R140_U23 ; R140_U196
g7295 or SI_5_ U93 ; R140_U197
g7296 nand U93 SI_5_ ; R140_U198
g7297 or SI_6_ U92 ; R140_U199
g7298 nand U92 SI_6_ ; R140_U200
g7299 or SI_7_ U91 ; R140_U201
g7300 not R140_U16 ; R140_U202
g7301 or SI_8_ U90 ; R140_U203
g7302 nand U90 SI_8_ ; R140_U204
g7303 or SI_9_ U89 ; R140_U205
g7304 nand SI_9_ U89 ; R140_U206
g7305 or SI_10_ U118 ; R140_U207
g7306 nand U118 SI_10_ ; R140_U208
g7307 or SI_11_ U117 ; R140_U209
g7308 nand R140_U209 R140_U183 ; R140_U210
g7309 not R140_U46 ; R140_U211
g7310 not R140_U181 ; R140_U212
g7311 or SI_12_ U116 ; R140_U213
g7312 nand U116 SI_12_ ; R140_U214
g7313 not R140_U179 ; R140_U215
g7314 or SI_13_ U115 ; R140_U216
g7315 nand U115 SI_13_ ; R140_U217
g7316 not R140_U177 ; R140_U218
g7317 or SI_14_ U114 ; R140_U219
g7318 nand U114 SI_14_ ; R140_U220
g7319 not R140_U175 ; R140_U221
g7320 or SI_15_ U113 ; R140_U222
g7321 nand R140_U222 R140_U175 ; R140_U223
g7322 nand U113 SI_15_ ; R140_U224
g7323 not R140_U173 ; R140_U225
g7324 or SI_16_ U112 ; R140_U226
g7325 nand R140_U226 R140_U173 ; R140_U227
g7326 nand U112 SI_16_ ; R140_U228
g7327 not R140_U171 ; R140_U229
g7328 or SI_17_ U111 ; R140_U230
g7329 nand R140_U230 R140_U171 ; R140_U231
g7330 nand U111 SI_17_ ; R140_U232
g7331 not R140_U169 ; R140_U233
g7332 or SI_18_ U110 ; R140_U234
g7333 nand R140_U234 R140_U169 ; R140_U235
g7334 nand U110 SI_18_ ; R140_U236
g7335 not R140_U167 ; R140_U237
g7336 or SI_19_ U109 ; R140_U238
g7337 nand R140_U238 R140_U167 ; R140_U239
g7338 nand U109 SI_19_ ; R140_U240
g7339 not R140_U164 ; R140_U241
g7340 or SI_20_ U107 ; R140_U242
g7341 nand R140_U242 R140_U164 ; R140_U243
g7342 nand U107 SI_20_ ; R140_U244
g7343 not R140_U162 ; R140_U245
g7344 or SI_21_ U106 ; R140_U246
g7345 nand R140_U246 R140_U162 ; R140_U247
g7346 nand U106 SI_21_ ; R140_U248
g7347 not R140_U160 ; R140_U249
g7348 or SI_22_ U105 ; R140_U250
g7349 nand R140_U250 R140_U160 ; R140_U251
g7350 nand U105 SI_22_ ; R140_U252
g7351 not R140_U158 ; R140_U253
g7352 or SI_23_ U104 ; R140_U254
g7353 nand R140_U254 R140_U158 ; R140_U255
g7354 nand U104 SI_23_ ; R140_U256
g7355 not R140_U156 ; R140_U257
g7356 or SI_24_ U103 ; R140_U258
g7357 nand R140_U258 R140_U156 ; R140_U259
g7358 nand U103 SI_24_ ; R140_U260
g7359 not R140_U154 ; R140_U261
g7360 or SI_25_ U102 ; R140_U262
g7361 nand R140_U262 R140_U154 ; R140_U263
g7362 nand U102 SI_25_ ; R140_U264
g7363 not R140_U152 ; R140_U265
g7364 or SI_26_ U101 ; R140_U266
g7365 nand R140_U266 R140_U152 ; R140_U267
g7366 nand U101 SI_26_ ; R140_U268
g7367 not R140_U150 ; R140_U269
g7368 or SI_27_ U100 ; R140_U270
g7369 nand R140_U270 R140_U150 ; R140_U271
g7370 nand U100 SI_27_ ; R140_U272
g7371 not R140_U148 ; R140_U273
g7372 or SI_28_ U99 ; R140_U274
g7373 nand R140_U274 R140_U148 ; R140_U275
g7374 nand U99 SI_28_ ; R140_U276
g7375 not R140_U146 ; R140_U277
g7376 or SI_29_ U98 ; R140_U278
g7377 nand R140_U278 R140_U146 ; R140_U279
g7378 nand U98 SI_29_ ; R140_U280
g7379 not R140_U143 ; R140_U281
g7380 nand U96 SI_30_ ; R140_U282
g7381 or U96 SI_30_ ; R140_U283
g7382 nand R140_U279 R140_U122 ; R140_U284
g7383 nand U120 SI_0_ U119 ; R140_U285
g7384 nand U119 SI_1_ ; R140_U286
g7385 nand R140_U191 R140_U193 ; R140_U287
g7386 nand R140_U196 R140_U197 ; R140_U288
g7387 not R140_U35 ; R140_U289
g7388 nand R140_U35 R140_U199 ; R140_U290
g7389 nand R140_U202 R140_U203 ; R140_U291
g7390 nand R140_U291 R140_U204 ; R140_U292
g7391 nand R140_U292 R140_U205 ; R140_U293
g7392 not R140_U82 ; R140_U294
g7393 nand R140_U82 R140_U207 ; R140_U295
g7394 nand R140_U7 R140_U183 ; R140_U296
g7395 nand R140_U211 R140_U213 ; R140_U297
g7396 not R140_U81 ; R140_U298
g7397 nand R140_U8 R140_U183 ; R140_U299
g7398 nand R140_U81 R140_U216 ; R140_U300
g7399 not R140_U80 ; R140_U301
g7400 nand R140_U120 R140_U183 ; R140_U302
g7401 nand R140_U80 R140_U219 ; R140_U303
g7402 nand R140_U306 R140_U286 R140_U305 ; R140_U304
g7403 nand U120 SI_0_ U119 ; R140_U305
g7404 nand SI_0_ SI_1_ U120 ; R140_U306
g7405 nand R140_U201 R140_U130 ; R140_U307
g7406 not R140_U128 ; R140_U308
g7407 nand R140_U5 R140_U130 ; R140_U309
g7408 not R140_U126 ; R140_U310
g7409 nand R140_U6 R140_U130 ; R140_U311
g7410 not R140_U185 ; R140_U312
g7411 nand R140_U118 R140_U130 ; R140_U313
g7412 not R140_U183 ; R140_U314
g7413 nand R140_U195 R140_U136 ; R140_U315
g7414 not R140_U134 ; R140_U316
g7415 nand R140_U4 R140_U136 ; R140_U317
g7416 not R140_U132 ; R140_U318
g7417 nand R140_U115 R140_U136 ; R140_U319
g7418 not R140_U130 ; R140_U320
g7419 nand R140_U113 R140_U144 ; R140_U321
g7420 not R140_U136 ; R140_U322
g7421 nand R140_U123 R140_U143 ; R140_U323
g7422 nand R140_U186 U119 ; R140_U324
g7423 nand U89 R140_U34 ; R140_U325
g7424 nand SI_9_ R140_U33 ; R140_U326
g7425 nand U89 R140_U34 ; R140_U327
g7426 nand SI_9_ R140_U33 ; R140_U328
g7427 nand R140_U328 R140_U327 ; R140_U329
g7428 nand R140_U125 R140_U126 ; R140_U330
g7429 nand R140_U310 R140_U329 ; R140_U331
g7430 nand U90 R140_U12 ; R140_U332
g7431 nand SI_8_ R140_U13 ; R140_U333
g7432 nand U90 R140_U12 ; R140_U334
g7433 nand SI_8_ R140_U13 ; R140_U335
g7434 nand R140_U335 R140_U334 ; R140_U336
g7435 nand R140_U127 R140_U128 ; R140_U337
g7436 nand R140_U308 R140_U336 ; R140_U338
g7437 nand U91 R140_U14 ; R140_U339
g7438 nand SI_7_ R140_U15 ; R140_U340
g7439 nand U91 R140_U14 ; R140_U341
g7440 nand SI_7_ R140_U15 ; R140_U342
g7441 nand R140_U342 R140_U341 ; R140_U343
g7442 nand R140_U129 R140_U130 ; R140_U344
g7443 nand R140_U320 R140_U343 ; R140_U345
g7444 nand U92 R140_U17 ; R140_U346
g7445 nand SI_6_ R140_U18 ; R140_U347
g7446 nand U92 R140_U17 ; R140_U348
g7447 nand SI_6_ R140_U18 ; R140_U349
g7448 nand R140_U349 R140_U348 ; R140_U350
g7449 nand R140_U131 R140_U132 ; R140_U351
g7450 nand R140_U318 R140_U350 ; R140_U352
g7451 nand U93 R140_U19 ; R140_U353
g7452 nand SI_5_ R140_U20 ; R140_U354
g7453 nand U93 R140_U19 ; R140_U355
g7454 nand SI_5_ R140_U20 ; R140_U356
g7455 nand R140_U356 R140_U355 ; R140_U357
g7456 nand R140_U133 R140_U134 ; R140_U358
g7457 nand R140_U316 R140_U357 ; R140_U359
g7458 nand U94 R140_U21 ; R140_U360
g7459 nand SI_4_ R140_U22 ; R140_U361
g7460 nand U94 R140_U21 ; R140_U362
g7461 nand SI_4_ R140_U22 ; R140_U363
g7462 nand R140_U363 R140_U362 ; R140_U364
g7463 nand R140_U135 R140_U136 ; R140_U365
g7464 nand R140_U322 R140_U364 ; R140_U366
g7465 nand U97 R140_U24 ; R140_U367
g7466 nand SI_3_ R140_U25 ; R140_U368
g7467 nand U97 R140_U24 ; R140_U369
g7468 nand SI_3_ R140_U25 ; R140_U370
g7469 nand R140_U370 R140_U369 ; R140_U371
g7470 nand R140_U137 R140_U138 ; R140_U372
g7471 nand R140_U192 R140_U371 ; R140_U373
g7472 nand U95 R140_U140 ; R140_U374
g7473 nand SI_31_ R140_U139 ; R140_U375
g7474 nand R140_U375 R140_U374 ; R140_U376
g7475 nand U95 R140_U140 ; R140_U377
g7476 nand SI_31_ R140_U139 ; R140_U378
g7477 nand R140_U9 R140_U77 R140_U78 ; R140_U379
g7478 nand SI_30_ R140_U376 U96 ; R140_U380
g7479 nand U96 R140_U77 ; R140_U381
g7480 nand SI_30_ R140_U78 ; R140_U382
g7481 nand U96 R140_U77 ; R140_U383
g7482 nand SI_30_ R140_U78 ; R140_U384
g7483 nand R140_U384 R140_U383 ; R140_U385
g7484 nand R140_U142 R140_U143 ; R140_U386
g7485 nand R140_U281 R140_U385 ; R140_U387
g7486 nand U108 R140_U26 ; R140_U388
g7487 nand SI_2_ R140_U27 ; R140_U389
g7488 nand U108 R140_U26 ; R140_U390
g7489 nand SI_2_ R140_U27 ; R140_U391
g7490 nand R140_U391 R140_U390 ; R140_U392
g7491 nand R140_U389 R140_U388 R140_U144 ; R140_U393
g7492 nand R140_U188 R140_U392 ; R140_U394
g7493 nand U98 R140_U75 ; R140_U395
g7494 nand SI_29_ R140_U76 ; R140_U396
g7495 nand U98 R140_U75 ; R140_U397
g7496 nand SI_29_ R140_U76 ; R140_U398
g7497 nand R140_U398 R140_U397 ; R140_U399
g7498 nand R140_U145 R140_U146 ; R140_U400
g7499 nand R140_U277 R140_U399 ; R140_U401
g7500 nand U99 R140_U73 ; R140_U402
g7501 nand SI_28_ R140_U74 ; R140_U403
g7502 nand U99 R140_U73 ; R140_U404
g7503 nand SI_28_ R140_U74 ; R140_U405
g7504 nand R140_U405 R140_U404 ; R140_U406
g7505 nand R140_U147 R140_U148 ; R140_U407
g7506 nand R140_U273 R140_U406 ; R140_U408
g7507 nand U100 R140_U71 ; R140_U409
g7508 nand SI_27_ R140_U72 ; R140_U410
g7509 nand U100 R140_U71 ; R140_U411
g7510 nand SI_27_ R140_U72 ; R140_U412
g7511 nand R140_U412 R140_U411 ; R140_U413
g7512 nand R140_U149 R140_U150 ; R140_U414
g7513 nand R140_U269 R140_U413 ; R140_U415
g7514 nand U101 R140_U69 ; R140_U416
g7515 nand SI_26_ R140_U70 ; R140_U417
g7516 nand U101 R140_U69 ; R140_U418
g7517 nand SI_26_ R140_U70 ; R140_U419
g7518 nand R140_U419 R140_U418 ; R140_U420
g7519 nand R140_U151 R140_U152 ; R140_U421
g7520 nand R140_U265 R140_U420 ; R140_U422
g7521 nand U102 R140_U67 ; R140_U423
g7522 nand SI_25_ R140_U68 ; R140_U424
g7523 nand U102 R140_U67 ; R140_U425
g7524 nand SI_25_ R140_U68 ; R140_U426
g7525 nand R140_U426 R140_U425 ; R140_U427
g7526 nand R140_U153 R140_U154 ; R140_U428
g7527 nand R140_U261 R140_U427 ; R140_U429
g7528 nand U103 R140_U65 ; R140_U430
g7529 nand SI_24_ R140_U66 ; R140_U431
g7530 nand U103 R140_U65 ; R140_U432
g7531 nand SI_24_ R140_U66 ; R140_U433
g7532 nand R140_U433 R140_U432 ; R140_U434
g7533 nand R140_U155 R140_U156 ; R140_U435
g7534 nand R140_U257 R140_U434 ; R140_U436
g7535 nand U104 R140_U63 ; R140_U437
g7536 nand SI_23_ R140_U64 ; R140_U438
g7537 nand U104 R140_U63 ; R140_U439
g7538 nand SI_23_ R140_U64 ; R140_U440
g7539 nand R140_U440 R140_U439 ; R140_U441
g7540 nand R140_U157 R140_U158 ; R140_U442
g7541 nand R140_U253 R140_U441 ; R140_U443
g7542 nand U105 R140_U61 ; R140_U444
g7543 nand SI_22_ R140_U62 ; R140_U445
g7544 nand U105 R140_U61 ; R140_U446
g7545 nand SI_22_ R140_U62 ; R140_U447
g7546 nand R140_U447 R140_U446 ; R140_U448
g7547 nand R140_U159 R140_U160 ; R140_U449
g7548 nand R140_U249 R140_U448 ; R140_U450
g7549 nand U106 R140_U59 ; R140_U451
g7550 nand SI_21_ R140_U60 ; R140_U452
g7551 nand U106 R140_U59 ; R140_U453
g7552 nand SI_21_ R140_U60 ; R140_U454
g7553 nand R140_U454 R140_U453 ; R140_U455
g7554 nand R140_U161 R140_U162 ; R140_U456
g7555 nand R140_U245 R140_U455 ; R140_U457
g7556 nand U107 R140_U57 ; R140_U458
g7557 nand SI_20_ R140_U58 ; R140_U459
g7558 nand U107 R140_U57 ; R140_U460
g7559 nand SI_20_ R140_U58 ; R140_U461
g7560 nand R140_U461 R140_U460 ; R140_U462
g7561 nand R140_U163 R140_U164 ; R140_U463
g7562 nand R140_U241 R140_U462 ; R140_U464
g7563 nand U119 R140_U165 ; R140_U465
g7564 nand R140_U187 R140_U32 ; R140_U466
g7565 nand R140_U466 R140_U465 ; R140_U467
g7566 nand R140_U165 R140_U32 SI_1_ ; R140_U468
g7567 nand R140_U467 R140_U29 ; R140_U469
g7568 nand U109 R140_U55 ; R140_U470
g7569 nand SI_19_ R140_U56 ; R140_U471
g7570 nand U109 R140_U55 ; R140_U472
g7571 nand SI_19_ R140_U56 ; R140_U473
g7572 nand R140_U473 R140_U472 ; R140_U474
g7573 nand R140_U166 R140_U167 ; R140_U475
g7574 nand R140_U237 R140_U474 ; R140_U476
g7575 nand U110 R140_U53 ; R140_U477
g7576 nand SI_18_ R140_U54 ; R140_U478
g7577 nand U110 R140_U53 ; R140_U479
g7578 nand SI_18_ R140_U54 ; R140_U480
g7579 nand R140_U480 R140_U479 ; R140_U481
g7580 nand R140_U168 R140_U169 ; R140_U482
g7581 nand R140_U233 R140_U481 ; R140_U483
g7582 nand U111 R140_U51 ; R140_U484
g7583 nand SI_17_ R140_U52 ; R140_U485
g7584 nand U111 R140_U51 ; R140_U486
g7585 nand SI_17_ R140_U52 ; R140_U487
g7586 nand R140_U487 R140_U486 ; R140_U488
g7587 nand R140_U170 R140_U171 ; R140_U489
g7588 nand R140_U229 R140_U488 ; R140_U490
g7589 nand U112 R140_U49 ; R140_U491
g7590 nand SI_16_ R140_U50 ; R140_U492
g7591 nand U112 R140_U49 ; R140_U493
g7592 nand SI_16_ R140_U50 ; R140_U494
g7593 nand R140_U494 R140_U493 ; R140_U495
g7594 nand R140_U172 R140_U173 ; R140_U496
g7595 nand R140_U225 R140_U495 ; R140_U497
g7596 nand U113 R140_U47 ; R140_U498
g7597 nand SI_15_ R140_U48 ; R140_U499
g7598 nand U113 R140_U47 ; R140_U500
g7599 nand SI_15_ R140_U48 ; R140_U501
g7600 nand R140_U501 R140_U500 ; R140_U502
g7601 nand R140_U174 R140_U175 ; R140_U503
g7602 nand R140_U221 R140_U502 ; R140_U504
g7603 nand U114 R140_U36 ; R140_U505
g7604 nand SI_14_ R140_U37 ; R140_U506
g7605 nand U114 R140_U36 ; R140_U507
g7606 nand SI_14_ R140_U37 ; R140_U508
g7607 nand R140_U508 R140_U507 ; R140_U509
g7608 nand R140_U176 R140_U177 ; R140_U510
g7609 nand R140_U218 R140_U509 ; R140_U511
g7610 nand U115 R140_U40 ; R140_U512
g7611 nand SI_13_ R140_U41 ; R140_U513
g7612 nand U115 R140_U40 ; R140_U514
g7613 nand SI_13_ R140_U41 ; R140_U515
g7614 nand R140_U515 R140_U514 ; R140_U516
g7615 nand R140_U178 R140_U179 ; R140_U517
g7616 nand R140_U215 R140_U516 ; R140_U518
g7617 nand U116 R140_U42 ; R140_U519
g7618 nand SI_12_ R140_U43 ; R140_U520
g7619 nand U116 R140_U42 ; R140_U521
g7620 nand SI_12_ R140_U43 ; R140_U522
g7621 nand R140_U522 R140_U521 ; R140_U523
g7622 nand R140_U180 R140_U181 ; R140_U524
g7623 nand R140_U212 R140_U523 ; R140_U525
g7624 nand U117 R140_U44 ; R140_U526
g7625 nand SI_11_ R140_U45 ; R140_U527
g7626 nand U117 R140_U44 ; R140_U528
g7627 nand SI_11_ R140_U45 ; R140_U529
g7628 nand R140_U529 R140_U528 ; R140_U530
g7629 nand R140_U182 R140_U183 ; R140_U531
g7630 nand R140_U314 R140_U530 ; R140_U532
g7631 nand U118 R140_U38 ; R140_U533
g7632 nand SI_10_ R140_U39 ; R140_U534
g7633 nand U118 R140_U38 ; R140_U535
g7634 nand SI_10_ R140_U39 ; R140_U536
g7635 nand R140_U536 R140_U535 ; R140_U537
g7636 nand R140_U184 R140_U185 ; R140_U538
g7637 nand R140_U312 R140_U537 ; R140_U539
g7638 nand U120 R140_U30 ; R140_U540
g7639 nand SI_0_ R140_U31 ; R140_U541
g7640 not P2_ADDR_REG_19__SCAN_IN ; LT_1079_19_U6
g7641 not P1_REG3_REG_3__SCAN_IN ; P1_ADD_99_U4
g7642 and P1_ADD_99_U102 P1_REG3_REG_28__SCAN_IN P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U5
g7643 not P1_REG3_REG_4__SCAN_IN ; P1_ADD_99_U6
g7644 nand P1_REG3_REG_4__SCAN_IN P1_REG3_REG_3__SCAN_IN ; P1_ADD_99_U7
g7645 not P1_REG3_REG_5__SCAN_IN ; P1_ADD_99_U8
g7646 nand P1_ADD_99_U80 P1_REG3_REG_5__SCAN_IN ; P1_ADD_99_U9
g7647 not P1_REG3_REG_6__SCAN_IN ; P1_ADD_99_U10
g7648 nand P1_ADD_99_U81 P1_REG3_REG_6__SCAN_IN ; P1_ADD_99_U11
g7649 not P1_REG3_REG_7__SCAN_IN ; P1_ADD_99_U12
g7650 nand P1_ADD_99_U82 P1_REG3_REG_7__SCAN_IN ; P1_ADD_99_U13
g7651 not P1_REG3_REG_8__SCAN_IN ; P1_ADD_99_U14
g7652 not P1_REG3_REG_9__SCAN_IN ; P1_ADD_99_U15
g7653 nand P1_ADD_99_U83 P1_REG3_REG_8__SCAN_IN ; P1_ADD_99_U16
g7654 nand P1_ADD_99_U84 P1_REG3_REG_9__SCAN_IN ; P1_ADD_99_U17
g7655 not P1_REG3_REG_10__SCAN_IN ; P1_ADD_99_U18
g7656 nand P1_ADD_99_U85 P1_REG3_REG_10__SCAN_IN ; P1_ADD_99_U19
g7657 not P1_REG3_REG_11__SCAN_IN ; P1_ADD_99_U20
g7658 nand P1_ADD_99_U86 P1_REG3_REG_11__SCAN_IN ; P1_ADD_99_U21
g7659 not P1_REG3_REG_12__SCAN_IN ; P1_ADD_99_U22
g7660 nand P1_ADD_99_U87 P1_REG3_REG_12__SCAN_IN ; P1_ADD_99_U23
g7661 not P1_REG3_REG_13__SCAN_IN ; P1_ADD_99_U24
g7662 nand P1_ADD_99_U88 P1_REG3_REG_13__SCAN_IN ; P1_ADD_99_U25
g7663 not P1_REG3_REG_14__SCAN_IN ; P1_ADD_99_U26
g7664 nand P1_ADD_99_U89 P1_REG3_REG_14__SCAN_IN ; P1_ADD_99_U27
g7665 not P1_REG3_REG_15__SCAN_IN ; P1_ADD_99_U28
g7666 nand P1_ADD_99_U90 P1_REG3_REG_15__SCAN_IN ; P1_ADD_99_U29
g7667 not P1_REG3_REG_16__SCAN_IN ; P1_ADD_99_U30
g7668 nand P1_ADD_99_U91 P1_REG3_REG_16__SCAN_IN ; P1_ADD_99_U31
g7669 not P1_REG3_REG_17__SCAN_IN ; P1_ADD_99_U32
g7670 nand P1_ADD_99_U92 P1_REG3_REG_17__SCAN_IN ; P1_ADD_99_U33
g7671 not P1_REG3_REG_18__SCAN_IN ; P1_ADD_99_U34
g7672 nand P1_ADD_99_U93 P1_REG3_REG_18__SCAN_IN ; P1_ADD_99_U35
g7673 not P1_REG3_REG_19__SCAN_IN ; P1_ADD_99_U36
g7674 nand P1_ADD_99_U94 P1_REG3_REG_19__SCAN_IN ; P1_ADD_99_U37
g7675 not P1_REG3_REG_20__SCAN_IN ; P1_ADD_99_U38
g7676 nand P1_ADD_99_U95 P1_REG3_REG_20__SCAN_IN ; P1_ADD_99_U39
g7677 not P1_REG3_REG_21__SCAN_IN ; P1_ADD_99_U40
g7678 nand P1_ADD_99_U96 P1_REG3_REG_21__SCAN_IN ; P1_ADD_99_U41
g7679 not P1_REG3_REG_22__SCAN_IN ; P1_ADD_99_U42
g7680 nand P1_ADD_99_U97 P1_REG3_REG_22__SCAN_IN ; P1_ADD_99_U43
g7681 not P1_REG3_REG_23__SCAN_IN ; P1_ADD_99_U44
g7682 nand P1_ADD_99_U98 P1_REG3_REG_23__SCAN_IN ; P1_ADD_99_U45
g7683 not P1_REG3_REG_24__SCAN_IN ; P1_ADD_99_U46
g7684 nand P1_ADD_99_U99 P1_REG3_REG_24__SCAN_IN ; P1_ADD_99_U47
g7685 not P1_REG3_REG_25__SCAN_IN ; P1_ADD_99_U48
g7686 nand P1_ADD_99_U100 P1_REG3_REG_25__SCAN_IN ; P1_ADD_99_U49
g7687 not P1_REG3_REG_26__SCAN_IN ; P1_ADD_99_U50
g7688 nand P1_ADD_99_U101 P1_REG3_REG_26__SCAN_IN ; P1_ADD_99_U51
g7689 not P1_REG3_REG_28__SCAN_IN ; P1_ADD_99_U52
g7690 not P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U53
g7691 nand P1_ADD_99_U105 P1_ADD_99_U104 ; P1_ADD_99_U54
g7692 nand P1_ADD_99_U107 P1_ADD_99_U106 ; P1_ADD_99_U55
g7693 nand P1_ADD_99_U109 P1_ADD_99_U108 ; P1_ADD_99_U56
g7694 nand P1_ADD_99_U111 P1_ADD_99_U110 ; P1_ADD_99_U57
g7695 nand P1_ADD_99_U113 P1_ADD_99_U112 ; P1_ADD_99_U58
g7696 nand P1_ADD_99_U115 P1_ADD_99_U114 ; P1_ADD_99_U59
g7697 nand P1_ADD_99_U117 P1_ADD_99_U116 ; P1_ADD_99_U60
g7698 nand P1_ADD_99_U119 P1_ADD_99_U118 ; P1_ADD_99_U61
g7699 nand P1_ADD_99_U121 P1_ADD_99_U120 ; P1_ADD_99_U62
g7700 nand P1_ADD_99_U123 P1_ADD_99_U122 ; P1_ADD_99_U63
g7701 nand P1_ADD_99_U125 P1_ADD_99_U124 ; P1_ADD_99_U64
g7702 nand P1_ADD_99_U127 P1_ADD_99_U126 ; P1_ADD_99_U65
g7703 nand P1_ADD_99_U129 P1_ADD_99_U128 ; P1_ADD_99_U66
g7704 nand P1_ADD_99_U131 P1_ADD_99_U130 ; P1_ADD_99_U67
g7705 nand P1_ADD_99_U133 P1_ADD_99_U132 ; P1_ADD_99_U68
g7706 nand P1_ADD_99_U135 P1_ADD_99_U134 ; P1_ADD_99_U69
g7707 nand P1_ADD_99_U137 P1_ADD_99_U136 ; P1_ADD_99_U70
g7708 nand P1_ADD_99_U139 P1_ADD_99_U138 ; P1_ADD_99_U71
g7709 nand P1_ADD_99_U141 P1_ADD_99_U140 ; P1_ADD_99_U72
g7710 nand P1_ADD_99_U143 P1_ADD_99_U142 ; P1_ADD_99_U73
g7711 nand P1_ADD_99_U145 P1_ADD_99_U144 ; P1_ADD_99_U74
g7712 nand P1_ADD_99_U147 P1_ADD_99_U146 ; P1_ADD_99_U75
g7713 nand P1_ADD_99_U149 P1_ADD_99_U148 ; P1_ADD_99_U76
g7714 nand P1_ADD_99_U151 P1_ADD_99_U150 ; P1_ADD_99_U77
g7715 nand P1_ADD_99_U153 P1_ADD_99_U152 ; P1_ADD_99_U78
g7716 nand P1_ADD_99_U102 P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U79
g7717 not P1_ADD_99_U7 ; P1_ADD_99_U80
g7718 not P1_ADD_99_U9 ; P1_ADD_99_U81
g7719 not P1_ADD_99_U11 ; P1_ADD_99_U82
g7720 not P1_ADD_99_U13 ; P1_ADD_99_U83
g7721 not P1_ADD_99_U16 ; P1_ADD_99_U84
g7722 not P1_ADD_99_U17 ; P1_ADD_99_U85
g7723 not P1_ADD_99_U19 ; P1_ADD_99_U86
g7724 not P1_ADD_99_U21 ; P1_ADD_99_U87
g7725 not P1_ADD_99_U23 ; P1_ADD_99_U88
g7726 not P1_ADD_99_U25 ; P1_ADD_99_U89
g7727 not P1_ADD_99_U27 ; P1_ADD_99_U90
g7728 not P1_ADD_99_U29 ; P1_ADD_99_U91
g7729 not P1_ADD_99_U31 ; P1_ADD_99_U92
g7730 not P1_ADD_99_U33 ; P1_ADD_99_U93
g7731 not P1_ADD_99_U35 ; P1_ADD_99_U94
g7732 not P1_ADD_99_U37 ; P1_ADD_99_U95
g7733 not P1_ADD_99_U39 ; P1_ADD_99_U96
g7734 not P1_ADD_99_U41 ; P1_ADD_99_U97
g7735 not P1_ADD_99_U43 ; P1_ADD_99_U98
g7736 not P1_ADD_99_U45 ; P1_ADD_99_U99
g7737 not P1_ADD_99_U47 ; P1_ADD_99_U100
g7738 not P1_ADD_99_U49 ; P1_ADD_99_U101
g7739 not P1_ADD_99_U51 ; P1_ADD_99_U102
g7740 not P1_ADD_99_U79 ; P1_ADD_99_U103
g7741 nand P1_ADD_99_U16 P1_REG3_REG_9__SCAN_IN ; P1_ADD_99_U104
g7742 nand P1_ADD_99_U84 P1_ADD_99_U15 ; P1_ADD_99_U105
g7743 nand P1_ADD_99_U13 P1_REG3_REG_8__SCAN_IN ; P1_ADD_99_U106
g7744 nand P1_ADD_99_U83 P1_ADD_99_U14 ; P1_ADD_99_U107
g7745 nand P1_ADD_99_U11 P1_REG3_REG_7__SCAN_IN ; P1_ADD_99_U108
g7746 nand P1_ADD_99_U82 P1_ADD_99_U12 ; P1_ADD_99_U109
g7747 nand P1_ADD_99_U9 P1_REG3_REG_6__SCAN_IN ; P1_ADD_99_U110
g7748 nand P1_ADD_99_U81 P1_ADD_99_U10 ; P1_ADD_99_U111
g7749 nand P1_ADD_99_U7 P1_REG3_REG_5__SCAN_IN ; P1_ADD_99_U112
g7750 nand P1_ADD_99_U80 P1_ADD_99_U8 ; P1_ADD_99_U113
g7751 nand P1_ADD_99_U4 P1_REG3_REG_4__SCAN_IN ; P1_ADD_99_U114
g7752 nand P1_ADD_99_U6 P1_REG3_REG_3__SCAN_IN ; P1_ADD_99_U115
g7753 nand P1_ADD_99_U79 P1_REG3_REG_28__SCAN_IN ; P1_ADD_99_U116
g7754 nand P1_ADD_99_U103 P1_ADD_99_U52 ; P1_ADD_99_U117
g7755 nand P1_ADD_99_U51 P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U118
g7756 nand P1_ADD_99_U102 P1_ADD_99_U53 ; P1_ADD_99_U119
g7757 nand P1_ADD_99_U49 P1_REG3_REG_26__SCAN_IN ; P1_ADD_99_U120
g7758 nand P1_ADD_99_U101 P1_ADD_99_U50 ; P1_ADD_99_U121
g7759 nand P1_ADD_99_U47 P1_REG3_REG_25__SCAN_IN ; P1_ADD_99_U122
g7760 nand P1_ADD_99_U100 P1_ADD_99_U48 ; P1_ADD_99_U123
g7761 nand P1_ADD_99_U45 P1_REG3_REG_24__SCAN_IN ; P1_ADD_99_U124
g7762 nand P1_ADD_99_U99 P1_ADD_99_U46 ; P1_ADD_99_U125
g7763 nand P1_ADD_99_U43 P1_REG3_REG_23__SCAN_IN ; P1_ADD_99_U126
g7764 nand P1_ADD_99_U98 P1_ADD_99_U44 ; P1_ADD_99_U127
g7765 nand P1_ADD_99_U41 P1_REG3_REG_22__SCAN_IN ; P1_ADD_99_U128
g7766 nand P1_ADD_99_U97 P1_ADD_99_U42 ; P1_ADD_99_U129
g7767 nand P1_ADD_99_U39 P1_REG3_REG_21__SCAN_IN ; P1_ADD_99_U130
g7768 nand P1_ADD_99_U96 P1_ADD_99_U40 ; P1_ADD_99_U131
g7769 nand P1_ADD_99_U37 P1_REG3_REG_20__SCAN_IN ; P1_ADD_99_U132
g7770 nand P1_ADD_99_U95 P1_ADD_99_U38 ; P1_ADD_99_U133
g7771 nand P1_ADD_99_U35 P1_REG3_REG_19__SCAN_IN ; P1_ADD_99_U134
g7772 nand P1_ADD_99_U94 P1_ADD_99_U36 ; P1_ADD_99_U135
g7773 nand P1_ADD_99_U33 P1_REG3_REG_18__SCAN_IN ; P1_ADD_99_U136
g7774 nand P1_ADD_99_U93 P1_ADD_99_U34 ; P1_ADD_99_U137
g7775 nand P1_ADD_99_U31 P1_REG3_REG_17__SCAN_IN ; P1_ADD_99_U138
g7776 nand P1_ADD_99_U92 P1_ADD_99_U32 ; P1_ADD_99_U139
g7777 nand P1_ADD_99_U29 P1_REG3_REG_16__SCAN_IN ; P1_ADD_99_U140
g7778 nand P1_ADD_99_U91 P1_ADD_99_U30 ; P1_ADD_99_U141
g7779 nand P1_ADD_99_U27 P1_REG3_REG_15__SCAN_IN ; P1_ADD_99_U142
g7780 nand P1_ADD_99_U90 P1_ADD_99_U28 ; P1_ADD_99_U143
g7781 nand P1_ADD_99_U25 P1_REG3_REG_14__SCAN_IN ; P1_ADD_99_U144
g7782 nand P1_ADD_99_U89 P1_ADD_99_U26 ; P1_ADD_99_U145
g7783 nand P1_ADD_99_U23 P1_REG3_REG_13__SCAN_IN ; P1_ADD_99_U146
g7784 nand P1_ADD_99_U88 P1_ADD_99_U24 ; P1_ADD_99_U147
g7785 nand P1_ADD_99_U21 P1_REG3_REG_12__SCAN_IN ; P1_ADD_99_U148
g7786 nand P1_ADD_99_U87 P1_ADD_99_U22 ; P1_ADD_99_U149
g7787 nand P1_ADD_99_U19 P1_REG3_REG_11__SCAN_IN ; P1_ADD_99_U150
g7788 nand P1_ADD_99_U86 P1_ADD_99_U20 ; P1_ADD_99_U151
g7789 nand P1_ADD_99_U17 P1_REG3_REG_10__SCAN_IN ; P1_ADD_99_U152
g7790 nand P1_ADD_99_U85 P1_ADD_99_U18 ; P1_ADD_99_U153
g7791 and P1_R1105_U95 P1_R1105_U94 ; P1_R1105_U4
g7792 and P1_R1105_U96 P1_R1105_U97 ; P1_R1105_U5
g7793 and P1_R1105_U113 P1_R1105_U112 ; P1_R1105_U6
g7794 and P1_R1105_U155 P1_R1105_U154 ; P1_R1105_U7
g7795 and P1_R1105_U164 P1_R1105_U163 ; P1_R1105_U8
g7796 and P1_R1105_U182 P1_R1105_U181 ; P1_R1105_U9
g7797 and P1_R1105_U218 P1_R1105_U215 ; P1_R1105_U10
g7798 and P1_R1105_U211 P1_R1105_U208 ; P1_R1105_U11
g7799 and P1_R1105_U202 P1_R1105_U199 ; P1_R1105_U12
g7800 and P1_R1105_U196 P1_R1105_U192 ; P1_R1105_U13
g7801 and P1_R1105_U151 P1_R1105_U148 ; P1_R1105_U14
g7802 and P1_R1105_U143 P1_R1105_U140 ; P1_R1105_U15
g7803 and P1_R1105_U129 P1_R1105_U126 ; P1_R1105_U16
g7804 not P1_REG2_REG_6__SCAN_IN ; P1_R1105_U17
g7805 not P1_U3470 ; P1_R1105_U18
g7806 not P1_U3473 ; P1_R1105_U19
g7807 nand P1_U3470 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U20
g7808 not P1_REG2_REG_7__SCAN_IN ; P1_R1105_U21
g7809 not P1_REG2_REG_4__SCAN_IN ; P1_R1105_U22
g7810 not P1_U3464 ; P1_R1105_U23
g7811 not P1_U3467 ; P1_R1105_U24
g7812 not P1_REG2_REG_2__SCAN_IN ; P1_R1105_U25
g7813 not P1_U3458 ; P1_R1105_U26
g7814 not P1_REG2_REG_0__SCAN_IN ; P1_R1105_U27
g7815 not P1_U3449 ; P1_R1105_U28
g7816 nand P1_U3449 P1_REG2_REG_0__SCAN_IN ; P1_R1105_U29
g7817 not P1_REG2_REG_3__SCAN_IN ; P1_R1105_U30
g7818 not P1_U3461 ; P1_R1105_U31
g7819 nand P1_U3464 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U32
g7820 not P1_REG2_REG_5__SCAN_IN ; P1_R1105_U33
g7821 not P1_REG2_REG_8__SCAN_IN ; P1_R1105_U34
g7822 not P1_U3476 ; P1_R1105_U35
g7823 not P1_U3479 ; P1_R1105_U36
g7824 not P1_REG2_REG_9__SCAN_IN ; P1_R1105_U37
g7825 nand P1_R1105_U49 P1_R1105_U121 ; P1_R1105_U38
g7826 nand P1_R1105_U110 P1_R1105_U108 P1_R1105_U109 ; P1_R1105_U39
g7827 nand P1_R1105_U98 P1_R1105_U99 ; P1_R1105_U40
g7828 nand P1_U3455 P1_REG2_REG_1__SCAN_IN ; P1_R1105_U41
g7829 nand P1_R1105_U136 P1_R1105_U134 P1_R1105_U135 ; P1_R1105_U42
g7830 nand P1_R1105_U132 P1_R1105_U131 ; P1_R1105_U43
g7831 not P1_REG2_REG_16__SCAN_IN ; P1_R1105_U44
g7832 not P1_U3500 ; P1_R1105_U45
g7833 not P1_U3503 ; P1_R1105_U46
g7834 nand P1_U3500 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U47
g7835 not P1_REG2_REG_17__SCAN_IN ; P1_R1105_U48
g7836 nand P1_U3476 P1_REG2_REG_8__SCAN_IN ; P1_R1105_U49
g7837 not P1_REG2_REG_10__SCAN_IN ; P1_R1105_U50
g7838 not P1_U3482 ; P1_R1105_U51
g7839 not P1_REG2_REG_12__SCAN_IN ; P1_R1105_U52
g7840 not P1_U3488 ; P1_R1105_U53
g7841 not P1_REG2_REG_11__SCAN_IN ; P1_R1105_U54
g7842 not P1_U3485 ; P1_R1105_U55
g7843 nand P1_U3485 P1_REG2_REG_11__SCAN_IN ; P1_R1105_U56
g7844 not P1_REG2_REG_13__SCAN_IN ; P1_R1105_U57
g7845 not P1_U3491 ; P1_R1105_U58
g7846 not P1_REG2_REG_14__SCAN_IN ; P1_R1105_U59
g7847 not P1_U3494 ; P1_R1105_U60
g7848 not P1_REG2_REG_15__SCAN_IN ; P1_R1105_U61
g7849 not P1_U3497 ; P1_R1105_U62
g7850 not P1_REG2_REG_18__SCAN_IN ; P1_R1105_U63
g7851 not P1_U3506 ; P1_R1105_U64
g7852 nand P1_R1105_U186 P1_R1105_U185 P1_R1105_U187 ; P1_R1105_U65
g7853 nand P1_R1105_U179 P1_R1105_U178 ; P1_R1105_U66
g7854 nand P1_R1105_U56 P1_R1105_U204 ; P1_R1105_U67
g7855 nand P1_R1105_U259 P1_R1105_U258 ; P1_R1105_U68
g7856 nand P1_R1105_U308 P1_R1105_U307 ; P1_R1105_U69
g7857 nand P1_R1105_U231 P1_R1105_U230 ; P1_R1105_U70
g7858 nand P1_R1105_U236 P1_R1105_U235 ; P1_R1105_U71
g7859 nand P1_R1105_U243 P1_R1105_U242 ; P1_R1105_U72
g7860 nand P1_R1105_U250 P1_R1105_U249 ; P1_R1105_U73
g7861 nand P1_R1105_U255 P1_R1105_U254 ; P1_R1105_U74
g7862 nand P1_R1105_U271 P1_R1105_U270 ; P1_R1105_U75
g7863 nand P1_R1105_U278 P1_R1105_U277 ; P1_R1105_U76
g7864 nand P1_R1105_U285 P1_R1105_U284 ; P1_R1105_U77
g7865 nand P1_R1105_U292 P1_R1105_U291 ; P1_R1105_U78
g7866 nand P1_R1105_U299 P1_R1105_U298 ; P1_R1105_U79
g7867 nand P1_R1105_U304 P1_R1105_U303 ; P1_R1105_U80
g7868 nand P1_R1105_U117 P1_R1105_U116 P1_R1105_U118 ; P1_R1105_U81
g7869 nand P1_R1105_U133 P1_R1105_U145 ; P1_R1105_U82
g7870 nand P1_R1105_U41 P1_R1105_U152 ; P1_R1105_U83
g7871 not P1_U3443 ; P1_R1105_U84
g7872 not P1_REG2_REG_19__SCAN_IN ; P1_R1105_U85
g7873 nand P1_R1105_U175 P1_R1105_U174 ; P1_R1105_U86
g7874 nand P1_R1105_U171 P1_R1105_U170 ; P1_R1105_U87
g7875 nand P1_R1105_U161 P1_R1105_U160 ; P1_R1105_U88
g7876 not P1_R1105_U32 ; P1_R1105_U89
g7877 nand P1_U3479 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U90
g7878 nand P1_U3488 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U91
g7879 not P1_R1105_U56 ; P1_R1105_U92
g7880 not P1_R1105_U49 ; P1_R1105_U93
g7881 or P1_U3467 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U94
g7882 or P1_U3464 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U95
g7883 or P1_U3461 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U96
g7884 or P1_U3458 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U97
g7885 not P1_R1105_U29 ; P1_R1105_U98
g7886 or P1_U3455 P1_REG2_REG_1__SCAN_IN ; P1_R1105_U99
g7887 not P1_R1105_U40 ; P1_R1105_U100
g7888 not P1_R1105_U41 ; P1_R1105_U101
g7889 nand P1_R1105_U40 P1_R1105_U41 ; P1_R1105_U102
g7890 nand P1_U3458 P1_R1105_U96 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U103
g7891 nand P1_R1105_U5 P1_R1105_U102 ; P1_R1105_U104
g7892 nand P1_U3461 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U105
g7893 nand P1_R1105_U105 P1_R1105_U103 P1_R1105_U104 ; P1_R1105_U106
g7894 nand P1_R1105_U33 P1_R1105_U32 ; P1_R1105_U107
g7895 nand P1_U3467 P1_R1105_U107 ; P1_R1105_U108
g7896 nand P1_R1105_U4 P1_R1105_U106 ; P1_R1105_U109
g7897 nand P1_R1105_U89 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U110
g7898 not P1_R1105_U39 ; P1_R1105_U111
g7899 or P1_U3473 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U112
g7900 or P1_U3470 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U113
g7901 not P1_R1105_U20 ; P1_R1105_U114
g7902 nand P1_R1105_U21 P1_R1105_U20 ; P1_R1105_U115
g7903 nand P1_U3473 P1_R1105_U115 ; P1_R1105_U116
g7904 nand P1_R1105_U114 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U117
g7905 nand P1_R1105_U6 P1_R1105_U39 ; P1_R1105_U118
g7906 not P1_R1105_U81 ; P1_R1105_U119
g7907 or P1_U3476 P1_REG2_REG_8__SCAN_IN ; P1_R1105_U120
g7908 nand P1_R1105_U120 P1_R1105_U81 ; P1_R1105_U121
g7909 not P1_R1105_U38 ; P1_R1105_U122
g7910 or P1_U3479 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U123
g7911 or P1_U3470 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U124
g7912 nand P1_R1105_U124 P1_R1105_U39 ; P1_R1105_U125
g7913 nand P1_R1105_U238 P1_R1105_U237 P1_R1105_U20 P1_R1105_U125 ; P1_R1105_U126
g7914 nand P1_R1105_U111 P1_R1105_U20 ; P1_R1105_U127
g7915 nand P1_U3473 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U128
g7916 nand P1_R1105_U128 P1_R1105_U6 P1_R1105_U127 ; P1_R1105_U129
g7917 or P1_U3470 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U130
g7918 nand P1_R1105_U101 P1_R1105_U97 ; P1_R1105_U131
g7919 nand P1_U3458 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U132
g7920 not P1_R1105_U43 ; P1_R1105_U133
g7921 nand P1_R1105_U100 P1_R1105_U5 ; P1_R1105_U134
g7922 nand P1_R1105_U43 P1_R1105_U96 ; P1_R1105_U135
g7923 nand P1_U3461 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U136
g7924 not P1_R1105_U42 ; P1_R1105_U137
g7925 or P1_U3464 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U138
g7926 nand P1_R1105_U138 P1_R1105_U42 ; P1_R1105_U139
g7927 nand P1_R1105_U245 P1_R1105_U244 P1_R1105_U32 P1_R1105_U139 ; P1_R1105_U140
g7928 nand P1_R1105_U137 P1_R1105_U32 ; P1_R1105_U141
g7929 nand P1_U3467 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U142
g7930 nand P1_R1105_U142 P1_R1105_U4 P1_R1105_U141 ; P1_R1105_U143
g7931 or P1_U3464 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U144
g7932 nand P1_R1105_U100 P1_R1105_U97 ; P1_R1105_U145
g7933 not P1_R1105_U82 ; P1_R1105_U146
g7934 nand P1_U3461 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U147
g7935 nand P1_R1105_U41 P1_R1105_U40 P1_R1105_U257 P1_R1105_U256 ; P1_R1105_U148
g7936 nand P1_R1105_U41 P1_R1105_U40 ; P1_R1105_U149
g7937 nand P1_U3458 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U150
g7938 nand P1_R1105_U150 P1_R1105_U97 P1_R1105_U149 ; P1_R1105_U151
g7939 or P1_U3455 P1_REG2_REG_1__SCAN_IN ; P1_R1105_U152
g7940 not P1_R1105_U83 ; P1_R1105_U153
g7941 or P1_U3479 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U154
g7942 or P1_U3482 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U155
g7943 nand P1_R1105_U93 P1_R1105_U7 ; P1_R1105_U156
g7944 nand P1_U3482 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U157
g7945 nand P1_R1105_U157 P1_R1105_U90 P1_R1105_U156 ; P1_R1105_U158
g7946 or P1_U3482 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U159
g7947 nand P1_R1105_U120 P1_R1105_U7 P1_R1105_U81 ; P1_R1105_U160
g7948 nand P1_R1105_U159 P1_R1105_U158 ; P1_R1105_U161
g7949 not P1_R1105_U88 ; P1_R1105_U162
g7950 or P1_U3491 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U163
g7951 or P1_U3488 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U164
g7952 nand P1_R1105_U92 P1_R1105_U8 ; P1_R1105_U165
g7953 nand P1_U3491 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U166
g7954 nand P1_R1105_U166 P1_R1105_U91 P1_R1105_U165 ; P1_R1105_U167
g7955 or P1_U3485 P1_REG2_REG_11__SCAN_IN ; P1_R1105_U168
g7956 or P1_U3491 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U169
g7957 nand P1_R1105_U168 P1_R1105_U8 P1_R1105_U88 ; P1_R1105_U170
g7958 nand P1_R1105_U169 P1_R1105_U167 ; P1_R1105_U171
g7959 not P1_R1105_U87 ; P1_R1105_U172
g7960 or P1_U3494 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U173
g7961 nand P1_R1105_U173 P1_R1105_U87 ; P1_R1105_U174
g7962 nand P1_U3494 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U175
g7963 not P1_R1105_U86 ; P1_R1105_U176
g7964 or P1_U3497 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U177
g7965 nand P1_R1105_U177 P1_R1105_U86 ; P1_R1105_U178
g7966 nand P1_U3497 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U179
g7967 not P1_R1105_U66 ; P1_R1105_U180
g7968 or P1_U3503 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U181
g7969 or P1_U3500 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U182
g7970 not P1_R1105_U47 ; P1_R1105_U183
g7971 nand P1_R1105_U48 P1_R1105_U47 ; P1_R1105_U184
g7972 nand P1_U3503 P1_R1105_U184 ; P1_R1105_U185
g7973 nand P1_R1105_U183 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U186
g7974 nand P1_R1105_U9 P1_R1105_U66 ; P1_R1105_U187
g7975 not P1_R1105_U65 ; P1_R1105_U188
g7976 or P1_U3506 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U189
g7977 nand P1_R1105_U189 P1_R1105_U65 ; P1_R1105_U190
g7978 nand P1_U3506 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U191
g7979 nand P1_R1105_U261 P1_R1105_U260 P1_R1105_U191 P1_R1105_U190 ; P1_R1105_U192
g7980 nand P1_U3506 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U193
g7981 nand P1_R1105_U188 P1_R1105_U193 ; P1_R1105_U194
g7982 or P1_U3506 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U195
g7983 nand P1_R1105_U195 P1_R1105_U264 P1_R1105_U194 ; P1_R1105_U196
g7984 or P1_U3500 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U197
g7985 nand P1_R1105_U197 P1_R1105_U66 ; P1_R1105_U198
g7986 nand P1_R1105_U273 P1_R1105_U272 P1_R1105_U47 P1_R1105_U198 ; P1_R1105_U199
g7987 nand P1_R1105_U180 P1_R1105_U47 ; P1_R1105_U200
g7988 nand P1_U3503 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U201
g7989 nand P1_R1105_U201 P1_R1105_U9 P1_R1105_U200 ; P1_R1105_U202
g7990 or P1_U3500 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U203
g7991 nand P1_R1105_U168 P1_R1105_U88 ; P1_R1105_U204
g7992 not P1_R1105_U67 ; P1_R1105_U205
g7993 or P1_U3488 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U206
g7994 nand P1_R1105_U206 P1_R1105_U67 ; P1_R1105_U207
g7995 nand P1_R1105_U294 P1_R1105_U293 P1_R1105_U91 P1_R1105_U207 ; P1_R1105_U208
g7996 nand P1_R1105_U205 P1_R1105_U91 ; P1_R1105_U209
g7997 nand P1_U3491 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U210
g7998 nand P1_R1105_U210 P1_R1105_U8 P1_R1105_U209 ; P1_R1105_U211
g7999 or P1_U3488 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U212
g8000 or P1_U3479 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U213
g8001 nand P1_R1105_U213 P1_R1105_U38 ; P1_R1105_U214
g8002 nand P1_R1105_U306 P1_R1105_U305 P1_R1105_U90 P1_R1105_U214 ; P1_R1105_U215
g8003 nand P1_R1105_U122 P1_R1105_U90 ; P1_R1105_U216
g8004 nand P1_U3482 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U217
g8005 nand P1_R1105_U217 P1_R1105_U7 P1_R1105_U216 ; P1_R1105_U218
g8006 nand P1_R1105_U123 P1_R1105_U90 ; P1_R1105_U219
g8007 nand P1_R1105_U120 P1_R1105_U49 ; P1_R1105_U220
g8008 nand P1_R1105_U130 P1_R1105_U20 ; P1_R1105_U221
g8009 nand P1_R1105_U144 P1_R1105_U32 ; P1_R1105_U222
g8010 nand P1_R1105_U147 P1_R1105_U96 ; P1_R1105_U223
g8011 nand P1_R1105_U203 P1_R1105_U47 ; P1_R1105_U224
g8012 nand P1_R1105_U212 P1_R1105_U91 ; P1_R1105_U225
g8013 nand P1_R1105_U168 P1_R1105_U56 ; P1_R1105_U226
g8014 nand P1_U3479 P1_R1105_U37 ; P1_R1105_U227
g8015 nand P1_R1105_U36 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U228
g8016 nand P1_R1105_U228 P1_R1105_U227 ; P1_R1105_U229
g8017 nand P1_R1105_U219 P1_R1105_U38 ; P1_R1105_U230
g8018 nand P1_R1105_U229 P1_R1105_U122 ; P1_R1105_U231
g8019 nand P1_U3476 P1_R1105_U34 ; P1_R1105_U232
g8020 nand P1_R1105_U35 P1_REG2_REG_8__SCAN_IN ; P1_R1105_U233
g8021 nand P1_R1105_U233 P1_R1105_U232 ; P1_R1105_U234
g8022 nand P1_R1105_U220 P1_R1105_U81 ; P1_R1105_U235
g8023 nand P1_R1105_U119 P1_R1105_U234 ; P1_R1105_U236
g8024 nand P1_U3473 P1_R1105_U21 ; P1_R1105_U237
g8025 nand P1_R1105_U19 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U238
g8026 nand P1_U3470 P1_R1105_U17 ; P1_R1105_U239
g8027 nand P1_R1105_U18 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U240
g8028 nand P1_R1105_U240 P1_R1105_U239 ; P1_R1105_U241
g8029 nand P1_R1105_U221 P1_R1105_U39 ; P1_R1105_U242
g8030 nand P1_R1105_U241 P1_R1105_U111 ; P1_R1105_U243
g8031 nand P1_U3467 P1_R1105_U33 ; P1_R1105_U244
g8032 nand P1_R1105_U24 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U245
g8033 nand P1_U3464 P1_R1105_U22 ; P1_R1105_U246
g8034 nand P1_R1105_U23 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U247
g8035 nand P1_R1105_U247 P1_R1105_U246 ; P1_R1105_U248
g8036 nand P1_R1105_U222 P1_R1105_U42 ; P1_R1105_U249
g8037 nand P1_R1105_U248 P1_R1105_U137 ; P1_R1105_U250
g8038 nand P1_U3461 P1_R1105_U30 ; P1_R1105_U251
g8039 nand P1_R1105_U31 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U252
g8040 nand P1_R1105_U252 P1_R1105_U251 ; P1_R1105_U253
g8041 nand P1_R1105_U223 P1_R1105_U82 ; P1_R1105_U254
g8042 nand P1_R1105_U146 P1_R1105_U253 ; P1_R1105_U255
g8043 nand P1_U3458 P1_R1105_U25 ; P1_R1105_U256
g8044 nand P1_R1105_U26 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U257
g8045 nand P1_R1105_U98 P1_R1105_U83 ; P1_R1105_U258
g8046 nand P1_R1105_U153 P1_R1105_U29 ; P1_R1105_U259
g8047 nand P1_U3443 P1_R1105_U85 ; P1_R1105_U260
g8048 nand P1_R1105_U84 P1_REG2_REG_19__SCAN_IN ; P1_R1105_U261
g8049 nand P1_U3443 P1_R1105_U85 ; P1_R1105_U262
g8050 nand P1_R1105_U84 P1_REG2_REG_19__SCAN_IN ; P1_R1105_U263
g8051 nand P1_R1105_U263 P1_R1105_U262 ; P1_R1105_U264
g8052 nand P1_U3506 P1_R1105_U63 ; P1_R1105_U265
g8053 nand P1_R1105_U64 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U266
g8054 nand P1_U3506 P1_R1105_U63 ; P1_R1105_U267
g8055 nand P1_R1105_U64 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U268
g8056 nand P1_R1105_U268 P1_R1105_U267 ; P1_R1105_U269
g8057 nand P1_R1105_U266 P1_R1105_U265 P1_R1105_U65 ; P1_R1105_U270
g8058 nand P1_R1105_U269 P1_R1105_U188 ; P1_R1105_U271
g8059 nand P1_U3503 P1_R1105_U48 ; P1_R1105_U272
g8060 nand P1_R1105_U46 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U273
g8061 nand P1_U3500 P1_R1105_U44 ; P1_R1105_U274
g8062 nand P1_R1105_U45 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U275
g8063 nand P1_R1105_U275 P1_R1105_U274 ; P1_R1105_U276
g8064 nand P1_R1105_U224 P1_R1105_U66 ; P1_R1105_U277
g8065 nand P1_R1105_U276 P1_R1105_U180 ; P1_R1105_U278
g8066 nand P1_U3497 P1_R1105_U61 ; P1_R1105_U279
g8067 nand P1_R1105_U62 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U280
g8068 nand P1_U3497 P1_R1105_U61 ; P1_R1105_U281
g8069 nand P1_R1105_U62 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U282
g8070 nand P1_R1105_U282 P1_R1105_U281 ; P1_R1105_U283
g8071 nand P1_R1105_U280 P1_R1105_U279 P1_R1105_U86 ; P1_R1105_U284
g8072 nand P1_R1105_U176 P1_R1105_U283 ; P1_R1105_U285
g8073 nand P1_U3494 P1_R1105_U59 ; P1_R1105_U286
g8074 nand P1_R1105_U60 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U287
g8075 nand P1_U3494 P1_R1105_U59 ; P1_R1105_U288
g8076 nand P1_R1105_U60 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U289
g8077 nand P1_R1105_U289 P1_R1105_U288 ; P1_R1105_U290
g8078 nand P1_R1105_U287 P1_R1105_U286 P1_R1105_U87 ; P1_R1105_U291
g8079 nand P1_R1105_U172 P1_R1105_U290 ; P1_R1105_U292
g8080 nand P1_U3491 P1_R1105_U57 ; P1_R1105_U293
g8081 nand P1_R1105_U58 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U294
g8082 nand P1_U3488 P1_R1105_U52 ; P1_R1105_U295
g8083 nand P1_R1105_U53 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U296
g8084 nand P1_R1105_U296 P1_R1105_U295 ; P1_R1105_U297
g8085 nand P1_R1105_U225 P1_R1105_U67 ; P1_R1105_U298
g8086 nand P1_R1105_U297 P1_R1105_U205 ; P1_R1105_U299
g8087 nand P1_U3485 P1_R1105_U54 ; P1_R1105_U300
g8088 nand P1_R1105_U55 P1_REG2_REG_11__SCAN_IN ; P1_R1105_U301
g8089 nand P1_R1105_U301 P1_R1105_U300 ; P1_R1105_U302
g8090 nand P1_R1105_U226 P1_R1105_U88 ; P1_R1105_U303
g8091 nand P1_R1105_U162 P1_R1105_U302 ; P1_R1105_U304
g8092 nand P1_U3482 P1_R1105_U50 ; P1_R1105_U305
g8093 nand P1_R1105_U51 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U306
g8094 nand P1_U3449 P1_R1105_U27 ; P1_R1105_U307
g8095 nand P1_R1105_U28 P1_REG2_REG_0__SCAN_IN ; P1_R1105_U308
g8096 and P1_SUB_88_U227 P1_SUB_88_U38 ; P1_SUB_88_U6
g8097 and P1_SUB_88_U225 P1_SUB_88_U192 ; P1_SUB_88_U7
g8098 and P1_SUB_88_U224 P1_SUB_88_U35 ; P1_SUB_88_U8
g8099 and P1_SUB_88_U223 P1_SUB_88_U36 ; P1_SUB_88_U9
g8100 and P1_SUB_88_U221 P1_SUB_88_U195 ; P1_SUB_88_U10
g8101 and P1_SUB_88_U220 P1_SUB_88_U34 ; P1_SUB_88_U11
g8102 and P1_SUB_88_U219 P1_SUB_88_U197 ; P1_SUB_88_U12
g8103 and P1_SUB_88_U217 P1_SUB_88_U198 ; P1_SUB_88_U13
g8104 and P1_SUB_88_U216 P1_SUB_88_U172 ; P1_SUB_88_U14
g8105 and P1_SUB_88_U215 P1_SUB_88_U200 ; P1_SUB_88_U15
g8106 and P1_SUB_88_U213 P1_SUB_88_U201 ; P1_SUB_88_U16
g8107 and P1_SUB_88_U212 P1_SUB_88_U169 ; P1_SUB_88_U17
g8108 and P1_SUB_88_U211 P1_SUB_88_U167 ; P1_SUB_88_U18
g8109 and P1_SUB_88_U209 P1_SUB_88_U204 ; P1_SUB_88_U19
g8110 and P1_SUB_88_U208 P1_SUB_88_U33 ; P1_SUB_88_U20
g8111 and P1_SUB_88_U207 P1_SUB_88_U27 ; P1_SUB_88_U21
g8112 and P1_SUB_88_U190 P1_SUB_88_U180 ; P1_SUB_88_U22
g8113 and P1_SUB_88_U189 P1_SUB_88_U29 ; P1_SUB_88_U23
g8114 and P1_SUB_88_U188 P1_SUB_88_U30 ; P1_SUB_88_U24
g8115 and P1_SUB_88_U186 P1_SUB_88_U183 ; P1_SUB_88_U25
g8116 and P1_SUB_88_U185 P1_SUB_88_U28 ; P1_SUB_88_U26
g8117 or P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_2__SCAN_IN ; P1_SUB_88_U27
g8118 nand P1_SUB_88_U44 P1_SUB_88_U230 P1_SUB_88_U43 ; P1_SUB_88_U28
g8119 nand P1_SUB_88_U45 P1_SUB_88_U230 ; P1_SUB_88_U29
g8120 nand P1_SUB_88_U46 P1_SUB_88_U181 ; P1_SUB_88_U30
g8121 not P1_IR_REG_7__SCAN_IN ; P1_SUB_88_U31
g8122 not P1_IR_REG_3__SCAN_IN ; P1_SUB_88_U32
g8123 nand P1_SUB_88_U56 P1_SUB_88_U51 ; P1_SUB_88_U33
g8124 nand P1_SUB_88_U130 P1_SUB_88_U129 P1_SUB_88_U128 P1_SUB_88_U127 ; P1_SUB_88_U34
g8125 nand P1_SUB_88_U156 P1_SUB_88_U184 ; P1_SUB_88_U35
g8126 nand P1_SUB_88_U157 P1_SUB_88_U193 ; P1_SUB_88_U36
g8127 not P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U37
g8128 nand P1_SUB_88_U158 P1_SUB_88_U184 ; P1_SUB_88_U38
g8129 not P1_IR_REG_11__SCAN_IN ; P1_SUB_88_U39
g8130 nand P1_SUB_88_U247 P1_SUB_88_U246 ; P1_SUB_88_U40
g8131 nand P1_SUB_88_U237 P1_SUB_88_U236 ; P1_SUB_88_U41
g8132 nand P1_SUB_88_U241 P1_SUB_88_U240 ; P1_SUB_88_U42
g8133 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U43
g8134 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN ; P1_SUB_88_U44
g8135 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U45
g8136 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U46
g8137 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U47
g8138 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U48
g8139 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U49
g8140 nor P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U50
g8141 and P1_SUB_88_U50 P1_SUB_88_U49 P1_SUB_88_U48 P1_SUB_88_U47 ; P1_SUB_88_U51
g8142 nor P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U52
g8143 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_27__SCAN_IN P1_IR_REG_28__SCAN_IN P1_IR_REG_29__SCAN_IN ; P1_SUB_88_U53
g8144 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U54
g8145 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U55
g8146 and P1_SUB_88_U55 P1_SUB_88_U54 P1_SUB_88_U53 P1_SUB_88_U52 ; P1_SUB_88_U56
g8147 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U57
g8148 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U58
g8149 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U59
g8150 nor P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U60
g8151 and P1_SUB_88_U60 P1_SUB_88_U59 P1_SUB_88_U58 P1_SUB_88_U57 ; P1_SUB_88_U61
g8152 nor P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U62
g8153 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_27__SCAN_IN P1_IR_REG_28__SCAN_IN ; P1_SUB_88_U63
g8154 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U64
g8155 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U65
g8156 and P1_SUB_88_U65 P1_SUB_88_U64 P1_SUB_88_U63 P1_SUB_88_U62 ; P1_SUB_88_U66
g8157 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U67
g8158 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U68
g8159 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U69
g8160 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U70
g8161 and P1_SUB_88_U70 P1_SUB_88_U69 P1_SUB_88_U68 P1_SUB_88_U67 ; P1_SUB_88_U71
g8162 nor P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U72
g8163 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_26__SCAN_IN P1_IR_REG_27__SCAN_IN ; P1_SUB_88_U73
g8164 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U74
g8165 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U75
g8166 and P1_SUB_88_U75 P1_SUB_88_U74 P1_SUB_88_U73 P1_SUB_88_U72 ; P1_SUB_88_U76
g8167 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U77
g8168 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U78
g8169 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U79
g8170 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U80
g8171 and P1_SUB_88_U80 P1_SUB_88_U79 P1_SUB_88_U78 P1_SUB_88_U77 ; P1_SUB_88_U81
g8172 nor P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U82
g8173 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U83
g8174 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U84
g8175 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U85
g8176 and P1_SUB_88_U85 P1_SUB_88_U84 P1_SUB_88_U83 P1_SUB_88_U82 ; P1_SUB_88_U86
g8177 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U87
g8178 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U88
g8179 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U89
g8180 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U90
g8181 and P1_SUB_88_U90 P1_SUB_88_U89 P1_SUB_88_U88 P1_SUB_88_U87 ; P1_SUB_88_U91
g8182 nor P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U92
g8183 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U93
g8184 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U94
g8185 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U95
g8186 and P1_SUB_88_U95 P1_SUB_88_U94 P1_SUB_88_U93 P1_SUB_88_U92 ; P1_SUB_88_U96
g8187 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U97
g8188 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U98
g8189 nor P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U99
g8190 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U100
g8191 and P1_SUB_88_U100 P1_SUB_88_U99 P1_SUB_88_U98 P1_SUB_88_U97 ; P1_SUB_88_U101
g8192 nor P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN ; P1_SUB_88_U102
g8193 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U103
g8194 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U104
g8195 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U105
g8196 and P1_SUB_88_U105 P1_SUB_88_U104 P1_SUB_88_U103 P1_SUB_88_U102 ; P1_SUB_88_U106
g8197 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U107
g8198 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U108
g8199 nor P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U109
g8200 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U110
g8201 and P1_SUB_88_U110 P1_SUB_88_U109 P1_SUB_88_U108 P1_SUB_88_U107 ; P1_SUB_88_U111
g8202 nor P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN ; P1_SUB_88_U112
g8203 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_24__SCAN_IN ; P1_SUB_88_U113
g8204 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U114
g8205 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U115
g8206 and P1_SUB_88_U115 P1_SUB_88_U114 P1_SUB_88_U113 P1_SUB_88_U112 ; P1_SUB_88_U116
g8207 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U117
g8208 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U118
g8209 nor P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U119
g8210 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U120
g8211 and P1_SUB_88_U120 P1_SUB_88_U119 P1_SUB_88_U118 P1_SUB_88_U117 ; P1_SUB_88_U121
g8212 nor P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U122
g8213 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_23__SCAN_IN ; P1_SUB_88_U123
g8214 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U124
g8215 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U125
g8216 and P1_SUB_88_U125 P1_SUB_88_U124 P1_SUB_88_U123 P1_SUB_88_U122 ; P1_SUB_88_U126
g8217 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U127
g8218 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U128
g8219 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U129
g8220 nor P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U130
g8221 nor P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U131
g8222 nor P1_IR_REG_19__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U132
g8223 nor P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U133
g8224 and P1_SUB_88_U132 P1_SUB_88_U131 P1_SUB_88_U133 ; P1_SUB_88_U134
g8225 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U135
g8226 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U136
g8227 and P1_SUB_88_U136 P1_SUB_88_U135 ; P1_SUB_88_U137
g8228 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U138
g8229 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U139
g8230 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U140
g8231 and P1_SUB_88_U140 P1_SUB_88_U139 ; P1_SUB_88_U141
g8232 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U142
g8233 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U143
g8234 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U144
g8235 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U145
g8236 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U146
g8237 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U147
g8238 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U148
g8239 nor P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U149
g8240 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U150
g8241 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U151
g8242 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U152
g8243 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U153
g8244 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U154
g8245 nor P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U155
g8246 nor P1_IR_REG_9__SCAN_IN P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U156
g8247 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U157
g8248 nor P1_IR_REG_9__SCAN_IN P1_IR_REG_10__SCAN_IN ; P1_SUB_88_U158
g8249 not P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U159
g8250 and P1_SUB_88_U233 P1_SUB_88_U232 ; P1_SUB_88_U160
g8251 not P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U161
g8252 and P1_SUB_88_U235 P1_SUB_88_U234 ; P1_SUB_88_U162
g8253 not P1_IR_REG_31__SCAN_IN ; P1_SUB_88_U163
g8254 not P1_IR_REG_30__SCAN_IN ; P1_SUB_88_U164
g8255 and P1_SUB_88_U239 P1_SUB_88_U238 ; P1_SUB_88_U165
g8256 not P1_IR_REG_27__SCAN_IN ; P1_SUB_88_U166
g8257 nand P1_SUB_88_U96 P1_SUB_88_U91 ; P1_SUB_88_U167
g8258 not P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U168
g8259 nand P1_SUB_88_U116 P1_SUB_88_U111 ; P1_SUB_88_U169
g8260 and P1_SUB_88_U243 P1_SUB_88_U242 ; P1_SUB_88_U170
g8261 not P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U171
g8262 nand P1_SUB_88_U144 P1_SUB_88_U143 P1_SUB_88_U145 P1_SUB_88_U147 P1_SUB_88_U146 ; P1_SUB_88_U172
g8263 and P1_SUB_88_U245 P1_SUB_88_U244 ; P1_SUB_88_U173
g8264 not P1_IR_REG_1__SCAN_IN ; P1_SUB_88_U174
g8265 not P1_IR_REG_0__SCAN_IN ; P1_SUB_88_U175
g8266 not P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U176
g8267 and P1_SUB_88_U249 P1_SUB_88_U248 ; P1_SUB_88_U177
g8268 not P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U178
g8269 and P1_SUB_88_U251 P1_SUB_88_U250 ; P1_SUB_88_U179
g8270 nand P1_SUB_88_U230 P1_SUB_88_U32 ; P1_SUB_88_U180
g8271 not P1_SUB_88_U29 ; P1_SUB_88_U181
g8272 not P1_SUB_88_U30 ; P1_SUB_88_U182
g8273 nand P1_SUB_88_U182 P1_SUB_88_U31 ; P1_SUB_88_U183
g8274 not P1_SUB_88_U28 ; P1_SUB_88_U184
g8275 nand P1_SUB_88_U183 P1_IR_REG_8__SCAN_IN ; P1_SUB_88_U185
g8276 nand P1_SUB_88_U30 P1_IR_REG_7__SCAN_IN ; P1_SUB_88_U186
g8277 nand P1_SUB_88_U181 P1_SUB_88_U161 ; P1_SUB_88_U187
g8278 nand P1_SUB_88_U187 P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U188
g8279 nand P1_SUB_88_U180 P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U189
g8280 nand P1_SUB_88_U27 P1_IR_REG_3__SCAN_IN ; P1_SUB_88_U190
g8281 not P1_SUB_88_U38 ; P1_SUB_88_U191
g8282 nand P1_SUB_88_U191 P1_SUB_88_U39 ; P1_SUB_88_U192
g8283 not P1_SUB_88_U35 ; P1_SUB_88_U193
g8284 not P1_SUB_88_U36 ; P1_SUB_88_U194
g8285 nand P1_SUB_88_U194 P1_SUB_88_U37 ; P1_SUB_88_U195
g8286 not P1_SUB_88_U34 ; P1_SUB_88_U196
g8287 nand P1_SUB_88_U155 P1_SUB_88_U154 P1_SUB_88_U153 P1_SUB_88_U152 ; P1_SUB_88_U197
g8288 nand P1_SUB_88_U151 P1_SUB_88_U150 P1_SUB_88_U149 P1_SUB_88_U148 ; P1_SUB_88_U198
g8289 not P1_SUB_88_U172 ; P1_SUB_88_U199
g8290 nand P1_SUB_88_U134 P1_SUB_88_U196 ; P1_SUB_88_U200
g8291 nand P1_SUB_88_U126 P1_SUB_88_U121 ; P1_SUB_88_U201
g8292 not P1_SUB_88_U169 ; P1_SUB_88_U202
g8293 not P1_SUB_88_U167 ; P1_SUB_88_U203
g8294 nand P1_SUB_88_U66 P1_SUB_88_U61 ; P1_SUB_88_U204
g8295 not P1_SUB_88_U33 ; P1_SUB_88_U205
g8296 or P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN ; P1_SUB_88_U206
g8297 nand P1_SUB_88_U206 P1_IR_REG_2__SCAN_IN ; P1_SUB_88_U207
g8298 nand P1_SUB_88_U204 P1_IR_REG_29__SCAN_IN ; P1_SUB_88_U208
g8299 nand P1_SUB_88_U229 P1_IR_REG_28__SCAN_IN ; P1_SUB_88_U209
g8300 nand P1_SUB_88_U106 P1_SUB_88_U101 ; P1_SUB_88_U210
g8301 nand P1_SUB_88_U210 P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U211
g8302 nand P1_SUB_88_U201 P1_IR_REG_24__SCAN_IN ; P1_SUB_88_U212
g8303 nand P1_SUB_88_U200 P1_IR_REG_23__SCAN_IN ; P1_SUB_88_U213
g8304 nand P1_SUB_88_U142 P1_SUB_88_U141 P1_SUB_88_U138 P1_SUB_88_U137 ; P1_SUB_88_U214
g8305 nand P1_SUB_88_U214 P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U215
g8306 nand P1_SUB_88_U198 P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U216
g8307 nand P1_SUB_88_U197 P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U217
g8308 nand P1_SUB_88_U196 P1_SUB_88_U176 ; P1_SUB_88_U218
g8309 nand P1_SUB_88_U218 P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U219
g8310 nand P1_SUB_88_U195 P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U220
g8311 nand P1_SUB_88_U36 P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U221
g8312 nand P1_SUB_88_U193 P1_SUB_88_U178 ; P1_SUB_88_U222
g8313 nand P1_SUB_88_U222 P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U223
g8314 nand P1_SUB_88_U192 P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U224
g8315 nand P1_SUB_88_U38 P1_IR_REG_11__SCAN_IN ; P1_SUB_88_U225
g8316 nand P1_SUB_88_U184 P1_SUB_88_U159 ; P1_SUB_88_U226
g8317 nand P1_SUB_88_U226 P1_IR_REG_10__SCAN_IN ; P1_SUB_88_U227
g8318 nand P1_SUB_88_U205 P1_SUB_88_U164 ; P1_SUB_88_U228
g8319 nand P1_SUB_88_U76 P1_SUB_88_U71 ; P1_SUB_88_U229
g8320 not P1_SUB_88_U27 ; P1_SUB_88_U230
g8321 nand P1_SUB_88_U86 P1_SUB_88_U81 ; P1_SUB_88_U231
g8322 nand P1_SUB_88_U28 P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U232
g8323 nand P1_SUB_88_U184 P1_SUB_88_U159 ; P1_SUB_88_U233
g8324 nand P1_SUB_88_U29 P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U234
g8325 nand P1_SUB_88_U181 P1_SUB_88_U161 ; P1_SUB_88_U235
g8326 nand P1_SUB_88_U228 P1_SUB_88_U163 ; P1_SUB_88_U236
g8327 nand P1_SUB_88_U205 P1_SUB_88_U164 P1_IR_REG_31__SCAN_IN ; P1_SUB_88_U237
g8328 nand P1_SUB_88_U33 P1_IR_REG_30__SCAN_IN ; P1_SUB_88_U238
g8329 nand P1_SUB_88_U205 P1_SUB_88_U164 ; P1_SUB_88_U239
g8330 nand P1_SUB_88_U203 P1_IR_REG_27__SCAN_IN ; P1_SUB_88_U240
g8331 nand P1_SUB_88_U231 P1_SUB_88_U166 ; P1_SUB_88_U241
g8332 nand P1_SUB_88_U169 P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U242
g8333 nand P1_SUB_88_U202 P1_SUB_88_U168 ; P1_SUB_88_U243
g8334 nand P1_SUB_88_U172 P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U244
g8335 nand P1_SUB_88_U199 P1_SUB_88_U171 ; P1_SUB_88_U245
g8336 nand P1_SUB_88_U175 P1_IR_REG_1__SCAN_IN ; P1_SUB_88_U246
g8337 nand P1_SUB_88_U174 P1_IR_REG_0__SCAN_IN ; P1_SUB_88_U247
g8338 nand P1_SUB_88_U34 P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U248
g8339 nand P1_SUB_88_U196 P1_SUB_88_U176 ; P1_SUB_88_U249
g8340 nand P1_SUB_88_U35 P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U250
g8341 nand P1_SUB_88_U193 P1_SUB_88_U178 ; P1_SUB_88_U251
g8342 not P1_U3057 ; P1_R1309_U6
g8343 not P1_U3054 ; P1_R1309_U7
g8344 and P1_R1309_U10 P1_R1309_U9 ; P1_R1309_U8
g8345 nand P1_U3054 P1_R1309_U6 ; P1_R1309_U9
g8346 nand P1_U3057 P1_R1309_U7 ; P1_R1309_U10
g8347 and P1_R1282_U135 P1_R1282_U35 ; P1_R1282_U6
g8348 and P1_R1282_U133 P1_R1282_U36 ; P1_R1282_U7
g8349 and P1_R1282_U132 P1_R1282_U37 ; P1_R1282_U8
g8350 and P1_R1282_U131 P1_R1282_U38 ; P1_R1282_U9
g8351 and P1_R1282_U129 P1_R1282_U39 ; P1_R1282_U10
g8352 and P1_R1282_U128 P1_R1282_U40 ; P1_R1282_U11
g8353 and P1_R1282_U127 P1_R1282_U41 ; P1_R1282_U12
g8354 and P1_R1282_U125 P1_R1282_U42 ; P1_R1282_U13
g8355 and P1_R1282_U123 P1_R1282_U43 ; P1_R1282_U14
g8356 and P1_R1282_U121 P1_R1282_U44 ; P1_R1282_U15
g8357 and P1_R1282_U119 P1_R1282_U45 ; P1_R1282_U16
g8358 and P1_R1282_U117 P1_R1282_U46 ; P1_R1282_U17
g8359 and P1_R1282_U115 P1_R1282_U25 ; P1_R1282_U18
g8360 and P1_R1282_U113 P1_R1282_U67 ; P1_R1282_U19
g8361 and P1_R1282_U98 P1_R1282_U26 ; P1_R1282_U20
g8362 and P1_R1282_U97 P1_R1282_U27 ; P1_R1282_U21
g8363 and P1_R1282_U96 P1_R1282_U28 ; P1_R1282_U22
g8364 and P1_R1282_U94 P1_R1282_U29 ; P1_R1282_U23
g8365 and P1_R1282_U93 P1_R1282_U30 ; P1_R1282_U24
g8366 or P1_U3456 P1_U3451 P1_U3459 ; P1_R1282_U25
g8367 nand P1_R1282_U87 P1_R1282_U34 ; P1_R1282_U26
g8368 nand P1_R1282_U88 P1_R1282_U33 ; P1_R1282_U27
g8369 nand P1_R1282_U58 P1_R1282_U89 ; P1_R1282_U28
g8370 nand P1_R1282_U90 P1_R1282_U32 ; P1_R1282_U29
g8371 nand P1_R1282_U91 P1_R1282_U31 ; P1_R1282_U30
g8372 not P1_U3477 ; P1_R1282_U31
g8373 not P1_U3474 ; P1_R1282_U32
g8374 not P1_U3465 ; P1_R1282_U33
g8375 not P1_U3462 ; P1_R1282_U34
g8376 nand P1_R1282_U59 P1_R1282_U92 ; P1_R1282_U35
g8377 nand P1_R1282_U99 P1_R1282_U56 ; P1_R1282_U36
g8378 nand P1_R1282_U100 P1_R1282_U55 ; P1_R1282_U37
g8379 nand P1_R1282_U60 P1_R1282_U101 ; P1_R1282_U38
g8380 nand P1_R1282_U102 P1_R1282_U54 ; P1_R1282_U39
g8381 nand P1_R1282_U103 P1_R1282_U53 ; P1_R1282_U40
g8382 nand P1_R1282_U61 P1_R1282_U104 ; P1_R1282_U41
g8383 nand P1_R1282_U105 P1_R1282_U81 P1_R1282_U52 ; P1_R1282_U42
g8384 nand P1_R1282_U106 P1_R1282_U77 P1_R1282_U51 ; P1_R1282_U43
g8385 nand P1_R1282_U107 P1_R1282_U75 P1_R1282_U50 ; P1_R1282_U44
g8386 nand P1_R1282_U108 P1_R1282_U73 P1_R1282_U49 ; P1_R1282_U45
g8387 nand P1_R1282_U109 P1_R1282_U71 P1_R1282_U48 ; P1_R1282_U46
g8388 not P1_U4017 ; P1_R1282_U47
g8389 not P1_U4007 ; P1_R1282_U48
g8390 not P1_U4009 ; P1_R1282_U49
g8391 not P1_U4011 ; P1_R1282_U50
g8392 not P1_U4013 ; P1_R1282_U51
g8393 not P1_U4015 ; P1_R1282_U52
g8394 not P1_U3501 ; P1_R1282_U53
g8395 not P1_U3498 ; P1_R1282_U54
g8396 not P1_U3489 ; P1_R1282_U55
g8397 not P1_U3486 ; P1_R1282_U56
g8398 nand P1_R1282_U153 P1_R1282_U152 ; P1_R1282_U57
g8399 nor P1_U3468 P1_U3471 ; P1_R1282_U58
g8400 nor P1_U3483 P1_U3480 ; P1_R1282_U59
g8401 nor P1_U3492 P1_U3495 ; P1_R1282_U60
g8402 nor P1_U3504 P1_U3507 ; P1_R1282_U61
g8403 not P1_U3480 ; P1_R1282_U62
g8404 and P1_R1282_U137 P1_R1282_U136 ; P1_R1282_U63
g8405 not P1_U3468 ; P1_R1282_U64
g8406 and P1_R1282_U139 P1_R1282_U138 ; P1_R1282_U65
g8407 not P1_U4016 ; P1_R1282_U66
g8408 nand P1_R1282_U110 P1_R1282_U69 P1_R1282_U47 ; P1_R1282_U67
g8409 and P1_R1282_U141 P1_R1282_U140 ; P1_R1282_U68
g8410 not P1_U4018 ; P1_R1282_U69
g8411 and P1_R1282_U143 P1_R1282_U142 ; P1_R1282_U70
g8412 not P1_U4008 ; P1_R1282_U71
g8413 and P1_R1282_U145 P1_R1282_U144 ; P1_R1282_U72
g8414 not P1_U4010 ; P1_R1282_U73
g8415 and P1_R1282_U147 P1_R1282_U146 ; P1_R1282_U74
g8416 not P1_U4012 ; P1_R1282_U75
g8417 and P1_R1282_U149 P1_R1282_U148 ; P1_R1282_U76
g8418 not P1_U4014 ; P1_R1282_U77
g8419 and P1_R1282_U151 P1_R1282_U150 ; P1_R1282_U78
g8420 not P1_U3456 ; P1_R1282_U79
g8421 not P1_U3451 ; P1_R1282_U80
g8422 not P1_U3509 ; P1_R1282_U81
g8423 and P1_R1282_U155 P1_R1282_U154 ; P1_R1282_U82
g8424 not P1_U3504 ; P1_R1282_U83
g8425 and P1_R1282_U157 P1_R1282_U156 ; P1_R1282_U84
g8426 not P1_U3492 ; P1_R1282_U85
g8427 and P1_R1282_U159 P1_R1282_U158 ; P1_R1282_U86
g8428 not P1_R1282_U25 ; P1_R1282_U87
g8429 not P1_R1282_U26 ; P1_R1282_U88
g8430 not P1_R1282_U27 ; P1_R1282_U89
g8431 not P1_R1282_U28 ; P1_R1282_U90
g8432 not P1_R1282_U29 ; P1_R1282_U91
g8433 not P1_R1282_U30 ; P1_R1282_U92
g8434 nand P1_U3477 P1_R1282_U29 ; P1_R1282_U93
g8435 nand P1_U3474 P1_R1282_U28 ; P1_R1282_U94
g8436 nand P1_R1282_U89 P1_R1282_U64 ; P1_R1282_U95
g8437 nand P1_U3471 P1_R1282_U95 ; P1_R1282_U96
g8438 nand P1_U3465 P1_R1282_U26 ; P1_R1282_U97
g8439 nand P1_U3462 P1_R1282_U25 ; P1_R1282_U98
g8440 not P1_R1282_U35 ; P1_R1282_U99
g8441 not P1_R1282_U36 ; P1_R1282_U100
g8442 not P1_R1282_U37 ; P1_R1282_U101
g8443 not P1_R1282_U38 ; P1_R1282_U102
g8444 not P1_R1282_U39 ; P1_R1282_U103
g8445 not P1_R1282_U40 ; P1_R1282_U104
g8446 not P1_R1282_U41 ; P1_R1282_U105
g8447 not P1_R1282_U42 ; P1_R1282_U106
g8448 not P1_R1282_U43 ; P1_R1282_U107
g8449 not P1_R1282_U44 ; P1_R1282_U108
g8450 not P1_R1282_U45 ; P1_R1282_U109
g8451 not P1_R1282_U46 ; P1_R1282_U110
g8452 not P1_R1282_U67 ; P1_R1282_U111
g8453 nand P1_R1282_U110 P1_R1282_U69 ; P1_R1282_U112
g8454 nand P1_U4017 P1_R1282_U112 ; P1_R1282_U113
g8455 or P1_U3456 P1_U3451 ; P1_R1282_U114
g8456 nand P1_U3459 P1_R1282_U114 ; P1_R1282_U115
g8457 nand P1_R1282_U109 P1_R1282_U71 ; P1_R1282_U116
g8458 nand P1_U4007 P1_R1282_U116 ; P1_R1282_U117
g8459 nand P1_R1282_U108 P1_R1282_U73 ; P1_R1282_U118
g8460 nand P1_U4009 P1_R1282_U118 ; P1_R1282_U119
g8461 nand P1_R1282_U107 P1_R1282_U75 ; P1_R1282_U120
g8462 nand P1_U4011 P1_R1282_U120 ; P1_R1282_U121
g8463 nand P1_R1282_U106 P1_R1282_U77 ; P1_R1282_U122
g8464 nand P1_U4013 P1_R1282_U122 ; P1_R1282_U123
g8465 nand P1_R1282_U105 P1_R1282_U81 ; P1_R1282_U124
g8466 nand P1_U4015 P1_R1282_U124 ; P1_R1282_U125
g8467 nand P1_R1282_U104 P1_R1282_U83 ; P1_R1282_U126
g8468 nand P1_U3507 P1_R1282_U126 ; P1_R1282_U127
g8469 nand P1_U3501 P1_R1282_U39 ; P1_R1282_U128
g8470 nand P1_U3498 P1_R1282_U38 ; P1_R1282_U129
g8471 nand P1_R1282_U101 P1_R1282_U85 ; P1_R1282_U130
g8472 nand P1_U3495 P1_R1282_U130 ; P1_R1282_U131
g8473 nand P1_U3489 P1_R1282_U36 ; P1_R1282_U132
g8474 nand P1_U3486 P1_R1282_U35 ; P1_R1282_U133
g8475 nand P1_R1282_U92 P1_R1282_U62 ; P1_R1282_U134
g8476 nand P1_U3483 P1_R1282_U134 ; P1_R1282_U135
g8477 nand P1_U3480 P1_R1282_U30 ; P1_R1282_U136
g8478 nand P1_R1282_U92 P1_R1282_U62 ; P1_R1282_U137
g8479 nand P1_U3468 P1_R1282_U27 ; P1_R1282_U138
g8480 nand P1_R1282_U89 P1_R1282_U64 ; P1_R1282_U139
g8481 nand P1_U4016 P1_R1282_U67 ; P1_R1282_U140
g8482 nand P1_R1282_U111 P1_R1282_U66 ; P1_R1282_U141
g8483 nand P1_U4018 P1_R1282_U46 ; P1_R1282_U142
g8484 nand P1_R1282_U110 P1_R1282_U69 ; P1_R1282_U143
g8485 nand P1_U4008 P1_R1282_U45 ; P1_R1282_U144
g8486 nand P1_R1282_U109 P1_R1282_U71 ; P1_R1282_U145
g8487 nand P1_U4010 P1_R1282_U44 ; P1_R1282_U146
g8488 nand P1_R1282_U108 P1_R1282_U73 ; P1_R1282_U147
g8489 nand P1_U4012 P1_R1282_U43 ; P1_R1282_U148
g8490 nand P1_R1282_U107 P1_R1282_U75 ; P1_R1282_U149
g8491 nand P1_U4014 P1_R1282_U42 ; P1_R1282_U150
g8492 nand P1_R1282_U106 P1_R1282_U77 ; P1_R1282_U151
g8493 nand P1_U3456 P1_R1282_U80 ; P1_R1282_U152
g8494 nand P1_U3451 P1_R1282_U79 ; P1_R1282_U153
g8495 nand P1_U3509 P1_R1282_U41 ; P1_R1282_U154
g8496 nand P1_R1282_U105 P1_R1282_U81 ; P1_R1282_U155
g8497 nand P1_U3504 P1_R1282_U40 ; P1_R1282_U156
g8498 nand P1_R1282_U104 P1_R1282_U83 ; P1_R1282_U157
g8499 nand P1_U3492 P1_R1282_U37 ; P1_R1282_U158
g8500 nand P1_R1282_U101 P1_R1282_U85 ; P1_R1282_U159
g8501 and P1_R1240_U176 P1_R1240_U175 ; P1_R1240_U4
g8502 and P1_R1240_U177 P1_R1240_U178 ; P1_R1240_U5
g8503 and P1_R1240_U194 P1_R1240_U193 ; P1_R1240_U6
g8504 and P1_R1240_U234 P1_R1240_U233 ; P1_R1240_U7
g8505 and P1_R1240_U243 P1_R1240_U242 ; P1_R1240_U8
g8506 and P1_R1240_U261 P1_R1240_U260 ; P1_R1240_U9
g8507 and P1_R1240_U269 P1_R1240_U268 ; P1_R1240_U10
g8508 and P1_R1240_U348 P1_R1240_U345 ; P1_R1240_U11
g8509 and P1_R1240_U341 P1_R1240_U338 ; P1_R1240_U12
g8510 and P1_R1240_U332 P1_R1240_U329 ; P1_R1240_U13
g8511 and P1_R1240_U323 P1_R1240_U320 ; P1_R1240_U14
g8512 and P1_R1240_U317 P1_R1240_U315 ; P1_R1240_U15
g8513 and P1_R1240_U310 P1_R1240_U307 ; P1_R1240_U16
g8514 and P1_R1240_U232 P1_R1240_U229 ; P1_R1240_U17
g8515 and P1_R1240_U224 P1_R1240_U221 ; P1_R1240_U18
g8516 and P1_R1240_U210 P1_R1240_U207 ; P1_R1240_U19
g8517 not P1_U3471 ; P1_R1240_U20
g8518 not P1_U3069 ; P1_R1240_U21
g8519 not P1_U3068 ; P1_R1240_U22
g8520 nand P1_U3069 P1_U3471 ; P1_R1240_U23
g8521 not P1_U3474 ; P1_R1240_U24
g8522 not P1_U3465 ; P1_R1240_U25
g8523 not P1_U3058 ; P1_R1240_U26
g8524 not P1_U3065 ; P1_R1240_U27
g8525 not P1_U3459 ; P1_R1240_U28
g8526 not P1_U3066 ; P1_R1240_U29
g8527 not P1_U3451 ; P1_R1240_U30
g8528 not P1_U3075 ; P1_R1240_U31
g8529 nand P1_U3075 P1_U3451 ; P1_R1240_U32
g8530 not P1_U3462 ; P1_R1240_U33
g8531 not P1_U3062 ; P1_R1240_U34
g8532 nand P1_U3058 P1_U3465 ; P1_R1240_U35
g8533 not P1_U3468 ; P1_R1240_U36
g8534 not P1_U3477 ; P1_R1240_U37
g8535 not P1_U3082 ; P1_R1240_U38
g8536 not P1_U3081 ; P1_R1240_U39
g8537 not P1_U3480 ; P1_R1240_U40
g8538 nand P1_R1240_U62 P1_R1240_U202 ; P1_R1240_U41
g8539 nand P1_R1240_U118 P1_R1240_U190 ; P1_R1240_U42
g8540 nand P1_R1240_U179 P1_R1240_U180 ; P1_R1240_U43
g8541 nand P1_U3456 P1_U3076 ; P1_R1240_U44
g8542 nand P1_R1240_U122 P1_R1240_U216 ; P1_R1240_U45
g8543 nand P1_R1240_U213 P1_R1240_U212 ; P1_R1240_U46
g8544 not P1_U4008 ; P1_R1240_U47
g8545 not P1_U3051 ; P1_R1240_U48
g8546 not P1_U3055 ; P1_R1240_U49
g8547 not P1_U4009 ; P1_R1240_U50
g8548 not P1_U4010 ; P1_R1240_U51
g8549 not P1_U3056 ; P1_R1240_U52
g8550 not P1_U4011 ; P1_R1240_U53
g8551 not P1_U3063 ; P1_R1240_U54
g8552 not P1_U4014 ; P1_R1240_U55
g8553 not P1_U3073 ; P1_R1240_U56
g8554 not P1_U3501 ; P1_R1240_U57
g8555 not P1_U3071 ; P1_R1240_U58
g8556 not P1_U3067 ; P1_R1240_U59
g8557 nand P1_U3071 P1_U3501 ; P1_R1240_U60
g8558 not P1_U3504 ; P1_R1240_U61
g8559 nand P1_U3082 P1_U3477 ; P1_R1240_U62
g8560 not P1_U3483 ; P1_R1240_U63
g8561 not P1_U3060 ; P1_R1240_U64
g8562 not P1_U3489 ; P1_R1240_U65
g8563 not P1_U3070 ; P1_R1240_U66
g8564 not P1_U3486 ; P1_R1240_U67
g8565 not P1_U3061 ; P1_R1240_U68
g8566 nand P1_U3061 P1_U3486 ; P1_R1240_U69
g8567 not P1_U3492 ; P1_R1240_U70
g8568 not P1_U3078 ; P1_R1240_U71
g8569 not P1_U3495 ; P1_R1240_U72
g8570 not P1_U3077 ; P1_R1240_U73
g8571 not P1_U3498 ; P1_R1240_U74
g8572 not P1_U3072 ; P1_R1240_U75
g8573 not P1_U3507 ; P1_R1240_U76
g8574 not P1_U3080 ; P1_R1240_U77
g8575 nand P1_U3080 P1_U3507 ; P1_R1240_U78
g8576 not P1_U3509 ; P1_R1240_U79
g8577 not P1_U3079 ; P1_R1240_U80
g8578 nand P1_U3079 P1_U3509 ; P1_R1240_U81
g8579 not P1_U4015 ; P1_R1240_U82
g8580 not P1_U4013 ; P1_R1240_U83
g8581 not P1_U3059 ; P1_R1240_U84
g8582 not P1_U4012 ; P1_R1240_U85
g8583 not P1_U3064 ; P1_R1240_U86
g8584 nand P1_U4009 P1_U3055 ; P1_R1240_U87
g8585 not P1_U3052 ; P1_R1240_U88
g8586 not P1_U4007 ; P1_R1240_U89
g8587 nand P1_R1240_U303 P1_R1240_U173 ; P1_R1240_U90
g8588 not P1_U3074 ; P1_R1240_U91
g8589 nand P1_R1240_U78 P1_R1240_U312 ; P1_R1240_U92
g8590 nand P1_R1240_U258 P1_R1240_U257 ; P1_R1240_U93
g8591 nand P1_R1240_U69 P1_R1240_U334 ; P1_R1240_U94
g8592 nand P1_R1240_U454 P1_R1240_U453 ; P1_R1240_U95
g8593 nand P1_R1240_U501 P1_R1240_U500 ; P1_R1240_U96
g8594 nand P1_R1240_U372 P1_R1240_U371 ; P1_R1240_U97
g8595 nand P1_R1240_U377 P1_R1240_U376 ; P1_R1240_U98
g8596 nand P1_R1240_U384 P1_R1240_U383 ; P1_R1240_U99
g8597 nand P1_R1240_U391 P1_R1240_U390 ; P1_R1240_U100
g8598 nand P1_R1240_U396 P1_R1240_U395 ; P1_R1240_U101
g8599 nand P1_R1240_U405 P1_R1240_U404 ; P1_R1240_U102
g8600 nand P1_R1240_U412 P1_R1240_U411 ; P1_R1240_U103
g8601 nand P1_R1240_U419 P1_R1240_U418 ; P1_R1240_U104
g8602 nand P1_R1240_U426 P1_R1240_U425 ; P1_R1240_U105
g8603 nand P1_R1240_U431 P1_R1240_U430 ; P1_R1240_U106
g8604 nand P1_R1240_U438 P1_R1240_U437 ; P1_R1240_U107
g8605 nand P1_R1240_U445 P1_R1240_U444 ; P1_R1240_U108
g8606 nand P1_R1240_U459 P1_R1240_U458 ; P1_R1240_U109
g8607 nand P1_R1240_U464 P1_R1240_U463 ; P1_R1240_U110
g8608 nand P1_R1240_U471 P1_R1240_U470 ; P1_R1240_U111
g8609 nand P1_R1240_U478 P1_R1240_U477 ; P1_R1240_U112
g8610 nand P1_R1240_U485 P1_R1240_U484 ; P1_R1240_U113
g8611 nand P1_R1240_U492 P1_R1240_U491 ; P1_R1240_U114
g8612 nand P1_R1240_U497 P1_R1240_U496 ; P1_R1240_U115
g8613 and P1_U3459 P1_U3066 ; P1_R1240_U116
g8614 and P1_R1240_U186 P1_R1240_U184 ; P1_R1240_U117
g8615 and P1_R1240_U191 P1_R1240_U189 ; P1_R1240_U118
g8616 and P1_R1240_U198 P1_R1240_U197 ; P1_R1240_U119
g8617 and P1_R1240_U379 P1_R1240_U378 P1_R1240_U23 ; P1_R1240_U120
g8618 and P1_R1240_U209 P1_R1240_U6 ; P1_R1240_U121
g8619 and P1_R1240_U217 P1_R1240_U215 ; P1_R1240_U122
g8620 and P1_R1240_U386 P1_R1240_U385 P1_R1240_U35 ; P1_R1240_U123
g8621 and P1_R1240_U223 P1_R1240_U4 ; P1_R1240_U124
g8622 and P1_R1240_U231 P1_R1240_U178 ; P1_R1240_U125
g8623 and P1_R1240_U201 P1_R1240_U7 ; P1_R1240_U126
g8624 and P1_R1240_U236 P1_R1240_U168 ; P1_R1240_U127
g8625 and P1_R1240_U245 P1_R1240_U169 ; P1_R1240_U128
g8626 and P1_R1240_U265 P1_R1240_U264 ; P1_R1240_U129
g8627 and P1_R1240_U10 P1_R1240_U279 ; P1_R1240_U130
g8628 and P1_R1240_U282 P1_R1240_U277 ; P1_R1240_U131
g8629 and P1_R1240_U298 P1_R1240_U295 ; P1_R1240_U132
g8630 and P1_R1240_U365 P1_R1240_U299 ; P1_R1240_U133
g8631 and P1_R1240_U156 P1_R1240_U275 ; P1_R1240_U134
g8632 and P1_R1240_U466 P1_R1240_U465 P1_R1240_U60 ; P1_R1240_U135
g8633 and P1_R1240_U487 P1_R1240_U486 P1_R1240_U169 ; P1_R1240_U136
g8634 and P1_R1240_U340 P1_R1240_U8 ; P1_R1240_U137
g8635 and P1_R1240_U499 P1_R1240_U498 P1_R1240_U168 ; P1_R1240_U138
g8636 and P1_R1240_U347 P1_R1240_U7 ; P1_R1240_U139
g8637 nand P1_R1240_U119 P1_R1240_U199 ; P1_R1240_U140
g8638 nand P1_R1240_U214 P1_R1240_U226 ; P1_R1240_U141
g8639 not P1_U3053 ; P1_R1240_U142
g8640 not P1_U4018 ; P1_R1240_U143
g8641 and P1_R1240_U400 P1_R1240_U399 ; P1_R1240_U144
g8642 nand P1_R1240_U301 P1_R1240_U166 P1_R1240_U361 ; P1_R1240_U145
g8643 and P1_R1240_U407 P1_R1240_U406 ; P1_R1240_U146
g8644 nand P1_R1240_U367 P1_R1240_U366 P1_R1240_U133 ; P1_R1240_U147
g8645 and P1_R1240_U414 P1_R1240_U413 ; P1_R1240_U148
g8646 nand P1_R1240_U362 P1_R1240_U296 P1_R1240_U87 ; P1_R1240_U149
g8647 and P1_R1240_U421 P1_R1240_U420 ; P1_R1240_U150
g8648 nand P1_R1240_U290 P1_R1240_U289 ; P1_R1240_U151
g8649 and P1_R1240_U433 P1_R1240_U432 ; P1_R1240_U152
g8650 nand P1_R1240_U286 P1_R1240_U285 ; P1_R1240_U153
g8651 and P1_R1240_U440 P1_R1240_U439 ; P1_R1240_U154
g8652 nand P1_R1240_U131 P1_R1240_U281 ; P1_R1240_U155
g8653 and P1_R1240_U447 P1_R1240_U446 ; P1_R1240_U156
g8654 and P1_R1240_U452 P1_R1240_U451 ; P1_R1240_U157
g8655 nand P1_R1240_U44 P1_R1240_U324 ; P1_R1240_U158
g8656 nand P1_R1240_U129 P1_R1240_U266 ; P1_R1240_U159
g8657 and P1_R1240_U473 P1_R1240_U472 ; P1_R1240_U160
g8658 nand P1_R1240_U254 P1_R1240_U253 ; P1_R1240_U161
g8659 and P1_R1240_U480 P1_R1240_U479 ; P1_R1240_U162
g8660 nand P1_R1240_U250 P1_R1240_U249 ; P1_R1240_U163
g8661 nand P1_R1240_U240 P1_R1240_U239 ; P1_R1240_U164
g8662 nand P1_R1240_U364 P1_R1240_U363 ; P1_R1240_U165
g8663 nand P1_U3052 P1_R1240_U147 ; P1_R1240_U166
g8664 not P1_R1240_U35 ; P1_R1240_U167
g8665 nand P1_U3480 P1_U3081 ; P1_R1240_U168
g8666 nand P1_U3070 P1_U3489 ; P1_R1240_U169
g8667 nand P1_U3056 P1_U4010 ; P1_R1240_U170
g8668 not P1_R1240_U69 ; P1_R1240_U171
g8669 not P1_R1240_U78 ; P1_R1240_U172
g8670 nand P1_U3063 P1_U4011 ; P1_R1240_U173
g8671 not P1_R1240_U62 ; P1_R1240_U174
g8672 or P1_U3065 P1_U3468 ; P1_R1240_U175
g8673 or P1_U3058 P1_U3465 ; P1_R1240_U176
g8674 or P1_U3462 P1_U3062 ; P1_R1240_U177
g8675 or P1_U3459 P1_U3066 ; P1_R1240_U178
g8676 not P1_R1240_U32 ; P1_R1240_U179
g8677 or P1_U3456 P1_U3076 ; P1_R1240_U180
g8678 not P1_R1240_U43 ; P1_R1240_U181
g8679 not P1_R1240_U44 ; P1_R1240_U182
g8680 nand P1_R1240_U43 P1_R1240_U44 ; P1_R1240_U183
g8681 nand P1_R1240_U116 P1_R1240_U177 ; P1_R1240_U184
g8682 nand P1_R1240_U5 P1_R1240_U183 ; P1_R1240_U185
g8683 nand P1_U3062 P1_U3462 ; P1_R1240_U186
g8684 nand P1_R1240_U117 P1_R1240_U185 ; P1_R1240_U187
g8685 nand P1_R1240_U36 P1_R1240_U35 ; P1_R1240_U188
g8686 nand P1_U3065 P1_R1240_U188 ; P1_R1240_U189
g8687 nand P1_R1240_U4 P1_R1240_U187 ; P1_R1240_U190
g8688 nand P1_U3468 P1_R1240_U167 ; P1_R1240_U191
g8689 not P1_R1240_U42 ; P1_R1240_U192
g8690 or P1_U3068 P1_U3474 ; P1_R1240_U193
g8691 or P1_U3069 P1_U3471 ; P1_R1240_U194
g8692 not P1_R1240_U23 ; P1_R1240_U195
g8693 nand P1_R1240_U24 P1_R1240_U23 ; P1_R1240_U196
g8694 nand P1_U3068 P1_R1240_U196 ; P1_R1240_U197
g8695 nand P1_U3474 P1_R1240_U195 ; P1_R1240_U198
g8696 nand P1_R1240_U6 P1_R1240_U42 ; P1_R1240_U199
g8697 not P1_R1240_U140 ; P1_R1240_U200
g8698 or P1_U3477 P1_U3082 ; P1_R1240_U201
g8699 nand P1_R1240_U201 P1_R1240_U140 ; P1_R1240_U202
g8700 not P1_R1240_U41 ; P1_R1240_U203
g8701 or P1_U3081 P1_U3480 ; P1_R1240_U204
g8702 or P1_U3471 P1_U3069 ; P1_R1240_U205
g8703 nand P1_R1240_U205 P1_R1240_U42 ; P1_R1240_U206
g8704 nand P1_R1240_U120 P1_R1240_U206 ; P1_R1240_U207
g8705 nand P1_R1240_U192 P1_R1240_U23 ; P1_R1240_U208
g8706 nand P1_U3474 P1_U3068 ; P1_R1240_U209
g8707 nand P1_R1240_U121 P1_R1240_U208 ; P1_R1240_U210
g8708 or P1_U3069 P1_U3471 ; P1_R1240_U211
g8709 nand P1_R1240_U182 P1_R1240_U178 ; P1_R1240_U212
g8710 nand P1_U3066 P1_U3459 ; P1_R1240_U213
g8711 not P1_R1240_U46 ; P1_R1240_U214
g8712 nand P1_R1240_U181 P1_R1240_U5 ; P1_R1240_U215
g8713 nand P1_R1240_U46 P1_R1240_U177 ; P1_R1240_U216
g8714 nand P1_U3062 P1_U3462 ; P1_R1240_U217
g8715 not P1_R1240_U45 ; P1_R1240_U218
g8716 or P1_U3465 P1_U3058 ; P1_R1240_U219
g8717 nand P1_R1240_U219 P1_R1240_U45 ; P1_R1240_U220
g8718 nand P1_R1240_U123 P1_R1240_U220 ; P1_R1240_U221
g8719 nand P1_R1240_U218 P1_R1240_U35 ; P1_R1240_U222
g8720 nand P1_U3468 P1_U3065 ; P1_R1240_U223
g8721 nand P1_R1240_U124 P1_R1240_U222 ; P1_R1240_U224
g8722 or P1_U3058 P1_U3465 ; P1_R1240_U225
g8723 nand P1_R1240_U181 P1_R1240_U178 ; P1_R1240_U226
g8724 not P1_R1240_U141 ; P1_R1240_U227
g8725 nand P1_U3062 P1_U3462 ; P1_R1240_U228
g8726 nand P1_R1240_U398 P1_R1240_U397 P1_R1240_U44 P1_R1240_U43 ; P1_R1240_U229
g8727 nand P1_R1240_U44 P1_R1240_U43 ; P1_R1240_U230
g8728 nand P1_U3066 P1_U3459 ; P1_R1240_U231
g8729 nand P1_R1240_U125 P1_R1240_U230 ; P1_R1240_U232
g8730 or P1_U3081 P1_U3480 ; P1_R1240_U233
g8731 or P1_U3060 P1_U3483 ; P1_R1240_U234
g8732 nand P1_R1240_U174 P1_R1240_U7 ; P1_R1240_U235
g8733 nand P1_U3060 P1_U3483 ; P1_R1240_U236
g8734 nand P1_R1240_U127 P1_R1240_U235 ; P1_R1240_U237
g8735 or P1_U3483 P1_U3060 ; P1_R1240_U238
g8736 nand P1_R1240_U126 P1_R1240_U140 ; P1_R1240_U239
g8737 nand P1_R1240_U238 P1_R1240_U237 ; P1_R1240_U240
g8738 not P1_R1240_U164 ; P1_R1240_U241
g8739 or P1_U3078 P1_U3492 ; P1_R1240_U242
g8740 or P1_U3070 P1_U3489 ; P1_R1240_U243
g8741 nand P1_R1240_U171 P1_R1240_U8 ; P1_R1240_U244
g8742 nand P1_U3078 P1_U3492 ; P1_R1240_U245
g8743 nand P1_R1240_U128 P1_R1240_U244 ; P1_R1240_U246
g8744 or P1_U3486 P1_U3061 ; P1_R1240_U247
g8745 or P1_U3492 P1_U3078 ; P1_R1240_U248
g8746 nand P1_R1240_U247 P1_R1240_U164 P1_R1240_U8 ; P1_R1240_U249
g8747 nand P1_R1240_U248 P1_R1240_U246 ; P1_R1240_U250
g8748 not P1_R1240_U163 ; P1_R1240_U251
g8749 or P1_U3495 P1_U3077 ; P1_R1240_U252
g8750 nand P1_R1240_U252 P1_R1240_U163 ; P1_R1240_U253
g8751 nand P1_U3077 P1_U3495 ; P1_R1240_U254
g8752 not P1_R1240_U161 ; P1_R1240_U255
g8753 or P1_U3498 P1_U3072 ; P1_R1240_U256
g8754 nand P1_R1240_U256 P1_R1240_U161 ; P1_R1240_U257
g8755 nand P1_U3072 P1_U3498 ; P1_R1240_U258
g8756 not P1_R1240_U93 ; P1_R1240_U259
g8757 or P1_U3067 P1_U3504 ; P1_R1240_U260
g8758 or P1_U3071 P1_U3501 ; P1_R1240_U261
g8759 not P1_R1240_U60 ; P1_R1240_U262
g8760 nand P1_R1240_U61 P1_R1240_U60 ; P1_R1240_U263
g8761 nand P1_U3067 P1_R1240_U263 ; P1_R1240_U264
g8762 nand P1_U3504 P1_R1240_U262 ; P1_R1240_U265
g8763 nand P1_R1240_U9 P1_R1240_U93 ; P1_R1240_U266
g8764 not P1_R1240_U159 ; P1_R1240_U267
g8765 or P1_U3074 P1_U4015 ; P1_R1240_U268
g8766 or P1_U3079 P1_U3509 ; P1_R1240_U269
g8767 or P1_U3073 P1_U4014 ; P1_R1240_U270
g8768 not P1_R1240_U81 ; P1_R1240_U271
g8769 nand P1_U4015 P1_R1240_U271 ; P1_R1240_U272
g8770 nand P1_R1240_U272 P1_R1240_U91 ; P1_R1240_U273
g8771 nand P1_R1240_U81 P1_R1240_U82 ; P1_R1240_U274
g8772 nand P1_R1240_U274 P1_R1240_U273 ; P1_R1240_U275
g8773 nand P1_R1240_U172 P1_R1240_U10 ; P1_R1240_U276
g8774 nand P1_U3073 P1_U4014 ; P1_R1240_U277
g8775 nand P1_R1240_U275 P1_R1240_U276 ; P1_R1240_U278
g8776 or P1_U3507 P1_U3080 ; P1_R1240_U279
g8777 or P1_U4014 P1_U3073 ; P1_R1240_U280
g8778 nand P1_R1240_U270 P1_R1240_U159 P1_R1240_U130 ; P1_R1240_U281
g8779 nand P1_R1240_U280 P1_R1240_U278 ; P1_R1240_U282
g8780 not P1_R1240_U155 ; P1_R1240_U283
g8781 or P1_U4013 P1_U3059 ; P1_R1240_U284
g8782 nand P1_R1240_U284 P1_R1240_U155 ; P1_R1240_U285
g8783 nand P1_U3059 P1_U4013 ; P1_R1240_U286
g8784 not P1_R1240_U153 ; P1_R1240_U287
g8785 or P1_U4012 P1_U3064 ; P1_R1240_U288
g8786 nand P1_R1240_U288 P1_R1240_U153 ; P1_R1240_U289
g8787 nand P1_U3064 P1_U4012 ; P1_R1240_U290
g8788 not P1_R1240_U151 ; P1_R1240_U291
g8789 or P1_U3056 P1_U4010 ; P1_R1240_U292
g8790 nand P1_R1240_U173 P1_R1240_U170 ; P1_R1240_U293
g8791 not P1_R1240_U87 ; P1_R1240_U294
g8792 or P1_U4011 P1_U3063 ; P1_R1240_U295
g8793 nand P1_R1240_U151 P1_R1240_U295 P1_R1240_U165 ; P1_R1240_U296
g8794 not P1_R1240_U149 ; P1_R1240_U297
g8795 or P1_U4008 P1_U3051 ; P1_R1240_U298
g8796 nand P1_U3051 P1_U4008 ; P1_R1240_U299
g8797 not P1_R1240_U147 ; P1_R1240_U300
g8798 nand P1_U4007 P1_R1240_U147 ; P1_R1240_U301
g8799 not P1_R1240_U145 ; P1_R1240_U302
g8800 nand P1_R1240_U295 P1_R1240_U151 ; P1_R1240_U303
g8801 not P1_R1240_U90 ; P1_R1240_U304
g8802 or P1_U4010 P1_U3056 ; P1_R1240_U305
g8803 nand P1_R1240_U305 P1_R1240_U90 ; P1_R1240_U306
g8804 nand P1_R1240_U306 P1_R1240_U170 P1_R1240_U150 ; P1_R1240_U307
g8805 nand P1_R1240_U304 P1_R1240_U170 ; P1_R1240_U308
g8806 nand P1_U4009 P1_U3055 ; P1_R1240_U309
g8807 nand P1_R1240_U308 P1_R1240_U309 P1_R1240_U165 ; P1_R1240_U310
g8808 or P1_U3056 P1_U4010 ; P1_R1240_U311
g8809 nand P1_R1240_U279 P1_R1240_U159 ; P1_R1240_U312
g8810 not P1_R1240_U92 ; P1_R1240_U313
g8811 nand P1_R1240_U10 P1_R1240_U92 ; P1_R1240_U314
g8812 nand P1_R1240_U134 P1_R1240_U314 ; P1_R1240_U315
g8813 nand P1_R1240_U314 P1_R1240_U275 ; P1_R1240_U316
g8814 nand P1_R1240_U450 P1_R1240_U316 ; P1_R1240_U317
g8815 or P1_U3509 P1_U3079 ; P1_R1240_U318
g8816 nand P1_R1240_U318 P1_R1240_U92 ; P1_R1240_U319
g8817 nand P1_R1240_U319 P1_R1240_U81 P1_R1240_U157 ; P1_R1240_U320
g8818 nand P1_R1240_U313 P1_R1240_U81 ; P1_R1240_U321
g8819 nand P1_U3074 P1_U4015 ; P1_R1240_U322
g8820 nand P1_R1240_U322 P1_R1240_U321 P1_R1240_U10 ; P1_R1240_U323
g8821 or P1_U3456 P1_U3076 ; P1_R1240_U324
g8822 not P1_R1240_U158 ; P1_R1240_U325
g8823 or P1_U3079 P1_U3509 ; P1_R1240_U326
g8824 or P1_U3501 P1_U3071 ; P1_R1240_U327
g8825 nand P1_R1240_U327 P1_R1240_U93 ; P1_R1240_U328
g8826 nand P1_R1240_U135 P1_R1240_U328 ; P1_R1240_U329
g8827 nand P1_R1240_U259 P1_R1240_U60 ; P1_R1240_U330
g8828 nand P1_U3504 P1_U3067 ; P1_R1240_U331
g8829 nand P1_R1240_U331 P1_R1240_U330 P1_R1240_U9 ; P1_R1240_U332
g8830 or P1_U3071 P1_U3501 ; P1_R1240_U333
g8831 nand P1_R1240_U247 P1_R1240_U164 ; P1_R1240_U334
g8832 not P1_R1240_U94 ; P1_R1240_U335
g8833 or P1_U3489 P1_U3070 ; P1_R1240_U336
g8834 nand P1_R1240_U336 P1_R1240_U94 ; P1_R1240_U337
g8835 nand P1_R1240_U136 P1_R1240_U337 ; P1_R1240_U338
g8836 nand P1_R1240_U335 P1_R1240_U169 ; P1_R1240_U339
g8837 nand P1_U3078 P1_U3492 ; P1_R1240_U340
g8838 nand P1_R1240_U137 P1_R1240_U339 ; P1_R1240_U341
g8839 or P1_U3070 P1_U3489 ; P1_R1240_U342
g8840 or P1_U3480 P1_U3081 ; P1_R1240_U343
g8841 nand P1_R1240_U343 P1_R1240_U41 ; P1_R1240_U344
g8842 nand P1_R1240_U138 P1_R1240_U344 ; P1_R1240_U345
g8843 nand P1_R1240_U203 P1_R1240_U168 ; P1_R1240_U346
g8844 nand P1_U3060 P1_U3483 ; P1_R1240_U347
g8845 nand P1_R1240_U139 P1_R1240_U346 ; P1_R1240_U348
g8846 nand P1_R1240_U204 P1_R1240_U168 ; P1_R1240_U349
g8847 nand P1_R1240_U201 P1_R1240_U62 ; P1_R1240_U350
g8848 nand P1_R1240_U211 P1_R1240_U23 ; P1_R1240_U351
g8849 nand P1_R1240_U225 P1_R1240_U35 ; P1_R1240_U352
g8850 nand P1_R1240_U228 P1_R1240_U177 ; P1_R1240_U353
g8851 nand P1_R1240_U311 P1_R1240_U170 ; P1_R1240_U354
g8852 nand P1_R1240_U295 P1_R1240_U173 ; P1_R1240_U355
g8853 nand P1_R1240_U326 P1_R1240_U81 ; P1_R1240_U356
g8854 nand P1_R1240_U279 P1_R1240_U78 ; P1_R1240_U357
g8855 nand P1_R1240_U333 P1_R1240_U60 ; P1_R1240_U358
g8856 nand P1_R1240_U342 P1_R1240_U169 ; P1_R1240_U359
g8857 nand P1_R1240_U247 P1_R1240_U69 ; P1_R1240_U360
g8858 nand P1_U4007 P1_U3052 ; P1_R1240_U361
g8859 nand P1_R1240_U293 P1_R1240_U165 ; P1_R1240_U362
g8860 nand P1_U3055 P1_R1240_U292 ; P1_R1240_U363
g8861 nand P1_U4009 P1_R1240_U292 ; P1_R1240_U364
g8862 nand P1_R1240_U293 P1_R1240_U165 P1_R1240_U298 ; P1_R1240_U365
g8863 nand P1_R1240_U151 P1_R1240_U165 P1_R1240_U132 ; P1_R1240_U366
g8864 nand P1_R1240_U294 P1_R1240_U298 ; P1_R1240_U367
g8865 nand P1_U3081 P1_R1240_U40 ; P1_R1240_U368
g8866 nand P1_U3480 P1_R1240_U39 ; P1_R1240_U369
g8867 nand P1_R1240_U369 P1_R1240_U368 ; P1_R1240_U370
g8868 nand P1_R1240_U349 P1_R1240_U41 ; P1_R1240_U371
g8869 nand P1_R1240_U370 P1_R1240_U203 ; P1_R1240_U372
g8870 nand P1_U3082 P1_R1240_U37 ; P1_R1240_U373
g8871 nand P1_U3477 P1_R1240_U38 ; P1_R1240_U374
g8872 nand P1_R1240_U374 P1_R1240_U373 ; P1_R1240_U375
g8873 nand P1_R1240_U350 P1_R1240_U140 ; P1_R1240_U376
g8874 nand P1_R1240_U200 P1_R1240_U375 ; P1_R1240_U377
g8875 nand P1_U3068 P1_R1240_U24 ; P1_R1240_U378
g8876 nand P1_U3474 P1_R1240_U22 ; P1_R1240_U379
g8877 nand P1_U3069 P1_R1240_U20 ; P1_R1240_U380
g8878 nand P1_U3471 P1_R1240_U21 ; P1_R1240_U381
g8879 nand P1_R1240_U381 P1_R1240_U380 ; P1_R1240_U382
g8880 nand P1_R1240_U351 P1_R1240_U42 ; P1_R1240_U383
g8881 nand P1_R1240_U382 P1_R1240_U192 ; P1_R1240_U384
g8882 nand P1_U3065 P1_R1240_U36 ; P1_R1240_U385
g8883 nand P1_U3468 P1_R1240_U27 ; P1_R1240_U386
g8884 nand P1_U3058 P1_R1240_U25 ; P1_R1240_U387
g8885 nand P1_U3465 P1_R1240_U26 ; P1_R1240_U388
g8886 nand P1_R1240_U388 P1_R1240_U387 ; P1_R1240_U389
g8887 nand P1_R1240_U352 P1_R1240_U45 ; P1_R1240_U390
g8888 nand P1_R1240_U389 P1_R1240_U218 ; P1_R1240_U391
g8889 nand P1_U3062 P1_R1240_U33 ; P1_R1240_U392
g8890 nand P1_U3462 P1_R1240_U34 ; P1_R1240_U393
g8891 nand P1_R1240_U393 P1_R1240_U392 ; P1_R1240_U394
g8892 nand P1_R1240_U353 P1_R1240_U141 ; P1_R1240_U395
g8893 nand P1_R1240_U227 P1_R1240_U394 ; P1_R1240_U396
g8894 nand P1_U3066 P1_R1240_U28 ; P1_R1240_U397
g8895 nand P1_U3459 P1_R1240_U29 ; P1_R1240_U398
g8896 nand P1_U3053 P1_R1240_U143 ; P1_R1240_U399
g8897 nand P1_U4018 P1_R1240_U142 ; P1_R1240_U400
g8898 nand P1_U3053 P1_R1240_U143 ; P1_R1240_U401
g8899 nand P1_U4018 P1_R1240_U142 ; P1_R1240_U402
g8900 nand P1_R1240_U402 P1_R1240_U401 ; P1_R1240_U403
g8901 nand P1_R1240_U144 P1_R1240_U145 ; P1_R1240_U404
g8902 nand P1_R1240_U302 P1_R1240_U403 ; P1_R1240_U405
g8903 nand P1_U3052 P1_R1240_U89 ; P1_R1240_U406
g8904 nand P1_U4007 P1_R1240_U88 ; P1_R1240_U407
g8905 nand P1_U3052 P1_R1240_U89 ; P1_R1240_U408
g8906 nand P1_U4007 P1_R1240_U88 ; P1_R1240_U409
g8907 nand P1_R1240_U409 P1_R1240_U408 ; P1_R1240_U410
g8908 nand P1_R1240_U146 P1_R1240_U147 ; P1_R1240_U411
g8909 nand P1_R1240_U300 P1_R1240_U410 ; P1_R1240_U412
g8910 nand P1_U3051 P1_R1240_U47 ; P1_R1240_U413
g8911 nand P1_U4008 P1_R1240_U48 ; P1_R1240_U414
g8912 nand P1_U3051 P1_R1240_U47 ; P1_R1240_U415
g8913 nand P1_U4008 P1_R1240_U48 ; P1_R1240_U416
g8914 nand P1_R1240_U416 P1_R1240_U415 ; P1_R1240_U417
g8915 nand P1_R1240_U148 P1_R1240_U149 ; P1_R1240_U418
g8916 nand P1_R1240_U297 P1_R1240_U417 ; P1_R1240_U419
g8917 nand P1_U3055 P1_R1240_U50 ; P1_R1240_U420
g8918 nand P1_U4009 P1_R1240_U49 ; P1_R1240_U421
g8919 nand P1_U3056 P1_R1240_U51 ; P1_R1240_U422
g8920 nand P1_U4010 P1_R1240_U52 ; P1_R1240_U423
g8921 nand P1_R1240_U423 P1_R1240_U422 ; P1_R1240_U424
g8922 nand P1_R1240_U354 P1_R1240_U90 ; P1_R1240_U425
g8923 nand P1_R1240_U424 P1_R1240_U304 ; P1_R1240_U426
g8924 nand P1_U3063 P1_R1240_U53 ; P1_R1240_U427
g8925 nand P1_U4011 P1_R1240_U54 ; P1_R1240_U428
g8926 nand P1_R1240_U428 P1_R1240_U427 ; P1_R1240_U429
g8927 nand P1_R1240_U355 P1_R1240_U151 ; P1_R1240_U430
g8928 nand P1_R1240_U291 P1_R1240_U429 ; P1_R1240_U431
g8929 nand P1_U3064 P1_R1240_U85 ; P1_R1240_U432
g8930 nand P1_U4012 P1_R1240_U86 ; P1_R1240_U433
g8931 nand P1_U3064 P1_R1240_U85 ; P1_R1240_U434
g8932 nand P1_U4012 P1_R1240_U86 ; P1_R1240_U435
g8933 nand P1_R1240_U435 P1_R1240_U434 ; P1_R1240_U436
g8934 nand P1_R1240_U152 P1_R1240_U153 ; P1_R1240_U437
g8935 nand P1_R1240_U287 P1_R1240_U436 ; P1_R1240_U438
g8936 nand P1_U3059 P1_R1240_U83 ; P1_R1240_U439
g8937 nand P1_U4013 P1_R1240_U84 ; P1_R1240_U440
g8938 nand P1_U3059 P1_R1240_U83 ; P1_R1240_U441
g8939 nand P1_U4013 P1_R1240_U84 ; P1_R1240_U442
g8940 nand P1_R1240_U442 P1_R1240_U441 ; P1_R1240_U443
g8941 nand P1_R1240_U154 P1_R1240_U155 ; P1_R1240_U444
g8942 nand P1_R1240_U283 P1_R1240_U443 ; P1_R1240_U445
g8943 nand P1_U3073 P1_R1240_U55 ; P1_R1240_U446
g8944 nand P1_U4014 P1_R1240_U56 ; P1_R1240_U447
g8945 nand P1_U3073 P1_R1240_U55 ; P1_R1240_U448
g8946 nand P1_U4014 P1_R1240_U56 ; P1_R1240_U449
g8947 nand P1_R1240_U449 P1_R1240_U448 ; P1_R1240_U450
g8948 nand P1_U3074 P1_R1240_U82 ; P1_R1240_U451
g8949 nand P1_U4015 P1_R1240_U91 ; P1_R1240_U452
g8950 nand P1_R1240_U179 P1_R1240_U158 ; P1_R1240_U453
g8951 nand P1_R1240_U325 P1_R1240_U32 ; P1_R1240_U454
g8952 nand P1_U3079 P1_R1240_U79 ; P1_R1240_U455
g8953 nand P1_U3509 P1_R1240_U80 ; P1_R1240_U456
g8954 nand P1_R1240_U456 P1_R1240_U455 ; P1_R1240_U457
g8955 nand P1_R1240_U356 P1_R1240_U92 ; P1_R1240_U458
g8956 nand P1_R1240_U457 P1_R1240_U313 ; P1_R1240_U459
g8957 nand P1_U3080 P1_R1240_U76 ; P1_R1240_U460
g8958 nand P1_U3507 P1_R1240_U77 ; P1_R1240_U461
g8959 nand P1_R1240_U461 P1_R1240_U460 ; P1_R1240_U462
g8960 nand P1_R1240_U357 P1_R1240_U159 ; P1_R1240_U463
g8961 nand P1_R1240_U267 P1_R1240_U462 ; P1_R1240_U464
g8962 nand P1_U3067 P1_R1240_U61 ; P1_R1240_U465
g8963 nand P1_U3504 P1_R1240_U59 ; P1_R1240_U466
g8964 nand P1_U3071 P1_R1240_U57 ; P1_R1240_U467
g8965 nand P1_U3501 P1_R1240_U58 ; P1_R1240_U468
g8966 nand P1_R1240_U468 P1_R1240_U467 ; P1_R1240_U469
g8967 nand P1_R1240_U358 P1_R1240_U93 ; P1_R1240_U470
g8968 nand P1_R1240_U469 P1_R1240_U259 ; P1_R1240_U471
g8969 nand P1_U3072 P1_R1240_U74 ; P1_R1240_U472
g8970 nand P1_U3498 P1_R1240_U75 ; P1_R1240_U473
g8971 nand P1_U3072 P1_R1240_U74 ; P1_R1240_U474
g8972 nand P1_U3498 P1_R1240_U75 ; P1_R1240_U475
g8973 nand P1_R1240_U475 P1_R1240_U474 ; P1_R1240_U476
g8974 nand P1_R1240_U160 P1_R1240_U161 ; P1_R1240_U477
g8975 nand P1_R1240_U255 P1_R1240_U476 ; P1_R1240_U478
g8976 nand P1_U3077 P1_R1240_U72 ; P1_R1240_U479
g8977 nand P1_U3495 P1_R1240_U73 ; P1_R1240_U480
g8978 nand P1_U3077 P1_R1240_U72 ; P1_R1240_U481
g8979 nand P1_U3495 P1_R1240_U73 ; P1_R1240_U482
g8980 nand P1_R1240_U482 P1_R1240_U481 ; P1_R1240_U483
g8981 nand P1_R1240_U162 P1_R1240_U163 ; P1_R1240_U484
g8982 nand P1_R1240_U251 P1_R1240_U483 ; P1_R1240_U485
g8983 nand P1_U3078 P1_R1240_U70 ; P1_R1240_U486
g8984 nand P1_U3492 P1_R1240_U71 ; P1_R1240_U487
g8985 nand P1_U3070 P1_R1240_U65 ; P1_R1240_U488
g8986 nand P1_U3489 P1_R1240_U66 ; P1_R1240_U489
g8987 nand P1_R1240_U489 P1_R1240_U488 ; P1_R1240_U490
g8988 nand P1_R1240_U359 P1_R1240_U94 ; P1_R1240_U491
g8989 nand P1_R1240_U490 P1_R1240_U335 ; P1_R1240_U492
g8990 nand P1_U3061 P1_R1240_U67 ; P1_R1240_U493
g8991 nand P1_U3486 P1_R1240_U68 ; P1_R1240_U494
g8992 nand P1_R1240_U494 P1_R1240_U493 ; P1_R1240_U495
g8993 nand P1_R1240_U360 P1_R1240_U164 ; P1_R1240_U496
g8994 nand P1_R1240_U241 P1_R1240_U495 ; P1_R1240_U497
g8995 nand P1_U3060 P1_R1240_U63 ; P1_R1240_U498
g8996 nand P1_U3483 P1_R1240_U64 ; P1_R1240_U499
g8997 nand P1_U3075 P1_R1240_U30 ; P1_R1240_U500
g8998 nand P1_U3451 P1_R1240_U31 ; P1_R1240_U501
g8999 and P1_R1162_U95 P1_R1162_U94 ; P1_R1162_U4
g9000 and P1_R1162_U96 P1_R1162_U97 ; P1_R1162_U5
g9001 and P1_R1162_U113 P1_R1162_U112 ; P1_R1162_U6
g9002 and P1_R1162_U155 P1_R1162_U154 ; P1_R1162_U7
g9003 and P1_R1162_U164 P1_R1162_U163 ; P1_R1162_U8
g9004 and P1_R1162_U182 P1_R1162_U181 ; P1_R1162_U9
g9005 and P1_R1162_U218 P1_R1162_U215 ; P1_R1162_U10
g9006 and P1_R1162_U211 P1_R1162_U208 ; P1_R1162_U11
g9007 and P1_R1162_U202 P1_R1162_U199 ; P1_R1162_U12
g9008 and P1_R1162_U196 P1_R1162_U192 ; P1_R1162_U13
g9009 and P1_R1162_U151 P1_R1162_U148 ; P1_R1162_U14
g9010 and P1_R1162_U143 P1_R1162_U140 ; P1_R1162_U15
g9011 and P1_R1162_U129 P1_R1162_U126 ; P1_R1162_U16
g9012 not P1_REG1_REG_6__SCAN_IN ; P1_R1162_U17
g9013 not P1_U3470 ; P1_R1162_U18
g9014 not P1_U3473 ; P1_R1162_U19
g9015 nand P1_U3470 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U20
g9016 not P1_REG1_REG_7__SCAN_IN ; P1_R1162_U21
g9017 not P1_REG1_REG_4__SCAN_IN ; P1_R1162_U22
g9018 not P1_U3464 ; P1_R1162_U23
g9019 not P1_U3467 ; P1_R1162_U24
g9020 not P1_REG1_REG_2__SCAN_IN ; P1_R1162_U25
g9021 not P1_U3458 ; P1_R1162_U26
g9022 not P1_REG1_REG_0__SCAN_IN ; P1_R1162_U27
g9023 not P1_U3449 ; P1_R1162_U28
g9024 nand P1_U3449 P1_REG1_REG_0__SCAN_IN ; P1_R1162_U29
g9025 not P1_REG1_REG_3__SCAN_IN ; P1_R1162_U30
g9026 not P1_U3461 ; P1_R1162_U31
g9027 nand P1_U3464 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U32
g9028 not P1_REG1_REG_5__SCAN_IN ; P1_R1162_U33
g9029 not P1_REG1_REG_8__SCAN_IN ; P1_R1162_U34
g9030 not P1_U3476 ; P1_R1162_U35
g9031 not P1_U3479 ; P1_R1162_U36
g9032 not P1_REG1_REG_9__SCAN_IN ; P1_R1162_U37
g9033 nand P1_R1162_U49 P1_R1162_U121 ; P1_R1162_U38
g9034 nand P1_R1162_U110 P1_R1162_U108 P1_R1162_U109 ; P1_R1162_U39
g9035 nand P1_R1162_U98 P1_R1162_U99 ; P1_R1162_U40
g9036 nand P1_U3455 P1_REG1_REG_1__SCAN_IN ; P1_R1162_U41
g9037 nand P1_R1162_U136 P1_R1162_U134 P1_R1162_U135 ; P1_R1162_U42
g9038 nand P1_R1162_U132 P1_R1162_U131 ; P1_R1162_U43
g9039 not P1_REG1_REG_16__SCAN_IN ; P1_R1162_U44
g9040 not P1_U3500 ; P1_R1162_U45
g9041 not P1_U3503 ; P1_R1162_U46
g9042 nand P1_U3500 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U47
g9043 not P1_REG1_REG_17__SCAN_IN ; P1_R1162_U48
g9044 nand P1_U3476 P1_REG1_REG_8__SCAN_IN ; P1_R1162_U49
g9045 not P1_REG1_REG_10__SCAN_IN ; P1_R1162_U50
g9046 not P1_U3482 ; P1_R1162_U51
g9047 not P1_REG1_REG_12__SCAN_IN ; P1_R1162_U52
g9048 not P1_U3488 ; P1_R1162_U53
g9049 not P1_REG1_REG_11__SCAN_IN ; P1_R1162_U54
g9050 not P1_U3485 ; P1_R1162_U55
g9051 nand P1_U3485 P1_REG1_REG_11__SCAN_IN ; P1_R1162_U56
g9052 not P1_REG1_REG_13__SCAN_IN ; P1_R1162_U57
g9053 not P1_U3491 ; P1_R1162_U58
g9054 not P1_REG1_REG_14__SCAN_IN ; P1_R1162_U59
g9055 not P1_U3494 ; P1_R1162_U60
g9056 not P1_REG1_REG_15__SCAN_IN ; P1_R1162_U61
g9057 not P1_U3497 ; P1_R1162_U62
g9058 not P1_REG1_REG_18__SCAN_IN ; P1_R1162_U63
g9059 not P1_U3506 ; P1_R1162_U64
g9060 nand P1_R1162_U186 P1_R1162_U185 P1_R1162_U187 ; P1_R1162_U65
g9061 nand P1_R1162_U179 P1_R1162_U178 ; P1_R1162_U66
g9062 nand P1_R1162_U56 P1_R1162_U204 ; P1_R1162_U67
g9063 nand P1_R1162_U259 P1_R1162_U258 ; P1_R1162_U68
g9064 nand P1_R1162_U308 P1_R1162_U307 ; P1_R1162_U69
g9065 nand P1_R1162_U231 P1_R1162_U230 ; P1_R1162_U70
g9066 nand P1_R1162_U236 P1_R1162_U235 ; P1_R1162_U71
g9067 nand P1_R1162_U243 P1_R1162_U242 ; P1_R1162_U72
g9068 nand P1_R1162_U250 P1_R1162_U249 ; P1_R1162_U73
g9069 nand P1_R1162_U255 P1_R1162_U254 ; P1_R1162_U74
g9070 nand P1_R1162_U271 P1_R1162_U270 ; P1_R1162_U75
g9071 nand P1_R1162_U278 P1_R1162_U277 ; P1_R1162_U76
g9072 nand P1_R1162_U285 P1_R1162_U284 ; P1_R1162_U77
g9073 nand P1_R1162_U292 P1_R1162_U291 ; P1_R1162_U78
g9074 nand P1_R1162_U299 P1_R1162_U298 ; P1_R1162_U79
g9075 nand P1_R1162_U304 P1_R1162_U303 ; P1_R1162_U80
g9076 nand P1_R1162_U117 P1_R1162_U116 P1_R1162_U118 ; P1_R1162_U81
g9077 nand P1_R1162_U133 P1_R1162_U145 ; P1_R1162_U82
g9078 nand P1_R1162_U41 P1_R1162_U152 ; P1_R1162_U83
g9079 not P1_U3443 ; P1_R1162_U84
g9080 not P1_REG1_REG_19__SCAN_IN ; P1_R1162_U85
g9081 nand P1_R1162_U175 P1_R1162_U174 ; P1_R1162_U86
g9082 nand P1_R1162_U171 P1_R1162_U170 ; P1_R1162_U87
g9083 nand P1_R1162_U161 P1_R1162_U160 ; P1_R1162_U88
g9084 not P1_R1162_U32 ; P1_R1162_U89
g9085 nand P1_U3479 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U90
g9086 nand P1_U3488 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U91
g9087 not P1_R1162_U56 ; P1_R1162_U92
g9088 not P1_R1162_U49 ; P1_R1162_U93
g9089 or P1_U3467 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U94
g9090 or P1_U3464 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U95
g9091 or P1_U3461 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U96
g9092 or P1_U3458 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U97
g9093 not P1_R1162_U29 ; P1_R1162_U98
g9094 or P1_U3455 P1_REG1_REG_1__SCAN_IN ; P1_R1162_U99
g9095 not P1_R1162_U40 ; P1_R1162_U100
g9096 not P1_R1162_U41 ; P1_R1162_U101
g9097 nand P1_R1162_U40 P1_R1162_U41 ; P1_R1162_U102
g9098 nand P1_U3458 P1_R1162_U96 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U103
g9099 nand P1_R1162_U5 P1_R1162_U102 ; P1_R1162_U104
g9100 nand P1_U3461 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U105
g9101 nand P1_R1162_U105 P1_R1162_U103 P1_R1162_U104 ; P1_R1162_U106
g9102 nand P1_R1162_U33 P1_R1162_U32 ; P1_R1162_U107
g9103 nand P1_U3467 P1_R1162_U107 ; P1_R1162_U108
g9104 nand P1_R1162_U4 P1_R1162_U106 ; P1_R1162_U109
g9105 nand P1_R1162_U89 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U110
g9106 not P1_R1162_U39 ; P1_R1162_U111
g9107 or P1_U3473 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U112
g9108 or P1_U3470 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U113
g9109 not P1_R1162_U20 ; P1_R1162_U114
g9110 nand P1_R1162_U21 P1_R1162_U20 ; P1_R1162_U115
g9111 nand P1_U3473 P1_R1162_U115 ; P1_R1162_U116
g9112 nand P1_R1162_U114 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U117
g9113 nand P1_R1162_U6 P1_R1162_U39 ; P1_R1162_U118
g9114 not P1_R1162_U81 ; P1_R1162_U119
g9115 or P1_U3476 P1_REG1_REG_8__SCAN_IN ; P1_R1162_U120
g9116 nand P1_R1162_U120 P1_R1162_U81 ; P1_R1162_U121
g9117 not P1_R1162_U38 ; P1_R1162_U122
g9118 or P1_U3479 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U123
g9119 or P1_U3470 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U124
g9120 nand P1_R1162_U124 P1_R1162_U39 ; P1_R1162_U125
g9121 nand P1_R1162_U238 P1_R1162_U237 P1_R1162_U20 P1_R1162_U125 ; P1_R1162_U126
g9122 nand P1_R1162_U111 P1_R1162_U20 ; P1_R1162_U127
g9123 nand P1_U3473 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U128
g9124 nand P1_R1162_U128 P1_R1162_U6 P1_R1162_U127 ; P1_R1162_U129
g9125 or P1_U3470 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U130
g9126 nand P1_R1162_U101 P1_R1162_U97 ; P1_R1162_U131
g9127 nand P1_U3458 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U132
g9128 not P1_R1162_U43 ; P1_R1162_U133
g9129 nand P1_R1162_U100 P1_R1162_U5 ; P1_R1162_U134
g9130 nand P1_R1162_U43 P1_R1162_U96 ; P1_R1162_U135
g9131 nand P1_U3461 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U136
g9132 not P1_R1162_U42 ; P1_R1162_U137
g9133 or P1_U3464 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U138
g9134 nand P1_R1162_U138 P1_R1162_U42 ; P1_R1162_U139
g9135 nand P1_R1162_U245 P1_R1162_U244 P1_R1162_U32 P1_R1162_U139 ; P1_R1162_U140
g9136 nand P1_R1162_U137 P1_R1162_U32 ; P1_R1162_U141
g9137 nand P1_U3467 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U142
g9138 nand P1_R1162_U142 P1_R1162_U4 P1_R1162_U141 ; P1_R1162_U143
g9139 or P1_U3464 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U144
g9140 nand P1_R1162_U100 P1_R1162_U97 ; P1_R1162_U145
g9141 not P1_R1162_U82 ; P1_R1162_U146
g9142 nand P1_U3461 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U147
g9143 nand P1_R1162_U257 P1_R1162_U256 P1_R1162_U41 P1_R1162_U40 ; P1_R1162_U148
g9144 nand P1_R1162_U41 P1_R1162_U40 ; P1_R1162_U149
g9145 nand P1_U3458 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U150
g9146 nand P1_R1162_U150 P1_R1162_U97 P1_R1162_U149 ; P1_R1162_U151
g9147 or P1_U3455 P1_REG1_REG_1__SCAN_IN ; P1_R1162_U152
g9148 not P1_R1162_U83 ; P1_R1162_U153
g9149 or P1_U3479 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U154
g9150 or P1_U3482 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U155
g9151 nand P1_R1162_U93 P1_R1162_U7 ; P1_R1162_U156
g9152 nand P1_U3482 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U157
g9153 nand P1_R1162_U157 P1_R1162_U90 P1_R1162_U156 ; P1_R1162_U158
g9154 or P1_U3482 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U159
g9155 nand P1_R1162_U120 P1_R1162_U7 P1_R1162_U81 ; P1_R1162_U160
g9156 nand P1_R1162_U159 P1_R1162_U158 ; P1_R1162_U161
g9157 not P1_R1162_U88 ; P1_R1162_U162
g9158 or P1_U3491 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U163
g9159 or P1_U3488 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U164
g9160 nand P1_R1162_U92 P1_R1162_U8 ; P1_R1162_U165
g9161 nand P1_U3491 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U166
g9162 nand P1_R1162_U166 P1_R1162_U91 P1_R1162_U165 ; P1_R1162_U167
g9163 or P1_U3485 P1_REG1_REG_11__SCAN_IN ; P1_R1162_U168
g9164 or P1_U3491 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U169
g9165 nand P1_R1162_U168 P1_R1162_U8 P1_R1162_U88 ; P1_R1162_U170
g9166 nand P1_R1162_U169 P1_R1162_U167 ; P1_R1162_U171
g9167 not P1_R1162_U87 ; P1_R1162_U172
g9168 or P1_U3494 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U173
g9169 nand P1_R1162_U173 P1_R1162_U87 ; P1_R1162_U174
g9170 nand P1_U3494 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U175
g9171 not P1_R1162_U86 ; P1_R1162_U176
g9172 or P1_U3497 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U177
g9173 nand P1_R1162_U177 P1_R1162_U86 ; P1_R1162_U178
g9174 nand P1_U3497 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U179
g9175 not P1_R1162_U66 ; P1_R1162_U180
g9176 or P1_U3503 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U181
g9177 or P1_U3500 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U182
g9178 not P1_R1162_U47 ; P1_R1162_U183
g9179 nand P1_R1162_U48 P1_R1162_U47 ; P1_R1162_U184
g9180 nand P1_U3503 P1_R1162_U184 ; P1_R1162_U185
g9181 nand P1_R1162_U183 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U186
g9182 nand P1_R1162_U9 P1_R1162_U66 ; P1_R1162_U187
g9183 not P1_R1162_U65 ; P1_R1162_U188
g9184 or P1_U3506 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U189
g9185 nand P1_R1162_U189 P1_R1162_U65 ; P1_R1162_U190
g9186 nand P1_U3506 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U191
g9187 nand P1_R1162_U261 P1_R1162_U260 P1_R1162_U191 P1_R1162_U190 ; P1_R1162_U192
g9188 nand P1_U3506 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U193
g9189 nand P1_R1162_U188 P1_R1162_U193 ; P1_R1162_U194
g9190 or P1_U3506 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U195
g9191 nand P1_R1162_U195 P1_R1162_U264 P1_R1162_U194 ; P1_R1162_U196
g9192 or P1_U3500 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U197
g9193 nand P1_R1162_U197 P1_R1162_U66 ; P1_R1162_U198
g9194 nand P1_R1162_U273 P1_R1162_U272 P1_R1162_U47 P1_R1162_U198 ; P1_R1162_U199
g9195 nand P1_R1162_U180 P1_R1162_U47 ; P1_R1162_U200
g9196 nand P1_U3503 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U201
g9197 nand P1_R1162_U201 P1_R1162_U9 P1_R1162_U200 ; P1_R1162_U202
g9198 or P1_U3500 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U203
g9199 nand P1_R1162_U168 P1_R1162_U88 ; P1_R1162_U204
g9200 not P1_R1162_U67 ; P1_R1162_U205
g9201 or P1_U3488 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U206
g9202 nand P1_R1162_U206 P1_R1162_U67 ; P1_R1162_U207
g9203 nand P1_R1162_U294 P1_R1162_U293 P1_R1162_U91 P1_R1162_U207 ; P1_R1162_U208
g9204 nand P1_R1162_U205 P1_R1162_U91 ; P1_R1162_U209
g9205 nand P1_U3491 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U210
g9206 nand P1_R1162_U210 P1_R1162_U8 P1_R1162_U209 ; P1_R1162_U211
g9207 or P1_U3488 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U212
g9208 or P1_U3479 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U213
g9209 nand P1_R1162_U213 P1_R1162_U38 ; P1_R1162_U214
g9210 nand P1_R1162_U306 P1_R1162_U305 P1_R1162_U90 P1_R1162_U214 ; P1_R1162_U215
g9211 nand P1_R1162_U122 P1_R1162_U90 ; P1_R1162_U216
g9212 nand P1_U3482 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U217
g9213 nand P1_R1162_U217 P1_R1162_U7 P1_R1162_U216 ; P1_R1162_U218
g9214 nand P1_R1162_U123 P1_R1162_U90 ; P1_R1162_U219
g9215 nand P1_R1162_U120 P1_R1162_U49 ; P1_R1162_U220
g9216 nand P1_R1162_U130 P1_R1162_U20 ; P1_R1162_U221
g9217 nand P1_R1162_U144 P1_R1162_U32 ; P1_R1162_U222
g9218 nand P1_R1162_U147 P1_R1162_U96 ; P1_R1162_U223
g9219 nand P1_R1162_U203 P1_R1162_U47 ; P1_R1162_U224
g9220 nand P1_R1162_U212 P1_R1162_U91 ; P1_R1162_U225
g9221 nand P1_R1162_U168 P1_R1162_U56 ; P1_R1162_U226
g9222 nand P1_U3479 P1_R1162_U37 ; P1_R1162_U227
g9223 nand P1_R1162_U36 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U228
g9224 nand P1_R1162_U228 P1_R1162_U227 ; P1_R1162_U229
g9225 nand P1_R1162_U219 P1_R1162_U38 ; P1_R1162_U230
g9226 nand P1_R1162_U229 P1_R1162_U122 ; P1_R1162_U231
g9227 nand P1_U3476 P1_R1162_U34 ; P1_R1162_U232
g9228 nand P1_R1162_U35 P1_REG1_REG_8__SCAN_IN ; P1_R1162_U233
g9229 nand P1_R1162_U233 P1_R1162_U232 ; P1_R1162_U234
g9230 nand P1_R1162_U220 P1_R1162_U81 ; P1_R1162_U235
g9231 nand P1_R1162_U119 P1_R1162_U234 ; P1_R1162_U236
g9232 nand P1_U3473 P1_R1162_U21 ; P1_R1162_U237
g9233 nand P1_R1162_U19 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U238
g9234 nand P1_U3470 P1_R1162_U17 ; P1_R1162_U239
g9235 nand P1_R1162_U18 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U240
g9236 nand P1_R1162_U240 P1_R1162_U239 ; P1_R1162_U241
g9237 nand P1_R1162_U221 P1_R1162_U39 ; P1_R1162_U242
g9238 nand P1_R1162_U241 P1_R1162_U111 ; P1_R1162_U243
g9239 nand P1_U3467 P1_R1162_U33 ; P1_R1162_U244
g9240 nand P1_R1162_U24 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U245
g9241 nand P1_U3464 P1_R1162_U22 ; P1_R1162_U246
g9242 nand P1_R1162_U23 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U247
g9243 nand P1_R1162_U247 P1_R1162_U246 ; P1_R1162_U248
g9244 nand P1_R1162_U222 P1_R1162_U42 ; P1_R1162_U249
g9245 nand P1_R1162_U248 P1_R1162_U137 ; P1_R1162_U250
g9246 nand P1_U3461 P1_R1162_U30 ; P1_R1162_U251
g9247 nand P1_R1162_U31 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U252
g9248 nand P1_R1162_U252 P1_R1162_U251 ; P1_R1162_U253
g9249 nand P1_R1162_U223 P1_R1162_U82 ; P1_R1162_U254
g9250 nand P1_R1162_U146 P1_R1162_U253 ; P1_R1162_U255
g9251 nand P1_U3458 P1_R1162_U25 ; P1_R1162_U256
g9252 nand P1_R1162_U26 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U257
g9253 nand P1_R1162_U98 P1_R1162_U83 ; P1_R1162_U258
g9254 nand P1_R1162_U153 P1_R1162_U29 ; P1_R1162_U259
g9255 nand P1_U3443 P1_R1162_U85 ; P1_R1162_U260
g9256 nand P1_R1162_U84 P1_REG1_REG_19__SCAN_IN ; P1_R1162_U261
g9257 nand P1_U3443 P1_R1162_U85 ; P1_R1162_U262
g9258 nand P1_R1162_U84 P1_REG1_REG_19__SCAN_IN ; P1_R1162_U263
g9259 nand P1_R1162_U263 P1_R1162_U262 ; P1_R1162_U264
g9260 nand P1_U3506 P1_R1162_U63 ; P1_R1162_U265
g9261 nand P1_R1162_U64 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U266
g9262 nand P1_U3506 P1_R1162_U63 ; P1_R1162_U267
g9263 nand P1_R1162_U64 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U268
g9264 nand P1_R1162_U268 P1_R1162_U267 ; P1_R1162_U269
g9265 nand P1_R1162_U266 P1_R1162_U265 P1_R1162_U65 ; P1_R1162_U270
g9266 nand P1_R1162_U269 P1_R1162_U188 ; P1_R1162_U271
g9267 nand P1_U3503 P1_R1162_U48 ; P1_R1162_U272
g9268 nand P1_R1162_U46 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U273
g9269 nand P1_U3500 P1_R1162_U44 ; P1_R1162_U274
g9270 nand P1_R1162_U45 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U275
g9271 nand P1_R1162_U275 P1_R1162_U274 ; P1_R1162_U276
g9272 nand P1_R1162_U224 P1_R1162_U66 ; P1_R1162_U277
g9273 nand P1_R1162_U276 P1_R1162_U180 ; P1_R1162_U278
g9274 nand P1_U3497 P1_R1162_U61 ; P1_R1162_U279
g9275 nand P1_R1162_U62 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U280
g9276 nand P1_U3497 P1_R1162_U61 ; P1_R1162_U281
g9277 nand P1_R1162_U62 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U282
g9278 nand P1_R1162_U282 P1_R1162_U281 ; P1_R1162_U283
g9279 nand P1_R1162_U280 P1_R1162_U279 P1_R1162_U86 ; P1_R1162_U284
g9280 nand P1_R1162_U176 P1_R1162_U283 ; P1_R1162_U285
g9281 nand P1_U3494 P1_R1162_U59 ; P1_R1162_U286
g9282 nand P1_R1162_U60 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U287
g9283 nand P1_U3494 P1_R1162_U59 ; P1_R1162_U288
g9284 nand P1_R1162_U60 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U289
g9285 nand P1_R1162_U289 P1_R1162_U288 ; P1_R1162_U290
g9286 nand P1_R1162_U287 P1_R1162_U286 P1_R1162_U87 ; P1_R1162_U291
g9287 nand P1_R1162_U172 P1_R1162_U290 ; P1_R1162_U292
g9288 nand P1_U3491 P1_R1162_U57 ; P1_R1162_U293
g9289 nand P1_R1162_U58 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U294
g9290 nand P1_U3488 P1_R1162_U52 ; P1_R1162_U295
g9291 nand P1_R1162_U53 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U296
g9292 nand P1_R1162_U296 P1_R1162_U295 ; P1_R1162_U297
g9293 nand P1_R1162_U225 P1_R1162_U67 ; P1_R1162_U298
g9294 nand P1_R1162_U297 P1_R1162_U205 ; P1_R1162_U299
g9295 nand P1_U3485 P1_R1162_U54 ; P1_R1162_U300
g9296 nand P1_R1162_U55 P1_REG1_REG_11__SCAN_IN ; P1_R1162_U301
g9297 nand P1_R1162_U301 P1_R1162_U300 ; P1_R1162_U302
g9298 nand P1_R1162_U226 P1_R1162_U88 ; P1_R1162_U303
g9299 nand P1_R1162_U162 P1_R1162_U302 ; P1_R1162_U304
g9300 nand P1_U3482 P1_R1162_U50 ; P1_R1162_U305
g9301 nand P1_R1162_U51 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U306
g9302 nand P1_U3449 P1_R1162_U27 ; P1_R1162_U307
g9303 nand P1_R1162_U28 P1_REG1_REG_0__SCAN_IN ; P1_R1162_U308
g9304 and P1_R1117_U184 P1_R1117_U201 ; P1_R1117_U6
g9305 and P1_R1117_U203 P1_R1117_U202 ; P1_R1117_U7
g9306 and P1_R1117_U179 P1_R1117_U240 ; P1_R1117_U8
g9307 and P1_R1117_U242 P1_R1117_U241 ; P1_R1117_U9
g9308 and P1_R1117_U259 P1_R1117_U258 ; P1_R1117_U10
g9309 and P1_R1117_U285 P1_R1117_U284 ; P1_R1117_U11
g9310 and P1_R1117_U383 P1_R1117_U382 ; P1_R1117_U12
g9311 nand P1_R1117_U340 P1_R1117_U343 ; P1_R1117_U13
g9312 nand P1_R1117_U329 P1_R1117_U332 ; P1_R1117_U14
g9313 nand P1_R1117_U318 P1_R1117_U321 ; P1_R1117_U15
g9314 nand P1_R1117_U310 P1_R1117_U312 ; P1_R1117_U16
g9315 nand P1_R1117_U156 P1_R1117_U175 P1_R1117_U348 ; P1_R1117_U17
g9316 nand P1_R1117_U236 P1_R1117_U238 ; P1_R1117_U18
g9317 nand P1_R1117_U228 P1_R1117_U231 ; P1_R1117_U19
g9318 nand P1_R1117_U220 P1_R1117_U222 ; P1_R1117_U20
g9319 nand P1_R1117_U25 P1_R1117_U346 ; P1_R1117_U21
g9320 not P1_U3474 ; P1_R1117_U22
g9321 not P1_U3459 ; P1_R1117_U23
g9322 not P1_U3451 ; P1_R1117_U24
g9323 nand P1_U3451 P1_R1117_U93 ; P1_R1117_U25
g9324 not P1_U3076 ; P1_R1117_U26
g9325 not P1_U3462 ; P1_R1117_U27
g9326 not P1_U3066 ; P1_R1117_U28
g9327 nand P1_U3066 P1_R1117_U23 ; P1_R1117_U29
g9328 not P1_U3062 ; P1_R1117_U30
g9329 not P1_U3471 ; P1_R1117_U31
g9330 not P1_U3468 ; P1_R1117_U32
g9331 not P1_U3465 ; P1_R1117_U33
g9332 not P1_U3069 ; P1_R1117_U34
g9333 not P1_U3065 ; P1_R1117_U35
g9334 not P1_U3058 ; P1_R1117_U36
g9335 nand P1_U3058 P1_R1117_U33 ; P1_R1117_U37
g9336 not P1_U3477 ; P1_R1117_U38
g9337 not P1_U3068 ; P1_R1117_U39
g9338 nand P1_U3068 P1_R1117_U22 ; P1_R1117_U40
g9339 not P1_U3082 ; P1_R1117_U41
g9340 not P1_U3480 ; P1_R1117_U42
g9341 not P1_U3081 ; P1_R1117_U43
g9342 nand P1_R1117_U209 P1_R1117_U208 ; P1_R1117_U44
g9343 nand P1_R1117_U37 P1_R1117_U224 ; P1_R1117_U45
g9344 nand P1_R1117_U193 P1_R1117_U192 ; P1_R1117_U46
g9345 not P1_U4009 ; P1_R1117_U47
g9346 not P1_U4013 ; P1_R1117_U48
g9347 not P1_U3498 ; P1_R1117_U49
g9348 not P1_U3486 ; P1_R1117_U50
g9349 not P1_U3483 ; P1_R1117_U51
g9350 not P1_U3061 ; P1_R1117_U52
g9351 not P1_U3060 ; P1_R1117_U53
g9352 nand P1_U3081 P1_R1117_U42 ; P1_R1117_U54
g9353 not P1_U3489 ; P1_R1117_U55
g9354 not P1_U3070 ; P1_R1117_U56
g9355 not P1_U3492 ; P1_R1117_U57
g9356 not P1_U3078 ; P1_R1117_U58
g9357 not P1_U3501 ; P1_R1117_U59
g9358 not P1_U3495 ; P1_R1117_U60
g9359 not P1_U3071 ; P1_R1117_U61
g9360 not P1_U3072 ; P1_R1117_U62
g9361 not P1_U3077 ; P1_R1117_U63
g9362 nand P1_U3077 P1_R1117_U60 ; P1_R1117_U64
g9363 not P1_U3504 ; P1_R1117_U65
g9364 not P1_U3067 ; P1_R1117_U66
g9365 nand P1_R1117_U269 P1_R1117_U268 ; P1_R1117_U67
g9366 not P1_U3080 ; P1_R1117_U68
g9367 not P1_U3509 ; P1_R1117_U69
g9368 not P1_U3079 ; P1_R1117_U70
g9369 not P1_U4015 ; P1_R1117_U71
g9370 not P1_U3074 ; P1_R1117_U72
g9371 not P1_U4012 ; P1_R1117_U73
g9372 not P1_U4014 ; P1_R1117_U74
g9373 not P1_U3064 ; P1_R1117_U75
g9374 not P1_U3059 ; P1_R1117_U76
g9375 not P1_U3073 ; P1_R1117_U77
g9376 nand P1_U3073 P1_R1117_U74 ; P1_R1117_U78
g9377 not P1_U4011 ; P1_R1117_U79
g9378 not P1_U3063 ; P1_R1117_U80
g9379 not P1_U4010 ; P1_R1117_U81
g9380 not P1_U3056 ; P1_R1117_U82
g9381 not P1_U4008 ; P1_R1117_U83
g9382 not P1_U3055 ; P1_R1117_U84
g9383 nand P1_U3055 P1_R1117_U47 ; P1_R1117_U85
g9384 not P1_U3051 ; P1_R1117_U86
g9385 not P1_U4007 ; P1_R1117_U87
g9386 not P1_U3052 ; P1_R1117_U88
g9387 nand P1_R1117_U299 P1_R1117_U298 ; P1_R1117_U89
g9388 nand P1_R1117_U78 P1_R1117_U314 ; P1_R1117_U90
g9389 nand P1_R1117_U64 P1_R1117_U325 ; P1_R1117_U91
g9390 nand P1_R1117_U54 P1_R1117_U336 ; P1_R1117_U92
g9391 not P1_U3075 ; P1_R1117_U93
g9392 nand P1_R1117_U393 P1_R1117_U392 ; P1_R1117_U94
g9393 nand P1_R1117_U407 P1_R1117_U406 ; P1_R1117_U95
g9394 nand P1_R1117_U412 P1_R1117_U411 ; P1_R1117_U96
g9395 nand P1_R1117_U428 P1_R1117_U427 ; P1_R1117_U97
g9396 nand P1_R1117_U433 P1_R1117_U432 ; P1_R1117_U98
g9397 nand P1_R1117_U438 P1_R1117_U437 ; P1_R1117_U99
g9398 nand P1_R1117_U443 P1_R1117_U442 ; P1_R1117_U100
g9399 nand P1_R1117_U448 P1_R1117_U447 ; P1_R1117_U101
g9400 nand P1_R1117_U464 P1_R1117_U463 ; P1_R1117_U102
g9401 nand P1_R1117_U469 P1_R1117_U468 ; P1_R1117_U103
g9402 nand P1_R1117_U352 P1_R1117_U351 ; P1_R1117_U104
g9403 nand P1_R1117_U361 P1_R1117_U360 ; P1_R1117_U105
g9404 nand P1_R1117_U368 P1_R1117_U367 ; P1_R1117_U106
g9405 nand P1_R1117_U372 P1_R1117_U371 ; P1_R1117_U107
g9406 nand P1_R1117_U381 P1_R1117_U380 ; P1_R1117_U108
g9407 nand P1_R1117_U402 P1_R1117_U401 ; P1_R1117_U109
g9408 nand P1_R1117_U419 P1_R1117_U418 ; P1_R1117_U110
g9409 nand P1_R1117_U423 P1_R1117_U422 ; P1_R1117_U111
g9410 nand P1_R1117_U455 P1_R1117_U454 ; P1_R1117_U112
g9411 nand P1_R1117_U459 P1_R1117_U458 ; P1_R1117_U113
g9412 nand P1_R1117_U476 P1_R1117_U475 ; P1_R1117_U114
g9413 and P1_R1117_U195 P1_R1117_U183 ; P1_R1117_U115
g9414 and P1_R1117_U198 P1_R1117_U199 ; P1_R1117_U116
g9415 and P1_R1117_U211 P1_R1117_U185 ; P1_R1117_U117
g9416 and P1_R1117_U214 P1_R1117_U215 ; P1_R1117_U118
g9417 and P1_R1117_U354 P1_R1117_U353 P1_R1117_U40 ; P1_R1117_U119
g9418 and P1_R1117_U357 P1_R1117_U185 ; P1_R1117_U120
g9419 and P1_R1117_U230 P1_R1117_U7 ; P1_R1117_U121
g9420 and P1_R1117_U364 P1_R1117_U184 ; P1_R1117_U122
g9421 and P1_R1117_U374 P1_R1117_U373 P1_R1117_U29 ; P1_R1117_U123
g9422 and P1_R1117_U377 P1_R1117_U183 ; P1_R1117_U124
g9423 and P1_R1117_U217 P1_R1117_U8 ; P1_R1117_U125
g9424 and P1_R1117_U262 P1_R1117_U180 ; P1_R1117_U126
g9425 and P1_R1117_U288 P1_R1117_U181 ; P1_R1117_U127
g9426 and P1_R1117_U304 P1_R1117_U305 ; P1_R1117_U128
g9427 and P1_R1117_U307 P1_R1117_U386 ; P1_R1117_U129
g9428 and P1_R1117_U305 P1_R1117_U304 P1_R1117_U308 ; P1_R1117_U130
g9429 nand P1_R1117_U390 P1_R1117_U389 ; P1_R1117_U131
g9430 and P1_R1117_U395 P1_R1117_U394 P1_R1117_U85 ; P1_R1117_U132
g9431 and P1_R1117_U398 P1_R1117_U182 ; P1_R1117_U133
g9432 nand P1_R1117_U404 P1_R1117_U403 ; P1_R1117_U134
g9433 nand P1_R1117_U409 P1_R1117_U408 ; P1_R1117_U135
g9434 and P1_R1117_U415 P1_R1117_U181 ; P1_R1117_U136
g9435 nand P1_R1117_U425 P1_R1117_U424 ; P1_R1117_U137
g9436 nand P1_R1117_U430 P1_R1117_U429 ; P1_R1117_U138
g9437 nand P1_R1117_U435 P1_R1117_U434 ; P1_R1117_U139
g9438 nand P1_R1117_U440 P1_R1117_U439 ; P1_R1117_U140
g9439 nand P1_R1117_U445 P1_R1117_U444 ; P1_R1117_U141
g9440 and P1_R1117_U451 P1_R1117_U180 ; P1_R1117_U142
g9441 nand P1_R1117_U461 P1_R1117_U460 ; P1_R1117_U143
g9442 nand P1_R1117_U466 P1_R1117_U465 ; P1_R1117_U144
g9443 and P1_R1117_U342 P1_R1117_U9 ; P1_R1117_U145
g9444 and P1_R1117_U472 P1_R1117_U179 ; P1_R1117_U146
g9445 and P1_R1117_U350 P1_R1117_U349 ; P1_R1117_U147
g9446 nand P1_R1117_U118 P1_R1117_U212 ; P1_R1117_U148
g9447 and P1_R1117_U359 P1_R1117_U358 ; P1_R1117_U149
g9448 and P1_R1117_U366 P1_R1117_U365 ; P1_R1117_U150
g9449 and P1_R1117_U370 P1_R1117_U369 ; P1_R1117_U151
g9450 nand P1_R1117_U116 P1_R1117_U196 ; P1_R1117_U152
g9451 and P1_R1117_U379 P1_R1117_U378 ; P1_R1117_U153
g9452 not P1_U4018 ; P1_R1117_U154
g9453 not P1_U3053 ; P1_R1117_U155
g9454 and P1_R1117_U388 P1_R1117_U387 ; P1_R1117_U156
g9455 nand P1_R1117_U128 P1_R1117_U302 ; P1_R1117_U157
g9456 and P1_R1117_U400 P1_R1117_U399 ; P1_R1117_U158
g9457 nand P1_R1117_U295 P1_R1117_U294 ; P1_R1117_U159
g9458 nand P1_R1117_U291 P1_R1117_U290 ; P1_R1117_U160
g9459 and P1_R1117_U417 P1_R1117_U416 ; P1_R1117_U161
g9460 and P1_R1117_U421 P1_R1117_U420 ; P1_R1117_U162
g9461 nand P1_R1117_U281 P1_R1117_U280 ; P1_R1117_U163
g9462 nand P1_R1117_U277 P1_R1117_U276 ; P1_R1117_U164
g9463 not P1_U3456 ; P1_R1117_U165
g9464 nand P1_R1117_U273 P1_R1117_U272 ; P1_R1117_U166
g9465 not P1_U3507 ; P1_R1117_U167
g9466 nand P1_R1117_U265 P1_R1117_U264 ; P1_R1117_U168
g9467 and P1_R1117_U453 P1_R1117_U452 ; P1_R1117_U169
g9468 and P1_R1117_U457 P1_R1117_U456 ; P1_R1117_U170
g9469 nand P1_R1117_U255 P1_R1117_U254 ; P1_R1117_U171
g9470 nand P1_R1117_U251 P1_R1117_U250 ; P1_R1117_U172
g9471 nand P1_R1117_U247 P1_R1117_U246 ; P1_R1117_U173
g9472 and P1_R1117_U474 P1_R1117_U473 ; P1_R1117_U174
g9473 nand P1_R1117_U129 P1_R1117_U157 ; P1_R1117_U175
g9474 not P1_R1117_U85 ; P1_R1117_U176
g9475 not P1_R1117_U29 ; P1_R1117_U177
g9476 not P1_R1117_U40 ; P1_R1117_U178
g9477 nand P1_U3483 P1_R1117_U53 ; P1_R1117_U179
g9478 nand P1_U3498 P1_R1117_U62 ; P1_R1117_U180
g9479 nand P1_U4013 P1_R1117_U76 ; P1_R1117_U181
g9480 nand P1_U4009 P1_R1117_U84 ; P1_R1117_U182
g9481 nand P1_U3459 P1_R1117_U28 ; P1_R1117_U183
g9482 nand P1_U3468 P1_R1117_U35 ; P1_R1117_U184
g9483 nand P1_U3474 P1_R1117_U39 ; P1_R1117_U185
g9484 not P1_R1117_U64 ; P1_R1117_U186
g9485 not P1_R1117_U78 ; P1_R1117_U187
g9486 not P1_R1117_U37 ; P1_R1117_U188
g9487 not P1_R1117_U54 ; P1_R1117_U189
g9488 not P1_R1117_U25 ; P1_R1117_U190
g9489 nand P1_R1117_U190 P1_R1117_U26 ; P1_R1117_U191
g9490 nand P1_R1117_U191 P1_R1117_U165 ; P1_R1117_U192
g9491 nand P1_U3076 P1_R1117_U25 ; P1_R1117_U193
g9492 not P1_R1117_U46 ; P1_R1117_U194
g9493 nand P1_U3462 P1_R1117_U30 ; P1_R1117_U195
g9494 nand P1_R1117_U115 P1_R1117_U46 ; P1_R1117_U196
g9495 nand P1_R1117_U30 P1_R1117_U29 ; P1_R1117_U197
g9496 nand P1_R1117_U197 P1_R1117_U27 ; P1_R1117_U198
g9497 nand P1_U3062 P1_R1117_U177 ; P1_R1117_U199
g9498 not P1_R1117_U152 ; P1_R1117_U200
g9499 nand P1_U3471 P1_R1117_U34 ; P1_R1117_U201
g9500 nand P1_U3069 P1_R1117_U31 ; P1_R1117_U202
g9501 nand P1_U3065 P1_R1117_U32 ; P1_R1117_U203
g9502 nand P1_R1117_U188 P1_R1117_U6 ; P1_R1117_U204
g9503 nand P1_R1117_U7 P1_R1117_U204 ; P1_R1117_U205
g9504 nand P1_U3465 P1_R1117_U36 ; P1_R1117_U206
g9505 nand P1_U3471 P1_R1117_U34 ; P1_R1117_U207
g9506 nand P1_R1117_U206 P1_R1117_U152 P1_R1117_U6 ; P1_R1117_U208
g9507 nand P1_R1117_U207 P1_R1117_U205 ; P1_R1117_U209
g9508 not P1_R1117_U44 ; P1_R1117_U210
g9509 nand P1_U3477 P1_R1117_U41 ; P1_R1117_U211
g9510 nand P1_R1117_U117 P1_R1117_U44 ; P1_R1117_U212
g9511 nand P1_R1117_U41 P1_R1117_U40 ; P1_R1117_U213
g9512 nand P1_R1117_U213 P1_R1117_U38 ; P1_R1117_U214
g9513 nand P1_U3082 P1_R1117_U178 ; P1_R1117_U215
g9514 not P1_R1117_U148 ; P1_R1117_U216
g9515 nand P1_U3480 P1_R1117_U43 ; P1_R1117_U217
g9516 nand P1_R1117_U217 P1_R1117_U54 ; P1_R1117_U218
g9517 nand P1_R1117_U210 P1_R1117_U40 ; P1_R1117_U219
g9518 nand P1_R1117_U120 P1_R1117_U219 ; P1_R1117_U220
g9519 nand P1_R1117_U44 P1_R1117_U185 ; P1_R1117_U221
g9520 nand P1_R1117_U119 P1_R1117_U221 ; P1_R1117_U222
g9521 nand P1_R1117_U40 P1_R1117_U185 ; P1_R1117_U223
g9522 nand P1_R1117_U206 P1_R1117_U152 ; P1_R1117_U224
g9523 not P1_R1117_U45 ; P1_R1117_U225
g9524 nand P1_U3065 P1_R1117_U32 ; P1_R1117_U226
g9525 nand P1_R1117_U225 P1_R1117_U226 ; P1_R1117_U227
g9526 nand P1_R1117_U122 P1_R1117_U227 ; P1_R1117_U228
g9527 nand P1_R1117_U45 P1_R1117_U184 ; P1_R1117_U229
g9528 nand P1_U3471 P1_R1117_U34 ; P1_R1117_U230
g9529 nand P1_R1117_U121 P1_R1117_U229 ; P1_R1117_U231
g9530 nand P1_U3065 P1_R1117_U32 ; P1_R1117_U232
g9531 nand P1_R1117_U184 P1_R1117_U232 ; P1_R1117_U233
g9532 nand P1_R1117_U206 P1_R1117_U37 ; P1_R1117_U234
g9533 nand P1_R1117_U194 P1_R1117_U29 ; P1_R1117_U235
g9534 nand P1_R1117_U124 P1_R1117_U235 ; P1_R1117_U236
g9535 nand P1_R1117_U46 P1_R1117_U183 ; P1_R1117_U237
g9536 nand P1_R1117_U123 P1_R1117_U237 ; P1_R1117_U238
g9537 nand P1_R1117_U29 P1_R1117_U183 ; P1_R1117_U239
g9538 nand P1_U3486 P1_R1117_U52 ; P1_R1117_U240
g9539 nand P1_U3061 P1_R1117_U50 ; P1_R1117_U241
g9540 nand P1_U3060 P1_R1117_U51 ; P1_R1117_U242
g9541 nand P1_R1117_U189 P1_R1117_U8 ; P1_R1117_U243
g9542 nand P1_R1117_U9 P1_R1117_U243 ; P1_R1117_U244
g9543 nand P1_U3486 P1_R1117_U52 ; P1_R1117_U245
g9544 nand P1_R1117_U125 P1_R1117_U148 ; P1_R1117_U246
g9545 nand P1_R1117_U245 P1_R1117_U244 ; P1_R1117_U247
g9546 not P1_R1117_U173 ; P1_R1117_U248
g9547 nand P1_U3489 P1_R1117_U56 ; P1_R1117_U249
g9548 nand P1_R1117_U249 P1_R1117_U173 ; P1_R1117_U250
g9549 nand P1_U3070 P1_R1117_U55 ; P1_R1117_U251
g9550 not P1_R1117_U172 ; P1_R1117_U252
g9551 nand P1_U3492 P1_R1117_U58 ; P1_R1117_U253
g9552 nand P1_R1117_U253 P1_R1117_U172 ; P1_R1117_U254
g9553 nand P1_U3078 P1_R1117_U57 ; P1_R1117_U255
g9554 not P1_R1117_U171 ; P1_R1117_U256
g9555 nand P1_U3501 P1_R1117_U61 ; P1_R1117_U257
g9556 nand P1_U3071 P1_R1117_U59 ; P1_R1117_U258
g9557 nand P1_U3072 P1_R1117_U49 ; P1_R1117_U259
g9558 nand P1_R1117_U186 P1_R1117_U180 ; P1_R1117_U260
g9559 nand P1_R1117_U10 P1_R1117_U260 ; P1_R1117_U261
g9560 nand P1_U3495 P1_R1117_U63 ; P1_R1117_U262
g9561 nand P1_U3501 P1_R1117_U61 ; P1_R1117_U263
g9562 nand P1_R1117_U171 P1_R1117_U126 P1_R1117_U257 ; P1_R1117_U264
g9563 nand P1_R1117_U263 P1_R1117_U261 ; P1_R1117_U265
g9564 not P1_R1117_U168 ; P1_R1117_U266
g9565 nand P1_U3504 P1_R1117_U66 ; P1_R1117_U267
g9566 nand P1_R1117_U267 P1_R1117_U168 ; P1_R1117_U268
g9567 nand P1_U3067 P1_R1117_U65 ; P1_R1117_U269
g9568 not P1_R1117_U67 ; P1_R1117_U270
g9569 nand P1_R1117_U270 P1_R1117_U68 ; P1_R1117_U271
g9570 nand P1_R1117_U271 P1_R1117_U167 ; P1_R1117_U272
g9571 nand P1_U3080 P1_R1117_U67 ; P1_R1117_U273
g9572 not P1_R1117_U166 ; P1_R1117_U274
g9573 nand P1_U3509 P1_R1117_U70 ; P1_R1117_U275
g9574 nand P1_R1117_U275 P1_R1117_U166 ; P1_R1117_U276
g9575 nand P1_U3079 P1_R1117_U69 ; P1_R1117_U277
g9576 not P1_R1117_U164 ; P1_R1117_U278
g9577 nand P1_U4015 P1_R1117_U72 ; P1_R1117_U279
g9578 nand P1_R1117_U279 P1_R1117_U164 ; P1_R1117_U280
g9579 nand P1_U3074 P1_R1117_U71 ; P1_R1117_U281
g9580 not P1_R1117_U163 ; P1_R1117_U282
g9581 nand P1_U4012 P1_R1117_U75 ; P1_R1117_U283
g9582 nand P1_U3064 P1_R1117_U73 ; P1_R1117_U284
g9583 nand P1_U3059 P1_R1117_U48 ; P1_R1117_U285
g9584 nand P1_R1117_U187 P1_R1117_U181 ; P1_R1117_U286
g9585 nand P1_R1117_U11 P1_R1117_U286 ; P1_R1117_U287
g9586 nand P1_U4014 P1_R1117_U77 ; P1_R1117_U288
g9587 nand P1_U4012 P1_R1117_U75 ; P1_R1117_U289
g9588 nand P1_R1117_U163 P1_R1117_U127 P1_R1117_U283 ; P1_R1117_U290
g9589 nand P1_R1117_U289 P1_R1117_U287 ; P1_R1117_U291
g9590 not P1_R1117_U160 ; P1_R1117_U292
g9591 nand P1_U4011 P1_R1117_U80 ; P1_R1117_U293
g9592 nand P1_R1117_U293 P1_R1117_U160 ; P1_R1117_U294
g9593 nand P1_U3063 P1_R1117_U79 ; P1_R1117_U295
g9594 not P1_R1117_U159 ; P1_R1117_U296
g9595 nand P1_U4010 P1_R1117_U82 ; P1_R1117_U297
g9596 nand P1_R1117_U297 P1_R1117_U159 ; P1_R1117_U298
g9597 nand P1_U3056 P1_R1117_U81 ; P1_R1117_U299
g9598 not P1_R1117_U89 ; P1_R1117_U300
g9599 nand P1_U4008 P1_R1117_U86 ; P1_R1117_U301
g9600 nand P1_R1117_U89 P1_R1117_U182 P1_R1117_U301 ; P1_R1117_U302
g9601 nand P1_R1117_U86 P1_R1117_U85 ; P1_R1117_U303
g9602 nand P1_R1117_U303 P1_R1117_U83 ; P1_R1117_U304
g9603 nand P1_U3051 P1_R1117_U176 ; P1_R1117_U305
g9604 not P1_R1117_U157 ; P1_R1117_U306
g9605 nand P1_U4007 P1_R1117_U88 ; P1_R1117_U307
g9606 nand P1_U3052 P1_R1117_U87 ; P1_R1117_U308
g9607 nand P1_R1117_U300 P1_R1117_U85 ; P1_R1117_U309
g9608 nand P1_R1117_U133 P1_R1117_U309 ; P1_R1117_U310
g9609 nand P1_R1117_U89 P1_R1117_U182 ; P1_R1117_U311
g9610 nand P1_R1117_U132 P1_R1117_U311 ; P1_R1117_U312
g9611 nand P1_R1117_U85 P1_R1117_U182 ; P1_R1117_U313
g9612 nand P1_R1117_U288 P1_R1117_U163 ; P1_R1117_U314
g9613 not P1_R1117_U90 ; P1_R1117_U315
g9614 nand P1_U3059 P1_R1117_U48 ; P1_R1117_U316
g9615 nand P1_R1117_U315 P1_R1117_U316 ; P1_R1117_U317
g9616 nand P1_R1117_U136 P1_R1117_U317 ; P1_R1117_U318
g9617 nand P1_R1117_U90 P1_R1117_U181 ; P1_R1117_U319
g9618 nand P1_U4012 P1_R1117_U75 ; P1_R1117_U320
g9619 nand P1_R1117_U320 P1_R1117_U319 P1_R1117_U11 ; P1_R1117_U321
g9620 nand P1_U3059 P1_R1117_U48 ; P1_R1117_U322
g9621 nand P1_R1117_U181 P1_R1117_U322 ; P1_R1117_U323
g9622 nand P1_R1117_U288 P1_R1117_U78 ; P1_R1117_U324
g9623 nand P1_R1117_U262 P1_R1117_U171 ; P1_R1117_U325
g9624 not P1_R1117_U91 ; P1_R1117_U326
g9625 nand P1_U3072 P1_R1117_U49 ; P1_R1117_U327
g9626 nand P1_R1117_U326 P1_R1117_U327 ; P1_R1117_U328
g9627 nand P1_R1117_U142 P1_R1117_U328 ; P1_R1117_U329
g9628 nand P1_R1117_U91 P1_R1117_U180 ; P1_R1117_U330
g9629 nand P1_U3501 P1_R1117_U61 ; P1_R1117_U331
g9630 nand P1_R1117_U331 P1_R1117_U330 P1_R1117_U10 ; P1_R1117_U332
g9631 nand P1_U3072 P1_R1117_U49 ; P1_R1117_U333
g9632 nand P1_R1117_U180 P1_R1117_U333 ; P1_R1117_U334
g9633 nand P1_R1117_U262 P1_R1117_U64 ; P1_R1117_U335
g9634 nand P1_R1117_U217 P1_R1117_U148 ; P1_R1117_U336
g9635 not P1_R1117_U92 ; P1_R1117_U337
g9636 nand P1_U3060 P1_R1117_U51 ; P1_R1117_U338
g9637 nand P1_R1117_U337 P1_R1117_U338 ; P1_R1117_U339
g9638 nand P1_R1117_U146 P1_R1117_U339 ; P1_R1117_U340
g9639 nand P1_R1117_U92 P1_R1117_U179 ; P1_R1117_U341
g9640 nand P1_U3486 P1_R1117_U52 ; P1_R1117_U342
g9641 nand P1_R1117_U145 P1_R1117_U341 ; P1_R1117_U343
g9642 nand P1_U3060 P1_R1117_U51 ; P1_R1117_U344
g9643 nand P1_R1117_U179 P1_R1117_U344 ; P1_R1117_U345
g9644 nand P1_U3075 P1_R1117_U24 ; P1_R1117_U346
g9645 nand P1_R1117_U89 P1_R1117_U182 P1_R1117_U301 ; P1_R1117_U347
g9646 nand P1_R1117_U12 P1_R1117_U347 P1_R1117_U130 ; P1_R1117_U348
g9647 nand P1_U3480 P1_R1117_U43 ; P1_R1117_U349
g9648 nand P1_U3081 P1_R1117_U42 ; P1_R1117_U350
g9649 nand P1_R1117_U218 P1_R1117_U148 ; P1_R1117_U351
g9650 nand P1_R1117_U216 P1_R1117_U147 ; P1_R1117_U352
g9651 nand P1_U3477 P1_R1117_U41 ; P1_R1117_U353
g9652 nand P1_U3082 P1_R1117_U38 ; P1_R1117_U354
g9653 nand P1_U3477 P1_R1117_U41 ; P1_R1117_U355
g9654 nand P1_U3082 P1_R1117_U38 ; P1_R1117_U356
g9655 nand P1_R1117_U356 P1_R1117_U355 ; P1_R1117_U357
g9656 nand P1_U3474 P1_R1117_U39 ; P1_R1117_U358
g9657 nand P1_U3068 P1_R1117_U22 ; P1_R1117_U359
g9658 nand P1_R1117_U223 P1_R1117_U44 ; P1_R1117_U360
g9659 nand P1_R1117_U149 P1_R1117_U210 ; P1_R1117_U361
g9660 nand P1_U3471 P1_R1117_U34 ; P1_R1117_U362
g9661 nand P1_U3069 P1_R1117_U31 ; P1_R1117_U363
g9662 nand P1_R1117_U363 P1_R1117_U362 ; P1_R1117_U364
g9663 nand P1_U3468 P1_R1117_U35 ; P1_R1117_U365
g9664 nand P1_U3065 P1_R1117_U32 ; P1_R1117_U366
g9665 nand P1_R1117_U233 P1_R1117_U45 ; P1_R1117_U367
g9666 nand P1_R1117_U150 P1_R1117_U225 ; P1_R1117_U368
g9667 nand P1_U3465 P1_R1117_U36 ; P1_R1117_U369
g9668 nand P1_U3058 P1_R1117_U33 ; P1_R1117_U370
g9669 nand P1_R1117_U234 P1_R1117_U152 ; P1_R1117_U371
g9670 nand P1_R1117_U200 P1_R1117_U151 ; P1_R1117_U372
g9671 nand P1_U3462 P1_R1117_U30 ; P1_R1117_U373
g9672 nand P1_U3062 P1_R1117_U27 ; P1_R1117_U374
g9673 nand P1_U3462 P1_R1117_U30 ; P1_R1117_U375
g9674 nand P1_U3062 P1_R1117_U27 ; P1_R1117_U376
g9675 nand P1_R1117_U376 P1_R1117_U375 ; P1_R1117_U377
g9676 nand P1_U3459 P1_R1117_U28 ; P1_R1117_U378
g9677 nand P1_U3066 P1_R1117_U23 ; P1_R1117_U379
g9678 nand P1_R1117_U239 P1_R1117_U46 ; P1_R1117_U380
g9679 nand P1_R1117_U153 P1_R1117_U194 ; P1_R1117_U381
g9680 nand P1_U4018 P1_R1117_U155 ; P1_R1117_U382
g9681 nand P1_U3053 P1_R1117_U154 ; P1_R1117_U383
g9682 nand P1_U4018 P1_R1117_U155 ; P1_R1117_U384
g9683 nand P1_U3053 P1_R1117_U154 ; P1_R1117_U385
g9684 nand P1_R1117_U385 P1_R1117_U384 ; P1_R1117_U386
g9685 nand P1_U3052 P1_R1117_U386 P1_R1117_U87 ; P1_R1117_U387
g9686 nand P1_R1117_U12 P1_R1117_U88 P1_U4007 ; P1_R1117_U388
g9687 nand P1_U4007 P1_R1117_U88 ; P1_R1117_U389
g9688 nand P1_U3052 P1_R1117_U87 ; P1_R1117_U390
g9689 not P1_R1117_U131 ; P1_R1117_U391
g9690 nand P1_R1117_U306 P1_R1117_U391 ; P1_R1117_U392
g9691 nand P1_R1117_U131 P1_R1117_U157 ; P1_R1117_U393
g9692 nand P1_U4008 P1_R1117_U86 ; P1_R1117_U394
g9693 nand P1_U3051 P1_R1117_U83 ; P1_R1117_U395
g9694 nand P1_U4008 P1_R1117_U86 ; P1_R1117_U396
g9695 nand P1_U3051 P1_R1117_U83 ; P1_R1117_U397
g9696 nand P1_R1117_U397 P1_R1117_U396 ; P1_R1117_U398
g9697 nand P1_U4009 P1_R1117_U84 ; P1_R1117_U399
g9698 nand P1_U3055 P1_R1117_U47 ; P1_R1117_U400
g9699 nand P1_R1117_U313 P1_R1117_U89 ; P1_R1117_U401
g9700 nand P1_R1117_U158 P1_R1117_U300 ; P1_R1117_U402
g9701 nand P1_U4010 P1_R1117_U82 ; P1_R1117_U403
g9702 nand P1_U3056 P1_R1117_U81 ; P1_R1117_U404
g9703 not P1_R1117_U134 ; P1_R1117_U405
g9704 nand P1_R1117_U296 P1_R1117_U405 ; P1_R1117_U406
g9705 nand P1_R1117_U134 P1_R1117_U159 ; P1_R1117_U407
g9706 nand P1_U4011 P1_R1117_U80 ; P1_R1117_U408
g9707 nand P1_U3063 P1_R1117_U79 ; P1_R1117_U409
g9708 not P1_R1117_U135 ; P1_R1117_U410
g9709 nand P1_R1117_U292 P1_R1117_U410 ; P1_R1117_U411
g9710 nand P1_R1117_U135 P1_R1117_U160 ; P1_R1117_U412
g9711 nand P1_U4012 P1_R1117_U75 ; P1_R1117_U413
g9712 nand P1_U3064 P1_R1117_U73 ; P1_R1117_U414
g9713 nand P1_R1117_U414 P1_R1117_U413 ; P1_R1117_U415
g9714 nand P1_U4013 P1_R1117_U76 ; P1_R1117_U416
g9715 nand P1_U3059 P1_R1117_U48 ; P1_R1117_U417
g9716 nand P1_R1117_U323 P1_R1117_U90 ; P1_R1117_U418
g9717 nand P1_R1117_U161 P1_R1117_U315 ; P1_R1117_U419
g9718 nand P1_U4014 P1_R1117_U77 ; P1_R1117_U420
g9719 nand P1_U3073 P1_R1117_U74 ; P1_R1117_U421
g9720 nand P1_R1117_U324 P1_R1117_U163 ; P1_R1117_U422
g9721 nand P1_R1117_U282 P1_R1117_U162 ; P1_R1117_U423
g9722 nand P1_U4015 P1_R1117_U72 ; P1_R1117_U424
g9723 nand P1_U3074 P1_R1117_U71 ; P1_R1117_U425
g9724 not P1_R1117_U137 ; P1_R1117_U426
g9725 nand P1_R1117_U278 P1_R1117_U426 ; P1_R1117_U427
g9726 nand P1_R1117_U137 P1_R1117_U164 ; P1_R1117_U428
g9727 nand P1_U3456 P1_R1117_U26 ; P1_R1117_U429
g9728 nand P1_U3076 P1_R1117_U165 ; P1_R1117_U430
g9729 not P1_R1117_U138 ; P1_R1117_U431
g9730 nand P1_R1117_U431 P1_R1117_U190 ; P1_R1117_U432
g9731 nand P1_R1117_U138 P1_R1117_U25 ; P1_R1117_U433
g9732 nand P1_U3509 P1_R1117_U70 ; P1_R1117_U434
g9733 nand P1_U3079 P1_R1117_U69 ; P1_R1117_U435
g9734 not P1_R1117_U139 ; P1_R1117_U436
g9735 nand P1_R1117_U274 P1_R1117_U436 ; P1_R1117_U437
g9736 nand P1_R1117_U139 P1_R1117_U166 ; P1_R1117_U438
g9737 nand P1_U3507 P1_R1117_U68 ; P1_R1117_U439
g9738 nand P1_U3080 P1_R1117_U167 ; P1_R1117_U440
g9739 not P1_R1117_U140 ; P1_R1117_U441
g9740 nand P1_R1117_U441 P1_R1117_U270 ; P1_R1117_U442
g9741 nand P1_R1117_U140 P1_R1117_U67 ; P1_R1117_U443
g9742 nand P1_U3504 P1_R1117_U66 ; P1_R1117_U444
g9743 nand P1_U3067 P1_R1117_U65 ; P1_R1117_U445
g9744 not P1_R1117_U141 ; P1_R1117_U446
g9745 nand P1_R1117_U266 P1_R1117_U446 ; P1_R1117_U447
g9746 nand P1_R1117_U141 P1_R1117_U168 ; P1_R1117_U448
g9747 nand P1_U3501 P1_R1117_U61 ; P1_R1117_U449
g9748 nand P1_U3071 P1_R1117_U59 ; P1_R1117_U450
g9749 nand P1_R1117_U450 P1_R1117_U449 ; P1_R1117_U451
g9750 nand P1_U3498 P1_R1117_U62 ; P1_R1117_U452
g9751 nand P1_U3072 P1_R1117_U49 ; P1_R1117_U453
g9752 nand P1_R1117_U334 P1_R1117_U91 ; P1_R1117_U454
g9753 nand P1_R1117_U169 P1_R1117_U326 ; P1_R1117_U455
g9754 nand P1_U3495 P1_R1117_U63 ; P1_R1117_U456
g9755 nand P1_U3077 P1_R1117_U60 ; P1_R1117_U457
g9756 nand P1_R1117_U335 P1_R1117_U171 ; P1_R1117_U458
g9757 nand P1_R1117_U256 P1_R1117_U170 ; P1_R1117_U459
g9758 nand P1_U3492 P1_R1117_U58 ; P1_R1117_U460
g9759 nand P1_U3078 P1_R1117_U57 ; P1_R1117_U461
g9760 not P1_R1117_U143 ; P1_R1117_U462
g9761 nand P1_R1117_U252 P1_R1117_U462 ; P1_R1117_U463
g9762 nand P1_R1117_U143 P1_R1117_U172 ; P1_R1117_U464
g9763 nand P1_U3489 P1_R1117_U56 ; P1_R1117_U465
g9764 nand P1_U3070 P1_R1117_U55 ; P1_R1117_U466
g9765 not P1_R1117_U144 ; P1_R1117_U467
g9766 nand P1_R1117_U248 P1_R1117_U467 ; P1_R1117_U468
g9767 nand P1_R1117_U144 P1_R1117_U173 ; P1_R1117_U469
g9768 nand P1_U3486 P1_R1117_U52 ; P1_R1117_U470
g9769 nand P1_U3061 P1_R1117_U50 ; P1_R1117_U471
g9770 nand P1_R1117_U471 P1_R1117_U470 ; P1_R1117_U472
g9771 nand P1_U3483 P1_R1117_U53 ; P1_R1117_U473
g9772 nand P1_U3060 P1_R1117_U51 ; P1_R1117_U474
g9773 nand P1_R1117_U345 P1_R1117_U92 ; P1_R1117_U475
g9774 nand P1_R1117_U174 P1_R1117_U337 ; P1_R1117_U476
g9775 and P1_R1375_U119 P1_R1375_U120 ; P1_R1375_U6
g9776 and P1_R1375_U137 P1_R1375_U136 ; P1_R1375_U7
g9777 and P1_R1375_U144 P1_R1375_U143 P1_R1375_U142 P1_R1375_U141 ; P1_R1375_U8
g9778 and P1_R1375_U164 P1_R1375_U163 ; P1_R1375_U9
g9779 and P1_R1375_U197 P1_R1375_U196 P1_R1375_U198 P1_R1375_U6 ; P1_R1375_U10
g9780 and P1_U4018 P1_R1375_U20 ; P1_R1375_U11
g9781 and P1_R1375_U207 P1_R1375_U206 P1_R1375_U118 P1_R1375_U117 ; P1_R1375_U12
g9782 and P1_U3451 P1_R1375_U48 ; P1_R1375_U13
g9783 and P1_R1375_U205 P1_R1375_U115 P1_R1375_U204 ; P1_R1375_U14
g9784 not P1_U4016 ; P1_R1375_U15
g9785 not P1_U4017 ; P1_R1375_U16
g9786 not P1_U3054 ; P1_R1375_U17
g9787 not P1_U4018 ; P1_R1375_U18
g9788 not P1_U3057 ; P1_R1375_U19
g9789 not P1_U3053 ; P1_R1375_U20
g9790 not P1_U3052 ; P1_R1375_U21
g9791 not P1_U4008 ; P1_R1375_U22
g9792 not P1_U3055 ; P1_R1375_U23
g9793 not P1_U4010 ; P1_R1375_U24
g9794 not P1_U4007 ; P1_R1375_U25
g9795 not P1_U4009 ; P1_R1375_U26
g9796 not P1_U4011 ; P1_R1375_U27
g9797 not P1_U3064 ; P1_R1375_U28
g9798 not P1_U4012 ; P1_R1375_U29
g9799 not P1_U3059 ; P1_R1375_U30
g9800 not P1_U3056 ; P1_R1375_U31
g9801 not P1_U3063 ; P1_R1375_U32
g9802 not P1_U3073 ; P1_R1375_U33
g9803 not P1_U3074 ; P1_R1375_U34
g9804 not P1_U3504 ; P1_R1375_U35
g9805 not P1_U3507 ; P1_R1375_U36
g9806 not P1_U3072 ; P1_R1375_U37
g9807 not P1_U3077 ; P1_R1375_U38
g9808 not P1_U3471 ; P1_R1375_U39
g9809 not P1_U3065 ; P1_R1375_U40
g9810 not P1_U3081 ; P1_R1375_U41
g9811 not P1_U3082 ; P1_R1375_U42
g9812 not P1_U3069 ; P1_R1375_U43
g9813 not P1_U3068 ; P1_R1375_U44
g9814 not P1_U3058 ; P1_R1375_U45
g9815 not P1_U3062 ; P1_R1375_U46
g9816 not P1_U3451 ; P1_R1375_U47
g9817 not P1_U3075 ; P1_R1375_U48
g9818 nand P1_R1375_U147 P1_R1375_U146 ; P1_R1375_U49
g9819 not P1_U3456 ; P1_R1375_U50
g9820 not P1_U3066 ; P1_R1375_U51
g9821 not P1_U3486 ; P1_R1375_U52
g9822 not P1_U3489 ; P1_R1375_U53
g9823 not P1_U3459 ; P1_R1375_U54
g9824 not P1_U3462 ; P1_R1375_U55
g9825 not P1_U3468 ; P1_R1375_U56
g9826 not P1_U3465 ; P1_R1375_U57
g9827 not P1_U3474 ; P1_R1375_U58
g9828 not P1_U3477 ; P1_R1375_U59
g9829 not P1_U3480 ; P1_R1375_U60
g9830 not P1_U3483 ; P1_R1375_U61
g9831 not P1_U3060 ; P1_R1375_U62
g9832 not P1_U3070 ; P1_R1375_U63
g9833 not P1_U3061 ; P1_R1375_U64
g9834 not P1_U3078 ; P1_R1375_U65
g9835 not P1_U3492 ; P1_R1375_U66
g9836 not P1_U3495 ; P1_R1375_U67
g9837 not P1_U3498 ; P1_R1375_U68
g9838 not P1_U3501 ; P1_R1375_U69
g9839 not P1_U3071 ; P1_R1375_U70
g9840 not P1_U3067 ; P1_R1375_U71
g9841 not P1_U3080 ; P1_R1375_U72
g9842 not P1_U3079 ; P1_R1375_U73
g9843 not P1_U3509 ; P1_R1375_U74
g9844 not P1_U4015 ; P1_R1375_U75
g9845 not P1_U4014 ; P1_R1375_U76
g9846 not P1_U4013 ; P1_R1375_U77
g9847 nand P1_R1375_U11 P1_R1375_U125 ; P1_R1375_U78
g9848 nand P1_R1375_U124 P1_R1375_U122 P1_R1375_U87 P1_R1375_U12 ; P1_R1375_U79
g9849 nand P1_R1375_U109 P1_R1375_U195 ; P1_R1375_U80
g9850 and P1_U4008 P1_R1375_U113 ; P1_R1375_U81
g9851 and P1_U4010 P1_R1375_U31 ; P1_R1375_U82
g9852 and P1_U4007 P1_R1375_U21 ; P1_R1375_U83
g9853 and P1_U4009 P1_R1375_U23 ; P1_R1375_U84
g9854 and P1_U3064 P1_R1375_U29 ; P1_R1375_U85
g9855 and P1_U3059 P1_R1375_U77 ; P1_R1375_U86
g9856 and P1_R1375_U123 P1_R1375_U121 ; P1_R1375_U87
g9857 and P1_R1375_U129 P1_R1375_U126 ; P1_R1375_U88
g9858 and P1_R1375_U131 P1_R1375_U201 P1_R1375_U128 ; P1_R1375_U89
g9859 and P1_U3065 P1_R1375_U56 ; P1_R1375_U90
g9860 and P1_R1375_U145 P1_R1375_U149 ; P1_R1375_U91
g9861 and P1_R1375_U91 P1_R1375_U140 ; P1_R1375_U92
g9862 and P1_R1375_U153 P1_R1375_U152 P1_R1375_U8 ; P1_R1375_U93
g9863 and P1_U3459 P1_R1375_U51 ; P1_R1375_U94
g9864 and P1_R1375_U161 P1_R1375_U160 P1_R1375_U159 ; P1_R1375_U95
g9865 and P1_U3474 P1_R1375_U44 ; P1_R1375_U96
g9866 and P1_R1375_U171 P1_R1375_U170 ; P1_R1375_U97
g9867 and P1_R1375_U97 P1_R1375_U9 ; P1_R1375_U98
g9868 and P1_U3060 P1_R1375_U61 ; P1_R1375_U99
g9869 and P1_U3061 P1_R1375_U52 ; P1_R1375_U100
g9870 and P1_R1375_U173 P1_R1375_U174 P1_R1375_U102 ; P1_R1375_U101
g9871 and P1_R1375_U177 P1_R1375_U176 ; P1_R1375_U102
g9872 and P1_R1375_U7 P1_R1375_U104 ; P1_R1375_U103
g9873 and P1_R1375_U185 P1_R1375_U186 ; P1_R1375_U104
g9874 and P1_U3071 P1_R1375_U69 ; P1_R1375_U105
g9875 and P1_U3067 P1_R1375_U35 ; P1_R1375_U106
g9876 and P1_R1375_U188 P1_R1375_U190 P1_R1375_U108 ; P1_R1375_U107
g9877 and P1_R1375_U192 P1_R1375_U191 ; P1_R1375_U108
g9878 and P1_R1375_U134 P1_R1375_U133 ; P1_R1375_U109
g9879 and P1_U4015 P1_R1375_U34 ; P1_R1375_U110
g9880 and P1_R1375_U128 P1_R1375_U127 ; P1_R1375_U111
g9881 and P1_R1375_U10 P1_R1375_U131 P1_R1375_U129 P1_R1375_U130 ; P1_R1375_U112
g9882 not P1_U3051 ; P1_R1375_U113
g9883 nand P1_R1375_U200 P1_R1375_U199 ; P1_R1375_U114
g9884 nand P1_U4016 P1_R1375_U17 ; P1_R1375_U115
g9885 nand P1_U3053 P1_R1375_U18 ; P1_R1375_U116
g9886 nand P1_U3052 P1_R1375_U25 ; P1_R1375_U117
g9887 nand P1_U3055 P1_R1375_U26 ; P1_R1375_U118
g9888 nand P1_U4011 P1_R1375_U32 ; P1_R1375_U119
g9889 nand P1_U4012 P1_R1375_U28 ; P1_R1375_U120
g9890 nand P1_R1375_U85 P1_R1375_U119 ; P1_R1375_U121
g9891 nand P1_R1375_U86 P1_R1375_U6 ; P1_R1375_U122
g9892 nand P1_U3056 P1_R1375_U24 ; P1_R1375_U123
g9893 nand P1_U3063 P1_R1375_U27 ; P1_R1375_U124
g9894 nand P1_U3057 P1_R1375_U16 ; P1_R1375_U125
g9895 nand P1_R1375_U81 P1_R1375_U117 P1_R1375_U115 ; P1_R1375_U126
g9896 nand P1_R1375_U82 P1_R1375_U12 P1_R1375_U115 ; P1_R1375_U127
g9897 nand P1_R1375_U115 P1_R1375_U19 P1_U4017 ; P1_R1375_U128
g9898 nand P1_R1375_U83 P1_R1375_U115 ; P1_R1375_U129
g9899 nand P1_R1375_U84 P1_R1375_U12 P1_R1375_U115 ; P1_R1375_U130
g9900 nand P1_U3054 P1_R1375_U15 ; P1_R1375_U131
g9901 nand P1_R1375_U79 P1_R1375_U130 P1_R1375_U88 P1_R1375_U127 ; P1_R1375_U132
g9902 nand P1_U3073 P1_R1375_U76 ; P1_R1375_U133
g9903 nand P1_U3074 P1_R1375_U75 ; P1_R1375_U134
g9904 nand P1_U3072 P1_R1375_U68 ; P1_R1375_U135
g9905 nand P1_U3504 P1_R1375_U71 ; P1_R1375_U136
g9906 nand P1_U3507 P1_R1375_U72 ; P1_R1375_U137
g9907 nand P1_U3077 P1_R1375_U67 ; P1_R1375_U138
g9908 nand P1_U3471 P1_R1375_U43 ; P1_R1375_U139
g9909 nand P1_R1375_U90 P1_R1375_U139 ; P1_R1375_U140
g9910 nand P1_U3081 P1_R1375_U60 ; P1_R1375_U141
g9911 nand P1_U3082 P1_R1375_U59 ; P1_R1375_U142
g9912 nand P1_U3069 P1_R1375_U39 ; P1_R1375_U143
g9913 nand P1_U3068 P1_R1375_U58 ; P1_R1375_U144
g9914 nand P1_U3058 P1_R1375_U57 ; P1_R1375_U145
g9915 or P1_U3448 P1_R1375_U13 ; P1_R1375_U146
g9916 nand P1_U3075 P1_R1375_U47 ; P1_R1375_U147
g9917 not P1_R1375_U49 ; P1_R1375_U148
g9918 nand P1_U3062 P1_R1375_U55 ; P1_R1375_U149
g9919 nand P1_U3456 P1_R1375_U148 ; P1_R1375_U150
g9920 nand P1_U3076 P1_R1375_U150 ; P1_R1375_U151
g9921 nand P1_R1375_U49 P1_R1375_U50 ; P1_R1375_U152
g9922 nand P1_U3066 P1_R1375_U54 ; P1_R1375_U153
g9923 nand P1_R1375_U92 P1_R1375_U151 P1_R1375_U93 ; P1_R1375_U154
g9924 nand P1_R1375_U94 P1_R1375_U149 ; P1_R1375_U155
g9925 nand P1_U3462 P1_R1375_U46 ; P1_R1375_U156
g9926 nand P1_R1375_U156 P1_R1375_U155 ; P1_R1375_U157
g9927 nand P1_R1375_U157 P1_R1375_U145 ; P1_R1375_U158
g9928 nand P1_U3468 P1_R1375_U40 ; P1_R1375_U159
g9929 nand P1_U3465 P1_R1375_U45 ; P1_R1375_U160
g9930 nand P1_U3471 P1_R1375_U43 ; P1_R1375_U161
g9931 nand P1_R1375_U158 P1_R1375_U95 ; P1_R1375_U162
g9932 nand P1_U3486 P1_R1375_U64 ; P1_R1375_U163
g9933 nand P1_U3489 P1_R1375_U63 ; P1_R1375_U164
g9934 nand P1_R1375_U96 P1_R1375_U142 ; P1_R1375_U165
g9935 nand P1_U3477 P1_R1375_U42 ; P1_R1375_U166
g9936 nand P1_R1375_U166 P1_R1375_U165 ; P1_R1375_U167
g9937 nand P1_R1375_U162 P1_R1375_U140 P1_R1375_U8 ; P1_R1375_U168
g9938 nand P1_R1375_U167 P1_R1375_U141 ; P1_R1375_U169
g9939 nand P1_U3480 P1_R1375_U41 ; P1_R1375_U170
g9940 nand P1_U3483 P1_R1375_U62 ; P1_R1375_U171
g9941 nand P1_R1375_U168 P1_R1375_U169 P1_R1375_U98 P1_R1375_U154 ; P1_R1375_U172
g9942 nand P1_R1375_U99 P1_R1375_U9 ; P1_R1375_U173
g9943 nand P1_U3070 P1_R1375_U53 ; P1_R1375_U174
g9944 nand P1_U3489 P1_R1375_U63 ; P1_R1375_U175
g9945 nand P1_R1375_U100 P1_R1375_U175 ; P1_R1375_U176
g9946 nand P1_U3078 P1_R1375_U66 ; P1_R1375_U177
g9947 nand P1_R1375_U172 P1_R1375_U101 ; P1_R1375_U178
g9948 nand P1_U3492 P1_R1375_U65 ; P1_R1375_U179
g9949 nand P1_R1375_U179 P1_R1375_U178 ; P1_R1375_U180
g9950 nand P1_R1375_U180 P1_R1375_U138 ; P1_R1375_U181
g9951 nand P1_U3495 P1_R1375_U38 ; P1_R1375_U182
g9952 nand P1_R1375_U182 P1_R1375_U181 ; P1_R1375_U183
g9953 nand P1_R1375_U183 P1_R1375_U135 ; P1_R1375_U184
g9954 nand P1_U3498 P1_R1375_U37 ; P1_R1375_U185
g9955 nand P1_U3501 P1_R1375_U70 ; P1_R1375_U186
g9956 nand P1_R1375_U184 P1_R1375_U103 ; P1_R1375_U187
g9957 nand P1_R1375_U105 P1_R1375_U7 ; P1_R1375_U188
g9958 nand P1_U3507 P1_R1375_U72 ; P1_R1375_U189
g9959 nand P1_R1375_U106 P1_R1375_U189 ; P1_R1375_U190
g9960 nand P1_U3080 P1_R1375_U36 ; P1_R1375_U191
g9961 nand P1_U3079 P1_R1375_U74 ; P1_R1375_U192
g9962 nand P1_R1375_U187 P1_R1375_U107 ; P1_R1375_U193
g9963 nand P1_U3509 P1_R1375_U73 ; P1_R1375_U194
g9964 nand P1_R1375_U194 P1_R1375_U193 ; P1_R1375_U195
g9965 nand P1_R1375_U110 P1_R1375_U133 ; P1_R1375_U196
g9966 nand P1_U4014 P1_R1375_U33 ; P1_R1375_U197
g9967 nand P1_U4013 P1_R1375_U30 ; P1_R1375_U198
g9968 nand P1_U4017 P1_R1375_U116 ; P1_R1375_U199
g9969 nand P1_R1375_U19 P1_R1375_U116 ; P1_R1375_U200
g9970 nand P1_R1375_U11 P1_R1375_U202 ; P1_R1375_U201
g9971 nand P1_U3057 P1_R1375_U16 ; P1_R1375_U202
g9972 nand P1_R1375_U132 P1_R1375_U114 ; P1_R1375_U203
g9973 nand P1_R1375_U89 P1_R1375_U203 ; P1_R1375_U204
g9974 nand P1_R1375_U126 P1_R1375_U80 P1_R1375_U78 P1_R1375_U111 P1_R1375_U112 ; P1_R1375_U205
g9975 nand P1_U3051 P1_R1375_U22 ; P1_R1375_U206
g9976 nand P1_U4008 P1_R1375_U113 ; P1_R1375_U207
g9977 and P1_U3057 P1_R1352_U7 ; P1_R1352_U6
g9978 not P1_U3054 ; P1_R1352_U7
g9979 and P1_R1207_U184 P1_R1207_U201 ; P1_R1207_U6
g9980 and P1_R1207_U203 P1_R1207_U202 ; P1_R1207_U7
g9981 and P1_R1207_U179 P1_R1207_U240 ; P1_R1207_U8
g9982 and P1_R1207_U242 P1_R1207_U241 ; P1_R1207_U9
g9983 and P1_R1207_U259 P1_R1207_U258 ; P1_R1207_U10
g9984 and P1_R1207_U285 P1_R1207_U284 ; P1_R1207_U11
g9985 and P1_R1207_U383 P1_R1207_U382 ; P1_R1207_U12
g9986 nand P1_R1207_U340 P1_R1207_U343 ; P1_R1207_U13
g9987 nand P1_R1207_U329 P1_R1207_U332 ; P1_R1207_U14
g9988 nand P1_R1207_U318 P1_R1207_U321 ; P1_R1207_U15
g9989 nand P1_R1207_U310 P1_R1207_U312 ; P1_R1207_U16
g9990 nand P1_R1207_U156 P1_R1207_U175 P1_R1207_U348 ; P1_R1207_U17
g9991 nand P1_R1207_U236 P1_R1207_U238 ; P1_R1207_U18
g9992 nand P1_R1207_U228 P1_R1207_U231 ; P1_R1207_U19
g9993 nand P1_R1207_U220 P1_R1207_U222 ; P1_R1207_U20
g9994 nand P1_R1207_U25 P1_R1207_U346 ; P1_R1207_U21
g9995 not P1_U3474 ; P1_R1207_U22
g9996 not P1_U3459 ; P1_R1207_U23
g9997 not P1_U3451 ; P1_R1207_U24
g9998 nand P1_U3451 P1_R1207_U93 ; P1_R1207_U25
g9999 not P1_U3076 ; P1_R1207_U26
g10000 not P1_U3462 ; P1_R1207_U27
g10001 not P1_U3066 ; P1_R1207_U28
g10002 nand P1_U3066 P1_R1207_U23 ; P1_R1207_U29
g10003 not P1_U3062 ; P1_R1207_U30
g10004 not P1_U3471 ; P1_R1207_U31
g10005 not P1_U3468 ; P1_R1207_U32
g10006 not P1_U3465 ; P1_R1207_U33
g10007 not P1_U3069 ; P1_R1207_U34
g10008 not P1_U3065 ; P1_R1207_U35
g10009 not P1_U3058 ; P1_R1207_U36
g10010 nand P1_U3058 P1_R1207_U33 ; P1_R1207_U37
g10011 not P1_U3477 ; P1_R1207_U38
g10012 not P1_U3068 ; P1_R1207_U39
g10013 nand P1_U3068 P1_R1207_U22 ; P1_R1207_U40
g10014 not P1_U3082 ; P1_R1207_U41
g10015 not P1_U3480 ; P1_R1207_U42
g10016 not P1_U3081 ; P1_R1207_U43
g10017 nand P1_R1207_U209 P1_R1207_U208 ; P1_R1207_U44
g10018 nand P1_R1207_U37 P1_R1207_U224 ; P1_R1207_U45
g10019 nand P1_R1207_U193 P1_R1207_U192 ; P1_R1207_U46
g10020 not P1_U4009 ; P1_R1207_U47
g10021 not P1_U4013 ; P1_R1207_U48
g10022 not P1_U3498 ; P1_R1207_U49
g10023 not P1_U3486 ; P1_R1207_U50
g10024 not P1_U3483 ; P1_R1207_U51
g10025 not P1_U3061 ; P1_R1207_U52
g10026 not P1_U3060 ; P1_R1207_U53
g10027 nand P1_U3081 P1_R1207_U42 ; P1_R1207_U54
g10028 not P1_U3489 ; P1_R1207_U55
g10029 not P1_U3070 ; P1_R1207_U56
g10030 not P1_U3492 ; P1_R1207_U57
g10031 not P1_U3078 ; P1_R1207_U58
g10032 not P1_U3501 ; P1_R1207_U59
g10033 not P1_U3495 ; P1_R1207_U60
g10034 not P1_U3071 ; P1_R1207_U61
g10035 not P1_U3072 ; P1_R1207_U62
g10036 not P1_U3077 ; P1_R1207_U63
g10037 nand P1_U3077 P1_R1207_U60 ; P1_R1207_U64
g10038 not P1_U3504 ; P1_R1207_U65
g10039 not P1_U3067 ; P1_R1207_U66
g10040 nand P1_R1207_U269 P1_R1207_U268 ; P1_R1207_U67
g10041 not P1_U3080 ; P1_R1207_U68
g10042 not P1_U3509 ; P1_R1207_U69
g10043 not P1_U3079 ; P1_R1207_U70
g10044 not P1_U4015 ; P1_R1207_U71
g10045 not P1_U3074 ; P1_R1207_U72
g10046 not P1_U4012 ; P1_R1207_U73
g10047 not P1_U4014 ; P1_R1207_U74
g10048 not P1_U3064 ; P1_R1207_U75
g10049 not P1_U3059 ; P1_R1207_U76
g10050 not P1_U3073 ; P1_R1207_U77
g10051 nand P1_U3073 P1_R1207_U74 ; P1_R1207_U78
g10052 not P1_U4011 ; P1_R1207_U79
g10053 not P1_U3063 ; P1_R1207_U80
g10054 not P1_U4010 ; P1_R1207_U81
g10055 not P1_U3056 ; P1_R1207_U82
g10056 not P1_U4008 ; P1_R1207_U83
g10057 not P1_U3055 ; P1_R1207_U84
g10058 nand P1_U3055 P1_R1207_U47 ; P1_R1207_U85
g10059 not P1_U3051 ; P1_R1207_U86
g10060 not P1_U4007 ; P1_R1207_U87
g10061 not P1_U3052 ; P1_R1207_U88
g10062 nand P1_R1207_U299 P1_R1207_U298 ; P1_R1207_U89
g10063 nand P1_R1207_U78 P1_R1207_U314 ; P1_R1207_U90
g10064 nand P1_R1207_U64 P1_R1207_U325 ; P1_R1207_U91
g10065 nand P1_R1207_U54 P1_R1207_U336 ; P1_R1207_U92
g10066 not P1_U3075 ; P1_R1207_U93
g10067 nand P1_R1207_U393 P1_R1207_U392 ; P1_R1207_U94
g10068 nand P1_R1207_U407 P1_R1207_U406 ; P1_R1207_U95
g10069 nand P1_R1207_U412 P1_R1207_U411 ; P1_R1207_U96
g10070 nand P1_R1207_U428 P1_R1207_U427 ; P1_R1207_U97
g10071 nand P1_R1207_U433 P1_R1207_U432 ; P1_R1207_U98
g10072 nand P1_R1207_U438 P1_R1207_U437 ; P1_R1207_U99
g10073 nand P1_R1207_U443 P1_R1207_U442 ; P1_R1207_U100
g10074 nand P1_R1207_U448 P1_R1207_U447 ; P1_R1207_U101
g10075 nand P1_R1207_U464 P1_R1207_U463 ; P1_R1207_U102
g10076 nand P1_R1207_U469 P1_R1207_U468 ; P1_R1207_U103
g10077 nand P1_R1207_U352 P1_R1207_U351 ; P1_R1207_U104
g10078 nand P1_R1207_U361 P1_R1207_U360 ; P1_R1207_U105
g10079 nand P1_R1207_U368 P1_R1207_U367 ; P1_R1207_U106
g10080 nand P1_R1207_U372 P1_R1207_U371 ; P1_R1207_U107
g10081 nand P1_R1207_U381 P1_R1207_U380 ; P1_R1207_U108
g10082 nand P1_R1207_U402 P1_R1207_U401 ; P1_R1207_U109
g10083 nand P1_R1207_U419 P1_R1207_U418 ; P1_R1207_U110
g10084 nand P1_R1207_U423 P1_R1207_U422 ; P1_R1207_U111
g10085 nand P1_R1207_U455 P1_R1207_U454 ; P1_R1207_U112
g10086 nand P1_R1207_U459 P1_R1207_U458 ; P1_R1207_U113
g10087 nand P1_R1207_U476 P1_R1207_U475 ; P1_R1207_U114
g10088 and P1_R1207_U195 P1_R1207_U183 ; P1_R1207_U115
g10089 and P1_R1207_U198 P1_R1207_U199 ; P1_R1207_U116
g10090 and P1_R1207_U211 P1_R1207_U185 ; P1_R1207_U117
g10091 and P1_R1207_U214 P1_R1207_U215 ; P1_R1207_U118
g10092 and P1_R1207_U354 P1_R1207_U353 P1_R1207_U40 ; P1_R1207_U119
g10093 and P1_R1207_U357 P1_R1207_U185 ; P1_R1207_U120
g10094 and P1_R1207_U230 P1_R1207_U7 ; P1_R1207_U121
g10095 and P1_R1207_U364 P1_R1207_U184 ; P1_R1207_U122
g10096 and P1_R1207_U374 P1_R1207_U373 P1_R1207_U29 ; P1_R1207_U123
g10097 and P1_R1207_U377 P1_R1207_U183 ; P1_R1207_U124
g10098 and P1_R1207_U217 P1_R1207_U8 ; P1_R1207_U125
g10099 and P1_R1207_U262 P1_R1207_U180 ; P1_R1207_U126
g10100 and P1_R1207_U288 P1_R1207_U181 ; P1_R1207_U127
g10101 and P1_R1207_U304 P1_R1207_U305 ; P1_R1207_U128
g10102 and P1_R1207_U307 P1_R1207_U386 ; P1_R1207_U129
g10103 and P1_R1207_U305 P1_R1207_U304 P1_R1207_U308 ; P1_R1207_U130
g10104 nand P1_R1207_U390 P1_R1207_U389 ; P1_R1207_U131
g10105 and P1_R1207_U395 P1_R1207_U394 P1_R1207_U85 ; P1_R1207_U132
g10106 and P1_R1207_U398 P1_R1207_U182 ; P1_R1207_U133
g10107 nand P1_R1207_U404 P1_R1207_U403 ; P1_R1207_U134
g10108 nand P1_R1207_U409 P1_R1207_U408 ; P1_R1207_U135
g10109 and P1_R1207_U415 P1_R1207_U181 ; P1_R1207_U136
g10110 nand P1_R1207_U425 P1_R1207_U424 ; P1_R1207_U137
g10111 nand P1_R1207_U430 P1_R1207_U429 ; P1_R1207_U138
g10112 nand P1_R1207_U435 P1_R1207_U434 ; P1_R1207_U139
g10113 nand P1_R1207_U440 P1_R1207_U439 ; P1_R1207_U140
g10114 nand P1_R1207_U445 P1_R1207_U444 ; P1_R1207_U141
g10115 and P1_R1207_U451 P1_R1207_U180 ; P1_R1207_U142
g10116 nand P1_R1207_U461 P1_R1207_U460 ; P1_R1207_U143
g10117 nand P1_R1207_U466 P1_R1207_U465 ; P1_R1207_U144
g10118 and P1_R1207_U342 P1_R1207_U9 ; P1_R1207_U145
g10119 and P1_R1207_U472 P1_R1207_U179 ; P1_R1207_U146
g10120 and P1_R1207_U350 P1_R1207_U349 ; P1_R1207_U147
g10121 nand P1_R1207_U118 P1_R1207_U212 ; P1_R1207_U148
g10122 and P1_R1207_U359 P1_R1207_U358 ; P1_R1207_U149
g10123 and P1_R1207_U366 P1_R1207_U365 ; P1_R1207_U150
g10124 and P1_R1207_U370 P1_R1207_U369 ; P1_R1207_U151
g10125 nand P1_R1207_U116 P1_R1207_U196 ; P1_R1207_U152
g10126 and P1_R1207_U379 P1_R1207_U378 ; P1_R1207_U153
g10127 not P1_U4018 ; P1_R1207_U154
g10128 not P1_U3053 ; P1_R1207_U155
g10129 and P1_R1207_U388 P1_R1207_U387 ; P1_R1207_U156
g10130 nand P1_R1207_U128 P1_R1207_U302 ; P1_R1207_U157
g10131 and P1_R1207_U400 P1_R1207_U399 ; P1_R1207_U158
g10132 nand P1_R1207_U295 P1_R1207_U294 ; P1_R1207_U159
g10133 nand P1_R1207_U291 P1_R1207_U290 ; P1_R1207_U160
g10134 and P1_R1207_U417 P1_R1207_U416 ; P1_R1207_U161
g10135 and P1_R1207_U421 P1_R1207_U420 ; P1_R1207_U162
g10136 nand P1_R1207_U281 P1_R1207_U280 ; P1_R1207_U163
g10137 nand P1_R1207_U277 P1_R1207_U276 ; P1_R1207_U164
g10138 not P1_U3456 ; P1_R1207_U165
g10139 nand P1_R1207_U273 P1_R1207_U272 ; P1_R1207_U166
g10140 not P1_U3507 ; P1_R1207_U167
g10141 nand P1_R1207_U265 P1_R1207_U264 ; P1_R1207_U168
g10142 and P1_R1207_U453 P1_R1207_U452 ; P1_R1207_U169
g10143 and P1_R1207_U457 P1_R1207_U456 ; P1_R1207_U170
g10144 nand P1_R1207_U255 P1_R1207_U254 ; P1_R1207_U171
g10145 nand P1_R1207_U251 P1_R1207_U250 ; P1_R1207_U172
g10146 nand P1_R1207_U247 P1_R1207_U246 ; P1_R1207_U173
g10147 and P1_R1207_U474 P1_R1207_U473 ; P1_R1207_U174
g10148 nand P1_R1207_U129 P1_R1207_U157 ; P1_R1207_U175
g10149 not P1_R1207_U85 ; P1_R1207_U176
g10150 not P1_R1207_U29 ; P1_R1207_U177
g10151 not P1_R1207_U40 ; P1_R1207_U178
g10152 nand P1_U3483 P1_R1207_U53 ; P1_R1207_U179
g10153 nand P1_U3498 P1_R1207_U62 ; P1_R1207_U180
g10154 nand P1_U4013 P1_R1207_U76 ; P1_R1207_U181
g10155 nand P1_U4009 P1_R1207_U84 ; P1_R1207_U182
g10156 nand P1_U3459 P1_R1207_U28 ; P1_R1207_U183
g10157 nand P1_U3468 P1_R1207_U35 ; P1_R1207_U184
g10158 nand P1_U3474 P1_R1207_U39 ; P1_R1207_U185
g10159 not P1_R1207_U64 ; P1_R1207_U186
g10160 not P1_R1207_U78 ; P1_R1207_U187
g10161 not P1_R1207_U37 ; P1_R1207_U188
g10162 not P1_R1207_U54 ; P1_R1207_U189
g10163 not P1_R1207_U25 ; P1_R1207_U190
g10164 nand P1_R1207_U190 P1_R1207_U26 ; P1_R1207_U191
g10165 nand P1_R1207_U191 P1_R1207_U165 ; P1_R1207_U192
g10166 nand P1_U3076 P1_R1207_U25 ; P1_R1207_U193
g10167 not P1_R1207_U46 ; P1_R1207_U194
g10168 nand P1_U3462 P1_R1207_U30 ; P1_R1207_U195
g10169 nand P1_R1207_U115 P1_R1207_U46 ; P1_R1207_U196
g10170 nand P1_R1207_U30 P1_R1207_U29 ; P1_R1207_U197
g10171 nand P1_R1207_U197 P1_R1207_U27 ; P1_R1207_U198
g10172 nand P1_U3062 P1_R1207_U177 ; P1_R1207_U199
g10173 not P1_R1207_U152 ; P1_R1207_U200
g10174 nand P1_U3471 P1_R1207_U34 ; P1_R1207_U201
g10175 nand P1_U3069 P1_R1207_U31 ; P1_R1207_U202
g10176 nand P1_U3065 P1_R1207_U32 ; P1_R1207_U203
g10177 nand P1_R1207_U188 P1_R1207_U6 ; P1_R1207_U204
g10178 nand P1_R1207_U7 P1_R1207_U204 ; P1_R1207_U205
g10179 nand P1_U3465 P1_R1207_U36 ; P1_R1207_U206
g10180 nand P1_U3471 P1_R1207_U34 ; P1_R1207_U207
g10181 nand P1_R1207_U206 P1_R1207_U152 P1_R1207_U6 ; P1_R1207_U208
g10182 nand P1_R1207_U207 P1_R1207_U205 ; P1_R1207_U209
g10183 not P1_R1207_U44 ; P1_R1207_U210
g10184 nand P1_U3477 P1_R1207_U41 ; P1_R1207_U211
g10185 nand P1_R1207_U117 P1_R1207_U44 ; P1_R1207_U212
g10186 nand P1_R1207_U41 P1_R1207_U40 ; P1_R1207_U213
g10187 nand P1_R1207_U213 P1_R1207_U38 ; P1_R1207_U214
g10188 nand P1_U3082 P1_R1207_U178 ; P1_R1207_U215
g10189 not P1_R1207_U148 ; P1_R1207_U216
g10190 nand P1_U3480 P1_R1207_U43 ; P1_R1207_U217
g10191 nand P1_R1207_U217 P1_R1207_U54 ; P1_R1207_U218
g10192 nand P1_R1207_U210 P1_R1207_U40 ; P1_R1207_U219
g10193 nand P1_R1207_U120 P1_R1207_U219 ; P1_R1207_U220
g10194 nand P1_R1207_U44 P1_R1207_U185 ; P1_R1207_U221
g10195 nand P1_R1207_U119 P1_R1207_U221 ; P1_R1207_U222
g10196 nand P1_R1207_U40 P1_R1207_U185 ; P1_R1207_U223
g10197 nand P1_R1207_U206 P1_R1207_U152 ; P1_R1207_U224
g10198 not P1_R1207_U45 ; P1_R1207_U225
g10199 nand P1_U3065 P1_R1207_U32 ; P1_R1207_U226
g10200 nand P1_R1207_U225 P1_R1207_U226 ; P1_R1207_U227
g10201 nand P1_R1207_U122 P1_R1207_U227 ; P1_R1207_U228
g10202 nand P1_R1207_U45 P1_R1207_U184 ; P1_R1207_U229
g10203 nand P1_U3471 P1_R1207_U34 ; P1_R1207_U230
g10204 nand P1_R1207_U121 P1_R1207_U229 ; P1_R1207_U231
g10205 nand P1_U3065 P1_R1207_U32 ; P1_R1207_U232
g10206 nand P1_R1207_U184 P1_R1207_U232 ; P1_R1207_U233
g10207 nand P1_R1207_U206 P1_R1207_U37 ; P1_R1207_U234
g10208 nand P1_R1207_U194 P1_R1207_U29 ; P1_R1207_U235
g10209 nand P1_R1207_U124 P1_R1207_U235 ; P1_R1207_U236
g10210 nand P1_R1207_U46 P1_R1207_U183 ; P1_R1207_U237
g10211 nand P1_R1207_U123 P1_R1207_U237 ; P1_R1207_U238
g10212 nand P1_R1207_U29 P1_R1207_U183 ; P1_R1207_U239
g10213 nand P1_U3486 P1_R1207_U52 ; P1_R1207_U240
g10214 nand P1_U3061 P1_R1207_U50 ; P1_R1207_U241
g10215 nand P1_U3060 P1_R1207_U51 ; P1_R1207_U242
g10216 nand P1_R1207_U189 P1_R1207_U8 ; P1_R1207_U243
g10217 nand P1_R1207_U9 P1_R1207_U243 ; P1_R1207_U244
g10218 nand P1_U3486 P1_R1207_U52 ; P1_R1207_U245
g10219 nand P1_R1207_U125 P1_R1207_U148 ; P1_R1207_U246
g10220 nand P1_R1207_U245 P1_R1207_U244 ; P1_R1207_U247
g10221 not P1_R1207_U173 ; P1_R1207_U248
g10222 nand P1_U3489 P1_R1207_U56 ; P1_R1207_U249
g10223 nand P1_R1207_U249 P1_R1207_U173 ; P1_R1207_U250
g10224 nand P1_U3070 P1_R1207_U55 ; P1_R1207_U251
g10225 not P1_R1207_U172 ; P1_R1207_U252
g10226 nand P1_U3492 P1_R1207_U58 ; P1_R1207_U253
g10227 nand P1_R1207_U253 P1_R1207_U172 ; P1_R1207_U254
g10228 nand P1_U3078 P1_R1207_U57 ; P1_R1207_U255
g10229 not P1_R1207_U171 ; P1_R1207_U256
g10230 nand P1_U3501 P1_R1207_U61 ; P1_R1207_U257
g10231 nand P1_U3071 P1_R1207_U59 ; P1_R1207_U258
g10232 nand P1_U3072 P1_R1207_U49 ; P1_R1207_U259
g10233 nand P1_R1207_U186 P1_R1207_U180 ; P1_R1207_U260
g10234 nand P1_R1207_U10 P1_R1207_U260 ; P1_R1207_U261
g10235 nand P1_U3495 P1_R1207_U63 ; P1_R1207_U262
g10236 nand P1_U3501 P1_R1207_U61 ; P1_R1207_U263
g10237 nand P1_R1207_U171 P1_R1207_U126 P1_R1207_U257 ; P1_R1207_U264
g10238 nand P1_R1207_U263 P1_R1207_U261 ; P1_R1207_U265
g10239 not P1_R1207_U168 ; P1_R1207_U266
g10240 nand P1_U3504 P1_R1207_U66 ; P1_R1207_U267
g10241 nand P1_R1207_U267 P1_R1207_U168 ; P1_R1207_U268
g10242 nand P1_U3067 P1_R1207_U65 ; P1_R1207_U269
g10243 not P1_R1207_U67 ; P1_R1207_U270
g10244 nand P1_R1207_U270 P1_R1207_U68 ; P1_R1207_U271
g10245 nand P1_R1207_U271 P1_R1207_U167 ; P1_R1207_U272
g10246 nand P1_U3080 P1_R1207_U67 ; P1_R1207_U273
g10247 not P1_R1207_U166 ; P1_R1207_U274
g10248 nand P1_U3509 P1_R1207_U70 ; P1_R1207_U275
g10249 nand P1_R1207_U275 P1_R1207_U166 ; P1_R1207_U276
g10250 nand P1_U3079 P1_R1207_U69 ; P1_R1207_U277
g10251 not P1_R1207_U164 ; P1_R1207_U278
g10252 nand P1_U4015 P1_R1207_U72 ; P1_R1207_U279
g10253 nand P1_R1207_U279 P1_R1207_U164 ; P1_R1207_U280
g10254 nand P1_U3074 P1_R1207_U71 ; P1_R1207_U281
g10255 not P1_R1207_U163 ; P1_R1207_U282
g10256 nand P1_U4012 P1_R1207_U75 ; P1_R1207_U283
g10257 nand P1_U3064 P1_R1207_U73 ; P1_R1207_U284
g10258 nand P1_U3059 P1_R1207_U48 ; P1_R1207_U285
g10259 nand P1_R1207_U187 P1_R1207_U181 ; P1_R1207_U286
g10260 nand P1_R1207_U11 P1_R1207_U286 ; P1_R1207_U287
g10261 nand P1_U4014 P1_R1207_U77 ; P1_R1207_U288
g10262 nand P1_U4012 P1_R1207_U75 ; P1_R1207_U289
g10263 nand P1_R1207_U163 P1_R1207_U127 P1_R1207_U283 ; P1_R1207_U290
g10264 nand P1_R1207_U289 P1_R1207_U287 ; P1_R1207_U291
g10265 not P1_R1207_U160 ; P1_R1207_U292
g10266 nand P1_U4011 P1_R1207_U80 ; P1_R1207_U293
g10267 nand P1_R1207_U293 P1_R1207_U160 ; P1_R1207_U294
g10268 nand P1_U3063 P1_R1207_U79 ; P1_R1207_U295
g10269 not P1_R1207_U159 ; P1_R1207_U296
g10270 nand P1_U4010 P1_R1207_U82 ; P1_R1207_U297
g10271 nand P1_R1207_U297 P1_R1207_U159 ; P1_R1207_U298
g10272 nand P1_U3056 P1_R1207_U81 ; P1_R1207_U299
g10273 not P1_R1207_U89 ; P1_R1207_U300
g10274 nand P1_U4008 P1_R1207_U86 ; P1_R1207_U301
g10275 nand P1_R1207_U89 P1_R1207_U182 P1_R1207_U301 ; P1_R1207_U302
g10276 nand P1_R1207_U86 P1_R1207_U85 ; P1_R1207_U303
g10277 nand P1_R1207_U303 P1_R1207_U83 ; P1_R1207_U304
g10278 nand P1_U3051 P1_R1207_U176 ; P1_R1207_U305
g10279 not P1_R1207_U157 ; P1_R1207_U306
g10280 nand P1_U4007 P1_R1207_U88 ; P1_R1207_U307
g10281 nand P1_U3052 P1_R1207_U87 ; P1_R1207_U308
g10282 nand P1_R1207_U300 P1_R1207_U85 ; P1_R1207_U309
g10283 nand P1_R1207_U133 P1_R1207_U309 ; P1_R1207_U310
g10284 nand P1_R1207_U89 P1_R1207_U182 ; P1_R1207_U311
g10285 nand P1_R1207_U132 P1_R1207_U311 ; P1_R1207_U312
g10286 nand P1_R1207_U85 P1_R1207_U182 ; P1_R1207_U313
g10287 nand P1_R1207_U288 P1_R1207_U163 ; P1_R1207_U314
g10288 not P1_R1207_U90 ; P1_R1207_U315
g10289 nand P1_U3059 P1_R1207_U48 ; P1_R1207_U316
g10290 nand P1_R1207_U315 P1_R1207_U316 ; P1_R1207_U317
g10291 nand P1_R1207_U136 P1_R1207_U317 ; P1_R1207_U318
g10292 nand P1_R1207_U90 P1_R1207_U181 ; P1_R1207_U319
g10293 nand P1_U4012 P1_R1207_U75 ; P1_R1207_U320
g10294 nand P1_R1207_U320 P1_R1207_U319 P1_R1207_U11 ; P1_R1207_U321
g10295 nand P1_U3059 P1_R1207_U48 ; P1_R1207_U322
g10296 nand P1_R1207_U181 P1_R1207_U322 ; P1_R1207_U323
g10297 nand P1_R1207_U288 P1_R1207_U78 ; P1_R1207_U324
g10298 nand P1_R1207_U262 P1_R1207_U171 ; P1_R1207_U325
g10299 not P1_R1207_U91 ; P1_R1207_U326
g10300 nand P1_U3072 P1_R1207_U49 ; P1_R1207_U327
g10301 nand P1_R1207_U326 P1_R1207_U327 ; P1_R1207_U328
g10302 nand P1_R1207_U142 P1_R1207_U328 ; P1_R1207_U329
g10303 nand P1_R1207_U91 P1_R1207_U180 ; P1_R1207_U330
g10304 nand P1_U3501 P1_R1207_U61 ; P1_R1207_U331
g10305 nand P1_R1207_U331 P1_R1207_U330 P1_R1207_U10 ; P1_R1207_U332
g10306 nand P1_U3072 P1_R1207_U49 ; P1_R1207_U333
g10307 nand P1_R1207_U180 P1_R1207_U333 ; P1_R1207_U334
g10308 nand P1_R1207_U262 P1_R1207_U64 ; P1_R1207_U335
g10309 nand P1_R1207_U217 P1_R1207_U148 ; P1_R1207_U336
g10310 not P1_R1207_U92 ; P1_R1207_U337
g10311 nand P1_U3060 P1_R1207_U51 ; P1_R1207_U338
g10312 nand P1_R1207_U337 P1_R1207_U338 ; P1_R1207_U339
g10313 nand P1_R1207_U146 P1_R1207_U339 ; P1_R1207_U340
g10314 nand P1_R1207_U92 P1_R1207_U179 ; P1_R1207_U341
g10315 nand P1_U3486 P1_R1207_U52 ; P1_R1207_U342
g10316 nand P1_R1207_U145 P1_R1207_U341 ; P1_R1207_U343
g10317 nand P1_U3060 P1_R1207_U51 ; P1_R1207_U344
g10318 nand P1_R1207_U179 P1_R1207_U344 ; P1_R1207_U345
g10319 nand P1_U3075 P1_R1207_U24 ; P1_R1207_U346
g10320 nand P1_R1207_U89 P1_R1207_U182 P1_R1207_U301 ; P1_R1207_U347
g10321 nand P1_R1207_U12 P1_R1207_U347 P1_R1207_U130 ; P1_R1207_U348
g10322 nand P1_U3480 P1_R1207_U43 ; P1_R1207_U349
g10323 nand P1_U3081 P1_R1207_U42 ; P1_R1207_U350
g10324 nand P1_R1207_U218 P1_R1207_U148 ; P1_R1207_U351
g10325 nand P1_R1207_U216 P1_R1207_U147 ; P1_R1207_U352
g10326 nand P1_U3477 P1_R1207_U41 ; P1_R1207_U353
g10327 nand P1_U3082 P1_R1207_U38 ; P1_R1207_U354
g10328 nand P1_U3477 P1_R1207_U41 ; P1_R1207_U355
g10329 nand P1_U3082 P1_R1207_U38 ; P1_R1207_U356
g10330 nand P1_R1207_U356 P1_R1207_U355 ; P1_R1207_U357
g10331 nand P1_U3474 P1_R1207_U39 ; P1_R1207_U358
g10332 nand P1_U3068 P1_R1207_U22 ; P1_R1207_U359
g10333 nand P1_R1207_U223 P1_R1207_U44 ; P1_R1207_U360
g10334 nand P1_R1207_U149 P1_R1207_U210 ; P1_R1207_U361
g10335 nand P1_U3471 P1_R1207_U34 ; P1_R1207_U362
g10336 nand P1_U3069 P1_R1207_U31 ; P1_R1207_U363
g10337 nand P1_R1207_U363 P1_R1207_U362 ; P1_R1207_U364
g10338 nand P1_U3468 P1_R1207_U35 ; P1_R1207_U365
g10339 nand P1_U3065 P1_R1207_U32 ; P1_R1207_U366
g10340 nand P1_R1207_U233 P1_R1207_U45 ; P1_R1207_U367
g10341 nand P1_R1207_U150 P1_R1207_U225 ; P1_R1207_U368
g10342 nand P1_U3465 P1_R1207_U36 ; P1_R1207_U369
g10343 nand P1_U3058 P1_R1207_U33 ; P1_R1207_U370
g10344 nand P1_R1207_U234 P1_R1207_U152 ; P1_R1207_U371
g10345 nand P1_R1207_U200 P1_R1207_U151 ; P1_R1207_U372
g10346 nand P1_U3462 P1_R1207_U30 ; P1_R1207_U373
g10347 nand P1_U3062 P1_R1207_U27 ; P1_R1207_U374
g10348 nand P1_U3462 P1_R1207_U30 ; P1_R1207_U375
g10349 nand P1_U3062 P1_R1207_U27 ; P1_R1207_U376
g10350 nand P1_R1207_U376 P1_R1207_U375 ; P1_R1207_U377
g10351 nand P1_U3459 P1_R1207_U28 ; P1_R1207_U378
g10352 nand P1_U3066 P1_R1207_U23 ; P1_R1207_U379
g10353 nand P1_R1207_U239 P1_R1207_U46 ; P1_R1207_U380
g10354 nand P1_R1207_U153 P1_R1207_U194 ; P1_R1207_U381
g10355 nand P1_U4018 P1_R1207_U155 ; P1_R1207_U382
g10356 nand P1_U3053 P1_R1207_U154 ; P1_R1207_U383
g10357 nand P1_U4018 P1_R1207_U155 ; P1_R1207_U384
g10358 nand P1_U3053 P1_R1207_U154 ; P1_R1207_U385
g10359 nand P1_R1207_U385 P1_R1207_U384 ; P1_R1207_U386
g10360 nand P1_U3052 P1_R1207_U386 P1_R1207_U87 ; P1_R1207_U387
g10361 nand P1_R1207_U12 P1_R1207_U88 P1_U4007 ; P1_R1207_U388
g10362 nand P1_U4007 P1_R1207_U88 ; P1_R1207_U389
g10363 nand P1_U3052 P1_R1207_U87 ; P1_R1207_U390
g10364 not P1_R1207_U131 ; P1_R1207_U391
g10365 nand P1_R1207_U306 P1_R1207_U391 ; P1_R1207_U392
g10366 nand P1_R1207_U131 P1_R1207_U157 ; P1_R1207_U393
g10367 nand P1_U4008 P1_R1207_U86 ; P1_R1207_U394
g10368 nand P1_U3051 P1_R1207_U83 ; P1_R1207_U395
g10369 nand P1_U4008 P1_R1207_U86 ; P1_R1207_U396
g10370 nand P1_U3051 P1_R1207_U83 ; P1_R1207_U397
g10371 nand P1_R1207_U397 P1_R1207_U396 ; P1_R1207_U398
g10372 nand P1_U4009 P1_R1207_U84 ; P1_R1207_U399
g10373 nand P1_U3055 P1_R1207_U47 ; P1_R1207_U400
g10374 nand P1_R1207_U313 P1_R1207_U89 ; P1_R1207_U401
g10375 nand P1_R1207_U158 P1_R1207_U300 ; P1_R1207_U402
g10376 nand P1_U4010 P1_R1207_U82 ; P1_R1207_U403
g10377 nand P1_U3056 P1_R1207_U81 ; P1_R1207_U404
g10378 not P1_R1207_U134 ; P1_R1207_U405
g10379 nand P1_R1207_U296 P1_R1207_U405 ; P1_R1207_U406
g10380 nand P1_R1207_U134 P1_R1207_U159 ; P1_R1207_U407
g10381 nand P1_U4011 P1_R1207_U80 ; P1_R1207_U408
g10382 nand P1_U3063 P1_R1207_U79 ; P1_R1207_U409
g10383 not P1_R1207_U135 ; P1_R1207_U410
g10384 nand P1_R1207_U292 P1_R1207_U410 ; P1_R1207_U411
g10385 nand P1_R1207_U135 P1_R1207_U160 ; P1_R1207_U412
g10386 nand P1_U4012 P1_R1207_U75 ; P1_R1207_U413
g10387 nand P1_U3064 P1_R1207_U73 ; P1_R1207_U414
g10388 nand P1_R1207_U414 P1_R1207_U413 ; P1_R1207_U415
g10389 nand P1_U4013 P1_R1207_U76 ; P1_R1207_U416
g10390 nand P1_U3059 P1_R1207_U48 ; P1_R1207_U417
g10391 nand P1_R1207_U323 P1_R1207_U90 ; P1_R1207_U418
g10392 nand P1_R1207_U161 P1_R1207_U315 ; P1_R1207_U419
g10393 nand P1_U4014 P1_R1207_U77 ; P1_R1207_U420
g10394 nand P1_U3073 P1_R1207_U74 ; P1_R1207_U421
g10395 nand P1_R1207_U324 P1_R1207_U163 ; P1_R1207_U422
g10396 nand P1_R1207_U282 P1_R1207_U162 ; P1_R1207_U423
g10397 nand P1_U4015 P1_R1207_U72 ; P1_R1207_U424
g10398 nand P1_U3074 P1_R1207_U71 ; P1_R1207_U425
g10399 not P1_R1207_U137 ; P1_R1207_U426
g10400 nand P1_R1207_U278 P1_R1207_U426 ; P1_R1207_U427
g10401 nand P1_R1207_U137 P1_R1207_U164 ; P1_R1207_U428
g10402 nand P1_U3456 P1_R1207_U26 ; P1_R1207_U429
g10403 nand P1_U3076 P1_R1207_U165 ; P1_R1207_U430
g10404 not P1_R1207_U138 ; P1_R1207_U431
g10405 nand P1_R1207_U431 P1_R1207_U190 ; P1_R1207_U432
g10406 nand P1_R1207_U138 P1_R1207_U25 ; P1_R1207_U433
g10407 nand P1_U3509 P1_R1207_U70 ; P1_R1207_U434
g10408 nand P1_U3079 P1_R1207_U69 ; P1_R1207_U435
g10409 not P1_R1207_U139 ; P1_R1207_U436
g10410 nand P1_R1207_U274 P1_R1207_U436 ; P1_R1207_U437
g10411 nand P1_R1207_U139 P1_R1207_U166 ; P1_R1207_U438
g10412 nand P1_U3507 P1_R1207_U68 ; P1_R1207_U439
g10413 nand P1_U3080 P1_R1207_U167 ; P1_R1207_U440
g10414 not P1_R1207_U140 ; P1_R1207_U441
g10415 nand P1_R1207_U441 P1_R1207_U270 ; P1_R1207_U442
g10416 nand P1_R1207_U140 P1_R1207_U67 ; P1_R1207_U443
g10417 nand P1_U3504 P1_R1207_U66 ; P1_R1207_U444
g10418 nand P1_U3067 P1_R1207_U65 ; P1_R1207_U445
g10419 not P1_R1207_U141 ; P1_R1207_U446
g10420 nand P1_R1207_U266 P1_R1207_U446 ; P1_R1207_U447
g10421 nand P1_R1207_U141 P1_R1207_U168 ; P1_R1207_U448
g10422 nand P1_U3501 P1_R1207_U61 ; P1_R1207_U449
g10423 nand P1_U3071 P1_R1207_U59 ; P1_R1207_U450
g10424 nand P1_R1207_U450 P1_R1207_U449 ; P1_R1207_U451
g10425 nand P1_U3498 P1_R1207_U62 ; P1_R1207_U452
g10426 nand P1_U3072 P1_R1207_U49 ; P1_R1207_U453
g10427 nand P1_R1207_U334 P1_R1207_U91 ; P1_R1207_U454
g10428 nand P1_R1207_U169 P1_R1207_U326 ; P1_R1207_U455
g10429 nand P1_U3495 P1_R1207_U63 ; P1_R1207_U456
g10430 nand P1_U3077 P1_R1207_U60 ; P1_R1207_U457
g10431 nand P1_R1207_U335 P1_R1207_U171 ; P1_R1207_U458
g10432 nand P1_R1207_U256 P1_R1207_U170 ; P1_R1207_U459
g10433 nand P1_U3492 P1_R1207_U58 ; P1_R1207_U460
g10434 nand P1_U3078 P1_R1207_U57 ; P1_R1207_U461
g10435 not P1_R1207_U143 ; P1_R1207_U462
g10436 nand P1_R1207_U252 P1_R1207_U462 ; P1_R1207_U463
g10437 nand P1_R1207_U143 P1_R1207_U172 ; P1_R1207_U464
g10438 nand P1_U3489 P1_R1207_U56 ; P1_R1207_U465
g10439 nand P1_U3070 P1_R1207_U55 ; P1_R1207_U466
g10440 not P1_R1207_U144 ; P1_R1207_U467
g10441 nand P1_R1207_U248 P1_R1207_U467 ; P1_R1207_U468
g10442 nand P1_R1207_U144 P1_R1207_U173 ; P1_R1207_U469
g10443 nand P1_U3486 P1_R1207_U52 ; P1_R1207_U470
g10444 nand P1_U3061 P1_R1207_U50 ; P1_R1207_U471
g10445 nand P1_R1207_U471 P1_R1207_U470 ; P1_R1207_U472
g10446 nand P1_U3483 P1_R1207_U53 ; P1_R1207_U473
g10447 nand P1_U3060 P1_R1207_U51 ; P1_R1207_U474
g10448 nand P1_R1207_U345 P1_R1207_U92 ; P1_R1207_U475
g10449 nand P1_R1207_U174 P1_R1207_U337 ; P1_R1207_U476
g10450 and P1_R1165_U210 P1_R1165_U209 ; P1_R1165_U4
g10451 and P1_R1165_U222 P1_R1165_U221 ; P1_R1165_U5
g10452 and P1_R1165_U253 P1_R1165_U252 ; P1_R1165_U6
g10453 and P1_R1165_U271 P1_R1165_U270 ; P1_R1165_U7
g10454 and P1_R1165_U283 P1_R1165_U282 ; P1_R1165_U8
g10455 and P1_R1165_U507 P1_R1165_U506 ; P1_R1165_U9
g10456 and P1_R1165_U339 P1_R1165_U336 ; P1_R1165_U10
g10457 and P1_R1165_U330 P1_R1165_U327 ; P1_R1165_U11
g10458 and P1_R1165_U323 P1_R1165_U320 ; P1_R1165_U12
g10459 and P1_R1165_U360 P1_R1165_U311 P1_R1165_U314 ; P1_R1165_U13
g10460 and P1_R1165_U245 P1_R1165_U242 ; P1_R1165_U14
g10461 and P1_R1165_U238 P1_R1165_U235 ; P1_R1165_U15
g10462 not P1_U3209 ; P1_R1165_U16
g10463 not P1_U3173 ; P1_R1165_U17
g10464 nand P1_U3173 P1_R1165_U58 ; P1_R1165_U18
g10465 not P1_U3172 ; P1_R1165_U19
g10466 not P1_U3175 ; P1_R1165_U20
g10467 not P1_U3177 ; P1_R1165_U21
g10468 nand P1_U3177 P1_R1165_U61 ; P1_R1165_U22
g10469 not P1_U3176 ; P1_R1165_U23
g10470 not P1_U3179 ; P1_R1165_U24
g10471 not P1_U3178 ; P1_R1165_U25
g10472 not P1_U3174 ; P1_R1165_U26
g10473 not P1_U3171 ; P1_R1165_U27
g10474 not P1_U3170 ; P1_R1165_U28
g10475 nand P1_R1165_U219 P1_R1165_U218 ; P1_R1165_U29
g10476 nand P1_R1165_U207 P1_R1165_U206 ; P1_R1165_U30
g10477 not P1_U3152 ; P1_R1165_U31
g10478 not P1_U3153 ; P1_R1165_U32
g10479 not P1_U3154 ; P1_R1165_U33
g10480 not P1_U3155 ; P1_R1165_U34
g10481 not P1_U3163 ; P1_R1165_U35
g10482 nand P1_U3163 P1_R1165_U71 ; P1_R1165_U36
g10483 not P1_U3162 ; P1_R1165_U37
g10484 not P1_U3169 ; P1_R1165_U38
g10485 not P1_U3167 ; P1_R1165_U39
g10486 not P1_U3168 ; P1_R1165_U40
g10487 nand P1_U3168 P1_R1165_U74 ; P1_R1165_U41
g10488 not P1_U3166 ; P1_R1165_U42
g10489 not P1_U3165 ; P1_R1165_U43
g10490 not P1_U3164 ; P1_R1165_U44
g10491 not P1_U3161 ; P1_R1165_U45
g10492 not P1_U3159 ; P1_R1165_U46
g10493 not P1_U3160 ; P1_R1165_U47
g10494 nand P1_U3160 P1_R1165_U80 ; P1_R1165_U48
g10495 not P1_U3158 ; P1_R1165_U49
g10496 not P1_U3157 ; P1_R1165_U50
g10497 not P1_U3156 ; P1_R1165_U51
g10498 nand P1_U3153 P1_R1165_U69 ; P1_R1165_U52
g10499 nand P1_R1165_U200 P1_R1165_U309 ; P1_R1165_U53
g10500 nand P1_R1165_U48 P1_R1165_U316 ; P1_R1165_U54
g10501 nand P1_R1165_U268 P1_R1165_U267 ; P1_R1165_U55
g10502 nand P1_R1165_U41 P1_R1165_U332 ; P1_R1165_U56
g10503 nand P1_R1165_U366 P1_R1165_U365 ; P1_R1165_U57
g10504 nand P1_R1165_U395 P1_R1165_U394 ; P1_R1165_U58
g10505 nand P1_R1165_U392 P1_R1165_U391 ; P1_R1165_U59
g10506 nand P1_R1165_U374 P1_R1165_U373 ; P1_R1165_U60
g10507 nand P1_R1165_U386 P1_R1165_U385 ; P1_R1165_U61
g10508 nand P1_R1165_U383 P1_R1165_U382 ; P1_R1165_U62
g10509 nand P1_R1165_U377 P1_R1165_U376 ; P1_R1165_U63
g10510 nand P1_R1165_U380 P1_R1165_U379 ; P1_R1165_U64
g10511 nand P1_R1165_U389 P1_R1165_U388 ; P1_R1165_U65
g10512 nand P1_R1165_U398 P1_R1165_U397 ; P1_R1165_U66
g10513 nand P1_R1165_U438 P1_R1165_U437 ; P1_R1165_U67
g10514 nand P1_R1165_U441 P1_R1165_U440 ; P1_R1165_U68
g10515 nand P1_R1165_U444 P1_R1165_U443 ; P1_R1165_U69
g10516 nand P1_R1165_U447 P1_R1165_U446 ; P1_R1165_U70
g10517 nand P1_R1165_U471 P1_R1165_U470 ; P1_R1165_U71
g10518 nand P1_R1165_U468 P1_R1165_U467 ; P1_R1165_U72
g10519 nand P1_R1165_U450 P1_R1165_U449 ; P1_R1165_U73
g10520 nand P1_R1165_U459 P1_R1165_U458 ; P1_R1165_U74
g10521 nand P1_R1165_U453 P1_R1165_U452 ; P1_R1165_U75
g10522 nand P1_R1165_U456 P1_R1165_U455 ; P1_R1165_U76
g10523 nand P1_R1165_U462 P1_R1165_U461 ; P1_R1165_U77
g10524 nand P1_R1165_U465 P1_R1165_U464 ; P1_R1165_U78
g10525 nand P1_R1165_U474 P1_R1165_U473 ; P1_R1165_U79
g10526 nand P1_R1165_U483 P1_R1165_U482 ; P1_R1165_U80
g10527 nand P1_R1165_U477 P1_R1165_U476 ; P1_R1165_U81
g10528 nand P1_R1165_U480 P1_R1165_U479 ; P1_R1165_U82
g10529 nand P1_R1165_U486 P1_R1165_U485 ; P1_R1165_U83
g10530 nand P1_R1165_U489 P1_R1165_U488 ; P1_R1165_U84
g10531 nand P1_R1165_U495 P1_R1165_U494 ; P1_R1165_U85
g10532 nand P1_R1165_U602 P1_R1165_U601 ; P1_R1165_U86
g10533 nand P1_R1165_U401 P1_R1165_U400 ; P1_R1165_U87
g10534 nand P1_R1165_U408 P1_R1165_U407 ; P1_R1165_U88
g10535 nand P1_R1165_U415 P1_R1165_U414 ; P1_R1165_U89
g10536 nand P1_R1165_U422 P1_R1165_U421 ; P1_R1165_U90
g10537 nand P1_R1165_U429 P1_R1165_U428 ; P1_R1165_U91
g10538 nand P1_R1165_U436 P1_R1165_U435 ; P1_R1165_U92
g10539 nand P1_R1165_U498 P1_R1165_U497 ; P1_R1165_U93
g10540 nand P1_R1165_U505 P1_R1165_U504 ; P1_R1165_U94
g10541 nand P1_R1165_U512 P1_R1165_U511 ; P1_R1165_U95
g10542 nand P1_R1165_U517 P1_R1165_U516 ; P1_R1165_U96
g10543 nand P1_R1165_U524 P1_R1165_U523 ; P1_R1165_U97
g10544 nand P1_R1165_U531 P1_R1165_U530 ; P1_R1165_U98
g10545 nand P1_R1165_U538 P1_R1165_U537 ; P1_R1165_U99
g10546 nand P1_R1165_U545 P1_R1165_U544 ; P1_R1165_U100
g10547 nand P1_R1165_U550 P1_R1165_U549 ; P1_R1165_U101
g10548 nand P1_R1165_U557 P1_R1165_U556 ; P1_R1165_U102
g10549 nand P1_R1165_U564 P1_R1165_U563 ; P1_R1165_U103
g10550 nand P1_R1165_U571 P1_R1165_U570 ; P1_R1165_U104
g10551 nand P1_R1165_U578 P1_R1165_U577 ; P1_R1165_U105
g10552 nand P1_R1165_U585 P1_R1165_U584 ; P1_R1165_U106
g10553 nand P1_R1165_U590 P1_R1165_U589 ; P1_R1165_U107
g10554 nand P1_R1165_U597 P1_R1165_U596 ; P1_R1165_U108
g10555 and P1_R1165_U213 P1_R1165_U212 ; P1_R1165_U109
g10556 and P1_R1165_U226 P1_R1165_U225 ; P1_R1165_U110
g10557 and P1_R1165_U410 P1_R1165_U409 P1_R1165_U18 ; P1_R1165_U111
g10558 and P1_R1165_U237 P1_R1165_U5 ; P1_R1165_U112
g10559 and P1_R1165_U431 P1_R1165_U430 P1_R1165_U22 ; P1_R1165_U113
g10560 and P1_R1165_U244 P1_R1165_U4 ; P1_R1165_U114
g10561 and P1_R1165_U257 P1_R1165_U6 ; P1_R1165_U115
g10562 and P1_R1165_U255 P1_R1165_U195 ; P1_R1165_U116
g10563 and P1_R1165_U275 P1_R1165_U274 ; P1_R1165_U117
g10564 and P1_R1165_U287 P1_R1165_U8 ; P1_R1165_U118
g10565 and P1_R1165_U285 P1_R1165_U196 ; P1_R1165_U119
g10566 and P1_R1165_U359 P1_R1165_U52 ; P1_R1165_U120
g10567 and P1_R1165_U308 P1_R1165_U303 ; P1_R1165_U121
g10568 and P1_R1165_U356 P1_R1165_U307 ; P1_R1165_U122
g10569 nand P1_R1165_U492 P1_R1165_U491 ; P1_R1165_U123
g10570 and P1_R1165_U352 P1_R1165_U52 ; P1_R1165_U124
g10571 and P1_R1165_U442 P1_R1165_U33 ; P1_R1165_U125
g10572 and P1_R1165_U200 P1_R1165_U197 ; P1_R1165_U126
g10573 and P1_R1165_U313 P1_R1165_U193 ; P1_R1165_U127
g10574 and P1_R1165_U9 P1_R1165_U197 ; P1_R1165_U128
g10575 and P1_R1165_U533 P1_R1165_U532 P1_R1165_U196 ; P1_R1165_U129
g10576 and P1_R1165_U322 P1_R1165_U8 ; P1_R1165_U130
g10577 and P1_R1165_U559 P1_R1165_U558 P1_R1165_U36 ; P1_R1165_U131
g10578 and P1_R1165_U329 P1_R1165_U7 ; P1_R1165_U132
g10579 and P1_R1165_U580 P1_R1165_U579 P1_R1165_U195 ; P1_R1165_U133
g10580 and P1_R1165_U338 P1_R1165_U6 ; P1_R1165_U134
g10581 nand P1_R1165_U599 P1_R1165_U598 ; P1_R1165_U135
g10582 not P1_U3199 ; P1_R1165_U136
g10583 and P1_R1165_U369 P1_R1165_U368 ; P1_R1165_U137
g10584 not P1_U3204 ; P1_R1165_U138
g10585 not P1_U3208 ; P1_R1165_U139
g10586 not P1_U3207 ; P1_R1165_U140
g10587 not P1_U3205 ; P1_R1165_U141
g10588 not P1_U3206 ; P1_R1165_U142
g10589 not P1_U3203 ; P1_R1165_U143
g10590 not P1_U3201 ; P1_R1165_U144
g10591 not P1_U3202 ; P1_R1165_U145
g10592 not P1_U3200 ; P1_R1165_U146
g10593 nand P1_R1165_U231 P1_R1165_U230 ; P1_R1165_U147
g10594 and P1_R1165_U403 P1_R1165_U402 ; P1_R1165_U148
g10595 nand P1_R1165_U110 P1_R1165_U227 ; P1_R1165_U149
g10596 and P1_R1165_U417 P1_R1165_U416 ; P1_R1165_U150
g10597 nand P1_R1165_U361 P1_R1165_U350 ; P1_R1165_U151
g10598 and P1_R1165_U424 P1_R1165_U423 ; P1_R1165_U152
g10599 nand P1_R1165_U109 P1_R1165_U214 ; P1_R1165_U153
g10600 not P1_U3181 ; P1_R1165_U154
g10601 not P1_U3183 ; P1_R1165_U155
g10602 not P1_U3182 ; P1_R1165_U156
g10603 not P1_U3184 ; P1_R1165_U157
g10604 not P1_U3198 ; P1_R1165_U158
g10605 not P1_U3195 ; P1_R1165_U159
g10606 not P1_U3196 ; P1_R1165_U160
g10607 not P1_U3197 ; P1_R1165_U161
g10608 not P1_U3194 ; P1_R1165_U162
g10609 not P1_U3193 ; P1_R1165_U163
g10610 not P1_U3191 ; P1_R1165_U164
g10611 not P1_U3192 ; P1_R1165_U165
g10612 not P1_U3190 ; P1_R1165_U166
g10613 not P1_U3187 ; P1_R1165_U167
g10614 not P1_U3188 ; P1_R1165_U168
g10615 not P1_U3189 ; P1_R1165_U169
g10616 not P1_U3186 ; P1_R1165_U170
g10617 not P1_U3185 ; P1_R1165_U171
g10618 not P1_U3151 ; P1_R1165_U172
g10619 not P1_U3180 ; P1_R1165_U173
g10620 and P1_R1165_U500 P1_R1165_U499 ; P1_R1165_U174
g10621 nand P1_R1165_U124 P1_R1165_U304 ; P1_R1165_U175
g10622 nand P1_R1165_U298 P1_R1165_U297 ; P1_R1165_U176
g10623 and P1_R1165_U519 P1_R1165_U518 ; P1_R1165_U177
g10624 nand P1_R1165_U294 P1_R1165_U293 ; P1_R1165_U178
g10625 and P1_R1165_U526 P1_R1165_U525 ; P1_R1165_U179
g10626 nand P1_R1165_U290 P1_R1165_U289 ; P1_R1165_U180
g10627 and P1_R1165_U540 P1_R1165_U539 ; P1_R1165_U181
g10628 nand P1_R1165_U203 P1_R1165_U202 ; P1_R1165_U182
g10629 nand P1_R1165_U280 P1_R1165_U279 ; P1_R1165_U183
g10630 and P1_R1165_U552 P1_R1165_U551 ; P1_R1165_U184
g10631 nand P1_R1165_U117 P1_R1165_U276 ; P1_R1165_U185
g10632 and P1_R1165_U566 P1_R1165_U565 ; P1_R1165_U186
g10633 nand P1_R1165_U264 P1_R1165_U263 ; P1_R1165_U187
g10634 and P1_R1165_U573 P1_R1165_U572 ; P1_R1165_U188
g10635 nand P1_R1165_U260 P1_R1165_U259 ; P1_R1165_U189
g10636 nand P1_R1165_U250 P1_R1165_U249 ; P1_R1165_U190
g10637 and P1_R1165_U592 P1_R1165_U591 ; P1_R1165_U191
g10638 nand P1_R1165_U363 P1_R1165_U353 ; P1_R1165_U192
g10639 nand P1_R1165_U355 P1_R1165_U354 ; P1_R1165_U193
g10640 not P1_R1165_U22 ; P1_R1165_U194
g10641 nand P1_U3167 P1_R1165_U76 ; P1_R1165_U195
g10642 nand P1_U3159 P1_R1165_U82 ; P1_R1165_U196
g10643 nand P1_U3154 P1_R1165_U68 ; P1_R1165_U197
g10644 not P1_R1165_U41 ; P1_R1165_U198
g10645 not P1_R1165_U48 ; P1_R1165_U199
g10646 nand P1_U3155 P1_R1165_U70 ; P1_R1165_U200
g10647 or P1_U3209 P1_U3179 ; P1_R1165_U201
g10648 nand P1_R1165_U63 P1_R1165_U201 ; P1_R1165_U202
g10649 nand P1_U3179 P1_U3209 ; P1_R1165_U203
g10650 not P1_R1165_U182 ; P1_R1165_U204
g10651 nand P1_R1165_U381 P1_R1165_U25 ; P1_R1165_U205
g10652 nand P1_R1165_U205 P1_R1165_U182 ; P1_R1165_U206
g10653 nand P1_U3178 P1_R1165_U64 ; P1_R1165_U207
g10654 not P1_R1165_U30 ; P1_R1165_U208
g10655 nand P1_R1165_U384 P1_R1165_U23 ; P1_R1165_U209
g10656 nand P1_R1165_U387 P1_R1165_U21 ; P1_R1165_U210
g10657 nand P1_R1165_U23 P1_R1165_U22 ; P1_R1165_U211
g10658 nand P1_R1165_U62 P1_R1165_U211 ; P1_R1165_U212
g10659 nand P1_U3176 P1_R1165_U194 ; P1_R1165_U213
g10660 nand P1_R1165_U4 P1_R1165_U30 ; P1_R1165_U214
g10661 not P1_R1165_U153 ; P1_R1165_U215
g10662 nand P1_R1165_U375 P1_R1165_U20 ; P1_R1165_U216
g10663 nand P1_R1165_U390 P1_R1165_U26 ; P1_R1165_U217
g10664 nand P1_R1165_U217 P1_R1165_U151 ; P1_R1165_U218
g10665 nand P1_U3174 P1_R1165_U65 ; P1_R1165_U219
g10666 not P1_R1165_U29 ; P1_R1165_U220
g10667 nand P1_R1165_U393 P1_R1165_U19 ; P1_R1165_U221
g10668 nand P1_R1165_U396 P1_R1165_U17 ; P1_R1165_U222
g10669 not P1_R1165_U18 ; P1_R1165_U223
g10670 nand P1_R1165_U19 P1_R1165_U18 ; P1_R1165_U224
g10671 nand P1_R1165_U59 P1_R1165_U224 ; P1_R1165_U225
g10672 nand P1_U3172 P1_R1165_U223 ; P1_R1165_U226
g10673 nand P1_R1165_U5 P1_R1165_U29 ; P1_R1165_U227
g10674 not P1_R1165_U149 ; P1_R1165_U228
g10675 nand P1_R1165_U399 P1_R1165_U27 ; P1_R1165_U229
g10676 nand P1_R1165_U229 P1_R1165_U149 ; P1_R1165_U230
g10677 nand P1_U3171 P1_R1165_U66 ; P1_R1165_U231
g10678 not P1_R1165_U147 ; P1_R1165_U232
g10679 nand P1_R1165_U396 P1_R1165_U17 ; P1_R1165_U233
g10680 nand P1_R1165_U233 P1_R1165_U29 ; P1_R1165_U234
g10681 nand P1_R1165_U111 P1_R1165_U234 ; P1_R1165_U235
g10682 nand P1_R1165_U220 P1_R1165_U18 ; P1_R1165_U236
g10683 nand P1_U3172 P1_R1165_U59 ; P1_R1165_U237
g10684 nand P1_R1165_U112 P1_R1165_U236 ; P1_R1165_U238
g10685 nand P1_R1165_U396 P1_R1165_U17 ; P1_R1165_U239
g10686 nand P1_R1165_U387 P1_R1165_U21 ; P1_R1165_U240
g10687 nand P1_R1165_U240 P1_R1165_U30 ; P1_R1165_U241
g10688 nand P1_R1165_U113 P1_R1165_U241 ; P1_R1165_U242
g10689 nand P1_R1165_U208 P1_R1165_U22 ; P1_R1165_U243
g10690 nand P1_U3176 P1_R1165_U62 ; P1_R1165_U244
g10691 nand P1_R1165_U114 P1_R1165_U243 ; P1_R1165_U245
g10692 nand P1_R1165_U387 P1_R1165_U21 ; P1_R1165_U246
g10693 nand P1_R1165_U367 P1_R1165_U28 ; P1_R1165_U247
g10694 nand P1_R1165_U451 P1_R1165_U38 ; P1_R1165_U248
g10695 nand P1_R1165_U248 P1_R1165_U192 ; P1_R1165_U249
g10696 nand P1_U3169 P1_R1165_U73 ; P1_R1165_U250
g10697 not P1_R1165_U190 ; P1_R1165_U251
g10698 nand P1_R1165_U454 P1_R1165_U42 ; P1_R1165_U252
g10699 nand P1_R1165_U457 P1_R1165_U39 ; P1_R1165_U253
g10700 nand P1_R1165_U198 P1_R1165_U6 ; P1_R1165_U254
g10701 nand P1_U3166 P1_R1165_U75 ; P1_R1165_U255
g10702 nand P1_R1165_U116 P1_R1165_U254 ; P1_R1165_U256
g10703 nand P1_R1165_U460 P1_R1165_U40 ; P1_R1165_U257
g10704 nand P1_R1165_U454 P1_R1165_U42 ; P1_R1165_U258
g10705 nand P1_R1165_U115 P1_R1165_U190 ; P1_R1165_U259
g10706 nand P1_R1165_U258 P1_R1165_U256 ; P1_R1165_U260
g10707 not P1_R1165_U189 ; P1_R1165_U261
g10708 nand P1_R1165_U463 P1_R1165_U43 ; P1_R1165_U262
g10709 nand P1_R1165_U262 P1_R1165_U189 ; P1_R1165_U263
g10710 nand P1_U3165 P1_R1165_U77 ; P1_R1165_U264
g10711 not P1_R1165_U187 ; P1_R1165_U265
g10712 nand P1_R1165_U466 P1_R1165_U44 ; P1_R1165_U266
g10713 nand P1_R1165_U266 P1_R1165_U187 ; P1_R1165_U267
g10714 nand P1_U3164 P1_R1165_U78 ; P1_R1165_U268
g10715 not P1_R1165_U55 ; P1_R1165_U269
g10716 nand P1_R1165_U469 P1_R1165_U37 ; P1_R1165_U270
g10717 nand P1_R1165_U472 P1_R1165_U35 ; P1_R1165_U271
g10718 not P1_R1165_U36 ; P1_R1165_U272
g10719 nand P1_R1165_U37 P1_R1165_U36 ; P1_R1165_U273
g10720 nand P1_R1165_U72 P1_R1165_U273 ; P1_R1165_U274
g10721 nand P1_U3162 P1_R1165_U272 ; P1_R1165_U275
g10722 nand P1_R1165_U7 P1_R1165_U55 ; P1_R1165_U276
g10723 not P1_R1165_U185 ; P1_R1165_U277
g10724 nand P1_R1165_U475 P1_R1165_U45 ; P1_R1165_U278
g10725 nand P1_R1165_U278 P1_R1165_U185 ; P1_R1165_U279
g10726 nand P1_U3161 P1_R1165_U79 ; P1_R1165_U280
g10727 not P1_R1165_U183 ; P1_R1165_U281
g10728 nand P1_R1165_U478 P1_R1165_U49 ; P1_R1165_U282
g10729 nand P1_R1165_U481 P1_R1165_U46 ; P1_R1165_U283
g10730 nand P1_R1165_U199 P1_R1165_U8 ; P1_R1165_U284
g10731 nand P1_U3158 P1_R1165_U81 ; P1_R1165_U285
g10732 nand P1_R1165_U119 P1_R1165_U284 ; P1_R1165_U286
g10733 nand P1_R1165_U484 P1_R1165_U47 ; P1_R1165_U287
g10734 nand P1_R1165_U478 P1_R1165_U49 ; P1_R1165_U288
g10735 nand P1_R1165_U118 P1_R1165_U183 ; P1_R1165_U289
g10736 nand P1_R1165_U288 P1_R1165_U286 ; P1_R1165_U290
g10737 not P1_R1165_U180 ; P1_R1165_U291
g10738 nand P1_R1165_U487 P1_R1165_U50 ; P1_R1165_U292
g10739 nand P1_R1165_U292 P1_R1165_U180 ; P1_R1165_U293
g10740 nand P1_U3157 P1_R1165_U83 ; P1_R1165_U294
g10741 not P1_R1165_U178 ; P1_R1165_U295
g10742 nand P1_R1165_U490 P1_R1165_U51 ; P1_R1165_U296
g10743 nand P1_R1165_U296 P1_R1165_U178 ; P1_R1165_U297
g10744 nand P1_U3156 P1_R1165_U84 ; P1_R1165_U298
g10745 not P1_R1165_U176 ; P1_R1165_U299
g10746 nand P1_R1165_U442 P1_R1165_U33 ; P1_R1165_U300
g10747 nand P1_R1165_U200 P1_R1165_U197 ; P1_R1165_U301
g10748 not P1_R1165_U52 ; P1_R1165_U302
g10749 nand P1_R1165_U448 P1_R1165_U34 ; P1_R1165_U303
g10750 nand P1_R1165_U176 P1_R1165_U303 P1_R1165_U193 ; P1_R1165_U304
g10751 not P1_R1165_U175 ; P1_R1165_U305
g10752 nand P1_R1165_U439 P1_R1165_U31 ; P1_R1165_U306
g10753 nand P1_U3152 P1_R1165_U67 ; P1_R1165_U307
g10754 nand P1_R1165_U439 P1_R1165_U31 ; P1_R1165_U308
g10755 nand P1_R1165_U303 P1_R1165_U176 ; P1_R1165_U309
g10756 not P1_R1165_U53 ; P1_R1165_U310
g10757 nand P1_R1165_U125 P1_R1165_U9 ; P1_R1165_U311
g10758 nand P1_R1165_U126 P1_R1165_U309 ; P1_R1165_U312
g10759 nand P1_U3153 P1_R1165_U69 ; P1_R1165_U313
g10760 nand P1_R1165_U127 P1_R1165_U312 ; P1_R1165_U314
g10761 nand P1_R1165_U442 P1_R1165_U33 ; P1_R1165_U315
g10762 nand P1_R1165_U287 P1_R1165_U183 ; P1_R1165_U316
g10763 not P1_R1165_U54 ; P1_R1165_U317
g10764 nand P1_R1165_U481 P1_R1165_U46 ; P1_R1165_U318
g10765 nand P1_R1165_U318 P1_R1165_U54 ; P1_R1165_U319
g10766 nand P1_R1165_U129 P1_R1165_U319 ; P1_R1165_U320
g10767 nand P1_R1165_U317 P1_R1165_U196 ; P1_R1165_U321
g10768 nand P1_U3158 P1_R1165_U81 ; P1_R1165_U322
g10769 nand P1_R1165_U130 P1_R1165_U321 ; P1_R1165_U323
g10770 nand P1_R1165_U481 P1_R1165_U46 ; P1_R1165_U324
g10771 nand P1_R1165_U472 P1_R1165_U35 ; P1_R1165_U325
g10772 nand P1_R1165_U325 P1_R1165_U55 ; P1_R1165_U326
g10773 nand P1_R1165_U131 P1_R1165_U326 ; P1_R1165_U327
g10774 nand P1_R1165_U269 P1_R1165_U36 ; P1_R1165_U328
g10775 nand P1_U3162 P1_R1165_U72 ; P1_R1165_U329
g10776 nand P1_R1165_U132 P1_R1165_U328 ; P1_R1165_U330
g10777 nand P1_R1165_U472 P1_R1165_U35 ; P1_R1165_U331
g10778 nand P1_R1165_U257 P1_R1165_U190 ; P1_R1165_U332
g10779 not P1_R1165_U56 ; P1_R1165_U333
g10780 nand P1_R1165_U457 P1_R1165_U39 ; P1_R1165_U334
g10781 nand P1_R1165_U334 P1_R1165_U56 ; P1_R1165_U335
g10782 nand P1_R1165_U133 P1_R1165_U335 ; P1_R1165_U336
g10783 nand P1_R1165_U333 P1_R1165_U195 ; P1_R1165_U337
g10784 nand P1_U3166 P1_R1165_U75 ; P1_R1165_U338
g10785 nand P1_R1165_U134 P1_R1165_U337 ; P1_R1165_U339
g10786 nand P1_R1165_U457 P1_R1165_U39 ; P1_R1165_U340
g10787 nand P1_R1165_U239 P1_R1165_U18 ; P1_R1165_U341
g10788 nand P1_R1165_U246 P1_R1165_U22 ; P1_R1165_U342
g10789 nand P1_R1165_U315 P1_R1165_U197 ; P1_R1165_U343
g10790 nand P1_R1165_U303 P1_R1165_U200 ; P1_R1165_U344
g10791 nand P1_R1165_U324 P1_R1165_U196 ; P1_R1165_U345
g10792 nand P1_R1165_U287 P1_R1165_U48 ; P1_R1165_U346
g10793 nand P1_R1165_U331 P1_R1165_U36 ; P1_R1165_U347
g10794 nand P1_R1165_U340 P1_R1165_U195 ; P1_R1165_U348
g10795 nand P1_R1165_U257 P1_R1165_U41 ; P1_R1165_U349
g10796 nand P1_U3175 P1_R1165_U60 ; P1_R1165_U350
g10797 nand P1_R1165_U352 P1_R1165_U304 P1_R1165_U120 ; P1_R1165_U351
g10798 nand P1_R1165_U301 P1_R1165_U193 ; P1_R1165_U352
g10799 nand P1_U3170 P1_R1165_U57 ; P1_R1165_U353
g10800 nand P1_R1165_U69 P1_R1165_U300 ; P1_R1165_U354
g10801 nand P1_U3153 P1_R1165_U300 ; P1_R1165_U355
g10802 nand P1_R1165_U301 P1_R1165_U193 P1_R1165_U308 ; P1_R1165_U356
g10803 nand P1_R1165_U176 P1_R1165_U193 P1_R1165_U121 ; P1_R1165_U357
g10804 nand P1_R1165_U302 P1_R1165_U308 ; P1_R1165_U358
g10805 nand P1_U3152 P1_R1165_U67 ; P1_R1165_U359
g10806 nand P1_R1165_U128 P1_R1165_U310 ; P1_R1165_U360
g10807 nand P1_R1165_U216 P1_R1165_U153 ; P1_R1165_U361
g10808 not P1_R1165_U151 ; P1_R1165_U362
g10809 nand P1_R1165_U247 P1_R1165_U147 ; P1_R1165_U363
g10810 not P1_R1165_U192 ; P1_R1165_U364
g10811 nand P1_U3209 P1_R1165_U136 ; P1_R1165_U365
g10812 nand P1_U3199 P1_R1165_U16 ; P1_R1165_U366
g10813 not P1_R1165_U57 ; P1_R1165_U367
g10814 nand P1_R1165_U367 P1_U3170 ; P1_R1165_U368
g10815 nand P1_R1165_U57 P1_R1165_U28 ; P1_R1165_U369
g10816 nand P1_R1165_U367 P1_U3170 ; P1_R1165_U370
g10817 nand P1_R1165_U57 P1_R1165_U28 ; P1_R1165_U371
g10818 nand P1_R1165_U371 P1_R1165_U370 ; P1_R1165_U372
g10819 nand P1_U3209 P1_R1165_U138 ; P1_R1165_U373
g10820 nand P1_U3204 P1_R1165_U16 ; P1_R1165_U374
g10821 not P1_R1165_U60 ; P1_R1165_U375
g10822 nand P1_U3209 P1_R1165_U139 ; P1_R1165_U376
g10823 nand P1_U3208 P1_R1165_U16 ; P1_R1165_U377
g10824 not P1_R1165_U63 ; P1_R1165_U378
g10825 nand P1_U3209 P1_R1165_U140 ; P1_R1165_U379
g10826 nand P1_U3207 P1_R1165_U16 ; P1_R1165_U380
g10827 not P1_R1165_U64 ; P1_R1165_U381
g10828 nand P1_U3209 P1_R1165_U141 ; P1_R1165_U382
g10829 nand P1_U3205 P1_R1165_U16 ; P1_R1165_U383
g10830 not P1_R1165_U62 ; P1_R1165_U384
g10831 nand P1_U3209 P1_R1165_U142 ; P1_R1165_U385
g10832 nand P1_U3206 P1_R1165_U16 ; P1_R1165_U386
g10833 not P1_R1165_U61 ; P1_R1165_U387
g10834 nand P1_U3209 P1_R1165_U143 ; P1_R1165_U388
g10835 nand P1_U3203 P1_R1165_U16 ; P1_R1165_U389
g10836 not P1_R1165_U65 ; P1_R1165_U390
g10837 nand P1_U3209 P1_R1165_U144 ; P1_R1165_U391
g10838 nand P1_U3201 P1_R1165_U16 ; P1_R1165_U392
g10839 not P1_R1165_U59 ; P1_R1165_U393
g10840 nand P1_U3209 P1_R1165_U145 ; P1_R1165_U394
g10841 nand P1_U3202 P1_R1165_U16 ; P1_R1165_U395
g10842 not P1_R1165_U58 ; P1_R1165_U396
g10843 nand P1_U3209 P1_R1165_U146 ; P1_R1165_U397
g10844 nand P1_U3200 P1_R1165_U16 ; P1_R1165_U398
g10845 not P1_R1165_U66 ; P1_R1165_U399
g10846 nand P1_R1165_U137 P1_R1165_U147 ; P1_R1165_U400
g10847 nand P1_R1165_U232 P1_R1165_U372 ; P1_R1165_U401
g10848 nand P1_R1165_U399 P1_U3171 ; P1_R1165_U402
g10849 nand P1_R1165_U66 P1_R1165_U27 ; P1_R1165_U403
g10850 nand P1_R1165_U399 P1_U3171 ; P1_R1165_U404
g10851 nand P1_R1165_U66 P1_R1165_U27 ; P1_R1165_U405
g10852 nand P1_R1165_U405 P1_R1165_U404 ; P1_R1165_U406
g10853 nand P1_R1165_U148 P1_R1165_U149 ; P1_R1165_U407
g10854 nand P1_R1165_U228 P1_R1165_U406 ; P1_R1165_U408
g10855 nand P1_R1165_U393 P1_U3172 ; P1_R1165_U409
g10856 nand P1_R1165_U59 P1_R1165_U19 ; P1_R1165_U410
g10857 nand P1_R1165_U396 P1_U3173 ; P1_R1165_U411
g10858 nand P1_R1165_U58 P1_R1165_U17 ; P1_R1165_U412
g10859 nand P1_R1165_U412 P1_R1165_U411 ; P1_R1165_U413
g10860 nand P1_R1165_U341 P1_R1165_U29 ; P1_R1165_U414
g10861 nand P1_R1165_U413 P1_R1165_U220 ; P1_R1165_U415
g10862 nand P1_R1165_U390 P1_U3174 ; P1_R1165_U416
g10863 nand P1_R1165_U65 P1_R1165_U26 ; P1_R1165_U417
g10864 nand P1_R1165_U390 P1_U3174 ; P1_R1165_U418
g10865 nand P1_R1165_U65 P1_R1165_U26 ; P1_R1165_U419
g10866 nand P1_R1165_U419 P1_R1165_U418 ; P1_R1165_U420
g10867 nand P1_R1165_U150 P1_R1165_U151 ; P1_R1165_U421
g10868 nand P1_R1165_U362 P1_R1165_U420 ; P1_R1165_U422
g10869 nand P1_R1165_U375 P1_U3175 ; P1_R1165_U423
g10870 nand P1_R1165_U60 P1_R1165_U20 ; P1_R1165_U424
g10871 nand P1_R1165_U375 P1_U3175 ; P1_R1165_U425
g10872 nand P1_R1165_U60 P1_R1165_U20 ; P1_R1165_U426
g10873 nand P1_R1165_U426 P1_R1165_U425 ; P1_R1165_U427
g10874 nand P1_R1165_U152 P1_R1165_U153 ; P1_R1165_U428
g10875 nand P1_R1165_U215 P1_R1165_U427 ; P1_R1165_U429
g10876 nand P1_R1165_U384 P1_U3176 ; P1_R1165_U430
g10877 nand P1_R1165_U62 P1_R1165_U23 ; P1_R1165_U431
g10878 nand P1_R1165_U387 P1_U3177 ; P1_R1165_U432
g10879 nand P1_R1165_U61 P1_R1165_U21 ; P1_R1165_U433
g10880 nand P1_R1165_U433 P1_R1165_U432 ; P1_R1165_U434
g10881 nand P1_R1165_U342 P1_R1165_U30 ; P1_R1165_U435
g10882 nand P1_R1165_U434 P1_R1165_U208 ; P1_R1165_U436
g10883 nand P1_U3209 P1_R1165_U154 ; P1_R1165_U437
g10884 nand P1_U3181 P1_R1165_U16 ; P1_R1165_U438
g10885 not P1_R1165_U67 ; P1_R1165_U439
g10886 nand P1_U3209 P1_R1165_U155 ; P1_R1165_U440
g10887 nand P1_U3183 P1_R1165_U16 ; P1_R1165_U441
g10888 not P1_R1165_U68 ; P1_R1165_U442
g10889 nand P1_U3209 P1_R1165_U156 ; P1_R1165_U443
g10890 nand P1_U3182 P1_R1165_U16 ; P1_R1165_U444
g10891 not P1_R1165_U69 ; P1_R1165_U445
g10892 nand P1_U3209 P1_R1165_U157 ; P1_R1165_U446
g10893 nand P1_U3184 P1_R1165_U16 ; P1_R1165_U447
g10894 not P1_R1165_U70 ; P1_R1165_U448
g10895 nand P1_U3209 P1_R1165_U158 ; P1_R1165_U449
g10896 nand P1_U3198 P1_R1165_U16 ; P1_R1165_U450
g10897 not P1_R1165_U73 ; P1_R1165_U451
g10898 nand P1_U3209 P1_R1165_U159 ; P1_R1165_U452
g10899 nand P1_U3195 P1_R1165_U16 ; P1_R1165_U453
g10900 not P1_R1165_U75 ; P1_R1165_U454
g10901 nand P1_U3209 P1_R1165_U160 ; P1_R1165_U455
g10902 nand P1_U3196 P1_R1165_U16 ; P1_R1165_U456
g10903 not P1_R1165_U76 ; P1_R1165_U457
g10904 nand P1_U3209 P1_R1165_U161 ; P1_R1165_U458
g10905 nand P1_U3197 P1_R1165_U16 ; P1_R1165_U459
g10906 not P1_R1165_U74 ; P1_R1165_U460
g10907 nand P1_U3209 P1_R1165_U162 ; P1_R1165_U461
g10908 nand P1_U3194 P1_R1165_U16 ; P1_R1165_U462
g10909 not P1_R1165_U77 ; P1_R1165_U463
g10910 nand P1_U3209 P1_R1165_U163 ; P1_R1165_U464
g10911 nand P1_U3193 P1_R1165_U16 ; P1_R1165_U465
g10912 not P1_R1165_U78 ; P1_R1165_U466
g10913 nand P1_U3209 P1_R1165_U164 ; P1_R1165_U467
g10914 nand P1_U3191 P1_R1165_U16 ; P1_R1165_U468
g10915 not P1_R1165_U72 ; P1_R1165_U469
g10916 nand P1_U3209 P1_R1165_U165 ; P1_R1165_U470
g10917 nand P1_U3192 P1_R1165_U16 ; P1_R1165_U471
g10918 not P1_R1165_U71 ; P1_R1165_U472
g10919 nand P1_U3209 P1_R1165_U166 ; P1_R1165_U473
g10920 nand P1_U3190 P1_R1165_U16 ; P1_R1165_U474
g10921 not P1_R1165_U79 ; P1_R1165_U475
g10922 nand P1_U3209 P1_R1165_U167 ; P1_R1165_U476
g10923 nand P1_U3187 P1_R1165_U16 ; P1_R1165_U477
g10924 not P1_R1165_U81 ; P1_R1165_U478
g10925 nand P1_U3209 P1_R1165_U168 ; P1_R1165_U479
g10926 nand P1_U3188 P1_R1165_U16 ; P1_R1165_U480
g10927 not P1_R1165_U82 ; P1_R1165_U481
g10928 nand P1_U3209 P1_R1165_U169 ; P1_R1165_U482
g10929 nand P1_U3189 P1_R1165_U16 ; P1_R1165_U483
g10930 not P1_R1165_U80 ; P1_R1165_U484
g10931 nand P1_U3209 P1_R1165_U170 ; P1_R1165_U485
g10932 nand P1_U3186 P1_R1165_U16 ; P1_R1165_U486
g10933 not P1_R1165_U83 ; P1_R1165_U487
g10934 nand P1_U3209 P1_R1165_U171 ; P1_R1165_U488
g10935 nand P1_U3185 P1_R1165_U16 ; P1_R1165_U489
g10936 not P1_R1165_U84 ; P1_R1165_U490
g10937 nand P1_U3209 P1_R1165_U172 ; P1_R1165_U491
g10938 nand P1_U3151 P1_R1165_U16 ; P1_R1165_U492
g10939 not P1_R1165_U123 ; P1_R1165_U493
g10940 nand P1_U3180 P1_R1165_U493 ; P1_R1165_U494
g10941 nand P1_R1165_U123 P1_R1165_U173 ; P1_R1165_U495
g10942 not P1_R1165_U85 ; P1_R1165_U496
g10943 nand P1_R1165_U351 P1_R1165_U306 P1_R1165_U496 ; P1_R1165_U497
g10944 nand P1_R1165_U358 P1_R1165_U357 P1_R1165_U122 P1_R1165_U85 ; P1_R1165_U498
g10945 nand P1_R1165_U439 P1_U3152 ; P1_R1165_U499
g10946 nand P1_R1165_U67 P1_R1165_U31 ; P1_R1165_U500
g10947 nand P1_R1165_U439 P1_U3152 ; P1_R1165_U501
g10948 nand P1_R1165_U67 P1_R1165_U31 ; P1_R1165_U502
g10949 nand P1_R1165_U502 P1_R1165_U501 ; P1_R1165_U503
g10950 nand P1_R1165_U174 P1_R1165_U175 ; P1_R1165_U504
g10951 nand P1_R1165_U305 P1_R1165_U503 ; P1_R1165_U505
g10952 nand P1_R1165_U445 P1_U3153 ; P1_R1165_U506
g10953 nand P1_R1165_U69 P1_R1165_U32 ; P1_R1165_U507
g10954 nand P1_R1165_U442 P1_U3154 ; P1_R1165_U508
g10955 nand P1_R1165_U68 P1_R1165_U33 ; P1_R1165_U509
g10956 nand P1_R1165_U509 P1_R1165_U508 ; P1_R1165_U510
g10957 nand P1_R1165_U343 P1_R1165_U53 ; P1_R1165_U511
g10958 nand P1_R1165_U510 P1_R1165_U310 ; P1_R1165_U512
g10959 nand P1_R1165_U448 P1_U3155 ; P1_R1165_U513
g10960 nand P1_R1165_U70 P1_R1165_U34 ; P1_R1165_U514
g10961 nand P1_R1165_U514 P1_R1165_U513 ; P1_R1165_U515
g10962 nand P1_R1165_U344 P1_R1165_U176 ; P1_R1165_U516
g10963 nand P1_R1165_U299 P1_R1165_U515 ; P1_R1165_U517
g10964 nand P1_R1165_U490 P1_U3156 ; P1_R1165_U518
g10965 nand P1_R1165_U84 P1_R1165_U51 ; P1_R1165_U519
g10966 nand P1_R1165_U490 P1_U3156 ; P1_R1165_U520
g10967 nand P1_R1165_U84 P1_R1165_U51 ; P1_R1165_U521
g10968 nand P1_R1165_U521 P1_R1165_U520 ; P1_R1165_U522
g10969 nand P1_R1165_U177 P1_R1165_U178 ; P1_R1165_U523
g10970 nand P1_R1165_U295 P1_R1165_U522 ; P1_R1165_U524
g10971 nand P1_R1165_U487 P1_U3157 ; P1_R1165_U525
g10972 nand P1_R1165_U83 P1_R1165_U50 ; P1_R1165_U526
g10973 nand P1_R1165_U487 P1_U3157 ; P1_R1165_U527
g10974 nand P1_R1165_U83 P1_R1165_U50 ; P1_R1165_U528
g10975 nand P1_R1165_U528 P1_R1165_U527 ; P1_R1165_U529
g10976 nand P1_R1165_U179 P1_R1165_U180 ; P1_R1165_U530
g10977 nand P1_R1165_U291 P1_R1165_U529 ; P1_R1165_U531
g10978 nand P1_R1165_U478 P1_U3158 ; P1_R1165_U532
g10979 nand P1_R1165_U81 P1_R1165_U49 ; P1_R1165_U533
g10980 nand P1_R1165_U481 P1_U3159 ; P1_R1165_U534
g10981 nand P1_R1165_U82 P1_R1165_U46 ; P1_R1165_U535
g10982 nand P1_R1165_U535 P1_R1165_U534 ; P1_R1165_U536
g10983 nand P1_R1165_U345 P1_R1165_U54 ; P1_R1165_U537
g10984 nand P1_R1165_U536 P1_R1165_U317 ; P1_R1165_U538
g10985 nand P1_R1165_U381 P1_U3178 ; P1_R1165_U539
g10986 nand P1_R1165_U64 P1_R1165_U25 ; P1_R1165_U540
g10987 nand P1_R1165_U381 P1_U3178 ; P1_R1165_U541
g10988 nand P1_R1165_U64 P1_R1165_U25 ; P1_R1165_U542
g10989 nand P1_R1165_U542 P1_R1165_U541 ; P1_R1165_U543
g10990 nand P1_R1165_U181 P1_R1165_U182 ; P1_R1165_U544
g10991 nand P1_R1165_U204 P1_R1165_U543 ; P1_R1165_U545
g10992 nand P1_R1165_U484 P1_U3160 ; P1_R1165_U546
g10993 nand P1_R1165_U80 P1_R1165_U47 ; P1_R1165_U547
g10994 nand P1_R1165_U547 P1_R1165_U546 ; P1_R1165_U548
g10995 nand P1_R1165_U346 P1_R1165_U183 ; P1_R1165_U549
g10996 nand P1_R1165_U281 P1_R1165_U548 ; P1_R1165_U550
g10997 nand P1_R1165_U475 P1_U3161 ; P1_R1165_U551
g10998 nand P1_R1165_U79 P1_R1165_U45 ; P1_R1165_U552
g10999 nand P1_R1165_U475 P1_U3161 ; P1_R1165_U553
g11000 nand P1_R1165_U79 P1_R1165_U45 ; P1_R1165_U554
g11001 nand P1_R1165_U554 P1_R1165_U553 ; P1_R1165_U555
g11002 nand P1_R1165_U184 P1_R1165_U185 ; P1_R1165_U556
g11003 nand P1_R1165_U277 P1_R1165_U555 ; P1_R1165_U557
g11004 nand P1_R1165_U469 P1_U3162 ; P1_R1165_U558
g11005 nand P1_R1165_U72 P1_R1165_U37 ; P1_R1165_U559
g11006 nand P1_R1165_U472 P1_U3163 ; P1_R1165_U560
g11007 nand P1_R1165_U71 P1_R1165_U35 ; P1_R1165_U561
g11008 nand P1_R1165_U561 P1_R1165_U560 ; P1_R1165_U562
g11009 nand P1_R1165_U347 P1_R1165_U55 ; P1_R1165_U563
g11010 nand P1_R1165_U562 P1_R1165_U269 ; P1_R1165_U564
g11011 nand P1_R1165_U466 P1_U3164 ; P1_R1165_U565
g11012 nand P1_R1165_U78 P1_R1165_U44 ; P1_R1165_U566
g11013 nand P1_R1165_U466 P1_U3164 ; P1_R1165_U567
g11014 nand P1_R1165_U78 P1_R1165_U44 ; P1_R1165_U568
g11015 nand P1_R1165_U568 P1_R1165_U567 ; P1_R1165_U569
g11016 nand P1_R1165_U186 P1_R1165_U187 ; P1_R1165_U570
g11017 nand P1_R1165_U265 P1_R1165_U569 ; P1_R1165_U571
g11018 nand P1_R1165_U463 P1_U3165 ; P1_R1165_U572
g11019 nand P1_R1165_U77 P1_R1165_U43 ; P1_R1165_U573
g11020 nand P1_R1165_U463 P1_U3165 ; P1_R1165_U574
g11021 nand P1_R1165_U77 P1_R1165_U43 ; P1_R1165_U575
g11022 nand P1_R1165_U575 P1_R1165_U574 ; P1_R1165_U576
g11023 nand P1_R1165_U188 P1_R1165_U189 ; P1_R1165_U577
g11024 nand P1_R1165_U261 P1_R1165_U576 ; P1_R1165_U578
g11025 nand P1_R1165_U454 P1_U3166 ; P1_R1165_U579
g11026 nand P1_R1165_U75 P1_R1165_U42 ; P1_R1165_U580
g11027 nand P1_R1165_U457 P1_U3167 ; P1_R1165_U581
g11028 nand P1_R1165_U76 P1_R1165_U39 ; P1_R1165_U582
g11029 nand P1_R1165_U582 P1_R1165_U581 ; P1_R1165_U583
g11030 nand P1_R1165_U348 P1_R1165_U56 ; P1_R1165_U584
g11031 nand P1_R1165_U583 P1_R1165_U333 ; P1_R1165_U585
g11032 nand P1_R1165_U460 P1_U3168 ; P1_R1165_U586
g11033 nand P1_R1165_U74 P1_R1165_U40 ; P1_R1165_U587
g11034 nand P1_R1165_U587 P1_R1165_U586 ; P1_R1165_U588
g11035 nand P1_R1165_U349 P1_R1165_U190 ; P1_R1165_U589
g11036 nand P1_R1165_U251 P1_R1165_U588 ; P1_R1165_U590
g11037 nand P1_R1165_U451 P1_U3169 ; P1_R1165_U591
g11038 nand P1_R1165_U73 P1_R1165_U38 ; P1_R1165_U592
g11039 nand P1_R1165_U451 P1_U3169 ; P1_R1165_U593
g11040 nand P1_R1165_U73 P1_R1165_U38 ; P1_R1165_U594
g11041 nand P1_R1165_U594 P1_R1165_U593 ; P1_R1165_U595
g11042 nand P1_R1165_U191 P1_R1165_U192 ; P1_R1165_U596
g11043 nand P1_R1165_U364 P1_R1165_U595 ; P1_R1165_U597
g11044 nand P1_U3179 P1_R1165_U16 ; P1_R1165_U598
g11045 nand P1_U3209 P1_R1165_U24 ; P1_R1165_U599
g11046 not P1_R1165_U135 ; P1_R1165_U600
g11047 nand P1_R1165_U63 P1_R1165_U600 ; P1_R1165_U601
g11048 nand P1_R1165_U135 P1_R1165_U378 ; P1_R1165_U602
g11049 and P1_R1150_U184 P1_R1150_U201 ; P1_R1150_U6
g11050 and P1_R1150_U203 P1_R1150_U202 ; P1_R1150_U7
g11051 and P1_R1150_U179 P1_R1150_U240 ; P1_R1150_U8
g11052 and P1_R1150_U242 P1_R1150_U241 ; P1_R1150_U9
g11053 and P1_R1150_U259 P1_R1150_U258 ; P1_R1150_U10
g11054 and P1_R1150_U285 P1_R1150_U284 ; P1_R1150_U11
g11055 and P1_R1150_U383 P1_R1150_U382 ; P1_R1150_U12
g11056 nand P1_R1150_U340 P1_R1150_U343 ; P1_R1150_U13
g11057 nand P1_R1150_U329 P1_R1150_U332 ; P1_R1150_U14
g11058 nand P1_R1150_U318 P1_R1150_U321 ; P1_R1150_U15
g11059 nand P1_R1150_U310 P1_R1150_U312 ; P1_R1150_U16
g11060 nand P1_R1150_U156 P1_R1150_U175 P1_R1150_U348 ; P1_R1150_U17
g11061 nand P1_R1150_U236 P1_R1150_U238 ; P1_R1150_U18
g11062 nand P1_R1150_U228 P1_R1150_U231 ; P1_R1150_U19
g11063 nand P1_R1150_U220 P1_R1150_U222 ; P1_R1150_U20
g11064 nand P1_R1150_U25 P1_R1150_U346 ; P1_R1150_U21
g11065 not P1_U3474 ; P1_R1150_U22
g11066 not P1_U3459 ; P1_R1150_U23
g11067 not P1_U3451 ; P1_R1150_U24
g11068 nand P1_U3451 P1_R1150_U93 ; P1_R1150_U25
g11069 not P1_U3076 ; P1_R1150_U26
g11070 not P1_U3462 ; P1_R1150_U27
g11071 not P1_U3066 ; P1_R1150_U28
g11072 nand P1_U3066 P1_R1150_U23 ; P1_R1150_U29
g11073 not P1_U3062 ; P1_R1150_U30
g11074 not P1_U3471 ; P1_R1150_U31
g11075 not P1_U3468 ; P1_R1150_U32
g11076 not P1_U3465 ; P1_R1150_U33
g11077 not P1_U3069 ; P1_R1150_U34
g11078 not P1_U3065 ; P1_R1150_U35
g11079 not P1_U3058 ; P1_R1150_U36
g11080 nand P1_U3058 P1_R1150_U33 ; P1_R1150_U37
g11081 not P1_U3477 ; P1_R1150_U38
g11082 not P1_U3068 ; P1_R1150_U39
g11083 nand P1_U3068 P1_R1150_U22 ; P1_R1150_U40
g11084 not P1_U3082 ; P1_R1150_U41
g11085 not P1_U3480 ; P1_R1150_U42
g11086 not P1_U3081 ; P1_R1150_U43
g11087 nand P1_R1150_U209 P1_R1150_U208 ; P1_R1150_U44
g11088 nand P1_R1150_U37 P1_R1150_U224 ; P1_R1150_U45
g11089 nand P1_R1150_U193 P1_R1150_U192 ; P1_R1150_U46
g11090 not P1_U4009 ; P1_R1150_U47
g11091 not P1_U4013 ; P1_R1150_U48
g11092 not P1_U3498 ; P1_R1150_U49
g11093 not P1_U3486 ; P1_R1150_U50
g11094 not P1_U3483 ; P1_R1150_U51
g11095 not P1_U3061 ; P1_R1150_U52
g11096 not P1_U3060 ; P1_R1150_U53
g11097 nand P1_U3081 P1_R1150_U42 ; P1_R1150_U54
g11098 not P1_U3489 ; P1_R1150_U55
g11099 not P1_U3070 ; P1_R1150_U56
g11100 not P1_U3492 ; P1_R1150_U57
g11101 not P1_U3078 ; P1_R1150_U58
g11102 not P1_U3501 ; P1_R1150_U59
g11103 not P1_U3495 ; P1_R1150_U60
g11104 not P1_U3071 ; P1_R1150_U61
g11105 not P1_U3072 ; P1_R1150_U62
g11106 not P1_U3077 ; P1_R1150_U63
g11107 nand P1_U3077 P1_R1150_U60 ; P1_R1150_U64
g11108 not P1_U3504 ; P1_R1150_U65
g11109 not P1_U3067 ; P1_R1150_U66
g11110 nand P1_R1150_U269 P1_R1150_U268 ; P1_R1150_U67
g11111 not P1_U3080 ; P1_R1150_U68
g11112 not P1_U3509 ; P1_R1150_U69
g11113 not P1_U3079 ; P1_R1150_U70
g11114 not P1_U4015 ; P1_R1150_U71
g11115 not P1_U3074 ; P1_R1150_U72
g11116 not P1_U4012 ; P1_R1150_U73
g11117 not P1_U4014 ; P1_R1150_U74
g11118 not P1_U3064 ; P1_R1150_U75
g11119 not P1_U3059 ; P1_R1150_U76
g11120 not P1_U3073 ; P1_R1150_U77
g11121 nand P1_U3073 P1_R1150_U74 ; P1_R1150_U78
g11122 not P1_U4011 ; P1_R1150_U79
g11123 not P1_U3063 ; P1_R1150_U80
g11124 not P1_U4010 ; P1_R1150_U81
g11125 not P1_U3056 ; P1_R1150_U82
g11126 not P1_U4008 ; P1_R1150_U83
g11127 not P1_U3055 ; P1_R1150_U84
g11128 nand P1_U3055 P1_R1150_U47 ; P1_R1150_U85
g11129 not P1_U3051 ; P1_R1150_U86
g11130 not P1_U4007 ; P1_R1150_U87
g11131 not P1_U3052 ; P1_R1150_U88
g11132 nand P1_R1150_U299 P1_R1150_U298 ; P1_R1150_U89
g11133 nand P1_R1150_U78 P1_R1150_U314 ; P1_R1150_U90
g11134 nand P1_R1150_U64 P1_R1150_U325 ; P1_R1150_U91
g11135 nand P1_R1150_U54 P1_R1150_U336 ; P1_R1150_U92
g11136 not P1_U3075 ; P1_R1150_U93
g11137 nand P1_R1150_U393 P1_R1150_U392 ; P1_R1150_U94
g11138 nand P1_R1150_U407 P1_R1150_U406 ; P1_R1150_U95
g11139 nand P1_R1150_U412 P1_R1150_U411 ; P1_R1150_U96
g11140 nand P1_R1150_U428 P1_R1150_U427 ; P1_R1150_U97
g11141 nand P1_R1150_U433 P1_R1150_U432 ; P1_R1150_U98
g11142 nand P1_R1150_U438 P1_R1150_U437 ; P1_R1150_U99
g11143 nand P1_R1150_U443 P1_R1150_U442 ; P1_R1150_U100
g11144 nand P1_R1150_U448 P1_R1150_U447 ; P1_R1150_U101
g11145 nand P1_R1150_U464 P1_R1150_U463 ; P1_R1150_U102
g11146 nand P1_R1150_U469 P1_R1150_U468 ; P1_R1150_U103
g11147 nand P1_R1150_U352 P1_R1150_U351 ; P1_R1150_U104
g11148 nand P1_R1150_U361 P1_R1150_U360 ; P1_R1150_U105
g11149 nand P1_R1150_U368 P1_R1150_U367 ; P1_R1150_U106
g11150 nand P1_R1150_U372 P1_R1150_U371 ; P1_R1150_U107
g11151 nand P1_R1150_U381 P1_R1150_U380 ; P1_R1150_U108
g11152 nand P1_R1150_U402 P1_R1150_U401 ; P1_R1150_U109
g11153 nand P1_R1150_U419 P1_R1150_U418 ; P1_R1150_U110
g11154 nand P1_R1150_U423 P1_R1150_U422 ; P1_R1150_U111
g11155 nand P1_R1150_U455 P1_R1150_U454 ; P1_R1150_U112
g11156 nand P1_R1150_U459 P1_R1150_U458 ; P1_R1150_U113
g11157 nand P1_R1150_U476 P1_R1150_U475 ; P1_R1150_U114
g11158 and P1_R1150_U195 P1_R1150_U183 ; P1_R1150_U115
g11159 and P1_R1150_U198 P1_R1150_U199 ; P1_R1150_U116
g11160 and P1_R1150_U211 P1_R1150_U185 ; P1_R1150_U117
g11161 and P1_R1150_U214 P1_R1150_U215 ; P1_R1150_U118
g11162 and P1_R1150_U354 P1_R1150_U353 P1_R1150_U40 ; P1_R1150_U119
g11163 and P1_R1150_U357 P1_R1150_U185 ; P1_R1150_U120
g11164 and P1_R1150_U230 P1_R1150_U7 ; P1_R1150_U121
g11165 and P1_R1150_U364 P1_R1150_U184 ; P1_R1150_U122
g11166 and P1_R1150_U374 P1_R1150_U373 P1_R1150_U29 ; P1_R1150_U123
g11167 and P1_R1150_U377 P1_R1150_U183 ; P1_R1150_U124
g11168 and P1_R1150_U217 P1_R1150_U8 ; P1_R1150_U125
g11169 and P1_R1150_U262 P1_R1150_U180 ; P1_R1150_U126
g11170 and P1_R1150_U288 P1_R1150_U181 ; P1_R1150_U127
g11171 and P1_R1150_U304 P1_R1150_U305 ; P1_R1150_U128
g11172 and P1_R1150_U307 P1_R1150_U386 ; P1_R1150_U129
g11173 and P1_R1150_U305 P1_R1150_U304 P1_R1150_U308 ; P1_R1150_U130
g11174 nand P1_R1150_U390 P1_R1150_U389 ; P1_R1150_U131
g11175 and P1_R1150_U395 P1_R1150_U394 P1_R1150_U85 ; P1_R1150_U132
g11176 and P1_R1150_U398 P1_R1150_U182 ; P1_R1150_U133
g11177 nand P1_R1150_U404 P1_R1150_U403 ; P1_R1150_U134
g11178 nand P1_R1150_U409 P1_R1150_U408 ; P1_R1150_U135
g11179 and P1_R1150_U415 P1_R1150_U181 ; P1_R1150_U136
g11180 nand P1_R1150_U425 P1_R1150_U424 ; P1_R1150_U137
g11181 nand P1_R1150_U430 P1_R1150_U429 ; P1_R1150_U138
g11182 nand P1_R1150_U435 P1_R1150_U434 ; P1_R1150_U139
g11183 nand P1_R1150_U440 P1_R1150_U439 ; P1_R1150_U140
g11184 nand P1_R1150_U445 P1_R1150_U444 ; P1_R1150_U141
g11185 and P1_R1150_U451 P1_R1150_U180 ; P1_R1150_U142
g11186 nand P1_R1150_U461 P1_R1150_U460 ; P1_R1150_U143
g11187 nand P1_R1150_U466 P1_R1150_U465 ; P1_R1150_U144
g11188 and P1_R1150_U342 P1_R1150_U9 ; P1_R1150_U145
g11189 and P1_R1150_U472 P1_R1150_U179 ; P1_R1150_U146
g11190 and P1_R1150_U350 P1_R1150_U349 ; P1_R1150_U147
g11191 nand P1_R1150_U118 P1_R1150_U212 ; P1_R1150_U148
g11192 and P1_R1150_U359 P1_R1150_U358 ; P1_R1150_U149
g11193 and P1_R1150_U366 P1_R1150_U365 ; P1_R1150_U150
g11194 and P1_R1150_U370 P1_R1150_U369 ; P1_R1150_U151
g11195 nand P1_R1150_U116 P1_R1150_U196 ; P1_R1150_U152
g11196 and P1_R1150_U379 P1_R1150_U378 ; P1_R1150_U153
g11197 not P1_U4018 ; P1_R1150_U154
g11198 not P1_U3053 ; P1_R1150_U155
g11199 and P1_R1150_U388 P1_R1150_U387 ; P1_R1150_U156
g11200 nand P1_R1150_U128 P1_R1150_U302 ; P1_R1150_U157
g11201 and P1_R1150_U400 P1_R1150_U399 ; P1_R1150_U158
g11202 nand P1_R1150_U295 P1_R1150_U294 ; P1_R1150_U159
g11203 nand P1_R1150_U291 P1_R1150_U290 ; P1_R1150_U160
g11204 and P1_R1150_U417 P1_R1150_U416 ; P1_R1150_U161
g11205 and P1_R1150_U421 P1_R1150_U420 ; P1_R1150_U162
g11206 nand P1_R1150_U281 P1_R1150_U280 ; P1_R1150_U163
g11207 nand P1_R1150_U277 P1_R1150_U276 ; P1_R1150_U164
g11208 not P1_U3456 ; P1_R1150_U165
g11209 nand P1_R1150_U273 P1_R1150_U272 ; P1_R1150_U166
g11210 not P1_U3507 ; P1_R1150_U167
g11211 nand P1_R1150_U265 P1_R1150_U264 ; P1_R1150_U168
g11212 and P1_R1150_U453 P1_R1150_U452 ; P1_R1150_U169
g11213 and P1_R1150_U457 P1_R1150_U456 ; P1_R1150_U170
g11214 nand P1_R1150_U255 P1_R1150_U254 ; P1_R1150_U171
g11215 nand P1_R1150_U251 P1_R1150_U250 ; P1_R1150_U172
g11216 nand P1_R1150_U247 P1_R1150_U246 ; P1_R1150_U173
g11217 and P1_R1150_U474 P1_R1150_U473 ; P1_R1150_U174
g11218 nand P1_R1150_U129 P1_R1150_U157 ; P1_R1150_U175
g11219 not P1_R1150_U85 ; P1_R1150_U176
g11220 not P1_R1150_U29 ; P1_R1150_U177
g11221 not P1_R1150_U40 ; P1_R1150_U178
g11222 nand P1_U3483 P1_R1150_U53 ; P1_R1150_U179
g11223 nand P1_U3498 P1_R1150_U62 ; P1_R1150_U180
g11224 nand P1_U4013 P1_R1150_U76 ; P1_R1150_U181
g11225 nand P1_U4009 P1_R1150_U84 ; P1_R1150_U182
g11226 nand P1_U3459 P1_R1150_U28 ; P1_R1150_U183
g11227 nand P1_U3468 P1_R1150_U35 ; P1_R1150_U184
g11228 nand P1_U3474 P1_R1150_U39 ; P1_R1150_U185
g11229 not P1_R1150_U64 ; P1_R1150_U186
g11230 not P1_R1150_U78 ; P1_R1150_U187
g11231 not P1_R1150_U37 ; P1_R1150_U188
g11232 not P1_R1150_U54 ; P1_R1150_U189
g11233 not P1_R1150_U25 ; P1_R1150_U190
g11234 nand P1_R1150_U190 P1_R1150_U26 ; P1_R1150_U191
g11235 nand P1_R1150_U191 P1_R1150_U165 ; P1_R1150_U192
g11236 nand P1_U3076 P1_R1150_U25 ; P1_R1150_U193
g11237 not P1_R1150_U46 ; P1_R1150_U194
g11238 nand P1_U3462 P1_R1150_U30 ; P1_R1150_U195
g11239 nand P1_R1150_U115 P1_R1150_U46 ; P1_R1150_U196
g11240 nand P1_R1150_U30 P1_R1150_U29 ; P1_R1150_U197
g11241 nand P1_R1150_U197 P1_R1150_U27 ; P1_R1150_U198
g11242 nand P1_U3062 P1_R1150_U177 ; P1_R1150_U199
g11243 not P1_R1150_U152 ; P1_R1150_U200
g11244 nand P1_U3471 P1_R1150_U34 ; P1_R1150_U201
g11245 nand P1_U3069 P1_R1150_U31 ; P1_R1150_U202
g11246 nand P1_U3065 P1_R1150_U32 ; P1_R1150_U203
g11247 nand P1_R1150_U188 P1_R1150_U6 ; P1_R1150_U204
g11248 nand P1_R1150_U7 P1_R1150_U204 ; P1_R1150_U205
g11249 nand P1_U3465 P1_R1150_U36 ; P1_R1150_U206
g11250 nand P1_U3471 P1_R1150_U34 ; P1_R1150_U207
g11251 nand P1_R1150_U206 P1_R1150_U152 P1_R1150_U6 ; P1_R1150_U208
g11252 nand P1_R1150_U207 P1_R1150_U205 ; P1_R1150_U209
g11253 not P1_R1150_U44 ; P1_R1150_U210
g11254 nand P1_U3477 P1_R1150_U41 ; P1_R1150_U211
g11255 nand P1_R1150_U117 P1_R1150_U44 ; P1_R1150_U212
g11256 nand P1_R1150_U41 P1_R1150_U40 ; P1_R1150_U213
g11257 nand P1_R1150_U213 P1_R1150_U38 ; P1_R1150_U214
g11258 nand P1_U3082 P1_R1150_U178 ; P1_R1150_U215
g11259 not P1_R1150_U148 ; P1_R1150_U216
g11260 nand P1_U3480 P1_R1150_U43 ; P1_R1150_U217
g11261 nand P1_R1150_U217 P1_R1150_U54 ; P1_R1150_U218
g11262 nand P1_R1150_U210 P1_R1150_U40 ; P1_R1150_U219
g11263 nand P1_R1150_U120 P1_R1150_U219 ; P1_R1150_U220
g11264 nand P1_R1150_U44 P1_R1150_U185 ; P1_R1150_U221
g11265 nand P1_R1150_U119 P1_R1150_U221 ; P1_R1150_U222
g11266 nand P1_R1150_U40 P1_R1150_U185 ; P1_R1150_U223
g11267 nand P1_R1150_U206 P1_R1150_U152 ; P1_R1150_U224
g11268 not P1_R1150_U45 ; P1_R1150_U225
g11269 nand P1_U3065 P1_R1150_U32 ; P1_R1150_U226
g11270 nand P1_R1150_U225 P1_R1150_U226 ; P1_R1150_U227
g11271 nand P1_R1150_U122 P1_R1150_U227 ; P1_R1150_U228
g11272 nand P1_R1150_U45 P1_R1150_U184 ; P1_R1150_U229
g11273 nand P1_U3471 P1_R1150_U34 ; P1_R1150_U230
g11274 nand P1_R1150_U121 P1_R1150_U229 ; P1_R1150_U231
g11275 nand P1_U3065 P1_R1150_U32 ; P1_R1150_U232
g11276 nand P1_R1150_U184 P1_R1150_U232 ; P1_R1150_U233
g11277 nand P1_R1150_U206 P1_R1150_U37 ; P1_R1150_U234
g11278 nand P1_R1150_U194 P1_R1150_U29 ; P1_R1150_U235
g11279 nand P1_R1150_U124 P1_R1150_U235 ; P1_R1150_U236
g11280 nand P1_R1150_U46 P1_R1150_U183 ; P1_R1150_U237
g11281 nand P1_R1150_U123 P1_R1150_U237 ; P1_R1150_U238
g11282 nand P1_R1150_U29 P1_R1150_U183 ; P1_R1150_U239
g11283 nand P1_U3486 P1_R1150_U52 ; P1_R1150_U240
g11284 nand P1_U3061 P1_R1150_U50 ; P1_R1150_U241
g11285 nand P1_U3060 P1_R1150_U51 ; P1_R1150_U242
g11286 nand P1_R1150_U189 P1_R1150_U8 ; P1_R1150_U243
g11287 nand P1_R1150_U9 P1_R1150_U243 ; P1_R1150_U244
g11288 nand P1_U3486 P1_R1150_U52 ; P1_R1150_U245
g11289 nand P1_R1150_U125 P1_R1150_U148 ; P1_R1150_U246
g11290 nand P1_R1150_U245 P1_R1150_U244 ; P1_R1150_U247
g11291 not P1_R1150_U173 ; P1_R1150_U248
g11292 nand P1_U3489 P1_R1150_U56 ; P1_R1150_U249
g11293 nand P1_R1150_U249 P1_R1150_U173 ; P1_R1150_U250
g11294 nand P1_U3070 P1_R1150_U55 ; P1_R1150_U251
g11295 not P1_R1150_U172 ; P1_R1150_U252
g11296 nand P1_U3492 P1_R1150_U58 ; P1_R1150_U253
g11297 nand P1_R1150_U253 P1_R1150_U172 ; P1_R1150_U254
g11298 nand P1_U3078 P1_R1150_U57 ; P1_R1150_U255
g11299 not P1_R1150_U171 ; P1_R1150_U256
g11300 nand P1_U3501 P1_R1150_U61 ; P1_R1150_U257
g11301 nand P1_U3071 P1_R1150_U59 ; P1_R1150_U258
g11302 nand P1_U3072 P1_R1150_U49 ; P1_R1150_U259
g11303 nand P1_R1150_U186 P1_R1150_U180 ; P1_R1150_U260
g11304 nand P1_R1150_U10 P1_R1150_U260 ; P1_R1150_U261
g11305 nand P1_U3495 P1_R1150_U63 ; P1_R1150_U262
g11306 nand P1_U3501 P1_R1150_U61 ; P1_R1150_U263
g11307 nand P1_R1150_U171 P1_R1150_U126 P1_R1150_U257 ; P1_R1150_U264
g11308 nand P1_R1150_U263 P1_R1150_U261 ; P1_R1150_U265
g11309 not P1_R1150_U168 ; P1_R1150_U266
g11310 nand P1_U3504 P1_R1150_U66 ; P1_R1150_U267
g11311 nand P1_R1150_U267 P1_R1150_U168 ; P1_R1150_U268
g11312 nand P1_U3067 P1_R1150_U65 ; P1_R1150_U269
g11313 not P1_R1150_U67 ; P1_R1150_U270
g11314 nand P1_R1150_U270 P1_R1150_U68 ; P1_R1150_U271
g11315 nand P1_R1150_U271 P1_R1150_U167 ; P1_R1150_U272
g11316 nand P1_U3080 P1_R1150_U67 ; P1_R1150_U273
g11317 not P1_R1150_U166 ; P1_R1150_U274
g11318 nand P1_U3509 P1_R1150_U70 ; P1_R1150_U275
g11319 nand P1_R1150_U275 P1_R1150_U166 ; P1_R1150_U276
g11320 nand P1_U3079 P1_R1150_U69 ; P1_R1150_U277
g11321 not P1_R1150_U164 ; P1_R1150_U278
g11322 nand P1_U4015 P1_R1150_U72 ; P1_R1150_U279
g11323 nand P1_R1150_U279 P1_R1150_U164 ; P1_R1150_U280
g11324 nand P1_U3074 P1_R1150_U71 ; P1_R1150_U281
g11325 not P1_R1150_U163 ; P1_R1150_U282
g11326 nand P1_U4012 P1_R1150_U75 ; P1_R1150_U283
g11327 nand P1_U3064 P1_R1150_U73 ; P1_R1150_U284
g11328 nand P1_U3059 P1_R1150_U48 ; P1_R1150_U285
g11329 nand P1_R1150_U187 P1_R1150_U181 ; P1_R1150_U286
g11330 nand P1_R1150_U11 P1_R1150_U286 ; P1_R1150_U287
g11331 nand P1_U4014 P1_R1150_U77 ; P1_R1150_U288
g11332 nand P1_U4012 P1_R1150_U75 ; P1_R1150_U289
g11333 nand P1_R1150_U163 P1_R1150_U127 P1_R1150_U283 ; P1_R1150_U290
g11334 nand P1_R1150_U289 P1_R1150_U287 ; P1_R1150_U291
g11335 not P1_R1150_U160 ; P1_R1150_U292
g11336 nand P1_U4011 P1_R1150_U80 ; P1_R1150_U293
g11337 nand P1_R1150_U293 P1_R1150_U160 ; P1_R1150_U294
g11338 nand P1_U3063 P1_R1150_U79 ; P1_R1150_U295
g11339 not P1_R1150_U159 ; P1_R1150_U296
g11340 nand P1_U4010 P1_R1150_U82 ; P1_R1150_U297
g11341 nand P1_R1150_U297 P1_R1150_U159 ; P1_R1150_U298
g11342 nand P1_U3056 P1_R1150_U81 ; P1_R1150_U299
g11343 not P1_R1150_U89 ; P1_R1150_U300
g11344 nand P1_U4008 P1_R1150_U86 ; P1_R1150_U301
g11345 nand P1_R1150_U89 P1_R1150_U182 P1_R1150_U301 ; P1_R1150_U302
g11346 nand P1_R1150_U86 P1_R1150_U85 ; P1_R1150_U303
g11347 nand P1_R1150_U303 P1_R1150_U83 ; P1_R1150_U304
g11348 nand P1_U3051 P1_R1150_U176 ; P1_R1150_U305
g11349 not P1_R1150_U157 ; P1_R1150_U306
g11350 nand P1_U4007 P1_R1150_U88 ; P1_R1150_U307
g11351 nand P1_U3052 P1_R1150_U87 ; P1_R1150_U308
g11352 nand P1_R1150_U300 P1_R1150_U85 ; P1_R1150_U309
g11353 nand P1_R1150_U133 P1_R1150_U309 ; P1_R1150_U310
g11354 nand P1_R1150_U89 P1_R1150_U182 ; P1_R1150_U311
g11355 nand P1_R1150_U132 P1_R1150_U311 ; P1_R1150_U312
g11356 nand P1_R1150_U85 P1_R1150_U182 ; P1_R1150_U313
g11357 nand P1_R1150_U288 P1_R1150_U163 ; P1_R1150_U314
g11358 not P1_R1150_U90 ; P1_R1150_U315
g11359 nand P1_U3059 P1_R1150_U48 ; P1_R1150_U316
g11360 nand P1_R1150_U315 P1_R1150_U316 ; P1_R1150_U317
g11361 nand P1_R1150_U136 P1_R1150_U317 ; P1_R1150_U318
g11362 nand P1_R1150_U90 P1_R1150_U181 ; P1_R1150_U319
g11363 nand P1_U4012 P1_R1150_U75 ; P1_R1150_U320
g11364 nand P1_R1150_U320 P1_R1150_U319 P1_R1150_U11 ; P1_R1150_U321
g11365 nand P1_U3059 P1_R1150_U48 ; P1_R1150_U322
g11366 nand P1_R1150_U181 P1_R1150_U322 ; P1_R1150_U323
g11367 nand P1_R1150_U288 P1_R1150_U78 ; P1_R1150_U324
g11368 nand P1_R1150_U262 P1_R1150_U171 ; P1_R1150_U325
g11369 not P1_R1150_U91 ; P1_R1150_U326
g11370 nand P1_U3072 P1_R1150_U49 ; P1_R1150_U327
g11371 nand P1_R1150_U326 P1_R1150_U327 ; P1_R1150_U328
g11372 nand P1_R1150_U142 P1_R1150_U328 ; P1_R1150_U329
g11373 nand P1_R1150_U91 P1_R1150_U180 ; P1_R1150_U330
g11374 nand P1_U3501 P1_R1150_U61 ; P1_R1150_U331
g11375 nand P1_R1150_U331 P1_R1150_U330 P1_R1150_U10 ; P1_R1150_U332
g11376 nand P1_U3072 P1_R1150_U49 ; P1_R1150_U333
g11377 nand P1_R1150_U180 P1_R1150_U333 ; P1_R1150_U334
g11378 nand P1_R1150_U262 P1_R1150_U64 ; P1_R1150_U335
g11379 nand P1_R1150_U217 P1_R1150_U148 ; P1_R1150_U336
g11380 not P1_R1150_U92 ; P1_R1150_U337
g11381 nand P1_U3060 P1_R1150_U51 ; P1_R1150_U338
g11382 nand P1_R1150_U337 P1_R1150_U338 ; P1_R1150_U339
g11383 nand P1_R1150_U146 P1_R1150_U339 ; P1_R1150_U340
g11384 nand P1_R1150_U92 P1_R1150_U179 ; P1_R1150_U341
g11385 nand P1_U3486 P1_R1150_U52 ; P1_R1150_U342
g11386 nand P1_R1150_U145 P1_R1150_U341 ; P1_R1150_U343
g11387 nand P1_U3060 P1_R1150_U51 ; P1_R1150_U344
g11388 nand P1_R1150_U179 P1_R1150_U344 ; P1_R1150_U345
g11389 nand P1_U3075 P1_R1150_U24 ; P1_R1150_U346
g11390 nand P1_R1150_U89 P1_R1150_U182 P1_R1150_U301 ; P1_R1150_U347
g11391 nand P1_R1150_U12 P1_R1150_U347 P1_R1150_U130 ; P1_R1150_U348
g11392 nand P1_U3480 P1_R1150_U43 ; P1_R1150_U349
g11393 nand P1_U3081 P1_R1150_U42 ; P1_R1150_U350
g11394 nand P1_R1150_U218 P1_R1150_U148 ; P1_R1150_U351
g11395 nand P1_R1150_U216 P1_R1150_U147 ; P1_R1150_U352
g11396 nand P1_U3477 P1_R1150_U41 ; P1_R1150_U353
g11397 nand P1_U3082 P1_R1150_U38 ; P1_R1150_U354
g11398 nand P1_U3477 P1_R1150_U41 ; P1_R1150_U355
g11399 nand P1_U3082 P1_R1150_U38 ; P1_R1150_U356
g11400 nand P1_R1150_U356 P1_R1150_U355 ; P1_R1150_U357
g11401 nand P1_U3474 P1_R1150_U39 ; P1_R1150_U358
g11402 nand P1_U3068 P1_R1150_U22 ; P1_R1150_U359
g11403 nand P1_R1150_U223 P1_R1150_U44 ; P1_R1150_U360
g11404 nand P1_R1150_U149 P1_R1150_U210 ; P1_R1150_U361
g11405 nand P1_U3471 P1_R1150_U34 ; P1_R1150_U362
g11406 nand P1_U3069 P1_R1150_U31 ; P1_R1150_U363
g11407 nand P1_R1150_U363 P1_R1150_U362 ; P1_R1150_U364
g11408 nand P1_U3468 P1_R1150_U35 ; P1_R1150_U365
g11409 nand P1_U3065 P1_R1150_U32 ; P1_R1150_U366
g11410 nand P1_R1150_U233 P1_R1150_U45 ; P1_R1150_U367
g11411 nand P1_R1150_U150 P1_R1150_U225 ; P1_R1150_U368
g11412 nand P1_U3465 P1_R1150_U36 ; P1_R1150_U369
g11413 nand P1_U3058 P1_R1150_U33 ; P1_R1150_U370
g11414 nand P1_R1150_U234 P1_R1150_U152 ; P1_R1150_U371
g11415 nand P1_R1150_U200 P1_R1150_U151 ; P1_R1150_U372
g11416 nand P1_U3462 P1_R1150_U30 ; P1_R1150_U373
g11417 nand P1_U3062 P1_R1150_U27 ; P1_R1150_U374
g11418 nand P1_U3462 P1_R1150_U30 ; P1_R1150_U375
g11419 nand P1_U3062 P1_R1150_U27 ; P1_R1150_U376
g11420 nand P1_R1150_U376 P1_R1150_U375 ; P1_R1150_U377
g11421 nand P1_U3459 P1_R1150_U28 ; P1_R1150_U378
g11422 nand P1_U3066 P1_R1150_U23 ; P1_R1150_U379
g11423 nand P1_R1150_U239 P1_R1150_U46 ; P1_R1150_U380
g11424 nand P1_R1150_U153 P1_R1150_U194 ; P1_R1150_U381
g11425 nand P1_U4018 P1_R1150_U155 ; P1_R1150_U382
g11426 nand P1_U3053 P1_R1150_U154 ; P1_R1150_U383
g11427 nand P1_U4018 P1_R1150_U155 ; P1_R1150_U384
g11428 nand P1_U3053 P1_R1150_U154 ; P1_R1150_U385
g11429 nand P1_R1150_U385 P1_R1150_U384 ; P1_R1150_U386
g11430 nand P1_U3052 P1_R1150_U386 P1_R1150_U87 ; P1_R1150_U387
g11431 nand P1_R1150_U12 P1_R1150_U88 P1_U4007 ; P1_R1150_U388
g11432 nand P1_U4007 P1_R1150_U88 ; P1_R1150_U389
g11433 nand P1_U3052 P1_R1150_U87 ; P1_R1150_U390
g11434 not P1_R1150_U131 ; P1_R1150_U391
g11435 nand P1_R1150_U306 P1_R1150_U391 ; P1_R1150_U392
g11436 nand P1_R1150_U131 P1_R1150_U157 ; P1_R1150_U393
g11437 nand P1_U4008 P1_R1150_U86 ; P1_R1150_U394
g11438 nand P1_U3051 P1_R1150_U83 ; P1_R1150_U395
g11439 nand P1_U4008 P1_R1150_U86 ; P1_R1150_U396
g11440 nand P1_U3051 P1_R1150_U83 ; P1_R1150_U397
g11441 nand P1_R1150_U397 P1_R1150_U396 ; P1_R1150_U398
g11442 nand P1_U4009 P1_R1150_U84 ; P1_R1150_U399
g11443 nand P1_U3055 P1_R1150_U47 ; P1_R1150_U400
g11444 nand P1_R1150_U313 P1_R1150_U89 ; P1_R1150_U401
g11445 nand P1_R1150_U158 P1_R1150_U300 ; P1_R1150_U402
g11446 nand P1_U4010 P1_R1150_U82 ; P1_R1150_U403
g11447 nand P1_U3056 P1_R1150_U81 ; P1_R1150_U404
g11448 not P1_R1150_U134 ; P1_R1150_U405
g11449 nand P1_R1150_U296 P1_R1150_U405 ; P1_R1150_U406
g11450 nand P1_R1150_U134 P1_R1150_U159 ; P1_R1150_U407
g11451 nand P1_U4011 P1_R1150_U80 ; P1_R1150_U408
g11452 nand P1_U3063 P1_R1150_U79 ; P1_R1150_U409
g11453 not P1_R1150_U135 ; P1_R1150_U410
g11454 nand P1_R1150_U292 P1_R1150_U410 ; P1_R1150_U411
g11455 nand P1_R1150_U135 P1_R1150_U160 ; P1_R1150_U412
g11456 nand P1_U4012 P1_R1150_U75 ; P1_R1150_U413
g11457 nand P1_U3064 P1_R1150_U73 ; P1_R1150_U414
g11458 nand P1_R1150_U414 P1_R1150_U413 ; P1_R1150_U415
g11459 nand P1_U4013 P1_R1150_U76 ; P1_R1150_U416
g11460 nand P1_U3059 P1_R1150_U48 ; P1_R1150_U417
g11461 nand P1_R1150_U323 P1_R1150_U90 ; P1_R1150_U418
g11462 nand P1_R1150_U161 P1_R1150_U315 ; P1_R1150_U419
g11463 nand P1_U4014 P1_R1150_U77 ; P1_R1150_U420
g11464 nand P1_U3073 P1_R1150_U74 ; P1_R1150_U421
g11465 nand P1_R1150_U324 P1_R1150_U163 ; P1_R1150_U422
g11466 nand P1_R1150_U282 P1_R1150_U162 ; P1_R1150_U423
g11467 nand P1_U4015 P1_R1150_U72 ; P1_R1150_U424
g11468 nand P1_U3074 P1_R1150_U71 ; P1_R1150_U425
g11469 not P1_R1150_U137 ; P1_R1150_U426
g11470 nand P1_R1150_U278 P1_R1150_U426 ; P1_R1150_U427
g11471 nand P1_R1150_U137 P1_R1150_U164 ; P1_R1150_U428
g11472 nand P1_U3456 P1_R1150_U26 ; P1_R1150_U429
g11473 nand P1_U3076 P1_R1150_U165 ; P1_R1150_U430
g11474 not P1_R1150_U138 ; P1_R1150_U431
g11475 nand P1_R1150_U431 P1_R1150_U190 ; P1_R1150_U432
g11476 nand P1_R1150_U138 P1_R1150_U25 ; P1_R1150_U433
g11477 nand P1_U3509 P1_R1150_U70 ; P1_R1150_U434
g11478 nand P1_U3079 P1_R1150_U69 ; P1_R1150_U435
g11479 not P1_R1150_U139 ; P1_R1150_U436
g11480 nand P1_R1150_U274 P1_R1150_U436 ; P1_R1150_U437
g11481 nand P1_R1150_U139 P1_R1150_U166 ; P1_R1150_U438
g11482 nand P1_U3507 P1_R1150_U68 ; P1_R1150_U439
g11483 nand P1_U3080 P1_R1150_U167 ; P1_R1150_U440
g11484 not P1_R1150_U140 ; P1_R1150_U441
g11485 nand P1_R1150_U441 P1_R1150_U270 ; P1_R1150_U442
g11486 nand P1_R1150_U140 P1_R1150_U67 ; P1_R1150_U443
g11487 nand P1_U3504 P1_R1150_U66 ; P1_R1150_U444
g11488 nand P1_U3067 P1_R1150_U65 ; P1_R1150_U445
g11489 not P1_R1150_U141 ; P1_R1150_U446
g11490 nand P1_R1150_U266 P1_R1150_U446 ; P1_R1150_U447
g11491 nand P1_R1150_U141 P1_R1150_U168 ; P1_R1150_U448
g11492 nand P1_U3501 P1_R1150_U61 ; P1_R1150_U449
g11493 nand P1_U3071 P1_R1150_U59 ; P1_R1150_U450
g11494 nand P1_R1150_U450 P1_R1150_U449 ; P1_R1150_U451
g11495 nand P1_U3498 P1_R1150_U62 ; P1_R1150_U452
g11496 nand P1_U3072 P1_R1150_U49 ; P1_R1150_U453
g11497 nand P1_R1150_U334 P1_R1150_U91 ; P1_R1150_U454
g11498 nand P1_R1150_U169 P1_R1150_U326 ; P1_R1150_U455
g11499 nand P1_U3495 P1_R1150_U63 ; P1_R1150_U456
g11500 nand P1_U3077 P1_R1150_U60 ; P1_R1150_U457
g11501 nand P1_R1150_U335 P1_R1150_U171 ; P1_R1150_U458
g11502 nand P1_R1150_U256 P1_R1150_U170 ; P1_R1150_U459
g11503 nand P1_U3492 P1_R1150_U58 ; P1_R1150_U460
g11504 nand P1_U3078 P1_R1150_U57 ; P1_R1150_U461
g11505 not P1_R1150_U143 ; P1_R1150_U462
g11506 nand P1_R1150_U252 P1_R1150_U462 ; P1_R1150_U463
g11507 nand P1_R1150_U143 P1_R1150_U172 ; P1_R1150_U464
g11508 nand P1_U3489 P1_R1150_U56 ; P1_R1150_U465
g11509 nand P1_U3070 P1_R1150_U55 ; P1_R1150_U466
g11510 not P1_R1150_U144 ; P1_R1150_U467
g11511 nand P1_R1150_U248 P1_R1150_U467 ; P1_R1150_U468
g11512 nand P1_R1150_U144 P1_R1150_U173 ; P1_R1150_U469
g11513 nand P1_U3486 P1_R1150_U52 ; P1_R1150_U470
g11514 nand P1_U3061 P1_R1150_U50 ; P1_R1150_U471
g11515 nand P1_R1150_U471 P1_R1150_U470 ; P1_R1150_U472
g11516 nand P1_U3483 P1_R1150_U53 ; P1_R1150_U473
g11517 nand P1_U3060 P1_R1150_U51 ; P1_R1150_U474
g11518 nand P1_R1150_U345 P1_R1150_U92 ; P1_R1150_U475
g11519 nand P1_R1150_U174 P1_R1150_U337 ; P1_R1150_U476
g11520 and P1_R1192_U184 P1_R1192_U201 ; P1_R1192_U6
g11521 and P1_R1192_U203 P1_R1192_U202 ; P1_R1192_U7
g11522 and P1_R1192_U179 P1_R1192_U240 ; P1_R1192_U8
g11523 and P1_R1192_U242 P1_R1192_U241 ; P1_R1192_U9
g11524 and P1_R1192_U259 P1_R1192_U258 ; P1_R1192_U10
g11525 and P1_R1192_U285 P1_R1192_U284 ; P1_R1192_U11
g11526 and P1_R1192_U383 P1_R1192_U382 ; P1_R1192_U12
g11527 nand P1_R1192_U340 P1_R1192_U343 ; P1_R1192_U13
g11528 nand P1_R1192_U329 P1_R1192_U332 ; P1_R1192_U14
g11529 nand P1_R1192_U318 P1_R1192_U321 ; P1_R1192_U15
g11530 nand P1_R1192_U310 P1_R1192_U312 ; P1_R1192_U16
g11531 nand P1_R1192_U156 P1_R1192_U175 P1_R1192_U348 ; P1_R1192_U17
g11532 nand P1_R1192_U236 P1_R1192_U238 ; P1_R1192_U18
g11533 nand P1_R1192_U228 P1_R1192_U231 ; P1_R1192_U19
g11534 nand P1_R1192_U220 P1_R1192_U222 ; P1_R1192_U20
g11535 nand P1_R1192_U25 P1_R1192_U346 ; P1_R1192_U21
g11536 not P1_U3474 ; P1_R1192_U22
g11537 not P1_U3459 ; P1_R1192_U23
g11538 not P1_U3451 ; P1_R1192_U24
g11539 nand P1_U3451 P1_R1192_U93 ; P1_R1192_U25
g11540 not P1_U3076 ; P1_R1192_U26
g11541 not P1_U3462 ; P1_R1192_U27
g11542 not P1_U3066 ; P1_R1192_U28
g11543 nand P1_U3066 P1_R1192_U23 ; P1_R1192_U29
g11544 not P1_U3062 ; P1_R1192_U30
g11545 not P1_U3471 ; P1_R1192_U31
g11546 not P1_U3468 ; P1_R1192_U32
g11547 not P1_U3465 ; P1_R1192_U33
g11548 not P1_U3069 ; P1_R1192_U34
g11549 not P1_U3065 ; P1_R1192_U35
g11550 not P1_U3058 ; P1_R1192_U36
g11551 nand P1_U3058 P1_R1192_U33 ; P1_R1192_U37
g11552 not P1_U3477 ; P1_R1192_U38
g11553 not P1_U3068 ; P1_R1192_U39
g11554 nand P1_U3068 P1_R1192_U22 ; P1_R1192_U40
g11555 not P1_U3082 ; P1_R1192_U41
g11556 not P1_U3480 ; P1_R1192_U42
g11557 not P1_U3081 ; P1_R1192_U43
g11558 nand P1_R1192_U209 P1_R1192_U208 ; P1_R1192_U44
g11559 nand P1_R1192_U37 P1_R1192_U224 ; P1_R1192_U45
g11560 nand P1_R1192_U193 P1_R1192_U192 ; P1_R1192_U46
g11561 not P1_U4009 ; P1_R1192_U47
g11562 not P1_U4013 ; P1_R1192_U48
g11563 not P1_U3498 ; P1_R1192_U49
g11564 not P1_U3486 ; P1_R1192_U50
g11565 not P1_U3483 ; P1_R1192_U51
g11566 not P1_U3061 ; P1_R1192_U52
g11567 not P1_U3060 ; P1_R1192_U53
g11568 nand P1_U3081 P1_R1192_U42 ; P1_R1192_U54
g11569 not P1_U3489 ; P1_R1192_U55
g11570 not P1_U3070 ; P1_R1192_U56
g11571 not P1_U3492 ; P1_R1192_U57
g11572 not P1_U3078 ; P1_R1192_U58
g11573 not P1_U3501 ; P1_R1192_U59
g11574 not P1_U3495 ; P1_R1192_U60
g11575 not P1_U3071 ; P1_R1192_U61
g11576 not P1_U3072 ; P1_R1192_U62
g11577 not P1_U3077 ; P1_R1192_U63
g11578 nand P1_U3077 P1_R1192_U60 ; P1_R1192_U64
g11579 not P1_U3504 ; P1_R1192_U65
g11580 not P1_U3067 ; P1_R1192_U66
g11581 nand P1_R1192_U269 P1_R1192_U268 ; P1_R1192_U67
g11582 not P1_U3080 ; P1_R1192_U68
g11583 not P1_U3509 ; P1_R1192_U69
g11584 not P1_U3079 ; P1_R1192_U70
g11585 not P1_U4015 ; P1_R1192_U71
g11586 not P1_U3074 ; P1_R1192_U72
g11587 not P1_U4012 ; P1_R1192_U73
g11588 not P1_U4014 ; P1_R1192_U74
g11589 not P1_U3064 ; P1_R1192_U75
g11590 not P1_U3059 ; P1_R1192_U76
g11591 not P1_U3073 ; P1_R1192_U77
g11592 nand P1_U3073 P1_R1192_U74 ; P1_R1192_U78
g11593 not P1_U4011 ; P1_R1192_U79
g11594 not P1_U3063 ; P1_R1192_U80
g11595 not P1_U4010 ; P1_R1192_U81
g11596 not P1_U3056 ; P1_R1192_U82
g11597 not P1_U4008 ; P1_R1192_U83
g11598 not P1_U3055 ; P1_R1192_U84
g11599 nand P1_U3055 P1_R1192_U47 ; P1_R1192_U85
g11600 not P1_U3051 ; P1_R1192_U86
g11601 not P1_U4007 ; P1_R1192_U87
g11602 not P1_U3052 ; P1_R1192_U88
g11603 nand P1_R1192_U299 P1_R1192_U298 ; P1_R1192_U89
g11604 nand P1_R1192_U78 P1_R1192_U314 ; P1_R1192_U90
g11605 nand P1_R1192_U64 P1_R1192_U325 ; P1_R1192_U91
g11606 nand P1_R1192_U54 P1_R1192_U336 ; P1_R1192_U92
g11607 not P1_U3075 ; P1_R1192_U93
g11608 nand P1_R1192_U393 P1_R1192_U392 ; P1_R1192_U94
g11609 nand P1_R1192_U407 P1_R1192_U406 ; P1_R1192_U95
g11610 nand P1_R1192_U412 P1_R1192_U411 ; P1_R1192_U96
g11611 nand P1_R1192_U428 P1_R1192_U427 ; P1_R1192_U97
g11612 nand P1_R1192_U433 P1_R1192_U432 ; P1_R1192_U98
g11613 nand P1_R1192_U438 P1_R1192_U437 ; P1_R1192_U99
g11614 nand P1_R1192_U443 P1_R1192_U442 ; P1_R1192_U100
g11615 nand P1_R1192_U448 P1_R1192_U447 ; P1_R1192_U101
g11616 nand P1_R1192_U464 P1_R1192_U463 ; P1_R1192_U102
g11617 nand P1_R1192_U469 P1_R1192_U468 ; P1_R1192_U103
g11618 nand P1_R1192_U352 P1_R1192_U351 ; P1_R1192_U104
g11619 nand P1_R1192_U361 P1_R1192_U360 ; P1_R1192_U105
g11620 nand P1_R1192_U368 P1_R1192_U367 ; P1_R1192_U106
g11621 nand P1_R1192_U372 P1_R1192_U371 ; P1_R1192_U107
g11622 nand P1_R1192_U381 P1_R1192_U380 ; P1_R1192_U108
g11623 nand P1_R1192_U402 P1_R1192_U401 ; P1_R1192_U109
g11624 nand P1_R1192_U419 P1_R1192_U418 ; P1_R1192_U110
g11625 nand P1_R1192_U423 P1_R1192_U422 ; P1_R1192_U111
g11626 nand P1_R1192_U455 P1_R1192_U454 ; P1_R1192_U112
g11627 nand P1_R1192_U459 P1_R1192_U458 ; P1_R1192_U113
g11628 nand P1_R1192_U476 P1_R1192_U475 ; P1_R1192_U114
g11629 and P1_R1192_U195 P1_R1192_U183 ; P1_R1192_U115
g11630 and P1_R1192_U198 P1_R1192_U199 ; P1_R1192_U116
g11631 and P1_R1192_U211 P1_R1192_U185 ; P1_R1192_U117
g11632 and P1_R1192_U214 P1_R1192_U215 ; P1_R1192_U118
g11633 and P1_R1192_U354 P1_R1192_U353 P1_R1192_U40 ; P1_R1192_U119
g11634 and P1_R1192_U357 P1_R1192_U185 ; P1_R1192_U120
g11635 and P1_R1192_U230 P1_R1192_U7 ; P1_R1192_U121
g11636 and P1_R1192_U364 P1_R1192_U184 ; P1_R1192_U122
g11637 and P1_R1192_U374 P1_R1192_U373 P1_R1192_U29 ; P1_R1192_U123
g11638 and P1_R1192_U377 P1_R1192_U183 ; P1_R1192_U124
g11639 and P1_R1192_U217 P1_R1192_U8 ; P1_R1192_U125
g11640 and P1_R1192_U262 P1_R1192_U180 ; P1_R1192_U126
g11641 and P1_R1192_U288 P1_R1192_U181 ; P1_R1192_U127
g11642 and P1_R1192_U304 P1_R1192_U305 ; P1_R1192_U128
g11643 and P1_R1192_U307 P1_R1192_U386 ; P1_R1192_U129
g11644 and P1_R1192_U305 P1_R1192_U304 P1_R1192_U308 ; P1_R1192_U130
g11645 nand P1_R1192_U390 P1_R1192_U389 ; P1_R1192_U131
g11646 and P1_R1192_U395 P1_R1192_U394 P1_R1192_U85 ; P1_R1192_U132
g11647 and P1_R1192_U398 P1_R1192_U182 ; P1_R1192_U133
g11648 nand P1_R1192_U404 P1_R1192_U403 ; P1_R1192_U134
g11649 nand P1_R1192_U409 P1_R1192_U408 ; P1_R1192_U135
g11650 and P1_R1192_U415 P1_R1192_U181 ; P1_R1192_U136
g11651 nand P1_R1192_U425 P1_R1192_U424 ; P1_R1192_U137
g11652 nand P1_R1192_U430 P1_R1192_U429 ; P1_R1192_U138
g11653 nand P1_R1192_U435 P1_R1192_U434 ; P1_R1192_U139
g11654 nand P1_R1192_U440 P1_R1192_U439 ; P1_R1192_U140
g11655 nand P1_R1192_U445 P1_R1192_U444 ; P1_R1192_U141
g11656 and P1_R1192_U451 P1_R1192_U180 ; P1_R1192_U142
g11657 nand P1_R1192_U461 P1_R1192_U460 ; P1_R1192_U143
g11658 nand P1_R1192_U466 P1_R1192_U465 ; P1_R1192_U144
g11659 and P1_R1192_U342 P1_R1192_U9 ; P1_R1192_U145
g11660 and P1_R1192_U472 P1_R1192_U179 ; P1_R1192_U146
g11661 and P1_R1192_U350 P1_R1192_U349 ; P1_R1192_U147
g11662 nand P1_R1192_U118 P1_R1192_U212 ; P1_R1192_U148
g11663 and P1_R1192_U359 P1_R1192_U358 ; P1_R1192_U149
g11664 and P1_R1192_U366 P1_R1192_U365 ; P1_R1192_U150
g11665 and P1_R1192_U370 P1_R1192_U369 ; P1_R1192_U151
g11666 nand P1_R1192_U116 P1_R1192_U196 ; P1_R1192_U152
g11667 and P1_R1192_U379 P1_R1192_U378 ; P1_R1192_U153
g11668 not P1_U4018 ; P1_R1192_U154
g11669 not P1_U3053 ; P1_R1192_U155
g11670 and P1_R1192_U388 P1_R1192_U387 ; P1_R1192_U156
g11671 nand P1_R1192_U128 P1_R1192_U302 ; P1_R1192_U157
g11672 and P1_R1192_U400 P1_R1192_U399 ; P1_R1192_U158
g11673 nand P1_R1192_U295 P1_R1192_U294 ; P1_R1192_U159
g11674 nand P1_R1192_U291 P1_R1192_U290 ; P1_R1192_U160
g11675 and P1_R1192_U417 P1_R1192_U416 ; P1_R1192_U161
g11676 and P1_R1192_U421 P1_R1192_U420 ; P1_R1192_U162
g11677 nand P1_R1192_U281 P1_R1192_U280 ; P1_R1192_U163
g11678 nand P1_R1192_U277 P1_R1192_U276 ; P1_R1192_U164
g11679 not P1_U3456 ; P1_R1192_U165
g11680 nand P1_R1192_U273 P1_R1192_U272 ; P1_R1192_U166
g11681 not P1_U3507 ; P1_R1192_U167
g11682 nand P1_R1192_U265 P1_R1192_U264 ; P1_R1192_U168
g11683 and P1_R1192_U453 P1_R1192_U452 ; P1_R1192_U169
g11684 and P1_R1192_U457 P1_R1192_U456 ; P1_R1192_U170
g11685 nand P1_R1192_U255 P1_R1192_U254 ; P1_R1192_U171
g11686 nand P1_R1192_U251 P1_R1192_U250 ; P1_R1192_U172
g11687 nand P1_R1192_U247 P1_R1192_U246 ; P1_R1192_U173
g11688 and P1_R1192_U474 P1_R1192_U473 ; P1_R1192_U174
g11689 nand P1_R1192_U129 P1_R1192_U157 ; P1_R1192_U175
g11690 not P1_R1192_U85 ; P1_R1192_U176
g11691 not P1_R1192_U29 ; P1_R1192_U177
g11692 not P1_R1192_U40 ; P1_R1192_U178
g11693 nand P1_U3483 P1_R1192_U53 ; P1_R1192_U179
g11694 nand P1_U3498 P1_R1192_U62 ; P1_R1192_U180
g11695 nand P1_U4013 P1_R1192_U76 ; P1_R1192_U181
g11696 nand P1_U4009 P1_R1192_U84 ; P1_R1192_U182
g11697 nand P1_U3459 P1_R1192_U28 ; P1_R1192_U183
g11698 nand P1_U3468 P1_R1192_U35 ; P1_R1192_U184
g11699 nand P1_U3474 P1_R1192_U39 ; P1_R1192_U185
g11700 not P1_R1192_U64 ; P1_R1192_U186
g11701 not P1_R1192_U78 ; P1_R1192_U187
g11702 not P1_R1192_U37 ; P1_R1192_U188
g11703 not P1_R1192_U54 ; P1_R1192_U189
g11704 not P1_R1192_U25 ; P1_R1192_U190
g11705 nand P1_R1192_U190 P1_R1192_U26 ; P1_R1192_U191
g11706 nand P1_R1192_U191 P1_R1192_U165 ; P1_R1192_U192
g11707 nand P1_U3076 P1_R1192_U25 ; P1_R1192_U193
g11708 not P1_R1192_U46 ; P1_R1192_U194
g11709 nand P1_U3462 P1_R1192_U30 ; P1_R1192_U195
g11710 nand P1_R1192_U115 P1_R1192_U46 ; P1_R1192_U196
g11711 nand P1_R1192_U30 P1_R1192_U29 ; P1_R1192_U197
g11712 nand P1_R1192_U197 P1_R1192_U27 ; P1_R1192_U198
g11713 nand P1_U3062 P1_R1192_U177 ; P1_R1192_U199
g11714 not P1_R1192_U152 ; P1_R1192_U200
g11715 nand P1_U3471 P1_R1192_U34 ; P1_R1192_U201
g11716 nand P1_U3069 P1_R1192_U31 ; P1_R1192_U202
g11717 nand P1_U3065 P1_R1192_U32 ; P1_R1192_U203
g11718 nand P1_R1192_U188 P1_R1192_U6 ; P1_R1192_U204
g11719 nand P1_R1192_U7 P1_R1192_U204 ; P1_R1192_U205
g11720 nand P1_U3465 P1_R1192_U36 ; P1_R1192_U206
g11721 nand P1_U3471 P1_R1192_U34 ; P1_R1192_U207
g11722 nand P1_R1192_U206 P1_R1192_U152 P1_R1192_U6 ; P1_R1192_U208
g11723 nand P1_R1192_U207 P1_R1192_U205 ; P1_R1192_U209
g11724 not P1_R1192_U44 ; P1_R1192_U210
g11725 nand P1_U3477 P1_R1192_U41 ; P1_R1192_U211
g11726 nand P1_R1192_U117 P1_R1192_U44 ; P1_R1192_U212
g11727 nand P1_R1192_U41 P1_R1192_U40 ; P1_R1192_U213
g11728 nand P1_R1192_U213 P1_R1192_U38 ; P1_R1192_U214
g11729 nand P1_U3082 P1_R1192_U178 ; P1_R1192_U215
g11730 not P1_R1192_U148 ; P1_R1192_U216
g11731 nand P1_U3480 P1_R1192_U43 ; P1_R1192_U217
g11732 nand P1_R1192_U217 P1_R1192_U54 ; P1_R1192_U218
g11733 nand P1_R1192_U210 P1_R1192_U40 ; P1_R1192_U219
g11734 nand P1_R1192_U120 P1_R1192_U219 ; P1_R1192_U220
g11735 nand P1_R1192_U44 P1_R1192_U185 ; P1_R1192_U221
g11736 nand P1_R1192_U119 P1_R1192_U221 ; P1_R1192_U222
g11737 nand P1_R1192_U40 P1_R1192_U185 ; P1_R1192_U223
g11738 nand P1_R1192_U206 P1_R1192_U152 ; P1_R1192_U224
g11739 not P1_R1192_U45 ; P1_R1192_U225
g11740 nand P1_U3065 P1_R1192_U32 ; P1_R1192_U226
g11741 nand P1_R1192_U225 P1_R1192_U226 ; P1_R1192_U227
g11742 nand P1_R1192_U122 P1_R1192_U227 ; P1_R1192_U228
g11743 nand P1_R1192_U45 P1_R1192_U184 ; P1_R1192_U229
g11744 nand P1_U3471 P1_R1192_U34 ; P1_R1192_U230
g11745 nand P1_R1192_U121 P1_R1192_U229 ; P1_R1192_U231
g11746 nand P1_U3065 P1_R1192_U32 ; P1_R1192_U232
g11747 nand P1_R1192_U184 P1_R1192_U232 ; P1_R1192_U233
g11748 nand P1_R1192_U206 P1_R1192_U37 ; P1_R1192_U234
g11749 nand P1_R1192_U194 P1_R1192_U29 ; P1_R1192_U235
g11750 nand P1_R1192_U124 P1_R1192_U235 ; P1_R1192_U236
g11751 nand P1_R1192_U46 P1_R1192_U183 ; P1_R1192_U237
g11752 nand P1_R1192_U123 P1_R1192_U237 ; P1_R1192_U238
g11753 nand P1_R1192_U29 P1_R1192_U183 ; P1_R1192_U239
g11754 nand P1_U3486 P1_R1192_U52 ; P1_R1192_U240
g11755 nand P1_U3061 P1_R1192_U50 ; P1_R1192_U241
g11756 nand P1_U3060 P1_R1192_U51 ; P1_R1192_U242
g11757 nand P1_R1192_U189 P1_R1192_U8 ; P1_R1192_U243
g11758 nand P1_R1192_U9 P1_R1192_U243 ; P1_R1192_U244
g11759 nand P1_U3486 P1_R1192_U52 ; P1_R1192_U245
g11760 nand P1_R1192_U125 P1_R1192_U148 ; P1_R1192_U246
g11761 nand P1_R1192_U245 P1_R1192_U244 ; P1_R1192_U247
g11762 not P1_R1192_U173 ; P1_R1192_U248
g11763 nand P1_U3489 P1_R1192_U56 ; P1_R1192_U249
g11764 nand P1_R1192_U249 P1_R1192_U173 ; P1_R1192_U250
g11765 nand P1_U3070 P1_R1192_U55 ; P1_R1192_U251
g11766 not P1_R1192_U172 ; P1_R1192_U252
g11767 nand P1_U3492 P1_R1192_U58 ; P1_R1192_U253
g11768 nand P1_R1192_U253 P1_R1192_U172 ; P1_R1192_U254
g11769 nand P1_U3078 P1_R1192_U57 ; P1_R1192_U255
g11770 not P1_R1192_U171 ; P1_R1192_U256
g11771 nand P1_U3501 P1_R1192_U61 ; P1_R1192_U257
g11772 nand P1_U3071 P1_R1192_U59 ; P1_R1192_U258
g11773 nand P1_U3072 P1_R1192_U49 ; P1_R1192_U259
g11774 nand P1_R1192_U186 P1_R1192_U180 ; P1_R1192_U260
g11775 nand P1_R1192_U10 P1_R1192_U260 ; P1_R1192_U261
g11776 nand P1_U3495 P1_R1192_U63 ; P1_R1192_U262
g11777 nand P1_U3501 P1_R1192_U61 ; P1_R1192_U263
g11778 nand P1_R1192_U171 P1_R1192_U126 P1_R1192_U257 ; P1_R1192_U264
g11779 nand P1_R1192_U263 P1_R1192_U261 ; P1_R1192_U265
g11780 not P1_R1192_U168 ; P1_R1192_U266
g11781 nand P1_U3504 P1_R1192_U66 ; P1_R1192_U267
g11782 nand P1_R1192_U267 P1_R1192_U168 ; P1_R1192_U268
g11783 nand P1_U3067 P1_R1192_U65 ; P1_R1192_U269
g11784 not P1_R1192_U67 ; P1_R1192_U270
g11785 nand P1_R1192_U270 P1_R1192_U68 ; P1_R1192_U271
g11786 nand P1_R1192_U271 P1_R1192_U167 ; P1_R1192_U272
g11787 nand P1_U3080 P1_R1192_U67 ; P1_R1192_U273
g11788 not P1_R1192_U166 ; P1_R1192_U274
g11789 nand P1_U3509 P1_R1192_U70 ; P1_R1192_U275
g11790 nand P1_R1192_U275 P1_R1192_U166 ; P1_R1192_U276
g11791 nand P1_U3079 P1_R1192_U69 ; P1_R1192_U277
g11792 not P1_R1192_U164 ; P1_R1192_U278
g11793 nand P1_U4015 P1_R1192_U72 ; P1_R1192_U279
g11794 nand P1_R1192_U279 P1_R1192_U164 ; P1_R1192_U280
g11795 nand P1_U3074 P1_R1192_U71 ; P1_R1192_U281
g11796 not P1_R1192_U163 ; P1_R1192_U282
g11797 nand P1_U4012 P1_R1192_U75 ; P1_R1192_U283
g11798 nand P1_U3064 P1_R1192_U73 ; P1_R1192_U284
g11799 nand P1_U3059 P1_R1192_U48 ; P1_R1192_U285
g11800 nand P1_R1192_U187 P1_R1192_U181 ; P1_R1192_U286
g11801 nand P1_R1192_U11 P1_R1192_U286 ; P1_R1192_U287
g11802 nand P1_U4014 P1_R1192_U77 ; P1_R1192_U288
g11803 nand P1_U4012 P1_R1192_U75 ; P1_R1192_U289
g11804 nand P1_R1192_U163 P1_R1192_U127 P1_R1192_U283 ; P1_R1192_U290
g11805 nand P1_R1192_U289 P1_R1192_U287 ; P1_R1192_U291
g11806 not P1_R1192_U160 ; P1_R1192_U292
g11807 nand P1_U4011 P1_R1192_U80 ; P1_R1192_U293
g11808 nand P1_R1192_U293 P1_R1192_U160 ; P1_R1192_U294
g11809 nand P1_U3063 P1_R1192_U79 ; P1_R1192_U295
g11810 not P1_R1192_U159 ; P1_R1192_U296
g11811 nand P1_U4010 P1_R1192_U82 ; P1_R1192_U297
g11812 nand P1_R1192_U297 P1_R1192_U159 ; P1_R1192_U298
g11813 nand P1_U3056 P1_R1192_U81 ; P1_R1192_U299
g11814 not P1_R1192_U89 ; P1_R1192_U300
g11815 nand P1_U4008 P1_R1192_U86 ; P1_R1192_U301
g11816 nand P1_R1192_U89 P1_R1192_U182 P1_R1192_U301 ; P1_R1192_U302
g11817 nand P1_R1192_U86 P1_R1192_U85 ; P1_R1192_U303
g11818 nand P1_R1192_U303 P1_R1192_U83 ; P1_R1192_U304
g11819 nand P1_U3051 P1_R1192_U176 ; P1_R1192_U305
g11820 not P1_R1192_U157 ; P1_R1192_U306
g11821 nand P1_U4007 P1_R1192_U88 ; P1_R1192_U307
g11822 nand P1_U3052 P1_R1192_U87 ; P1_R1192_U308
g11823 nand P1_R1192_U300 P1_R1192_U85 ; P1_R1192_U309
g11824 nand P1_R1192_U133 P1_R1192_U309 ; P1_R1192_U310
g11825 nand P1_R1192_U89 P1_R1192_U182 ; P1_R1192_U311
g11826 nand P1_R1192_U132 P1_R1192_U311 ; P1_R1192_U312
g11827 nand P1_R1192_U85 P1_R1192_U182 ; P1_R1192_U313
g11828 nand P1_R1192_U288 P1_R1192_U163 ; P1_R1192_U314
g11829 not P1_R1192_U90 ; P1_R1192_U315
g11830 nand P1_U3059 P1_R1192_U48 ; P1_R1192_U316
g11831 nand P1_R1192_U315 P1_R1192_U316 ; P1_R1192_U317
g11832 nand P1_R1192_U136 P1_R1192_U317 ; P1_R1192_U318
g11833 nand P1_R1192_U90 P1_R1192_U181 ; P1_R1192_U319
g11834 nand P1_U4012 P1_R1192_U75 ; P1_R1192_U320
g11835 nand P1_R1192_U320 P1_R1192_U319 P1_R1192_U11 ; P1_R1192_U321
g11836 nand P1_U3059 P1_R1192_U48 ; P1_R1192_U322
g11837 nand P1_R1192_U181 P1_R1192_U322 ; P1_R1192_U323
g11838 nand P1_R1192_U288 P1_R1192_U78 ; P1_R1192_U324
g11839 nand P1_R1192_U262 P1_R1192_U171 ; P1_R1192_U325
g11840 not P1_R1192_U91 ; P1_R1192_U326
g11841 nand P1_U3072 P1_R1192_U49 ; P1_R1192_U327
g11842 nand P1_R1192_U326 P1_R1192_U327 ; P1_R1192_U328
g11843 nand P1_R1192_U142 P1_R1192_U328 ; P1_R1192_U329
g11844 nand P1_R1192_U91 P1_R1192_U180 ; P1_R1192_U330
g11845 nand P1_U3501 P1_R1192_U61 ; P1_R1192_U331
g11846 nand P1_R1192_U331 P1_R1192_U330 P1_R1192_U10 ; P1_R1192_U332
g11847 nand P1_U3072 P1_R1192_U49 ; P1_R1192_U333
g11848 nand P1_R1192_U180 P1_R1192_U333 ; P1_R1192_U334
g11849 nand P1_R1192_U262 P1_R1192_U64 ; P1_R1192_U335
g11850 nand P1_R1192_U217 P1_R1192_U148 ; P1_R1192_U336
g11851 not P1_R1192_U92 ; P1_R1192_U337
g11852 nand P1_U3060 P1_R1192_U51 ; P1_R1192_U338
g11853 nand P1_R1192_U337 P1_R1192_U338 ; P1_R1192_U339
g11854 nand P1_R1192_U146 P1_R1192_U339 ; P1_R1192_U340
g11855 nand P1_R1192_U92 P1_R1192_U179 ; P1_R1192_U341
g11856 nand P1_U3486 P1_R1192_U52 ; P1_R1192_U342
g11857 nand P1_R1192_U145 P1_R1192_U341 ; P1_R1192_U343
g11858 nand P1_U3060 P1_R1192_U51 ; P1_R1192_U344
g11859 nand P1_R1192_U179 P1_R1192_U344 ; P1_R1192_U345
g11860 nand P1_U3075 P1_R1192_U24 ; P1_R1192_U346
g11861 nand P1_R1192_U89 P1_R1192_U182 P1_R1192_U301 ; P1_R1192_U347
g11862 nand P1_R1192_U12 P1_R1192_U347 P1_R1192_U130 ; P1_R1192_U348
g11863 nand P1_U3480 P1_R1192_U43 ; P1_R1192_U349
g11864 nand P1_U3081 P1_R1192_U42 ; P1_R1192_U350
g11865 nand P1_R1192_U218 P1_R1192_U148 ; P1_R1192_U351
g11866 nand P1_R1192_U216 P1_R1192_U147 ; P1_R1192_U352
g11867 nand P1_U3477 P1_R1192_U41 ; P1_R1192_U353
g11868 nand P1_U3082 P1_R1192_U38 ; P1_R1192_U354
g11869 nand P1_U3477 P1_R1192_U41 ; P1_R1192_U355
g11870 nand P1_U3082 P1_R1192_U38 ; P1_R1192_U356
g11871 nand P1_R1192_U356 P1_R1192_U355 ; P1_R1192_U357
g11872 nand P1_U3474 P1_R1192_U39 ; P1_R1192_U358
g11873 nand P1_U3068 P1_R1192_U22 ; P1_R1192_U359
g11874 nand P1_R1192_U223 P1_R1192_U44 ; P1_R1192_U360
g11875 nand P1_R1192_U149 P1_R1192_U210 ; P1_R1192_U361
g11876 nand P1_U3471 P1_R1192_U34 ; P1_R1192_U362
g11877 nand P1_U3069 P1_R1192_U31 ; P1_R1192_U363
g11878 nand P1_R1192_U363 P1_R1192_U362 ; P1_R1192_U364
g11879 nand P1_U3468 P1_R1192_U35 ; P1_R1192_U365
g11880 nand P1_U3065 P1_R1192_U32 ; P1_R1192_U366
g11881 nand P1_R1192_U233 P1_R1192_U45 ; P1_R1192_U367
g11882 nand P1_R1192_U150 P1_R1192_U225 ; P1_R1192_U368
g11883 nand P1_U3465 P1_R1192_U36 ; P1_R1192_U369
g11884 nand P1_U3058 P1_R1192_U33 ; P1_R1192_U370
g11885 nand P1_R1192_U234 P1_R1192_U152 ; P1_R1192_U371
g11886 nand P1_R1192_U200 P1_R1192_U151 ; P1_R1192_U372
g11887 nand P1_U3462 P1_R1192_U30 ; P1_R1192_U373
g11888 nand P1_U3062 P1_R1192_U27 ; P1_R1192_U374
g11889 nand P1_U3462 P1_R1192_U30 ; P1_R1192_U375
g11890 nand P1_U3062 P1_R1192_U27 ; P1_R1192_U376
g11891 nand P1_R1192_U376 P1_R1192_U375 ; P1_R1192_U377
g11892 nand P1_U3459 P1_R1192_U28 ; P1_R1192_U378
g11893 nand P1_U3066 P1_R1192_U23 ; P1_R1192_U379
g11894 nand P1_R1192_U239 P1_R1192_U46 ; P1_R1192_U380
g11895 nand P1_R1192_U153 P1_R1192_U194 ; P1_R1192_U381
g11896 nand P1_U4018 P1_R1192_U155 ; P1_R1192_U382
g11897 nand P1_U3053 P1_R1192_U154 ; P1_R1192_U383
g11898 nand P1_U4018 P1_R1192_U155 ; P1_R1192_U384
g11899 nand P1_U3053 P1_R1192_U154 ; P1_R1192_U385
g11900 nand P1_R1192_U385 P1_R1192_U384 ; P1_R1192_U386
g11901 nand P1_U3052 P1_R1192_U386 P1_R1192_U87 ; P1_R1192_U387
g11902 nand P1_R1192_U12 P1_R1192_U88 P1_U4007 ; P1_R1192_U388
g11903 nand P1_U4007 P1_R1192_U88 ; P1_R1192_U389
g11904 nand P1_U3052 P1_R1192_U87 ; P1_R1192_U390
g11905 not P1_R1192_U131 ; P1_R1192_U391
g11906 nand P1_R1192_U306 P1_R1192_U391 ; P1_R1192_U392
g11907 nand P1_R1192_U131 P1_R1192_U157 ; P1_R1192_U393
g11908 nand P1_U4008 P1_R1192_U86 ; P1_R1192_U394
g11909 nand P1_U3051 P1_R1192_U83 ; P1_R1192_U395
g11910 nand P1_U4008 P1_R1192_U86 ; P1_R1192_U396
g11911 nand P1_U3051 P1_R1192_U83 ; P1_R1192_U397
g11912 nand P1_R1192_U397 P1_R1192_U396 ; P1_R1192_U398
g11913 nand P1_U4009 P1_R1192_U84 ; P1_R1192_U399
g11914 nand P1_U3055 P1_R1192_U47 ; P1_R1192_U400
g11915 nand P1_R1192_U313 P1_R1192_U89 ; P1_R1192_U401
g11916 nand P1_R1192_U158 P1_R1192_U300 ; P1_R1192_U402
g11917 nand P1_U4010 P1_R1192_U82 ; P1_R1192_U403
g11918 nand P1_U3056 P1_R1192_U81 ; P1_R1192_U404
g11919 not P1_R1192_U134 ; P1_R1192_U405
g11920 nand P1_R1192_U296 P1_R1192_U405 ; P1_R1192_U406
g11921 nand P1_R1192_U134 P1_R1192_U159 ; P1_R1192_U407
g11922 nand P1_U4011 P1_R1192_U80 ; P1_R1192_U408
g11923 nand P1_U3063 P1_R1192_U79 ; P1_R1192_U409
g11924 not P1_R1192_U135 ; P1_R1192_U410
g11925 nand P1_R1192_U292 P1_R1192_U410 ; P1_R1192_U411
g11926 nand P1_R1192_U135 P1_R1192_U160 ; P1_R1192_U412
g11927 nand P1_U4012 P1_R1192_U75 ; P1_R1192_U413
g11928 nand P1_U3064 P1_R1192_U73 ; P1_R1192_U414
g11929 nand P1_R1192_U414 P1_R1192_U413 ; P1_R1192_U415
g11930 nand P1_U4013 P1_R1192_U76 ; P1_R1192_U416
g11931 nand P1_U3059 P1_R1192_U48 ; P1_R1192_U417
g11932 nand P1_R1192_U323 P1_R1192_U90 ; P1_R1192_U418
g11933 nand P1_R1192_U161 P1_R1192_U315 ; P1_R1192_U419
g11934 nand P1_U4014 P1_R1192_U77 ; P1_R1192_U420
g11935 nand P1_U3073 P1_R1192_U74 ; P1_R1192_U421
g11936 nand P1_R1192_U324 P1_R1192_U163 ; P1_R1192_U422
g11937 nand P1_R1192_U282 P1_R1192_U162 ; P1_R1192_U423
g11938 nand P1_U4015 P1_R1192_U72 ; P1_R1192_U424
g11939 nand P1_U3074 P1_R1192_U71 ; P1_R1192_U425
g11940 not P1_R1192_U137 ; P1_R1192_U426
g11941 nand P1_R1192_U278 P1_R1192_U426 ; P1_R1192_U427
g11942 nand P1_R1192_U137 P1_R1192_U164 ; P1_R1192_U428
g11943 nand P1_U3456 P1_R1192_U26 ; P1_R1192_U429
g11944 nand P1_U3076 P1_R1192_U165 ; P1_R1192_U430
g11945 not P1_R1192_U138 ; P1_R1192_U431
g11946 nand P1_R1192_U431 P1_R1192_U190 ; P1_R1192_U432
g11947 nand P1_R1192_U138 P1_R1192_U25 ; P1_R1192_U433
g11948 nand P1_U3509 P1_R1192_U70 ; P1_R1192_U434
g11949 nand P1_U3079 P1_R1192_U69 ; P1_R1192_U435
g11950 not P1_R1192_U139 ; P1_R1192_U436
g11951 nand P1_R1192_U274 P1_R1192_U436 ; P1_R1192_U437
g11952 nand P1_R1192_U139 P1_R1192_U166 ; P1_R1192_U438
g11953 nand P1_U3507 P1_R1192_U68 ; P1_R1192_U439
g11954 nand P1_U3080 P1_R1192_U167 ; P1_R1192_U440
g11955 not P1_R1192_U140 ; P1_R1192_U441
g11956 nand P1_R1192_U441 P1_R1192_U270 ; P1_R1192_U442
g11957 nand P1_R1192_U140 P1_R1192_U67 ; P1_R1192_U443
g11958 nand P1_U3504 P1_R1192_U66 ; P1_R1192_U444
g11959 nand P1_U3067 P1_R1192_U65 ; P1_R1192_U445
g11960 not P1_R1192_U141 ; P1_R1192_U446
g11961 nand P1_R1192_U266 P1_R1192_U446 ; P1_R1192_U447
g11962 nand P1_R1192_U141 P1_R1192_U168 ; P1_R1192_U448
g11963 nand P1_U3501 P1_R1192_U61 ; P1_R1192_U449
g11964 nand P1_U3071 P1_R1192_U59 ; P1_R1192_U450
g11965 nand P1_R1192_U450 P1_R1192_U449 ; P1_R1192_U451
g11966 nand P1_U3498 P1_R1192_U62 ; P1_R1192_U452
g11967 nand P1_U3072 P1_R1192_U49 ; P1_R1192_U453
g11968 nand P1_R1192_U334 P1_R1192_U91 ; P1_R1192_U454
g11969 nand P1_R1192_U169 P1_R1192_U326 ; P1_R1192_U455
g11970 nand P1_U3495 P1_R1192_U63 ; P1_R1192_U456
g11971 nand P1_U3077 P1_R1192_U60 ; P1_R1192_U457
g11972 nand P1_R1192_U335 P1_R1192_U171 ; P1_R1192_U458
g11973 nand P1_R1192_U256 P1_R1192_U170 ; P1_R1192_U459
g11974 nand P1_U3492 P1_R1192_U58 ; P1_R1192_U460
g11975 nand P1_U3078 P1_R1192_U57 ; P1_R1192_U461
g11976 not P1_R1192_U143 ; P1_R1192_U462
g11977 nand P1_R1192_U252 P1_R1192_U462 ; P1_R1192_U463
g11978 nand P1_R1192_U143 P1_R1192_U172 ; P1_R1192_U464
g11979 nand P1_U3489 P1_R1192_U56 ; P1_R1192_U465
g11980 nand P1_U3070 P1_R1192_U55 ; P1_R1192_U466
g11981 not P1_R1192_U144 ; P1_R1192_U467
g11982 nand P1_R1192_U248 P1_R1192_U467 ; P1_R1192_U468
g11983 nand P1_R1192_U144 P1_R1192_U173 ; P1_R1192_U469
g11984 nand P1_U3486 P1_R1192_U52 ; P1_R1192_U470
g11985 nand P1_U3061 P1_R1192_U50 ; P1_R1192_U471
g11986 nand P1_R1192_U471 P1_R1192_U470 ; P1_R1192_U472
g11987 nand P1_U3483 P1_R1192_U53 ; P1_R1192_U473
g11988 nand P1_U3060 P1_R1192_U51 ; P1_R1192_U474
g11989 nand P1_R1192_U345 P1_R1192_U92 ; P1_R1192_U475
g11990 nand P1_R1192_U174 P1_R1192_U337 ; P1_R1192_U476
g11991 and P1_LT_201_U109 P1_LT_201_U108 ; P1_LT_201_U6
g11992 and P1_LT_201_U111 P1_LT_201_U112 ; P1_LT_201_U7
g11993 and P1_LT_201_U113 P1_LT_201_U114 ; P1_LT_201_U8
g11994 and P1_LT_201_U81 P1_LT_201_U116 P1_LT_201_U118 P1_LT_201_U8 ; P1_LT_201_U9
g11995 and P1_LT_201_U126 P1_LT_201_U125 ; P1_LT_201_U10
g11996 and P1_LT_201_U127 P1_LT_201_U124 P1_LT_201_U84 P1_LT_201_U85 ; P1_LT_201_U11
g11997 and P1_LT_201_U141 P1_LT_201_U140 ; P1_LT_201_U12
g11998 and P1_LT_201_U102 P1_LT_201_U193 ; P1_LT_201_U13
g11999 and P1_LT_201_U189 P1_LT_201_U104 ; P1_LT_201_U14
g12000 not P1_U3594 ; P1_LT_201_U15
g12001 not P1_U3595 ; P1_LT_201_U16
g12002 not P1_U4017 ; P1_LT_201_U17
g12003 not P1_U4018 ; P1_LT_201_U18
g12004 not P1_U3599 ; P1_LT_201_U19
g12005 not P1_U4011 ; P1_LT_201_U20
g12006 not P1_U4010 ; P1_LT_201_U21
g12007 not P1_U3604 ; P1_LT_201_U22
g12008 not P1_U4014 ; P1_LT_201_U23
g12009 not P1_U3605 ; P1_LT_201_U24
g12010 not P1_U4015 ; P1_LT_201_U25
g12011 not P1_U3509 ; P1_LT_201_U26
g12012 not P1_U3609 ; P1_LT_201_U27
g12013 not P1_U3507 ; P1_LT_201_U28
g12014 not P1_U3610 ; P1_LT_201_U29
g12015 not P1_U3608 ; P1_LT_201_U30
g12016 not P1_U3606 ; P1_LT_201_U31
g12017 not P1_U3504 ; P1_LT_201_U32
g12018 not P1_U3501 ; P1_LT_201_U33
g12019 not P1_U3611 ; P1_LT_201_U34
g12020 not P1_U3612 ; P1_LT_201_U35
g12021 not P1_U3474 ; P1_LT_201_U36
g12022 not P1_U3590 ; P1_LT_201_U37
g12023 not P1_U3471 ; P1_LT_201_U38
g12024 not P1_U3591 ; P1_LT_201_U39
g12025 not P1_U3587 ; P1_LT_201_U40
g12026 not P1_U3617 ; P1_LT_201_U41
g12027 not P1_U3588 ; P1_LT_201_U42
g12028 not P1_U3589 ; P1_LT_201_U43
g12029 not P1_U3592 ; P1_LT_201_U44
g12030 not P1_U3593 ; P1_LT_201_U45
g12031 nand P1_U3451 P1_LT_201_U105 ; P1_LT_201_U46
g12032 not P1_U3456 ; P1_LT_201_U47
g12033 not P1_U3596 ; P1_LT_201_U48
g12034 not P1_U3489 ; P1_LT_201_U49
g12035 not P1_U3492 ; P1_LT_201_U50
g12036 not P1_U3459 ; P1_LT_201_U51
g12037 not P1_U3462 ; P1_LT_201_U52
g12038 not P1_U3465 ; P1_LT_201_U53
g12039 not P1_U3468 ; P1_LT_201_U54
g12040 not P1_U3477 ; P1_LT_201_U55
g12041 not P1_U3480 ; P1_LT_201_U56
g12042 not P1_U3483 ; P1_LT_201_U57
g12043 not P1_U3486 ; P1_LT_201_U58
g12044 not P1_U3615 ; P1_LT_201_U59
g12045 not P1_U3616 ; P1_LT_201_U60
g12046 not P1_U3613 ; P1_LT_201_U61
g12047 not P1_U3614 ; P1_LT_201_U62
g12048 not P1_U3495 ; P1_LT_201_U63
g12049 not P1_U3498 ; P1_LT_201_U64
g12050 not P1_U4013 ; P1_LT_201_U65
g12051 not P1_U4012 ; P1_LT_201_U66
g12052 not P1_U3603 ; P1_LT_201_U67
g12053 not P1_U3600 ; P1_LT_201_U68
g12054 not P1_U3602 ; P1_LT_201_U69
g12055 not P1_U3601 ; P1_LT_201_U70
g12056 not P1_U4009 ; P1_LT_201_U71
g12057 not P1_U4008 ; P1_LT_201_U72
g12058 not P1_U4007 ; P1_LT_201_U73
g12059 not P1_U3597 ; P1_LT_201_U74
g12060 not P1_U4016 ; P1_LT_201_U75
g12061 and P1_U4014 P1_LT_201_U24 ; P1_LT_201_U76
g12062 and P1_U4015 P1_LT_201_U31 ; P1_LT_201_U77
g12063 and P1_LT_201_U171 P1_LT_201_U170 ; P1_LT_201_U78
g12064 and P1_U3609 P1_LT_201_U28 ; P1_LT_201_U79
g12065 and P1_U3610 P1_LT_201_U32 ; P1_LT_201_U80
g12066 and P1_LT_201_U117 P1_LT_201_U115 ; P1_LT_201_U81
g12067 and P1_U3590 P1_LT_201_U38 ; P1_LT_201_U82
g12068 and P1_U3591 P1_LT_201_U54 ; P1_LT_201_U83
g12069 and P1_LT_201_U129 P1_LT_201_U128 ; P1_LT_201_U84
g12070 and P1_LT_201_U133 P1_LT_201_U132 P1_LT_201_U131 P1_LT_201_U130 ; P1_LT_201_U85
g12071 and P1_LT_201_U137 P1_LT_201_U138 ; P1_LT_201_U86
g12072 and P1_LT_201_U86 P1_LT_201_U136 ; P1_LT_201_U87
g12073 and P1_U3459 P1_LT_201_U48 ; P1_LT_201_U88
g12074 and P1_U3462 P1_LT_201_U45 ; P1_LT_201_U89
g12075 and P1_LT_201_U131 P1_LT_201_U124 P1_LT_201_U130 ; P1_LT_201_U90
g12076 and P1_LT_201_U154 P1_LT_201_U139 ; P1_LT_201_U91
g12077 and P1_LT_201_U157 P1_LT_201_U156 ; P1_LT_201_U92
g12078 and P1_LT_201_U92 P1_LT_201_U12 ; P1_LT_201_U93
g12079 and P1_U3615 P1_LT_201_U49 ; P1_LT_201_U94
g12080 and P1_U3616 P1_LT_201_U58 ; P1_LT_201_U95
g12081 and P1_LT_201_U160 P1_LT_201_U161 ; P1_LT_201_U96
g12082 and P1_LT_201_U163 P1_LT_201_U162 ; P1_LT_201_U97
g12083 and P1_LT_201_U174 P1_LT_201_U173 P1_LT_201_U120 P1_LT_201_U121 ; P1_LT_201_U98
g12084 and P1_LT_201_U178 P1_LT_201_U177 ; P1_LT_201_U99
g12085 and P1_U3603 P1_LT_201_U66 ; P1_LT_201_U100
g12086 and P1_LT_201_U195 P1_LT_201_U184 ; P1_LT_201_U101
g12087 and P1_LT_201_U187 P1_LT_201_U73 ; P1_LT_201_U102
g12088 and P1_U3597 P1_LT_201_U18 ; P1_LT_201_U103
g12089 and P1_LT_201_U191 P1_LT_201_U107 P1_LT_201_U190 ; P1_LT_201_U104
g12090 not P1_U3618 ; P1_LT_201_U105
g12091 nand P1_U3594 P1_LT_201_U75 ; P1_LT_201_U106
g12092 nand P1_LT_201_U106 P1_U3595 P1_LT_201_U17 ; P1_LT_201_U107
g12093 nand P1_U4017 P1_LT_201_U16 ; P1_LT_201_U108
g12094 nand P1_U3594 P1_LT_201_U75 ; P1_LT_201_U109
g12095 nand P1_U3599 P1_LT_201_U72 ; P1_LT_201_U110
g12096 nand P1_U3509 P1_LT_201_U30 ; P1_LT_201_U111
g12097 nand P1_U3507 P1_LT_201_U27 ; P1_LT_201_U112
g12098 nand P1_U3604 P1_LT_201_U65 ; P1_LT_201_U113
g12099 nand P1_U3605 P1_LT_201_U23 ; P1_LT_201_U114
g12100 nand P1_LT_201_U79 P1_LT_201_U111 ; P1_LT_201_U115
g12101 nand P1_LT_201_U80 P1_LT_201_U7 ; P1_LT_201_U116
g12102 nand P1_U3608 P1_LT_201_U26 ; P1_LT_201_U117
g12103 nand P1_U3606 P1_LT_201_U25 ; P1_LT_201_U118
g12104 nand P1_U3611 P1_LT_201_U33 ; P1_LT_201_U119
g12105 nand P1_U4011 P1_LT_201_U69 ; P1_LT_201_U120
g12106 nand P1_U4010 P1_LT_201_U70 ; P1_LT_201_U121
g12107 nand P1_U3612 P1_LT_201_U64 ; P1_LT_201_U122
g12108 nand P1_U3474 P1_LT_201_U43 ; P1_LT_201_U123
g12109 nand P1_LT_201_U82 P1_LT_201_U123 ; P1_LT_201_U124
g12110 nand P1_U3471 P1_LT_201_U37 ; P1_LT_201_U125
g12111 nand P1_U3474 P1_LT_201_U43 ; P1_LT_201_U126
g12112 nand P1_LT_201_U83 P1_LT_201_U10 ; P1_LT_201_U127
g12113 nand P1_U3587 P1_LT_201_U56 ; P1_LT_201_U128
g12114 nand P1_U3617 P1_LT_201_U57 ; P1_LT_201_U129
g12115 nand P1_U3588 P1_LT_201_U55 ; P1_LT_201_U130
g12116 nand P1_U3589 P1_LT_201_U36 ; P1_LT_201_U131
g12117 nand P1_U3592 P1_LT_201_U53 ; P1_LT_201_U132
g12118 nand P1_U3593 P1_LT_201_U52 ; P1_LT_201_U133
g12119 not P1_LT_201_U46 ; P1_LT_201_U134
g12120 nand P1_U3456 P1_LT_201_U134 ; P1_LT_201_U135
g12121 nand P1_U3607 P1_LT_201_U135 ; P1_LT_201_U136
g12122 nand P1_LT_201_U46 P1_LT_201_U47 ; P1_LT_201_U137
g12123 nand P1_U3596 P1_LT_201_U51 ; P1_LT_201_U138
g12124 nand P1_LT_201_U87 P1_LT_201_U11 ; P1_LT_201_U139
g12125 nand P1_U3489 P1_LT_201_U59 ; P1_LT_201_U140
g12126 nand P1_U3492 P1_LT_201_U62 ; P1_LT_201_U141
g12127 nand P1_LT_201_U89 P1_LT_201_U132 ; P1_LT_201_U142
g12128 nand P1_U3465 P1_LT_201_U44 ; P1_LT_201_U143
g12129 nand P1_LT_201_U143 P1_LT_201_U142 P1_LT_201_U10 ; P1_LT_201_U144
g12130 nand P1_LT_201_U144 P1_LT_201_U127 ; P1_LT_201_U145
g12131 nand P1_U3468 P1_LT_201_U39 ; P1_LT_201_U146
g12132 nand P1_LT_201_U146 P1_LT_201_U145 ; P1_LT_201_U147
g12133 nand P1_LT_201_U90 P1_LT_201_U147 ; P1_LT_201_U148
g12134 nand P1_U3477 P1_LT_201_U42 ; P1_LT_201_U149
g12135 nand P1_LT_201_U149 P1_LT_201_U148 ; P1_LT_201_U150
g12136 nand P1_LT_201_U150 P1_LT_201_U128 ; P1_LT_201_U151
g12137 nand P1_U3480 P1_LT_201_U40 ; P1_LT_201_U152
g12138 nand P1_LT_201_U152 P1_LT_201_U151 ; P1_LT_201_U153
g12139 nand P1_LT_201_U88 P1_LT_201_U11 ; P1_LT_201_U154
g12140 nand P1_LT_201_U153 P1_LT_201_U129 ; P1_LT_201_U155
g12141 nand P1_U3483 P1_LT_201_U41 ; P1_LT_201_U156
g12142 nand P1_U3486 P1_LT_201_U60 ; P1_LT_201_U157
g12143 nand P1_LT_201_U91 P1_LT_201_U155 P1_LT_201_U93 ; P1_LT_201_U158
g12144 nand P1_U3492 P1_LT_201_U62 ; P1_LT_201_U159
g12145 nand P1_LT_201_U94 P1_LT_201_U159 ; P1_LT_201_U160
g12146 nand P1_LT_201_U95 P1_LT_201_U12 ; P1_LT_201_U161
g12147 nand P1_U3613 P1_LT_201_U63 ; P1_LT_201_U162
g12148 nand P1_U3614 P1_LT_201_U50 ; P1_LT_201_U163
g12149 nand P1_LT_201_U96 P1_LT_201_U158 P1_LT_201_U97 ; P1_LT_201_U164
g12150 nand P1_U3495 P1_LT_201_U61 ; P1_LT_201_U165
g12151 nand P1_LT_201_U165 P1_LT_201_U164 ; P1_LT_201_U166
g12152 nand P1_LT_201_U166 P1_LT_201_U122 ; P1_LT_201_U167
g12153 nand P1_U3498 P1_LT_201_U35 ; P1_LT_201_U168
g12154 nand P1_LT_201_U168 P1_LT_201_U167 ; P1_LT_201_U169
g12155 nand P1_U3504 P1_LT_201_U29 ; P1_LT_201_U170
g12156 nand P1_U3501 P1_LT_201_U34 ; P1_LT_201_U171
g12157 nand P1_LT_201_U78 P1_LT_201_U7 ; P1_LT_201_U172
g12158 nand P1_LT_201_U76 P1_LT_201_U113 ; P1_LT_201_U173
g12159 nand P1_LT_201_U77 P1_LT_201_U8 ; P1_LT_201_U174
g12160 nand P1_LT_201_U9 P1_LT_201_U172 ; P1_LT_201_U175
g12161 nand P1_LT_201_U169 P1_LT_201_U119 P1_LT_201_U9 ; P1_LT_201_U176
g12162 nand P1_U4013 P1_LT_201_U22 ; P1_LT_201_U177
g12163 nand P1_U4012 P1_LT_201_U67 ; P1_LT_201_U178
g12164 nand P1_LT_201_U176 P1_LT_201_U175 P1_LT_201_U99 P1_LT_201_U98 ; P1_LT_201_U179
g12165 nand P1_LT_201_U120 P1_LT_201_U100 P1_LT_201_U121 ; P1_LT_201_U180
g12166 nand P1_U4010 P1_LT_201_U70 ; P1_LT_201_U181
g12167 nand P1_U3602 P1_LT_201_U20 ; P1_LT_201_U182
g12168 nand P1_U3601 P1_LT_201_U21 ; P1_LT_201_U183
g12169 nand P1_U3600 P1_LT_201_U71 ; P1_LT_201_U184
g12170 nand P1_LT_201_U180 P1_LT_201_U179 P1_LT_201_U101 ; P1_LT_201_U185
g12171 nand P1_U4009 P1_LT_201_U68 ; P1_LT_201_U186
g12172 nand P1_U4008 P1_LT_201_U19 ; P1_LT_201_U187
g12173 nand P1_U4018 P1_LT_201_U74 ; P1_LT_201_U188
g12174 nand P1_LT_201_U6 P1_LT_201_U198 P1_LT_201_U196 P1_LT_201_U188 ; P1_LT_201_U189
g12175 nand P1_LT_201_U103 P1_LT_201_U6 ; P1_LT_201_U190
g12176 nand P1_U4016 P1_LT_201_U15 ; P1_LT_201_U191
g12177 nand P1_LT_201_U186 P1_LT_201_U185 ; P1_LT_201_U192
g12178 nand P1_LT_201_U192 P1_LT_201_U110 ; P1_LT_201_U193
g12179 nand P1_LT_201_U183 P1_LT_201_U182 ; P1_LT_201_U194
g12180 nand P1_LT_201_U194 P1_LT_201_U181 ; P1_LT_201_U195
g12181 or P1_U3598 P1_LT_201_U13 ; P1_LT_201_U196
g12182 nand P1_LT_201_U187 P1_LT_201_U193 ; P1_LT_201_U197
g12183 nand P1_U4007 P1_LT_201_U197 ; P1_LT_201_U198
g12184 and P1_R1360_U111 P1_R1360_U112 ; P1_R1360_U6
g12185 and P1_R1360_U116 P1_R1360_U115 ; P1_R1360_U7
g12186 and P1_R1360_U118 P1_R1360_U119 ; P1_R1360_U8
g12187 and P1_R1360_U123 P1_R1360_U122 ; P1_R1360_U9
g12188 and P1_R1360_U199 P1_R1360_U185 P1_R1360_U186 P1_R1360_U184 P1_R1360_U183 ; P1_R1360_U10
g12189 and P1_R1360_U183 P1_R1360_U104 ; P1_R1360_U11
g12190 and P1_R1360_U203 P1_R1360_U202 ; P1_R1360_U12
g12191 and P1_R1360_U205 P1_R1360_U204 ; P1_R1360_U13
g12192 nand P1_R1360_U108 P1_R1360_U200 P1_R1360_U107 ; P1_R1360_U14
g12193 not P1_U3086 ; P1_R1360_U15
g12194 not P1_U3085 ; P1_R1360_U16
g12195 not P1_U3119 ; P1_R1360_U17
g12196 not P1_U3087 ; P1_R1360_U18
g12197 not P1_U3088 ; P1_R1360_U19
g12198 not P1_U3121 ; P1_R1360_U20
g12199 not P1_U3120 ; P1_R1360_U21
g12200 not P1_U3118 ; P1_R1360_U22
g12201 not P1_U3125 ; P1_R1360_U23
g12202 not P1_U3124 ; P1_R1360_U24
g12203 not P1_U3095 ; P1_R1360_U25
g12204 not P1_U3096 ; P1_R1360_U26
g12205 not P1_U3131 ; P1_R1360_U27
g12206 not P1_U3130 ; P1_R1360_U28
g12207 not P1_U3101 ; P1_R1360_U29
g12208 not P1_U3102 ; P1_R1360_U30
g12209 not P1_U3137 ; P1_R1360_U31
g12210 not P1_U3136 ; P1_R1360_U32
g12211 not P1_U3107 ; P1_R1360_U33
g12212 not P1_U3140 ; P1_R1360_U34
g12213 not P1_U3108 ; P1_R1360_U35
g12214 not P1_U3141 ; P1_R1360_U36
g12215 not P1_U3110 ; P1_R1360_U37
g12216 not P1_U3109 ; P1_R1360_U38
g12217 not P1_U3112 ; P1_R1360_U39
g12218 not P1_U3111 ; P1_R1360_U40
g12219 not P1_U3114 ; P1_R1360_U41
g12220 not P1_U3113 ; P1_R1360_U42
g12221 not P1_U3115 ; P1_R1360_U43
g12222 not P1_U3147 ; P1_R1360_U44
g12223 not P1_U3146 ; P1_R1360_U45
g12224 not P1_U3145 ; P1_R1360_U46
g12225 not P1_U3144 ; P1_R1360_U47
g12226 not P1_U3143 ; P1_R1360_U48
g12227 not P1_U3142 ; P1_R1360_U49
g12228 not P1_U3139 ; P1_R1360_U50
g12229 not P1_U3138 ; P1_R1360_U51
g12230 not P1_U3106 ; P1_R1360_U52
g12231 not P1_U3104 ; P1_R1360_U53
g12232 not P1_U3105 ; P1_R1360_U54
g12233 not P1_U3103 ; P1_R1360_U55
g12234 not P1_U3135 ; P1_R1360_U56
g12235 not P1_U3134 ; P1_R1360_U57
g12236 not P1_U3133 ; P1_R1360_U58
g12237 not P1_U3132 ; P1_R1360_U59
g12238 not P1_U3100 ; P1_R1360_U60
g12239 not P1_U3099 ; P1_R1360_U61
g12240 not P1_U3098 ; P1_R1360_U62
g12241 not P1_U3097 ; P1_R1360_U63
g12242 not P1_U3129 ; P1_R1360_U64
g12243 not P1_U3128 ; P1_R1360_U65
g12244 not P1_U3127 ; P1_R1360_U66
g12245 not P1_U3126 ; P1_R1360_U67
g12246 not P1_U3090 ; P1_R1360_U68
g12247 not P1_U3089 ; P1_R1360_U69
g12248 not P1_U3093 ; P1_R1360_U70
g12249 not P1_U3094 ; P1_R1360_U71
g12250 not P1_U3091 ; P1_R1360_U72
g12251 not P1_U3092 ; P1_R1360_U73
g12252 not P1_U3122 ; P1_R1360_U74
g12253 not P1_U3123 ; P1_R1360_U75
g12254 not P1_U3150 ; P1_R1360_U76
g12255 and P1_R1360_U18 P1_U3119 ; P1_R1360_U77
g12256 and P1_R1360_U183 P1_R1360_U184 ; P1_R1360_U78
g12257 and P1_U3140 P1_R1360_U35 ; P1_R1360_U79
g12258 and P1_U3141 P1_R1360_U38 ; P1_R1360_U80
g12259 and P1_R1360_U127 P1_R1360_U126 P1_R1360_U125 P1_R1360_U124 ; P1_R1360_U81
g12260 and P1_R1360_U130 P1_R1360_U131 P1_R1360_U129 ; P1_R1360_U82
g12261 and P1_U3147 P1_R1360_U43 ; P1_R1360_U83
g12262 and P1_R1360_U85 P1_R1360_U132 ; P1_R1360_U84
g12263 and P1_R1360_U144 P1_R1360_U143 ; P1_R1360_U85
g12264 and P1_R1360_U121 P1_R1360_U120 ; P1_R1360_U86
g12265 and P1_R1360_U8 P1_R1360_U86 ; P1_R1360_U87
g12266 and P1_R1360_U147 P1_R1360_U146 P1_R1360_U90 ; P1_R1360_U88
g12267 and P1_R1360_U150 P1_R1360_U149 ; P1_R1360_U89
g12268 and P1_R1360_U89 P1_R1360_U9 ; P1_R1360_U90
g12269 and P1_U3106 P1_R1360_U51 ; P1_R1360_U91
g12270 and P1_U3105 P1_R1360_U31 ; P1_R1360_U92
g12271 and P1_R1360_U152 P1_R1360_U153 P1_R1360_U94 ; P1_R1360_U93
g12272 and P1_R1360_U156 P1_R1360_U155 ; P1_R1360_U94
g12273 and P1_R1360_U7 P1_R1360_U96 ; P1_R1360_U95
g12274 and P1_R1360_U164 P1_R1360_U165 ; P1_R1360_U96
g12275 and P1_U3100 P1_R1360_U59 ; P1_R1360_U97
g12276 and P1_U3099 P1_R1360_U27 ; P1_R1360_U98
g12277 and P1_R1360_U167 P1_R1360_U169 P1_R1360_U100 ; P1_R1360_U99
g12278 and P1_R1360_U171 P1_R1360_U170 ; P1_R1360_U100
g12279 and P1_R1360_U179 P1_R1360_U180 ; P1_R1360_U101
g12280 and P1_U3093 P1_R1360_U23 ; P1_R1360_U102
g12281 and P1_U3094 P1_R1360_U67 ; P1_R1360_U103
g12282 and P1_R1360_U181 P1_R1360_U185 P1_R1360_U186 P1_R1360_U106 P1_R1360_U184 ; P1_R1360_U104
g12283 and P1_R1360_U190 P1_R1360_U189 ; P1_R1360_U105
g12284 and P1_R1360_U188 P1_R1360_U187 P1_R1360_U105 ; P1_R1360_U106
g12285 and P1_R1360_U196 P1_R1360_U194 P1_R1360_U195 ; P1_R1360_U107
g12286 and P1_R1360_U201 P1_R1360_U13 ; P1_R1360_U108
g12287 not P1_U3117 ; P1_R1360_U109
g12288 nand P1_U3095 P1_R1360_U66 ; P1_R1360_U110
g12289 nand P1_U3124 P1_R1360_U73 ; P1_R1360_U111
g12290 nand P1_U3125 P1_R1360_U70 ; P1_R1360_U112
g12291 nand P1_U3096 P1_R1360_U65 ; P1_R1360_U113
g12292 nand P1_U3101 P1_R1360_U58 ; P1_R1360_U114
g12293 nand P1_U3131 P1_R1360_U61 ; P1_R1360_U115
g12294 nand P1_U3130 P1_R1360_U62 ; P1_R1360_U116
g12295 nand P1_U3102 P1_R1360_U57 ; P1_R1360_U117
g12296 nand P1_U3107 P1_R1360_U50 ; P1_R1360_U118
g12297 nand P1_U3108 P1_R1360_U34 ; P1_R1360_U119
g12298 nand P1_U3110 P1_R1360_U49 ; P1_R1360_U120
g12299 nand P1_U3109 P1_R1360_U36 ; P1_R1360_U121
g12300 nand P1_U3137 P1_R1360_U54 ; P1_R1360_U122
g12301 nand P1_U3136 P1_R1360_U53 ; P1_R1360_U123
g12302 nand P1_U3112 P1_R1360_U47 ; P1_R1360_U124
g12303 nand P1_U3111 P1_R1360_U48 ; P1_R1360_U125
g12304 nand P1_U3114 P1_R1360_U45 ; P1_R1360_U126
g12305 nand P1_U3113 P1_R1360_U46 ; P1_R1360_U127
g12306 nand P1_U3148 P1_U3149 ; P1_R1360_U128
g12307 nand P1_U3116 P1_R1360_U128 ; P1_R1360_U129
g12308 or P1_U3148 P1_U3149 ; P1_R1360_U130
g12309 nand P1_U3115 P1_R1360_U44 ; P1_R1360_U131
g12310 nand P1_R1360_U82 P1_R1360_U81 ; P1_R1360_U132
g12311 nand P1_R1360_U83 P1_R1360_U126 ; P1_R1360_U133
g12312 nand P1_U3146 P1_R1360_U41 ; P1_R1360_U134
g12313 nand P1_R1360_U134 P1_R1360_U133 ; P1_R1360_U135
g12314 nand P1_R1360_U135 P1_R1360_U127 ; P1_R1360_U136
g12315 nand P1_U3145 P1_R1360_U42 ; P1_R1360_U137
g12316 nand P1_R1360_U137 P1_R1360_U136 ; P1_R1360_U138
g12317 nand P1_R1360_U138 P1_R1360_U124 ; P1_R1360_U139
g12318 nand P1_U3144 P1_R1360_U39 ; P1_R1360_U140
g12319 nand P1_R1360_U140 P1_R1360_U139 ; P1_R1360_U141
g12320 nand P1_R1360_U141 P1_R1360_U125 ; P1_R1360_U142
g12321 nand P1_U3143 P1_R1360_U40 ; P1_R1360_U143
g12322 nand P1_U3142 P1_R1360_U37 ; P1_R1360_U144
g12323 nand P1_R1360_U142 P1_R1360_U84 ; P1_R1360_U145
g12324 nand P1_R1360_U79 P1_R1360_U118 ; P1_R1360_U146
g12325 nand P1_R1360_U80 P1_R1360_U8 ; P1_R1360_U147
g12326 nand P1_R1360_U87 P1_R1360_U145 ; P1_R1360_U148
g12327 nand P1_U3139 P1_R1360_U33 ; P1_R1360_U149
g12328 nand P1_U3138 P1_R1360_U52 ; P1_R1360_U150
g12329 nand P1_R1360_U148 P1_R1360_U88 ; P1_R1360_U151
g12330 nand P1_R1360_U91 P1_R1360_U9 ; P1_R1360_U152
g12331 nand P1_U3104 P1_R1360_U32 ; P1_R1360_U153
g12332 nand P1_U3136 P1_R1360_U53 ; P1_R1360_U154
g12333 nand P1_R1360_U92 P1_R1360_U154 ; P1_R1360_U155
g12334 nand P1_U3103 P1_R1360_U56 ; P1_R1360_U156
g12335 nand P1_R1360_U151 P1_R1360_U93 ; P1_R1360_U157
g12336 nand P1_U3135 P1_R1360_U55 ; P1_R1360_U158
g12337 nand P1_R1360_U158 P1_R1360_U157 ; P1_R1360_U159
g12338 nand P1_R1360_U159 P1_R1360_U117 ; P1_R1360_U160
g12339 nand P1_U3134 P1_R1360_U30 ; P1_R1360_U161
g12340 nand P1_R1360_U161 P1_R1360_U160 ; P1_R1360_U162
g12341 nand P1_R1360_U162 P1_R1360_U114 ; P1_R1360_U163
g12342 nand P1_U3133 P1_R1360_U29 ; P1_R1360_U164
g12343 nand P1_U3132 P1_R1360_U60 ; P1_R1360_U165
g12344 nand P1_R1360_U163 P1_R1360_U95 ; P1_R1360_U166
g12345 nand P1_R1360_U97 P1_R1360_U7 ; P1_R1360_U167
g12346 nand P1_U3130 P1_R1360_U62 ; P1_R1360_U168
g12347 nand P1_R1360_U98 P1_R1360_U168 ; P1_R1360_U169
g12348 nand P1_U3098 P1_R1360_U28 ; P1_R1360_U170
g12349 nand P1_U3097 P1_R1360_U64 ; P1_R1360_U171
g12350 nand P1_R1360_U166 P1_R1360_U99 ; P1_R1360_U172
g12351 nand P1_U3129 P1_R1360_U63 ; P1_R1360_U173
g12352 nand P1_R1360_U173 P1_R1360_U172 ; P1_R1360_U174
g12353 nand P1_R1360_U174 P1_R1360_U113 ; P1_R1360_U175
g12354 nand P1_U3128 P1_R1360_U26 ; P1_R1360_U176
g12355 nand P1_R1360_U176 P1_R1360_U175 ; P1_R1360_U177
g12356 nand P1_R1360_U177 P1_R1360_U110 ; P1_R1360_U178
g12357 nand P1_U3127 P1_R1360_U25 ; P1_R1360_U179
g12358 nand P1_U3126 P1_R1360_U71 ; P1_R1360_U180
g12359 nand P1_R1360_U101 P1_R1360_U178 P1_R1360_U6 ; P1_R1360_U181
g12360 nand P1_U3086 P1_R1360_U22 ; P1_R1360_U182
g12361 nand P1_U3087 P1_R1360_U17 ; P1_R1360_U183
g12362 nand P1_U3088 P1_R1360_U21 ; P1_R1360_U184
g12363 nand P1_U3090 P1_R1360_U74 ; P1_R1360_U185
g12364 nand P1_U3089 P1_R1360_U20 ; P1_R1360_U186
g12365 nand P1_R1360_U102 P1_R1360_U111 ; P1_R1360_U187
g12366 nand P1_R1360_U103 P1_R1360_U6 ; P1_R1360_U188
g12367 nand P1_U3091 P1_R1360_U75 ; P1_R1360_U189
g12368 nand P1_U3092 P1_R1360_U24 ; P1_R1360_U190
g12369 nand P1_U3121 P1_R1360_U69 ; P1_R1360_U191
g12370 nand P1_U3120 P1_R1360_U19 ; P1_R1360_U192
g12371 nand P1_R1360_U192 P1_R1360_U191 ; P1_R1360_U193
g12372 nand P1_R1360_U77 P1_R1360_U12 P1_R1360_U182 ; P1_R1360_U194
g12373 nand P1_R1360_U12 P1_R1360_U193 P1_R1360_U78 P1_R1360_U182 ; P1_R1360_U195
g12374 nand P1_R1360_U12 P1_R1360_U15 P1_U3118 ; P1_R1360_U196
g12375 nand P1_U3122 P1_R1360_U68 ; P1_R1360_U197
g12376 nand P1_U3123 P1_R1360_U72 ; P1_R1360_U198
g12377 nand P1_R1360_U198 P1_R1360_U197 ; P1_R1360_U199
g12378 nand P1_R1360_U12 P1_R1360_U11 P1_R1360_U182 ; P1_R1360_U200
g12379 nand P1_R1360_U12 P1_R1360_U10 P1_R1360_U182 ; P1_R1360_U201
g12380 nand P1_U3085 P1_R1360_U109 ; P1_R1360_U202
g12381 nand P1_U3117 P1_R1360_U16 ; P1_R1360_U203
g12382 nand P1_U3150 P1_U3085 P1_R1360_U109 ; P1_R1360_U204
g12383 nand P1_R1360_U76 P1_R1360_U16 P1_U3117 ; P1_R1360_U205
g12384 and P1_R1171_U176 P1_R1171_U175 ; P1_R1171_U4
g12385 and P1_R1171_U177 P1_R1171_U178 ; P1_R1171_U5
g12386 and P1_R1171_U194 P1_R1171_U193 ; P1_R1171_U6
g12387 and P1_R1171_U234 P1_R1171_U233 ; P1_R1171_U7
g12388 and P1_R1171_U243 P1_R1171_U242 ; P1_R1171_U8
g12389 and P1_R1171_U261 P1_R1171_U260 ; P1_R1171_U9
g12390 and P1_R1171_U269 P1_R1171_U268 ; P1_R1171_U10
g12391 and P1_R1171_U348 P1_R1171_U345 ; P1_R1171_U11
g12392 and P1_R1171_U341 P1_R1171_U338 ; P1_R1171_U12
g12393 and P1_R1171_U332 P1_R1171_U329 ; P1_R1171_U13
g12394 and P1_R1171_U323 P1_R1171_U320 ; P1_R1171_U14
g12395 and P1_R1171_U317 P1_R1171_U315 ; P1_R1171_U15
g12396 and P1_R1171_U310 P1_R1171_U307 ; P1_R1171_U16
g12397 and P1_R1171_U232 P1_R1171_U229 ; P1_R1171_U17
g12398 and P1_R1171_U224 P1_R1171_U221 ; P1_R1171_U18
g12399 and P1_R1171_U210 P1_R1171_U207 ; P1_R1171_U19
g12400 not P1_U3471 ; P1_R1171_U20
g12401 not P1_U3069 ; P1_R1171_U21
g12402 not P1_U3068 ; P1_R1171_U22
g12403 nand P1_U3069 P1_U3471 ; P1_R1171_U23
g12404 not P1_U3474 ; P1_R1171_U24
g12405 not P1_U3465 ; P1_R1171_U25
g12406 not P1_U3058 ; P1_R1171_U26
g12407 not P1_U3065 ; P1_R1171_U27
g12408 not P1_U3459 ; P1_R1171_U28
g12409 not P1_U3066 ; P1_R1171_U29
g12410 not P1_U3451 ; P1_R1171_U30
g12411 not P1_U3075 ; P1_R1171_U31
g12412 nand P1_U3075 P1_U3451 ; P1_R1171_U32
g12413 not P1_U3462 ; P1_R1171_U33
g12414 not P1_U3062 ; P1_R1171_U34
g12415 nand P1_U3058 P1_U3465 ; P1_R1171_U35
g12416 not P1_U3468 ; P1_R1171_U36
g12417 not P1_U3477 ; P1_R1171_U37
g12418 not P1_U3082 ; P1_R1171_U38
g12419 not P1_U3081 ; P1_R1171_U39
g12420 not P1_U3480 ; P1_R1171_U40
g12421 nand P1_R1171_U62 P1_R1171_U202 ; P1_R1171_U41
g12422 nand P1_R1171_U118 P1_R1171_U190 ; P1_R1171_U42
g12423 nand P1_R1171_U179 P1_R1171_U180 ; P1_R1171_U43
g12424 nand P1_U3456 P1_U3076 ; P1_R1171_U44
g12425 nand P1_R1171_U122 P1_R1171_U216 ; P1_R1171_U45
g12426 nand P1_R1171_U213 P1_R1171_U212 ; P1_R1171_U46
g12427 not P1_U4008 ; P1_R1171_U47
g12428 not P1_U3051 ; P1_R1171_U48
g12429 not P1_U3055 ; P1_R1171_U49
g12430 not P1_U4009 ; P1_R1171_U50
g12431 not P1_U4010 ; P1_R1171_U51
g12432 not P1_U3056 ; P1_R1171_U52
g12433 not P1_U4011 ; P1_R1171_U53
g12434 not P1_U3063 ; P1_R1171_U54
g12435 not P1_U4014 ; P1_R1171_U55
g12436 not P1_U3073 ; P1_R1171_U56
g12437 not P1_U3501 ; P1_R1171_U57
g12438 not P1_U3071 ; P1_R1171_U58
g12439 not P1_U3067 ; P1_R1171_U59
g12440 nand P1_U3071 P1_U3501 ; P1_R1171_U60
g12441 not P1_U3504 ; P1_R1171_U61
g12442 nand P1_U3082 P1_U3477 ; P1_R1171_U62
g12443 not P1_U3483 ; P1_R1171_U63
g12444 not P1_U3060 ; P1_R1171_U64
g12445 not P1_U3489 ; P1_R1171_U65
g12446 not P1_U3070 ; P1_R1171_U66
g12447 not P1_U3486 ; P1_R1171_U67
g12448 not P1_U3061 ; P1_R1171_U68
g12449 nand P1_U3061 P1_U3486 ; P1_R1171_U69
g12450 not P1_U3492 ; P1_R1171_U70
g12451 not P1_U3078 ; P1_R1171_U71
g12452 not P1_U3495 ; P1_R1171_U72
g12453 not P1_U3077 ; P1_R1171_U73
g12454 not P1_U3498 ; P1_R1171_U74
g12455 not P1_U3072 ; P1_R1171_U75
g12456 not P1_U3507 ; P1_R1171_U76
g12457 not P1_U3080 ; P1_R1171_U77
g12458 nand P1_U3080 P1_U3507 ; P1_R1171_U78
g12459 not P1_U3509 ; P1_R1171_U79
g12460 not P1_U3079 ; P1_R1171_U80
g12461 nand P1_U3079 P1_U3509 ; P1_R1171_U81
g12462 not P1_U4015 ; P1_R1171_U82
g12463 not P1_U4013 ; P1_R1171_U83
g12464 not P1_U3059 ; P1_R1171_U84
g12465 not P1_U4012 ; P1_R1171_U85
g12466 not P1_U3064 ; P1_R1171_U86
g12467 nand P1_U4009 P1_U3055 ; P1_R1171_U87
g12468 not P1_U3052 ; P1_R1171_U88
g12469 not P1_U4007 ; P1_R1171_U89
g12470 nand P1_R1171_U303 P1_R1171_U173 ; P1_R1171_U90
g12471 not P1_U3074 ; P1_R1171_U91
g12472 nand P1_R1171_U78 P1_R1171_U312 ; P1_R1171_U92
g12473 nand P1_R1171_U258 P1_R1171_U257 ; P1_R1171_U93
g12474 nand P1_R1171_U69 P1_R1171_U334 ; P1_R1171_U94
g12475 nand P1_R1171_U454 P1_R1171_U453 ; P1_R1171_U95
g12476 nand P1_R1171_U501 P1_R1171_U500 ; P1_R1171_U96
g12477 nand P1_R1171_U372 P1_R1171_U371 ; P1_R1171_U97
g12478 nand P1_R1171_U377 P1_R1171_U376 ; P1_R1171_U98
g12479 nand P1_R1171_U384 P1_R1171_U383 ; P1_R1171_U99
g12480 nand P1_R1171_U391 P1_R1171_U390 ; P1_R1171_U100
g12481 nand P1_R1171_U396 P1_R1171_U395 ; P1_R1171_U101
g12482 nand P1_R1171_U405 P1_R1171_U404 ; P1_R1171_U102
g12483 nand P1_R1171_U412 P1_R1171_U411 ; P1_R1171_U103
g12484 nand P1_R1171_U419 P1_R1171_U418 ; P1_R1171_U104
g12485 nand P1_R1171_U426 P1_R1171_U425 ; P1_R1171_U105
g12486 nand P1_R1171_U431 P1_R1171_U430 ; P1_R1171_U106
g12487 nand P1_R1171_U438 P1_R1171_U437 ; P1_R1171_U107
g12488 nand P1_R1171_U445 P1_R1171_U444 ; P1_R1171_U108
g12489 nand P1_R1171_U459 P1_R1171_U458 ; P1_R1171_U109
g12490 nand P1_R1171_U464 P1_R1171_U463 ; P1_R1171_U110
g12491 nand P1_R1171_U471 P1_R1171_U470 ; P1_R1171_U111
g12492 nand P1_R1171_U478 P1_R1171_U477 ; P1_R1171_U112
g12493 nand P1_R1171_U485 P1_R1171_U484 ; P1_R1171_U113
g12494 nand P1_R1171_U492 P1_R1171_U491 ; P1_R1171_U114
g12495 nand P1_R1171_U497 P1_R1171_U496 ; P1_R1171_U115
g12496 and P1_U3459 P1_U3066 ; P1_R1171_U116
g12497 and P1_R1171_U186 P1_R1171_U184 ; P1_R1171_U117
g12498 and P1_R1171_U191 P1_R1171_U189 ; P1_R1171_U118
g12499 and P1_R1171_U198 P1_R1171_U197 ; P1_R1171_U119
g12500 and P1_R1171_U379 P1_R1171_U378 P1_R1171_U23 ; P1_R1171_U120
g12501 and P1_R1171_U209 P1_R1171_U6 ; P1_R1171_U121
g12502 and P1_R1171_U217 P1_R1171_U215 ; P1_R1171_U122
g12503 and P1_R1171_U386 P1_R1171_U385 P1_R1171_U35 ; P1_R1171_U123
g12504 and P1_R1171_U223 P1_R1171_U4 ; P1_R1171_U124
g12505 and P1_R1171_U231 P1_R1171_U178 ; P1_R1171_U125
g12506 and P1_R1171_U201 P1_R1171_U7 ; P1_R1171_U126
g12507 and P1_R1171_U236 P1_R1171_U168 ; P1_R1171_U127
g12508 and P1_R1171_U245 P1_R1171_U169 ; P1_R1171_U128
g12509 and P1_R1171_U265 P1_R1171_U264 ; P1_R1171_U129
g12510 and P1_R1171_U10 P1_R1171_U279 ; P1_R1171_U130
g12511 and P1_R1171_U282 P1_R1171_U277 ; P1_R1171_U131
g12512 and P1_R1171_U298 P1_R1171_U295 ; P1_R1171_U132
g12513 and P1_R1171_U365 P1_R1171_U299 ; P1_R1171_U133
g12514 and P1_R1171_U156 P1_R1171_U275 ; P1_R1171_U134
g12515 and P1_R1171_U466 P1_R1171_U465 P1_R1171_U60 ; P1_R1171_U135
g12516 and P1_R1171_U487 P1_R1171_U486 P1_R1171_U169 ; P1_R1171_U136
g12517 and P1_R1171_U340 P1_R1171_U8 ; P1_R1171_U137
g12518 and P1_R1171_U499 P1_R1171_U498 P1_R1171_U168 ; P1_R1171_U138
g12519 and P1_R1171_U347 P1_R1171_U7 ; P1_R1171_U139
g12520 nand P1_R1171_U119 P1_R1171_U199 ; P1_R1171_U140
g12521 nand P1_R1171_U214 P1_R1171_U226 ; P1_R1171_U141
g12522 not P1_U3053 ; P1_R1171_U142
g12523 not P1_U4018 ; P1_R1171_U143
g12524 and P1_R1171_U400 P1_R1171_U399 ; P1_R1171_U144
g12525 nand P1_R1171_U301 P1_R1171_U166 P1_R1171_U361 ; P1_R1171_U145
g12526 and P1_R1171_U407 P1_R1171_U406 ; P1_R1171_U146
g12527 nand P1_R1171_U367 P1_R1171_U366 P1_R1171_U133 ; P1_R1171_U147
g12528 and P1_R1171_U414 P1_R1171_U413 ; P1_R1171_U148
g12529 nand P1_R1171_U362 P1_R1171_U296 P1_R1171_U87 ; P1_R1171_U149
g12530 and P1_R1171_U421 P1_R1171_U420 ; P1_R1171_U150
g12531 nand P1_R1171_U290 P1_R1171_U289 ; P1_R1171_U151
g12532 and P1_R1171_U433 P1_R1171_U432 ; P1_R1171_U152
g12533 nand P1_R1171_U286 P1_R1171_U285 ; P1_R1171_U153
g12534 and P1_R1171_U440 P1_R1171_U439 ; P1_R1171_U154
g12535 nand P1_R1171_U131 P1_R1171_U281 ; P1_R1171_U155
g12536 and P1_R1171_U447 P1_R1171_U446 ; P1_R1171_U156
g12537 and P1_R1171_U452 P1_R1171_U451 ; P1_R1171_U157
g12538 nand P1_R1171_U44 P1_R1171_U324 ; P1_R1171_U158
g12539 nand P1_R1171_U129 P1_R1171_U266 ; P1_R1171_U159
g12540 and P1_R1171_U473 P1_R1171_U472 ; P1_R1171_U160
g12541 nand P1_R1171_U254 P1_R1171_U253 ; P1_R1171_U161
g12542 and P1_R1171_U480 P1_R1171_U479 ; P1_R1171_U162
g12543 nand P1_R1171_U250 P1_R1171_U249 ; P1_R1171_U163
g12544 nand P1_R1171_U240 P1_R1171_U239 ; P1_R1171_U164
g12545 nand P1_R1171_U364 P1_R1171_U363 ; P1_R1171_U165
g12546 nand P1_U3052 P1_R1171_U147 ; P1_R1171_U166
g12547 not P1_R1171_U35 ; P1_R1171_U167
g12548 nand P1_U3480 P1_U3081 ; P1_R1171_U168
g12549 nand P1_U3070 P1_U3489 ; P1_R1171_U169
g12550 nand P1_U3056 P1_U4010 ; P1_R1171_U170
g12551 not P1_R1171_U69 ; P1_R1171_U171
g12552 not P1_R1171_U78 ; P1_R1171_U172
g12553 nand P1_U3063 P1_U4011 ; P1_R1171_U173
g12554 not P1_R1171_U62 ; P1_R1171_U174
g12555 or P1_U3065 P1_U3468 ; P1_R1171_U175
g12556 or P1_U3058 P1_U3465 ; P1_R1171_U176
g12557 or P1_U3462 P1_U3062 ; P1_R1171_U177
g12558 or P1_U3459 P1_U3066 ; P1_R1171_U178
g12559 not P1_R1171_U32 ; P1_R1171_U179
g12560 or P1_U3456 P1_U3076 ; P1_R1171_U180
g12561 not P1_R1171_U43 ; P1_R1171_U181
g12562 not P1_R1171_U44 ; P1_R1171_U182
g12563 nand P1_R1171_U43 P1_R1171_U44 ; P1_R1171_U183
g12564 nand P1_R1171_U116 P1_R1171_U177 ; P1_R1171_U184
g12565 nand P1_R1171_U5 P1_R1171_U183 ; P1_R1171_U185
g12566 nand P1_U3062 P1_U3462 ; P1_R1171_U186
g12567 nand P1_R1171_U117 P1_R1171_U185 ; P1_R1171_U187
g12568 nand P1_R1171_U36 P1_R1171_U35 ; P1_R1171_U188
g12569 nand P1_U3065 P1_R1171_U188 ; P1_R1171_U189
g12570 nand P1_R1171_U4 P1_R1171_U187 ; P1_R1171_U190
g12571 nand P1_U3468 P1_R1171_U167 ; P1_R1171_U191
g12572 not P1_R1171_U42 ; P1_R1171_U192
g12573 or P1_U3068 P1_U3474 ; P1_R1171_U193
g12574 or P1_U3069 P1_U3471 ; P1_R1171_U194
g12575 not P1_R1171_U23 ; P1_R1171_U195
g12576 nand P1_R1171_U24 P1_R1171_U23 ; P1_R1171_U196
g12577 nand P1_U3068 P1_R1171_U196 ; P1_R1171_U197
g12578 nand P1_U3474 P1_R1171_U195 ; P1_R1171_U198
g12579 nand P1_R1171_U6 P1_R1171_U42 ; P1_R1171_U199
g12580 not P1_R1171_U140 ; P1_R1171_U200
g12581 or P1_U3477 P1_U3082 ; P1_R1171_U201
g12582 nand P1_R1171_U201 P1_R1171_U140 ; P1_R1171_U202
g12583 not P1_R1171_U41 ; P1_R1171_U203
g12584 or P1_U3081 P1_U3480 ; P1_R1171_U204
g12585 or P1_U3471 P1_U3069 ; P1_R1171_U205
g12586 nand P1_R1171_U205 P1_R1171_U42 ; P1_R1171_U206
g12587 nand P1_R1171_U120 P1_R1171_U206 ; P1_R1171_U207
g12588 nand P1_R1171_U192 P1_R1171_U23 ; P1_R1171_U208
g12589 nand P1_U3474 P1_U3068 ; P1_R1171_U209
g12590 nand P1_R1171_U121 P1_R1171_U208 ; P1_R1171_U210
g12591 or P1_U3069 P1_U3471 ; P1_R1171_U211
g12592 nand P1_R1171_U182 P1_R1171_U178 ; P1_R1171_U212
g12593 nand P1_U3066 P1_U3459 ; P1_R1171_U213
g12594 not P1_R1171_U46 ; P1_R1171_U214
g12595 nand P1_R1171_U181 P1_R1171_U5 ; P1_R1171_U215
g12596 nand P1_R1171_U46 P1_R1171_U177 ; P1_R1171_U216
g12597 nand P1_U3062 P1_U3462 ; P1_R1171_U217
g12598 not P1_R1171_U45 ; P1_R1171_U218
g12599 or P1_U3465 P1_U3058 ; P1_R1171_U219
g12600 nand P1_R1171_U219 P1_R1171_U45 ; P1_R1171_U220
g12601 nand P1_R1171_U123 P1_R1171_U220 ; P1_R1171_U221
g12602 nand P1_R1171_U218 P1_R1171_U35 ; P1_R1171_U222
g12603 nand P1_U3468 P1_U3065 ; P1_R1171_U223
g12604 nand P1_R1171_U124 P1_R1171_U222 ; P1_R1171_U224
g12605 or P1_U3058 P1_U3465 ; P1_R1171_U225
g12606 nand P1_R1171_U181 P1_R1171_U178 ; P1_R1171_U226
g12607 not P1_R1171_U141 ; P1_R1171_U227
g12608 nand P1_U3062 P1_U3462 ; P1_R1171_U228
g12609 nand P1_R1171_U398 P1_R1171_U397 P1_R1171_U44 P1_R1171_U43 ; P1_R1171_U229
g12610 nand P1_R1171_U44 P1_R1171_U43 ; P1_R1171_U230
g12611 nand P1_U3066 P1_U3459 ; P1_R1171_U231
g12612 nand P1_R1171_U125 P1_R1171_U230 ; P1_R1171_U232
g12613 or P1_U3081 P1_U3480 ; P1_R1171_U233
g12614 or P1_U3060 P1_U3483 ; P1_R1171_U234
g12615 nand P1_R1171_U174 P1_R1171_U7 ; P1_R1171_U235
g12616 nand P1_U3060 P1_U3483 ; P1_R1171_U236
g12617 nand P1_R1171_U127 P1_R1171_U235 ; P1_R1171_U237
g12618 or P1_U3483 P1_U3060 ; P1_R1171_U238
g12619 nand P1_R1171_U126 P1_R1171_U140 ; P1_R1171_U239
g12620 nand P1_R1171_U238 P1_R1171_U237 ; P1_R1171_U240
g12621 not P1_R1171_U164 ; P1_R1171_U241
g12622 or P1_U3078 P1_U3492 ; P1_R1171_U242
g12623 or P1_U3070 P1_U3489 ; P1_R1171_U243
g12624 nand P1_R1171_U171 P1_R1171_U8 ; P1_R1171_U244
g12625 nand P1_U3078 P1_U3492 ; P1_R1171_U245
g12626 nand P1_R1171_U128 P1_R1171_U244 ; P1_R1171_U246
g12627 or P1_U3486 P1_U3061 ; P1_R1171_U247
g12628 or P1_U3492 P1_U3078 ; P1_R1171_U248
g12629 nand P1_R1171_U247 P1_R1171_U164 P1_R1171_U8 ; P1_R1171_U249
g12630 nand P1_R1171_U248 P1_R1171_U246 ; P1_R1171_U250
g12631 not P1_R1171_U163 ; P1_R1171_U251
g12632 or P1_U3495 P1_U3077 ; P1_R1171_U252
g12633 nand P1_R1171_U252 P1_R1171_U163 ; P1_R1171_U253
g12634 nand P1_U3077 P1_U3495 ; P1_R1171_U254
g12635 not P1_R1171_U161 ; P1_R1171_U255
g12636 or P1_U3498 P1_U3072 ; P1_R1171_U256
g12637 nand P1_R1171_U256 P1_R1171_U161 ; P1_R1171_U257
g12638 nand P1_U3072 P1_U3498 ; P1_R1171_U258
g12639 not P1_R1171_U93 ; P1_R1171_U259
g12640 or P1_U3067 P1_U3504 ; P1_R1171_U260
g12641 or P1_U3071 P1_U3501 ; P1_R1171_U261
g12642 not P1_R1171_U60 ; P1_R1171_U262
g12643 nand P1_R1171_U61 P1_R1171_U60 ; P1_R1171_U263
g12644 nand P1_U3067 P1_R1171_U263 ; P1_R1171_U264
g12645 nand P1_U3504 P1_R1171_U262 ; P1_R1171_U265
g12646 nand P1_R1171_U9 P1_R1171_U93 ; P1_R1171_U266
g12647 not P1_R1171_U159 ; P1_R1171_U267
g12648 or P1_U3074 P1_U4015 ; P1_R1171_U268
g12649 or P1_U3079 P1_U3509 ; P1_R1171_U269
g12650 or P1_U3073 P1_U4014 ; P1_R1171_U270
g12651 not P1_R1171_U81 ; P1_R1171_U271
g12652 nand P1_U4015 P1_R1171_U271 ; P1_R1171_U272
g12653 nand P1_R1171_U272 P1_R1171_U91 ; P1_R1171_U273
g12654 nand P1_R1171_U81 P1_R1171_U82 ; P1_R1171_U274
g12655 nand P1_R1171_U274 P1_R1171_U273 ; P1_R1171_U275
g12656 nand P1_R1171_U172 P1_R1171_U10 ; P1_R1171_U276
g12657 nand P1_U3073 P1_U4014 ; P1_R1171_U277
g12658 nand P1_R1171_U275 P1_R1171_U276 ; P1_R1171_U278
g12659 or P1_U3507 P1_U3080 ; P1_R1171_U279
g12660 or P1_U4014 P1_U3073 ; P1_R1171_U280
g12661 nand P1_R1171_U270 P1_R1171_U159 P1_R1171_U130 ; P1_R1171_U281
g12662 nand P1_R1171_U280 P1_R1171_U278 ; P1_R1171_U282
g12663 not P1_R1171_U155 ; P1_R1171_U283
g12664 or P1_U4013 P1_U3059 ; P1_R1171_U284
g12665 nand P1_R1171_U284 P1_R1171_U155 ; P1_R1171_U285
g12666 nand P1_U3059 P1_U4013 ; P1_R1171_U286
g12667 not P1_R1171_U153 ; P1_R1171_U287
g12668 or P1_U4012 P1_U3064 ; P1_R1171_U288
g12669 nand P1_R1171_U288 P1_R1171_U153 ; P1_R1171_U289
g12670 nand P1_U3064 P1_U4012 ; P1_R1171_U290
g12671 not P1_R1171_U151 ; P1_R1171_U291
g12672 or P1_U3056 P1_U4010 ; P1_R1171_U292
g12673 nand P1_R1171_U173 P1_R1171_U170 ; P1_R1171_U293
g12674 not P1_R1171_U87 ; P1_R1171_U294
g12675 or P1_U4011 P1_U3063 ; P1_R1171_U295
g12676 nand P1_R1171_U151 P1_R1171_U295 P1_R1171_U165 ; P1_R1171_U296
g12677 not P1_R1171_U149 ; P1_R1171_U297
g12678 or P1_U4008 P1_U3051 ; P1_R1171_U298
g12679 nand P1_U3051 P1_U4008 ; P1_R1171_U299
g12680 not P1_R1171_U147 ; P1_R1171_U300
g12681 nand P1_U4007 P1_R1171_U147 ; P1_R1171_U301
g12682 not P1_R1171_U145 ; P1_R1171_U302
g12683 nand P1_R1171_U295 P1_R1171_U151 ; P1_R1171_U303
g12684 not P1_R1171_U90 ; P1_R1171_U304
g12685 or P1_U4010 P1_U3056 ; P1_R1171_U305
g12686 nand P1_R1171_U305 P1_R1171_U90 ; P1_R1171_U306
g12687 nand P1_R1171_U306 P1_R1171_U170 P1_R1171_U150 ; P1_R1171_U307
g12688 nand P1_R1171_U304 P1_R1171_U170 ; P1_R1171_U308
g12689 nand P1_U4009 P1_U3055 ; P1_R1171_U309
g12690 nand P1_R1171_U308 P1_R1171_U309 P1_R1171_U165 ; P1_R1171_U310
g12691 or P1_U3056 P1_U4010 ; P1_R1171_U311
g12692 nand P1_R1171_U279 P1_R1171_U159 ; P1_R1171_U312
g12693 not P1_R1171_U92 ; P1_R1171_U313
g12694 nand P1_R1171_U10 P1_R1171_U92 ; P1_R1171_U314
g12695 nand P1_R1171_U134 P1_R1171_U314 ; P1_R1171_U315
g12696 nand P1_R1171_U314 P1_R1171_U275 ; P1_R1171_U316
g12697 nand P1_R1171_U450 P1_R1171_U316 ; P1_R1171_U317
g12698 or P1_U3509 P1_U3079 ; P1_R1171_U318
g12699 nand P1_R1171_U318 P1_R1171_U92 ; P1_R1171_U319
g12700 nand P1_R1171_U319 P1_R1171_U81 P1_R1171_U157 ; P1_R1171_U320
g12701 nand P1_R1171_U313 P1_R1171_U81 ; P1_R1171_U321
g12702 nand P1_U3074 P1_U4015 ; P1_R1171_U322
g12703 nand P1_R1171_U322 P1_R1171_U321 P1_R1171_U10 ; P1_R1171_U323
g12704 or P1_U3456 P1_U3076 ; P1_R1171_U324
g12705 not P1_R1171_U158 ; P1_R1171_U325
g12706 or P1_U3079 P1_U3509 ; P1_R1171_U326
g12707 or P1_U3501 P1_U3071 ; P1_R1171_U327
g12708 nand P1_R1171_U327 P1_R1171_U93 ; P1_R1171_U328
g12709 nand P1_R1171_U135 P1_R1171_U328 ; P1_R1171_U329
g12710 nand P1_R1171_U259 P1_R1171_U60 ; P1_R1171_U330
g12711 nand P1_U3504 P1_U3067 ; P1_R1171_U331
g12712 nand P1_R1171_U331 P1_R1171_U330 P1_R1171_U9 ; P1_R1171_U332
g12713 or P1_U3071 P1_U3501 ; P1_R1171_U333
g12714 nand P1_R1171_U247 P1_R1171_U164 ; P1_R1171_U334
g12715 not P1_R1171_U94 ; P1_R1171_U335
g12716 or P1_U3489 P1_U3070 ; P1_R1171_U336
g12717 nand P1_R1171_U336 P1_R1171_U94 ; P1_R1171_U337
g12718 nand P1_R1171_U136 P1_R1171_U337 ; P1_R1171_U338
g12719 nand P1_R1171_U335 P1_R1171_U169 ; P1_R1171_U339
g12720 nand P1_U3078 P1_U3492 ; P1_R1171_U340
g12721 nand P1_R1171_U137 P1_R1171_U339 ; P1_R1171_U341
g12722 or P1_U3070 P1_U3489 ; P1_R1171_U342
g12723 or P1_U3480 P1_U3081 ; P1_R1171_U343
g12724 nand P1_R1171_U343 P1_R1171_U41 ; P1_R1171_U344
g12725 nand P1_R1171_U138 P1_R1171_U344 ; P1_R1171_U345
g12726 nand P1_R1171_U203 P1_R1171_U168 ; P1_R1171_U346
g12727 nand P1_U3060 P1_U3483 ; P1_R1171_U347
g12728 nand P1_R1171_U139 P1_R1171_U346 ; P1_R1171_U348
g12729 nand P1_R1171_U204 P1_R1171_U168 ; P1_R1171_U349
g12730 nand P1_R1171_U201 P1_R1171_U62 ; P1_R1171_U350
g12731 nand P1_R1171_U211 P1_R1171_U23 ; P1_R1171_U351
g12732 nand P1_R1171_U225 P1_R1171_U35 ; P1_R1171_U352
g12733 nand P1_R1171_U228 P1_R1171_U177 ; P1_R1171_U353
g12734 nand P1_R1171_U311 P1_R1171_U170 ; P1_R1171_U354
g12735 nand P1_R1171_U295 P1_R1171_U173 ; P1_R1171_U355
g12736 nand P1_R1171_U326 P1_R1171_U81 ; P1_R1171_U356
g12737 nand P1_R1171_U279 P1_R1171_U78 ; P1_R1171_U357
g12738 nand P1_R1171_U333 P1_R1171_U60 ; P1_R1171_U358
g12739 nand P1_R1171_U342 P1_R1171_U169 ; P1_R1171_U359
g12740 nand P1_R1171_U247 P1_R1171_U69 ; P1_R1171_U360
g12741 nand P1_U4007 P1_U3052 ; P1_R1171_U361
g12742 nand P1_R1171_U293 P1_R1171_U165 ; P1_R1171_U362
g12743 nand P1_U3055 P1_R1171_U292 ; P1_R1171_U363
g12744 nand P1_U4009 P1_R1171_U292 ; P1_R1171_U364
g12745 nand P1_R1171_U293 P1_R1171_U165 P1_R1171_U298 ; P1_R1171_U365
g12746 nand P1_R1171_U151 P1_R1171_U165 P1_R1171_U132 ; P1_R1171_U366
g12747 nand P1_R1171_U294 P1_R1171_U298 ; P1_R1171_U367
g12748 nand P1_U3081 P1_R1171_U40 ; P1_R1171_U368
g12749 nand P1_U3480 P1_R1171_U39 ; P1_R1171_U369
g12750 nand P1_R1171_U369 P1_R1171_U368 ; P1_R1171_U370
g12751 nand P1_R1171_U349 P1_R1171_U41 ; P1_R1171_U371
g12752 nand P1_R1171_U370 P1_R1171_U203 ; P1_R1171_U372
g12753 nand P1_U3082 P1_R1171_U37 ; P1_R1171_U373
g12754 nand P1_U3477 P1_R1171_U38 ; P1_R1171_U374
g12755 nand P1_R1171_U374 P1_R1171_U373 ; P1_R1171_U375
g12756 nand P1_R1171_U350 P1_R1171_U140 ; P1_R1171_U376
g12757 nand P1_R1171_U200 P1_R1171_U375 ; P1_R1171_U377
g12758 nand P1_U3068 P1_R1171_U24 ; P1_R1171_U378
g12759 nand P1_U3474 P1_R1171_U22 ; P1_R1171_U379
g12760 nand P1_U3069 P1_R1171_U20 ; P1_R1171_U380
g12761 nand P1_U3471 P1_R1171_U21 ; P1_R1171_U381
g12762 nand P1_R1171_U381 P1_R1171_U380 ; P1_R1171_U382
g12763 nand P1_R1171_U351 P1_R1171_U42 ; P1_R1171_U383
g12764 nand P1_R1171_U382 P1_R1171_U192 ; P1_R1171_U384
g12765 nand P1_U3065 P1_R1171_U36 ; P1_R1171_U385
g12766 nand P1_U3468 P1_R1171_U27 ; P1_R1171_U386
g12767 nand P1_U3058 P1_R1171_U25 ; P1_R1171_U387
g12768 nand P1_U3465 P1_R1171_U26 ; P1_R1171_U388
g12769 nand P1_R1171_U388 P1_R1171_U387 ; P1_R1171_U389
g12770 nand P1_R1171_U352 P1_R1171_U45 ; P1_R1171_U390
g12771 nand P1_R1171_U389 P1_R1171_U218 ; P1_R1171_U391
g12772 nand P1_U3062 P1_R1171_U33 ; P1_R1171_U392
g12773 nand P1_U3462 P1_R1171_U34 ; P1_R1171_U393
g12774 nand P1_R1171_U393 P1_R1171_U392 ; P1_R1171_U394
g12775 nand P1_R1171_U353 P1_R1171_U141 ; P1_R1171_U395
g12776 nand P1_R1171_U227 P1_R1171_U394 ; P1_R1171_U396
g12777 nand P1_U3066 P1_R1171_U28 ; P1_R1171_U397
g12778 nand P1_U3459 P1_R1171_U29 ; P1_R1171_U398
g12779 nand P1_U3053 P1_R1171_U143 ; P1_R1171_U399
g12780 nand P1_U4018 P1_R1171_U142 ; P1_R1171_U400
g12781 nand P1_U3053 P1_R1171_U143 ; P1_R1171_U401
g12782 nand P1_U4018 P1_R1171_U142 ; P1_R1171_U402
g12783 nand P1_R1171_U402 P1_R1171_U401 ; P1_R1171_U403
g12784 nand P1_R1171_U144 P1_R1171_U145 ; P1_R1171_U404
g12785 nand P1_R1171_U302 P1_R1171_U403 ; P1_R1171_U405
g12786 nand P1_U3052 P1_R1171_U89 ; P1_R1171_U406
g12787 nand P1_U4007 P1_R1171_U88 ; P1_R1171_U407
g12788 nand P1_U3052 P1_R1171_U89 ; P1_R1171_U408
g12789 nand P1_U4007 P1_R1171_U88 ; P1_R1171_U409
g12790 nand P1_R1171_U409 P1_R1171_U408 ; P1_R1171_U410
g12791 nand P1_R1171_U146 P1_R1171_U147 ; P1_R1171_U411
g12792 nand P1_R1171_U300 P1_R1171_U410 ; P1_R1171_U412
g12793 nand P1_U3051 P1_R1171_U47 ; P1_R1171_U413
g12794 nand P1_U4008 P1_R1171_U48 ; P1_R1171_U414
g12795 nand P1_U3051 P1_R1171_U47 ; P1_R1171_U415
g12796 nand P1_U4008 P1_R1171_U48 ; P1_R1171_U416
g12797 nand P1_R1171_U416 P1_R1171_U415 ; P1_R1171_U417
g12798 nand P1_R1171_U148 P1_R1171_U149 ; P1_R1171_U418
g12799 nand P1_R1171_U297 P1_R1171_U417 ; P1_R1171_U419
g12800 nand P1_U3055 P1_R1171_U50 ; P1_R1171_U420
g12801 nand P1_U4009 P1_R1171_U49 ; P1_R1171_U421
g12802 nand P1_U3056 P1_R1171_U51 ; P1_R1171_U422
g12803 nand P1_U4010 P1_R1171_U52 ; P1_R1171_U423
g12804 nand P1_R1171_U423 P1_R1171_U422 ; P1_R1171_U424
g12805 nand P1_R1171_U354 P1_R1171_U90 ; P1_R1171_U425
g12806 nand P1_R1171_U424 P1_R1171_U304 ; P1_R1171_U426
g12807 nand P1_U3063 P1_R1171_U53 ; P1_R1171_U427
g12808 nand P1_U4011 P1_R1171_U54 ; P1_R1171_U428
g12809 nand P1_R1171_U428 P1_R1171_U427 ; P1_R1171_U429
g12810 nand P1_R1171_U355 P1_R1171_U151 ; P1_R1171_U430
g12811 nand P1_R1171_U291 P1_R1171_U429 ; P1_R1171_U431
g12812 nand P1_U3064 P1_R1171_U85 ; P1_R1171_U432
g12813 nand P1_U4012 P1_R1171_U86 ; P1_R1171_U433
g12814 nand P1_U3064 P1_R1171_U85 ; P1_R1171_U434
g12815 nand P1_U4012 P1_R1171_U86 ; P1_R1171_U435
g12816 nand P1_R1171_U435 P1_R1171_U434 ; P1_R1171_U436
g12817 nand P1_R1171_U152 P1_R1171_U153 ; P1_R1171_U437
g12818 nand P1_R1171_U287 P1_R1171_U436 ; P1_R1171_U438
g12819 nand P1_U3059 P1_R1171_U83 ; P1_R1171_U439
g12820 nand P1_U4013 P1_R1171_U84 ; P1_R1171_U440
g12821 nand P1_U3059 P1_R1171_U83 ; P1_R1171_U441
g12822 nand P1_U4013 P1_R1171_U84 ; P1_R1171_U442
g12823 nand P1_R1171_U442 P1_R1171_U441 ; P1_R1171_U443
g12824 nand P1_R1171_U154 P1_R1171_U155 ; P1_R1171_U444
g12825 nand P1_R1171_U283 P1_R1171_U443 ; P1_R1171_U445
g12826 nand P1_U3073 P1_R1171_U55 ; P1_R1171_U446
g12827 nand P1_U4014 P1_R1171_U56 ; P1_R1171_U447
g12828 nand P1_U3073 P1_R1171_U55 ; P1_R1171_U448
g12829 nand P1_U4014 P1_R1171_U56 ; P1_R1171_U449
g12830 nand P1_R1171_U449 P1_R1171_U448 ; P1_R1171_U450
g12831 nand P1_U3074 P1_R1171_U82 ; P1_R1171_U451
g12832 nand P1_U4015 P1_R1171_U91 ; P1_R1171_U452
g12833 nand P1_R1171_U179 P1_R1171_U158 ; P1_R1171_U453
g12834 nand P1_R1171_U325 P1_R1171_U32 ; P1_R1171_U454
g12835 nand P1_U3079 P1_R1171_U79 ; P1_R1171_U455
g12836 nand P1_U3509 P1_R1171_U80 ; P1_R1171_U456
g12837 nand P1_R1171_U456 P1_R1171_U455 ; P1_R1171_U457
g12838 nand P1_R1171_U356 P1_R1171_U92 ; P1_R1171_U458
g12839 nand P1_R1171_U457 P1_R1171_U313 ; P1_R1171_U459
g12840 nand P1_U3080 P1_R1171_U76 ; P1_R1171_U460
g12841 nand P1_U3507 P1_R1171_U77 ; P1_R1171_U461
g12842 nand P1_R1171_U461 P1_R1171_U460 ; P1_R1171_U462
g12843 nand P1_R1171_U357 P1_R1171_U159 ; P1_R1171_U463
g12844 nand P1_R1171_U267 P1_R1171_U462 ; P1_R1171_U464
g12845 nand P1_U3067 P1_R1171_U61 ; P1_R1171_U465
g12846 nand P1_U3504 P1_R1171_U59 ; P1_R1171_U466
g12847 nand P1_U3071 P1_R1171_U57 ; P1_R1171_U467
g12848 nand P1_U3501 P1_R1171_U58 ; P1_R1171_U468
g12849 nand P1_R1171_U468 P1_R1171_U467 ; P1_R1171_U469
g12850 nand P1_R1171_U358 P1_R1171_U93 ; P1_R1171_U470
g12851 nand P1_R1171_U469 P1_R1171_U259 ; P1_R1171_U471
g12852 nand P1_U3072 P1_R1171_U74 ; P1_R1171_U472
g12853 nand P1_U3498 P1_R1171_U75 ; P1_R1171_U473
g12854 nand P1_U3072 P1_R1171_U74 ; P1_R1171_U474
g12855 nand P1_U3498 P1_R1171_U75 ; P1_R1171_U475
g12856 nand P1_R1171_U475 P1_R1171_U474 ; P1_R1171_U476
g12857 nand P1_R1171_U160 P1_R1171_U161 ; P1_R1171_U477
g12858 nand P1_R1171_U255 P1_R1171_U476 ; P1_R1171_U478
g12859 nand P1_U3077 P1_R1171_U72 ; P1_R1171_U479
g12860 nand P1_U3495 P1_R1171_U73 ; P1_R1171_U480
g12861 nand P1_U3077 P1_R1171_U72 ; P1_R1171_U481
g12862 nand P1_U3495 P1_R1171_U73 ; P1_R1171_U482
g12863 nand P1_R1171_U482 P1_R1171_U481 ; P1_R1171_U483
g12864 nand P1_R1171_U162 P1_R1171_U163 ; P1_R1171_U484
g12865 nand P1_R1171_U251 P1_R1171_U483 ; P1_R1171_U485
g12866 nand P1_U3078 P1_R1171_U70 ; P1_R1171_U486
g12867 nand P1_U3492 P1_R1171_U71 ; P1_R1171_U487
g12868 nand P1_U3070 P1_R1171_U65 ; P1_R1171_U488
g12869 nand P1_U3489 P1_R1171_U66 ; P1_R1171_U489
g12870 nand P1_R1171_U489 P1_R1171_U488 ; P1_R1171_U490
g12871 nand P1_R1171_U359 P1_R1171_U94 ; P1_R1171_U491
g12872 nand P1_R1171_U490 P1_R1171_U335 ; P1_R1171_U492
g12873 nand P1_U3061 P1_R1171_U67 ; P1_R1171_U493
g12874 nand P1_U3486 P1_R1171_U68 ; P1_R1171_U494
g12875 nand P1_R1171_U494 P1_R1171_U493 ; P1_R1171_U495
g12876 nand P1_R1171_U360 P1_R1171_U164 ; P1_R1171_U496
g12877 nand P1_R1171_U241 P1_R1171_U495 ; P1_R1171_U497
g12878 nand P1_U3060 P1_R1171_U63 ; P1_R1171_U498
g12879 nand P1_U3483 P1_R1171_U64 ; P1_R1171_U499
g12880 nand P1_U3075 P1_R1171_U30 ; P1_R1171_U500
g12881 nand P1_U3451 P1_R1171_U31 ; P1_R1171_U501
g12882 and P1_R1138_U176 P1_R1138_U175 ; P1_R1138_U4
g12883 and P1_R1138_U177 P1_R1138_U178 ; P1_R1138_U5
g12884 and P1_R1138_U194 P1_R1138_U193 ; P1_R1138_U6
g12885 and P1_R1138_U234 P1_R1138_U233 ; P1_R1138_U7
g12886 and P1_R1138_U243 P1_R1138_U242 ; P1_R1138_U8
g12887 and P1_R1138_U261 P1_R1138_U260 ; P1_R1138_U9
g12888 and P1_R1138_U269 P1_R1138_U268 ; P1_R1138_U10
g12889 and P1_R1138_U348 P1_R1138_U345 ; P1_R1138_U11
g12890 and P1_R1138_U341 P1_R1138_U338 ; P1_R1138_U12
g12891 and P1_R1138_U332 P1_R1138_U329 ; P1_R1138_U13
g12892 and P1_R1138_U323 P1_R1138_U320 ; P1_R1138_U14
g12893 and P1_R1138_U317 P1_R1138_U315 ; P1_R1138_U15
g12894 and P1_R1138_U310 P1_R1138_U307 ; P1_R1138_U16
g12895 and P1_R1138_U232 P1_R1138_U229 ; P1_R1138_U17
g12896 and P1_R1138_U224 P1_R1138_U221 ; P1_R1138_U18
g12897 and P1_R1138_U210 P1_R1138_U207 ; P1_R1138_U19
g12898 not P1_U3471 ; P1_R1138_U20
g12899 not P1_U3069 ; P1_R1138_U21
g12900 not P1_U3068 ; P1_R1138_U22
g12901 nand P1_U3069 P1_U3471 ; P1_R1138_U23
g12902 not P1_U3474 ; P1_R1138_U24
g12903 not P1_U3465 ; P1_R1138_U25
g12904 not P1_U3058 ; P1_R1138_U26
g12905 not P1_U3065 ; P1_R1138_U27
g12906 not P1_U3459 ; P1_R1138_U28
g12907 not P1_U3066 ; P1_R1138_U29
g12908 not P1_U3451 ; P1_R1138_U30
g12909 not P1_U3075 ; P1_R1138_U31
g12910 nand P1_U3075 P1_U3451 ; P1_R1138_U32
g12911 not P1_U3462 ; P1_R1138_U33
g12912 not P1_U3062 ; P1_R1138_U34
g12913 nand P1_U3058 P1_U3465 ; P1_R1138_U35
g12914 not P1_U3468 ; P1_R1138_U36
g12915 not P1_U3477 ; P1_R1138_U37
g12916 not P1_U3082 ; P1_R1138_U38
g12917 not P1_U3081 ; P1_R1138_U39
g12918 not P1_U3480 ; P1_R1138_U40
g12919 nand P1_R1138_U62 P1_R1138_U202 ; P1_R1138_U41
g12920 nand P1_R1138_U118 P1_R1138_U190 ; P1_R1138_U42
g12921 nand P1_R1138_U179 P1_R1138_U180 ; P1_R1138_U43
g12922 nand P1_U3456 P1_U3076 ; P1_R1138_U44
g12923 nand P1_R1138_U122 P1_R1138_U216 ; P1_R1138_U45
g12924 nand P1_R1138_U213 P1_R1138_U212 ; P1_R1138_U46
g12925 not P1_U4008 ; P1_R1138_U47
g12926 not P1_U3051 ; P1_R1138_U48
g12927 not P1_U3055 ; P1_R1138_U49
g12928 not P1_U4009 ; P1_R1138_U50
g12929 not P1_U4010 ; P1_R1138_U51
g12930 not P1_U3056 ; P1_R1138_U52
g12931 not P1_U4011 ; P1_R1138_U53
g12932 not P1_U3063 ; P1_R1138_U54
g12933 not P1_U4014 ; P1_R1138_U55
g12934 not P1_U3073 ; P1_R1138_U56
g12935 not P1_U3501 ; P1_R1138_U57
g12936 not P1_U3071 ; P1_R1138_U58
g12937 not P1_U3067 ; P1_R1138_U59
g12938 nand P1_U3071 P1_U3501 ; P1_R1138_U60
g12939 not P1_U3504 ; P1_R1138_U61
g12940 nand P1_U3082 P1_U3477 ; P1_R1138_U62
g12941 not P1_U3483 ; P1_R1138_U63
g12942 not P1_U3060 ; P1_R1138_U64
g12943 not P1_U3489 ; P1_R1138_U65
g12944 not P1_U3070 ; P1_R1138_U66
g12945 not P1_U3486 ; P1_R1138_U67
g12946 not P1_U3061 ; P1_R1138_U68
g12947 nand P1_U3061 P1_U3486 ; P1_R1138_U69
g12948 not P1_U3492 ; P1_R1138_U70
g12949 not P1_U3078 ; P1_R1138_U71
g12950 not P1_U3495 ; P1_R1138_U72
g12951 not P1_U3077 ; P1_R1138_U73
g12952 not P1_U3498 ; P1_R1138_U74
g12953 not P1_U3072 ; P1_R1138_U75
g12954 not P1_U3507 ; P1_R1138_U76
g12955 not P1_U3080 ; P1_R1138_U77
g12956 nand P1_U3080 P1_U3507 ; P1_R1138_U78
g12957 not P1_U3509 ; P1_R1138_U79
g12958 not P1_U3079 ; P1_R1138_U80
g12959 nand P1_U3079 P1_U3509 ; P1_R1138_U81
g12960 not P1_U4015 ; P1_R1138_U82
g12961 not P1_U4013 ; P1_R1138_U83
g12962 not P1_U3059 ; P1_R1138_U84
g12963 not P1_U4012 ; P1_R1138_U85
g12964 not P1_U3064 ; P1_R1138_U86
g12965 nand P1_U4009 P1_U3055 ; P1_R1138_U87
g12966 not P1_U3052 ; P1_R1138_U88
g12967 not P1_U4007 ; P1_R1138_U89
g12968 nand P1_R1138_U303 P1_R1138_U173 ; P1_R1138_U90
g12969 not P1_U3074 ; P1_R1138_U91
g12970 nand P1_R1138_U78 P1_R1138_U312 ; P1_R1138_U92
g12971 nand P1_R1138_U258 P1_R1138_U257 ; P1_R1138_U93
g12972 nand P1_R1138_U69 P1_R1138_U334 ; P1_R1138_U94
g12973 nand P1_R1138_U454 P1_R1138_U453 ; P1_R1138_U95
g12974 nand P1_R1138_U501 P1_R1138_U500 ; P1_R1138_U96
g12975 nand P1_R1138_U372 P1_R1138_U371 ; P1_R1138_U97
g12976 nand P1_R1138_U377 P1_R1138_U376 ; P1_R1138_U98
g12977 nand P1_R1138_U384 P1_R1138_U383 ; P1_R1138_U99
g12978 nand P1_R1138_U391 P1_R1138_U390 ; P1_R1138_U100
g12979 nand P1_R1138_U396 P1_R1138_U395 ; P1_R1138_U101
g12980 nand P1_R1138_U405 P1_R1138_U404 ; P1_R1138_U102
g12981 nand P1_R1138_U412 P1_R1138_U411 ; P1_R1138_U103
g12982 nand P1_R1138_U419 P1_R1138_U418 ; P1_R1138_U104
g12983 nand P1_R1138_U426 P1_R1138_U425 ; P1_R1138_U105
g12984 nand P1_R1138_U431 P1_R1138_U430 ; P1_R1138_U106
g12985 nand P1_R1138_U438 P1_R1138_U437 ; P1_R1138_U107
g12986 nand P1_R1138_U445 P1_R1138_U444 ; P1_R1138_U108
g12987 nand P1_R1138_U459 P1_R1138_U458 ; P1_R1138_U109
g12988 nand P1_R1138_U464 P1_R1138_U463 ; P1_R1138_U110
g12989 nand P1_R1138_U471 P1_R1138_U470 ; P1_R1138_U111
g12990 nand P1_R1138_U478 P1_R1138_U477 ; P1_R1138_U112
g12991 nand P1_R1138_U485 P1_R1138_U484 ; P1_R1138_U113
g12992 nand P1_R1138_U492 P1_R1138_U491 ; P1_R1138_U114
g12993 nand P1_R1138_U497 P1_R1138_U496 ; P1_R1138_U115
g12994 and P1_U3459 P1_U3066 ; P1_R1138_U116
g12995 and P1_R1138_U186 P1_R1138_U184 ; P1_R1138_U117
g12996 and P1_R1138_U191 P1_R1138_U189 ; P1_R1138_U118
g12997 and P1_R1138_U198 P1_R1138_U197 ; P1_R1138_U119
g12998 and P1_R1138_U379 P1_R1138_U378 P1_R1138_U23 ; P1_R1138_U120
g12999 and P1_R1138_U209 P1_R1138_U6 ; P1_R1138_U121
g13000 and P1_R1138_U217 P1_R1138_U215 ; P1_R1138_U122
g13001 and P1_R1138_U386 P1_R1138_U385 P1_R1138_U35 ; P1_R1138_U123
g13002 and P1_R1138_U223 P1_R1138_U4 ; P1_R1138_U124
g13003 and P1_R1138_U231 P1_R1138_U178 ; P1_R1138_U125
g13004 and P1_R1138_U201 P1_R1138_U7 ; P1_R1138_U126
g13005 and P1_R1138_U236 P1_R1138_U168 ; P1_R1138_U127
g13006 and P1_R1138_U245 P1_R1138_U169 ; P1_R1138_U128
g13007 and P1_R1138_U265 P1_R1138_U264 ; P1_R1138_U129
g13008 and P1_R1138_U10 P1_R1138_U279 ; P1_R1138_U130
g13009 and P1_R1138_U282 P1_R1138_U277 ; P1_R1138_U131
g13010 and P1_R1138_U298 P1_R1138_U295 ; P1_R1138_U132
g13011 and P1_R1138_U365 P1_R1138_U299 ; P1_R1138_U133
g13012 and P1_R1138_U156 P1_R1138_U275 ; P1_R1138_U134
g13013 and P1_R1138_U466 P1_R1138_U465 P1_R1138_U60 ; P1_R1138_U135
g13014 and P1_R1138_U487 P1_R1138_U486 P1_R1138_U169 ; P1_R1138_U136
g13015 and P1_R1138_U340 P1_R1138_U8 ; P1_R1138_U137
g13016 and P1_R1138_U499 P1_R1138_U498 P1_R1138_U168 ; P1_R1138_U138
g13017 and P1_R1138_U347 P1_R1138_U7 ; P1_R1138_U139
g13018 nand P1_R1138_U119 P1_R1138_U199 ; P1_R1138_U140
g13019 nand P1_R1138_U214 P1_R1138_U226 ; P1_R1138_U141
g13020 not P1_U3053 ; P1_R1138_U142
g13021 not P1_U4018 ; P1_R1138_U143
g13022 and P1_R1138_U400 P1_R1138_U399 ; P1_R1138_U144
g13023 nand P1_R1138_U301 P1_R1138_U166 P1_R1138_U361 ; P1_R1138_U145
g13024 and P1_R1138_U407 P1_R1138_U406 ; P1_R1138_U146
g13025 nand P1_R1138_U367 P1_R1138_U366 P1_R1138_U133 ; P1_R1138_U147
g13026 and P1_R1138_U414 P1_R1138_U413 ; P1_R1138_U148
g13027 nand P1_R1138_U362 P1_R1138_U296 P1_R1138_U87 ; P1_R1138_U149
g13028 and P1_R1138_U421 P1_R1138_U420 ; P1_R1138_U150
g13029 nand P1_R1138_U290 P1_R1138_U289 ; P1_R1138_U151
g13030 and P1_R1138_U433 P1_R1138_U432 ; P1_R1138_U152
g13031 nand P1_R1138_U286 P1_R1138_U285 ; P1_R1138_U153
g13032 and P1_R1138_U440 P1_R1138_U439 ; P1_R1138_U154
g13033 nand P1_R1138_U131 P1_R1138_U281 ; P1_R1138_U155
g13034 and P1_R1138_U447 P1_R1138_U446 ; P1_R1138_U156
g13035 and P1_R1138_U452 P1_R1138_U451 ; P1_R1138_U157
g13036 nand P1_R1138_U44 P1_R1138_U324 ; P1_R1138_U158
g13037 nand P1_R1138_U129 P1_R1138_U266 ; P1_R1138_U159
g13038 and P1_R1138_U473 P1_R1138_U472 ; P1_R1138_U160
g13039 nand P1_R1138_U254 P1_R1138_U253 ; P1_R1138_U161
g13040 and P1_R1138_U480 P1_R1138_U479 ; P1_R1138_U162
g13041 nand P1_R1138_U250 P1_R1138_U249 ; P1_R1138_U163
g13042 nand P1_R1138_U240 P1_R1138_U239 ; P1_R1138_U164
g13043 nand P1_R1138_U364 P1_R1138_U363 ; P1_R1138_U165
g13044 nand P1_U3052 P1_R1138_U147 ; P1_R1138_U166
g13045 not P1_R1138_U35 ; P1_R1138_U167
g13046 nand P1_U3480 P1_U3081 ; P1_R1138_U168
g13047 nand P1_U3070 P1_U3489 ; P1_R1138_U169
g13048 nand P1_U3056 P1_U4010 ; P1_R1138_U170
g13049 not P1_R1138_U69 ; P1_R1138_U171
g13050 not P1_R1138_U78 ; P1_R1138_U172
g13051 nand P1_U3063 P1_U4011 ; P1_R1138_U173
g13052 not P1_R1138_U62 ; P1_R1138_U174
g13053 or P1_U3065 P1_U3468 ; P1_R1138_U175
g13054 or P1_U3058 P1_U3465 ; P1_R1138_U176
g13055 or P1_U3462 P1_U3062 ; P1_R1138_U177
g13056 or P1_U3459 P1_U3066 ; P1_R1138_U178
g13057 not P1_R1138_U32 ; P1_R1138_U179
g13058 or P1_U3456 P1_U3076 ; P1_R1138_U180
g13059 not P1_R1138_U43 ; P1_R1138_U181
g13060 not P1_R1138_U44 ; P1_R1138_U182
g13061 nand P1_R1138_U43 P1_R1138_U44 ; P1_R1138_U183
g13062 nand P1_R1138_U116 P1_R1138_U177 ; P1_R1138_U184
g13063 nand P1_R1138_U5 P1_R1138_U183 ; P1_R1138_U185
g13064 nand P1_U3062 P1_U3462 ; P1_R1138_U186
g13065 nand P1_R1138_U117 P1_R1138_U185 ; P1_R1138_U187
g13066 nand P1_R1138_U36 P1_R1138_U35 ; P1_R1138_U188
g13067 nand P1_U3065 P1_R1138_U188 ; P1_R1138_U189
g13068 nand P1_R1138_U4 P1_R1138_U187 ; P1_R1138_U190
g13069 nand P1_U3468 P1_R1138_U167 ; P1_R1138_U191
g13070 not P1_R1138_U42 ; P1_R1138_U192
g13071 or P1_U3068 P1_U3474 ; P1_R1138_U193
g13072 or P1_U3069 P1_U3471 ; P1_R1138_U194
g13073 not P1_R1138_U23 ; P1_R1138_U195
g13074 nand P1_R1138_U24 P1_R1138_U23 ; P1_R1138_U196
g13075 nand P1_U3068 P1_R1138_U196 ; P1_R1138_U197
g13076 nand P1_U3474 P1_R1138_U195 ; P1_R1138_U198
g13077 nand P1_R1138_U6 P1_R1138_U42 ; P1_R1138_U199
g13078 not P1_R1138_U140 ; P1_R1138_U200
g13079 or P1_U3477 P1_U3082 ; P1_R1138_U201
g13080 nand P1_R1138_U201 P1_R1138_U140 ; P1_R1138_U202
g13081 not P1_R1138_U41 ; P1_R1138_U203
g13082 or P1_U3081 P1_U3480 ; P1_R1138_U204
g13083 or P1_U3471 P1_U3069 ; P1_R1138_U205
g13084 nand P1_R1138_U205 P1_R1138_U42 ; P1_R1138_U206
g13085 nand P1_R1138_U120 P1_R1138_U206 ; P1_R1138_U207
g13086 nand P1_R1138_U192 P1_R1138_U23 ; P1_R1138_U208
g13087 nand P1_U3474 P1_U3068 ; P1_R1138_U209
g13088 nand P1_R1138_U121 P1_R1138_U208 ; P1_R1138_U210
g13089 or P1_U3069 P1_U3471 ; P1_R1138_U211
g13090 nand P1_R1138_U182 P1_R1138_U178 ; P1_R1138_U212
g13091 nand P1_U3066 P1_U3459 ; P1_R1138_U213
g13092 not P1_R1138_U46 ; P1_R1138_U214
g13093 nand P1_R1138_U181 P1_R1138_U5 ; P1_R1138_U215
g13094 nand P1_R1138_U46 P1_R1138_U177 ; P1_R1138_U216
g13095 nand P1_U3062 P1_U3462 ; P1_R1138_U217
g13096 not P1_R1138_U45 ; P1_R1138_U218
g13097 or P1_U3465 P1_U3058 ; P1_R1138_U219
g13098 nand P1_R1138_U219 P1_R1138_U45 ; P1_R1138_U220
g13099 nand P1_R1138_U123 P1_R1138_U220 ; P1_R1138_U221
g13100 nand P1_R1138_U218 P1_R1138_U35 ; P1_R1138_U222
g13101 nand P1_U3468 P1_U3065 ; P1_R1138_U223
g13102 nand P1_R1138_U124 P1_R1138_U222 ; P1_R1138_U224
g13103 or P1_U3058 P1_U3465 ; P1_R1138_U225
g13104 nand P1_R1138_U181 P1_R1138_U178 ; P1_R1138_U226
g13105 not P1_R1138_U141 ; P1_R1138_U227
g13106 nand P1_U3062 P1_U3462 ; P1_R1138_U228
g13107 nand P1_R1138_U398 P1_R1138_U397 P1_R1138_U44 P1_R1138_U43 ; P1_R1138_U229
g13108 nand P1_R1138_U44 P1_R1138_U43 ; P1_R1138_U230
g13109 nand P1_U3066 P1_U3459 ; P1_R1138_U231
g13110 nand P1_R1138_U125 P1_R1138_U230 ; P1_R1138_U232
g13111 or P1_U3081 P1_U3480 ; P1_R1138_U233
g13112 or P1_U3060 P1_U3483 ; P1_R1138_U234
g13113 nand P1_R1138_U174 P1_R1138_U7 ; P1_R1138_U235
g13114 nand P1_U3060 P1_U3483 ; P1_R1138_U236
g13115 nand P1_R1138_U127 P1_R1138_U235 ; P1_R1138_U237
g13116 or P1_U3483 P1_U3060 ; P1_R1138_U238
g13117 nand P1_R1138_U126 P1_R1138_U140 ; P1_R1138_U239
g13118 nand P1_R1138_U238 P1_R1138_U237 ; P1_R1138_U240
g13119 not P1_R1138_U164 ; P1_R1138_U241
g13120 or P1_U3078 P1_U3492 ; P1_R1138_U242
g13121 or P1_U3070 P1_U3489 ; P1_R1138_U243
g13122 nand P1_R1138_U171 P1_R1138_U8 ; P1_R1138_U244
g13123 nand P1_U3078 P1_U3492 ; P1_R1138_U245
g13124 nand P1_R1138_U128 P1_R1138_U244 ; P1_R1138_U246
g13125 or P1_U3486 P1_U3061 ; P1_R1138_U247
g13126 or P1_U3492 P1_U3078 ; P1_R1138_U248
g13127 nand P1_R1138_U247 P1_R1138_U164 P1_R1138_U8 ; P1_R1138_U249
g13128 nand P1_R1138_U248 P1_R1138_U246 ; P1_R1138_U250
g13129 not P1_R1138_U163 ; P1_R1138_U251
g13130 or P1_U3495 P1_U3077 ; P1_R1138_U252
g13131 nand P1_R1138_U252 P1_R1138_U163 ; P1_R1138_U253
g13132 nand P1_U3077 P1_U3495 ; P1_R1138_U254
g13133 not P1_R1138_U161 ; P1_R1138_U255
g13134 or P1_U3498 P1_U3072 ; P1_R1138_U256
g13135 nand P1_R1138_U256 P1_R1138_U161 ; P1_R1138_U257
g13136 nand P1_U3072 P1_U3498 ; P1_R1138_U258
g13137 not P1_R1138_U93 ; P1_R1138_U259
g13138 or P1_U3067 P1_U3504 ; P1_R1138_U260
g13139 or P1_U3071 P1_U3501 ; P1_R1138_U261
g13140 not P1_R1138_U60 ; P1_R1138_U262
g13141 nand P1_R1138_U61 P1_R1138_U60 ; P1_R1138_U263
g13142 nand P1_U3067 P1_R1138_U263 ; P1_R1138_U264
g13143 nand P1_U3504 P1_R1138_U262 ; P1_R1138_U265
g13144 nand P1_R1138_U9 P1_R1138_U93 ; P1_R1138_U266
g13145 not P1_R1138_U159 ; P1_R1138_U267
g13146 or P1_U3074 P1_U4015 ; P1_R1138_U268
g13147 or P1_U3079 P1_U3509 ; P1_R1138_U269
g13148 or P1_U3073 P1_U4014 ; P1_R1138_U270
g13149 not P1_R1138_U81 ; P1_R1138_U271
g13150 nand P1_U4015 P1_R1138_U271 ; P1_R1138_U272
g13151 nand P1_R1138_U272 P1_R1138_U91 ; P1_R1138_U273
g13152 nand P1_R1138_U81 P1_R1138_U82 ; P1_R1138_U274
g13153 nand P1_R1138_U274 P1_R1138_U273 ; P1_R1138_U275
g13154 nand P1_R1138_U172 P1_R1138_U10 ; P1_R1138_U276
g13155 nand P1_U3073 P1_U4014 ; P1_R1138_U277
g13156 nand P1_R1138_U275 P1_R1138_U276 ; P1_R1138_U278
g13157 or P1_U3507 P1_U3080 ; P1_R1138_U279
g13158 or P1_U4014 P1_U3073 ; P1_R1138_U280
g13159 nand P1_R1138_U270 P1_R1138_U159 P1_R1138_U130 ; P1_R1138_U281
g13160 nand P1_R1138_U280 P1_R1138_U278 ; P1_R1138_U282
g13161 not P1_R1138_U155 ; P1_R1138_U283
g13162 or P1_U4013 P1_U3059 ; P1_R1138_U284
g13163 nand P1_R1138_U284 P1_R1138_U155 ; P1_R1138_U285
g13164 nand P1_U3059 P1_U4013 ; P1_R1138_U286
g13165 not P1_R1138_U153 ; P1_R1138_U287
g13166 or P1_U4012 P1_U3064 ; P1_R1138_U288
g13167 nand P1_R1138_U288 P1_R1138_U153 ; P1_R1138_U289
g13168 nand P1_U3064 P1_U4012 ; P1_R1138_U290
g13169 not P1_R1138_U151 ; P1_R1138_U291
g13170 or P1_U3056 P1_U4010 ; P1_R1138_U292
g13171 nand P1_R1138_U173 P1_R1138_U170 ; P1_R1138_U293
g13172 not P1_R1138_U87 ; P1_R1138_U294
g13173 or P1_U4011 P1_U3063 ; P1_R1138_U295
g13174 nand P1_R1138_U151 P1_R1138_U295 P1_R1138_U165 ; P1_R1138_U296
g13175 not P1_R1138_U149 ; P1_R1138_U297
g13176 or P1_U4008 P1_U3051 ; P1_R1138_U298
g13177 nand P1_U3051 P1_U4008 ; P1_R1138_U299
g13178 not P1_R1138_U147 ; P1_R1138_U300
g13179 nand P1_U4007 P1_R1138_U147 ; P1_R1138_U301
g13180 not P1_R1138_U145 ; P1_R1138_U302
g13181 nand P1_R1138_U295 P1_R1138_U151 ; P1_R1138_U303
g13182 not P1_R1138_U90 ; P1_R1138_U304
g13183 or P1_U4010 P1_U3056 ; P1_R1138_U305
g13184 nand P1_R1138_U305 P1_R1138_U90 ; P1_R1138_U306
g13185 nand P1_R1138_U306 P1_R1138_U170 P1_R1138_U150 ; P1_R1138_U307
g13186 nand P1_R1138_U304 P1_R1138_U170 ; P1_R1138_U308
g13187 nand P1_U4009 P1_U3055 ; P1_R1138_U309
g13188 nand P1_R1138_U308 P1_R1138_U309 P1_R1138_U165 ; P1_R1138_U310
g13189 or P1_U3056 P1_U4010 ; P1_R1138_U311
g13190 nand P1_R1138_U279 P1_R1138_U159 ; P1_R1138_U312
g13191 not P1_R1138_U92 ; P1_R1138_U313
g13192 nand P1_R1138_U10 P1_R1138_U92 ; P1_R1138_U314
g13193 nand P1_R1138_U134 P1_R1138_U314 ; P1_R1138_U315
g13194 nand P1_R1138_U314 P1_R1138_U275 ; P1_R1138_U316
g13195 nand P1_R1138_U450 P1_R1138_U316 ; P1_R1138_U317
g13196 or P1_U3509 P1_U3079 ; P1_R1138_U318
g13197 nand P1_R1138_U318 P1_R1138_U92 ; P1_R1138_U319
g13198 nand P1_R1138_U319 P1_R1138_U81 P1_R1138_U157 ; P1_R1138_U320
g13199 nand P1_R1138_U313 P1_R1138_U81 ; P1_R1138_U321
g13200 nand P1_U3074 P1_U4015 ; P1_R1138_U322
g13201 nand P1_R1138_U322 P1_R1138_U321 P1_R1138_U10 ; P1_R1138_U323
g13202 or P1_U3456 P1_U3076 ; P1_R1138_U324
g13203 not P1_R1138_U158 ; P1_R1138_U325
g13204 or P1_U3079 P1_U3509 ; P1_R1138_U326
g13205 or P1_U3501 P1_U3071 ; P1_R1138_U327
g13206 nand P1_R1138_U327 P1_R1138_U93 ; P1_R1138_U328
g13207 nand P1_R1138_U135 P1_R1138_U328 ; P1_R1138_U329
g13208 nand P1_R1138_U259 P1_R1138_U60 ; P1_R1138_U330
g13209 nand P1_U3504 P1_U3067 ; P1_R1138_U331
g13210 nand P1_R1138_U331 P1_R1138_U330 P1_R1138_U9 ; P1_R1138_U332
g13211 or P1_U3071 P1_U3501 ; P1_R1138_U333
g13212 nand P1_R1138_U247 P1_R1138_U164 ; P1_R1138_U334
g13213 not P1_R1138_U94 ; P1_R1138_U335
g13214 or P1_U3489 P1_U3070 ; P1_R1138_U336
g13215 nand P1_R1138_U336 P1_R1138_U94 ; P1_R1138_U337
g13216 nand P1_R1138_U136 P1_R1138_U337 ; P1_R1138_U338
g13217 nand P1_R1138_U335 P1_R1138_U169 ; P1_R1138_U339
g13218 nand P1_U3078 P1_U3492 ; P1_R1138_U340
g13219 nand P1_R1138_U137 P1_R1138_U339 ; P1_R1138_U341
g13220 or P1_U3070 P1_U3489 ; P1_R1138_U342
g13221 or P1_U3480 P1_U3081 ; P1_R1138_U343
g13222 nand P1_R1138_U343 P1_R1138_U41 ; P1_R1138_U344
g13223 nand P1_R1138_U138 P1_R1138_U344 ; P1_R1138_U345
g13224 nand P1_R1138_U203 P1_R1138_U168 ; P1_R1138_U346
g13225 nand P1_U3060 P1_U3483 ; P1_R1138_U347
g13226 nand P1_R1138_U139 P1_R1138_U346 ; P1_R1138_U348
g13227 nand P1_R1138_U204 P1_R1138_U168 ; P1_R1138_U349
g13228 nand P1_R1138_U201 P1_R1138_U62 ; P1_R1138_U350
g13229 nand P1_R1138_U211 P1_R1138_U23 ; P1_R1138_U351
g13230 nand P1_R1138_U225 P1_R1138_U35 ; P1_R1138_U352
g13231 nand P1_R1138_U228 P1_R1138_U177 ; P1_R1138_U353
g13232 nand P1_R1138_U311 P1_R1138_U170 ; P1_R1138_U354
g13233 nand P1_R1138_U295 P1_R1138_U173 ; P1_R1138_U355
g13234 nand P1_R1138_U326 P1_R1138_U81 ; P1_R1138_U356
g13235 nand P1_R1138_U279 P1_R1138_U78 ; P1_R1138_U357
g13236 nand P1_R1138_U333 P1_R1138_U60 ; P1_R1138_U358
g13237 nand P1_R1138_U342 P1_R1138_U169 ; P1_R1138_U359
g13238 nand P1_R1138_U247 P1_R1138_U69 ; P1_R1138_U360
g13239 nand P1_U4007 P1_U3052 ; P1_R1138_U361
g13240 nand P1_R1138_U293 P1_R1138_U165 ; P1_R1138_U362
g13241 nand P1_U3055 P1_R1138_U292 ; P1_R1138_U363
g13242 nand P1_U4009 P1_R1138_U292 ; P1_R1138_U364
g13243 nand P1_R1138_U293 P1_R1138_U165 P1_R1138_U298 ; P1_R1138_U365
g13244 nand P1_R1138_U151 P1_R1138_U165 P1_R1138_U132 ; P1_R1138_U366
g13245 nand P1_R1138_U294 P1_R1138_U298 ; P1_R1138_U367
g13246 nand P1_U3081 P1_R1138_U40 ; P1_R1138_U368
g13247 nand P1_U3480 P1_R1138_U39 ; P1_R1138_U369
g13248 nand P1_R1138_U369 P1_R1138_U368 ; P1_R1138_U370
g13249 nand P1_R1138_U349 P1_R1138_U41 ; P1_R1138_U371
g13250 nand P1_R1138_U370 P1_R1138_U203 ; P1_R1138_U372
g13251 nand P1_U3082 P1_R1138_U37 ; P1_R1138_U373
g13252 nand P1_U3477 P1_R1138_U38 ; P1_R1138_U374
g13253 nand P1_R1138_U374 P1_R1138_U373 ; P1_R1138_U375
g13254 nand P1_R1138_U350 P1_R1138_U140 ; P1_R1138_U376
g13255 nand P1_R1138_U200 P1_R1138_U375 ; P1_R1138_U377
g13256 nand P1_U3068 P1_R1138_U24 ; P1_R1138_U378
g13257 nand P1_U3474 P1_R1138_U22 ; P1_R1138_U379
g13258 nand P1_U3069 P1_R1138_U20 ; P1_R1138_U380
g13259 nand P1_U3471 P1_R1138_U21 ; P1_R1138_U381
g13260 nand P1_R1138_U381 P1_R1138_U380 ; P1_R1138_U382
g13261 nand P1_R1138_U351 P1_R1138_U42 ; P1_R1138_U383
g13262 nand P1_R1138_U382 P1_R1138_U192 ; P1_R1138_U384
g13263 nand P1_U3065 P1_R1138_U36 ; P1_R1138_U385
g13264 nand P1_U3468 P1_R1138_U27 ; P1_R1138_U386
g13265 nand P1_U3058 P1_R1138_U25 ; P1_R1138_U387
g13266 nand P1_U3465 P1_R1138_U26 ; P1_R1138_U388
g13267 nand P1_R1138_U388 P1_R1138_U387 ; P1_R1138_U389
g13268 nand P1_R1138_U352 P1_R1138_U45 ; P1_R1138_U390
g13269 nand P1_R1138_U389 P1_R1138_U218 ; P1_R1138_U391
g13270 nand P1_U3062 P1_R1138_U33 ; P1_R1138_U392
g13271 nand P1_U3462 P1_R1138_U34 ; P1_R1138_U393
g13272 nand P1_R1138_U393 P1_R1138_U392 ; P1_R1138_U394
g13273 nand P1_R1138_U353 P1_R1138_U141 ; P1_R1138_U395
g13274 nand P1_R1138_U227 P1_R1138_U394 ; P1_R1138_U396
g13275 nand P1_U3066 P1_R1138_U28 ; P1_R1138_U397
g13276 nand P1_U3459 P1_R1138_U29 ; P1_R1138_U398
g13277 nand P1_U3053 P1_R1138_U143 ; P1_R1138_U399
g13278 nand P1_U4018 P1_R1138_U142 ; P1_R1138_U400
g13279 nand P1_U3053 P1_R1138_U143 ; P1_R1138_U401
g13280 nand P1_U4018 P1_R1138_U142 ; P1_R1138_U402
g13281 nand P1_R1138_U402 P1_R1138_U401 ; P1_R1138_U403
g13282 nand P1_R1138_U144 P1_R1138_U145 ; P1_R1138_U404
g13283 nand P1_R1138_U302 P1_R1138_U403 ; P1_R1138_U405
g13284 nand P1_U3052 P1_R1138_U89 ; P1_R1138_U406
g13285 nand P1_U4007 P1_R1138_U88 ; P1_R1138_U407
g13286 nand P1_U3052 P1_R1138_U89 ; P1_R1138_U408
g13287 nand P1_U4007 P1_R1138_U88 ; P1_R1138_U409
g13288 nand P1_R1138_U409 P1_R1138_U408 ; P1_R1138_U410
g13289 nand P1_R1138_U146 P1_R1138_U147 ; P1_R1138_U411
g13290 nand P1_R1138_U300 P1_R1138_U410 ; P1_R1138_U412
g13291 nand P1_U3051 P1_R1138_U47 ; P1_R1138_U413
g13292 nand P1_U4008 P1_R1138_U48 ; P1_R1138_U414
g13293 nand P1_U3051 P1_R1138_U47 ; P1_R1138_U415
g13294 nand P1_U4008 P1_R1138_U48 ; P1_R1138_U416
g13295 nand P1_R1138_U416 P1_R1138_U415 ; P1_R1138_U417
g13296 nand P1_R1138_U148 P1_R1138_U149 ; P1_R1138_U418
g13297 nand P1_R1138_U297 P1_R1138_U417 ; P1_R1138_U419
g13298 nand P1_U3055 P1_R1138_U50 ; P1_R1138_U420
g13299 nand P1_U4009 P1_R1138_U49 ; P1_R1138_U421
g13300 nand P1_U3056 P1_R1138_U51 ; P1_R1138_U422
g13301 nand P1_U4010 P1_R1138_U52 ; P1_R1138_U423
g13302 nand P1_R1138_U423 P1_R1138_U422 ; P1_R1138_U424
g13303 nand P1_R1138_U354 P1_R1138_U90 ; P1_R1138_U425
g13304 nand P1_R1138_U424 P1_R1138_U304 ; P1_R1138_U426
g13305 nand P1_U3063 P1_R1138_U53 ; P1_R1138_U427
g13306 nand P1_U4011 P1_R1138_U54 ; P1_R1138_U428
g13307 nand P1_R1138_U428 P1_R1138_U427 ; P1_R1138_U429
g13308 nand P1_R1138_U355 P1_R1138_U151 ; P1_R1138_U430
g13309 nand P1_R1138_U291 P1_R1138_U429 ; P1_R1138_U431
g13310 nand P1_U3064 P1_R1138_U85 ; P1_R1138_U432
g13311 nand P1_U4012 P1_R1138_U86 ; P1_R1138_U433
g13312 nand P1_U3064 P1_R1138_U85 ; P1_R1138_U434
g13313 nand P1_U4012 P1_R1138_U86 ; P1_R1138_U435
g13314 nand P1_R1138_U435 P1_R1138_U434 ; P1_R1138_U436
g13315 nand P1_R1138_U152 P1_R1138_U153 ; P1_R1138_U437
g13316 nand P1_R1138_U287 P1_R1138_U436 ; P1_R1138_U438
g13317 nand P1_U3059 P1_R1138_U83 ; P1_R1138_U439
g13318 nand P1_U4013 P1_R1138_U84 ; P1_R1138_U440
g13319 nand P1_U3059 P1_R1138_U83 ; P1_R1138_U441
g13320 nand P1_U4013 P1_R1138_U84 ; P1_R1138_U442
g13321 nand P1_R1138_U442 P1_R1138_U441 ; P1_R1138_U443
g13322 nand P1_R1138_U154 P1_R1138_U155 ; P1_R1138_U444
g13323 nand P1_R1138_U283 P1_R1138_U443 ; P1_R1138_U445
g13324 nand P1_U3073 P1_R1138_U55 ; P1_R1138_U446
g13325 nand P1_U4014 P1_R1138_U56 ; P1_R1138_U447
g13326 nand P1_U3073 P1_R1138_U55 ; P1_R1138_U448
g13327 nand P1_U4014 P1_R1138_U56 ; P1_R1138_U449
g13328 nand P1_R1138_U449 P1_R1138_U448 ; P1_R1138_U450
g13329 nand P1_U3074 P1_R1138_U82 ; P1_R1138_U451
g13330 nand P1_U4015 P1_R1138_U91 ; P1_R1138_U452
g13331 nand P1_R1138_U179 P1_R1138_U158 ; P1_R1138_U453
g13332 nand P1_R1138_U325 P1_R1138_U32 ; P1_R1138_U454
g13333 nand P1_U3079 P1_R1138_U79 ; P1_R1138_U455
g13334 nand P1_U3509 P1_R1138_U80 ; P1_R1138_U456
g13335 nand P1_R1138_U456 P1_R1138_U455 ; P1_R1138_U457
g13336 nand P1_R1138_U356 P1_R1138_U92 ; P1_R1138_U458
g13337 nand P1_R1138_U457 P1_R1138_U313 ; P1_R1138_U459
g13338 nand P1_U3080 P1_R1138_U76 ; P1_R1138_U460
g13339 nand P1_U3507 P1_R1138_U77 ; P1_R1138_U461
g13340 nand P1_R1138_U461 P1_R1138_U460 ; P1_R1138_U462
g13341 nand P1_R1138_U357 P1_R1138_U159 ; P1_R1138_U463
g13342 nand P1_R1138_U267 P1_R1138_U462 ; P1_R1138_U464
g13343 nand P1_U3067 P1_R1138_U61 ; P1_R1138_U465
g13344 nand P1_U3504 P1_R1138_U59 ; P1_R1138_U466
g13345 nand P1_U3071 P1_R1138_U57 ; P1_R1138_U467
g13346 nand P1_U3501 P1_R1138_U58 ; P1_R1138_U468
g13347 nand P1_R1138_U468 P1_R1138_U467 ; P1_R1138_U469
g13348 nand P1_R1138_U358 P1_R1138_U93 ; P1_R1138_U470
g13349 nand P1_R1138_U469 P1_R1138_U259 ; P1_R1138_U471
g13350 nand P1_U3072 P1_R1138_U74 ; P1_R1138_U472
g13351 nand P1_U3498 P1_R1138_U75 ; P1_R1138_U473
g13352 nand P1_U3072 P1_R1138_U74 ; P1_R1138_U474
g13353 nand P1_U3498 P1_R1138_U75 ; P1_R1138_U475
g13354 nand P1_R1138_U475 P1_R1138_U474 ; P1_R1138_U476
g13355 nand P1_R1138_U160 P1_R1138_U161 ; P1_R1138_U477
g13356 nand P1_R1138_U255 P1_R1138_U476 ; P1_R1138_U478
g13357 nand P1_U3077 P1_R1138_U72 ; P1_R1138_U479
g13358 nand P1_U3495 P1_R1138_U73 ; P1_R1138_U480
g13359 nand P1_U3077 P1_R1138_U72 ; P1_R1138_U481
g13360 nand P1_U3495 P1_R1138_U73 ; P1_R1138_U482
g13361 nand P1_R1138_U482 P1_R1138_U481 ; P1_R1138_U483
g13362 nand P1_R1138_U162 P1_R1138_U163 ; P1_R1138_U484
g13363 nand P1_R1138_U251 P1_R1138_U483 ; P1_R1138_U485
g13364 nand P1_U3078 P1_R1138_U70 ; P1_R1138_U486
g13365 nand P1_U3492 P1_R1138_U71 ; P1_R1138_U487
g13366 nand P1_U3070 P1_R1138_U65 ; P1_R1138_U488
g13367 nand P1_U3489 P1_R1138_U66 ; P1_R1138_U489
g13368 nand P1_R1138_U489 P1_R1138_U488 ; P1_R1138_U490
g13369 nand P1_R1138_U359 P1_R1138_U94 ; P1_R1138_U491
g13370 nand P1_R1138_U490 P1_R1138_U335 ; P1_R1138_U492
g13371 nand P1_U3061 P1_R1138_U67 ; P1_R1138_U493
g13372 nand P1_U3486 P1_R1138_U68 ; P1_R1138_U494
g13373 nand P1_R1138_U494 P1_R1138_U493 ; P1_R1138_U495
g13374 nand P1_R1138_U360 P1_R1138_U164 ; P1_R1138_U496
g13375 nand P1_R1138_U241 P1_R1138_U495 ; P1_R1138_U497
g13376 nand P1_U3060 P1_R1138_U63 ; P1_R1138_U498
g13377 nand P1_U3483 P1_R1138_U64 ; P1_R1138_U499
g13378 nand P1_U3075 P1_R1138_U30 ; P1_R1138_U500
g13379 nand P1_U3451 P1_R1138_U31 ; P1_R1138_U501
g13380 and P1_R1222_U176 P1_R1222_U175 ; P1_R1222_U4
g13381 and P1_R1222_U177 P1_R1222_U178 ; P1_R1222_U5
g13382 and P1_R1222_U194 P1_R1222_U193 ; P1_R1222_U6
g13383 and P1_R1222_U234 P1_R1222_U233 ; P1_R1222_U7
g13384 and P1_R1222_U243 P1_R1222_U242 ; P1_R1222_U8
g13385 and P1_R1222_U261 P1_R1222_U260 ; P1_R1222_U9
g13386 and P1_R1222_U269 P1_R1222_U268 ; P1_R1222_U10
g13387 and P1_R1222_U348 P1_R1222_U345 ; P1_R1222_U11
g13388 and P1_R1222_U341 P1_R1222_U338 ; P1_R1222_U12
g13389 and P1_R1222_U332 P1_R1222_U329 ; P1_R1222_U13
g13390 and P1_R1222_U323 P1_R1222_U320 ; P1_R1222_U14
g13391 and P1_R1222_U317 P1_R1222_U315 ; P1_R1222_U15
g13392 and P1_R1222_U310 P1_R1222_U307 ; P1_R1222_U16
g13393 and P1_R1222_U232 P1_R1222_U229 ; P1_R1222_U17
g13394 and P1_R1222_U224 P1_R1222_U221 ; P1_R1222_U18
g13395 and P1_R1222_U210 P1_R1222_U207 ; P1_R1222_U19
g13396 not P1_U3471 ; P1_R1222_U20
g13397 not P1_U3069 ; P1_R1222_U21
g13398 not P1_U3068 ; P1_R1222_U22
g13399 nand P1_U3069 P1_U3471 ; P1_R1222_U23
g13400 not P1_U3474 ; P1_R1222_U24
g13401 not P1_U3465 ; P1_R1222_U25
g13402 not P1_U3058 ; P1_R1222_U26
g13403 not P1_U3065 ; P1_R1222_U27
g13404 not P1_U3459 ; P1_R1222_U28
g13405 not P1_U3066 ; P1_R1222_U29
g13406 not P1_U3451 ; P1_R1222_U30
g13407 not P1_U3075 ; P1_R1222_U31
g13408 nand P1_U3075 P1_U3451 ; P1_R1222_U32
g13409 not P1_U3462 ; P1_R1222_U33
g13410 not P1_U3062 ; P1_R1222_U34
g13411 nand P1_U3058 P1_U3465 ; P1_R1222_U35
g13412 not P1_U3468 ; P1_R1222_U36
g13413 not P1_U3477 ; P1_R1222_U37
g13414 not P1_U3082 ; P1_R1222_U38
g13415 not P1_U3081 ; P1_R1222_U39
g13416 not P1_U3480 ; P1_R1222_U40
g13417 nand P1_R1222_U62 P1_R1222_U202 ; P1_R1222_U41
g13418 nand P1_R1222_U118 P1_R1222_U190 ; P1_R1222_U42
g13419 nand P1_R1222_U179 P1_R1222_U180 ; P1_R1222_U43
g13420 nand P1_U3456 P1_U3076 ; P1_R1222_U44
g13421 nand P1_R1222_U122 P1_R1222_U216 ; P1_R1222_U45
g13422 nand P1_R1222_U213 P1_R1222_U212 ; P1_R1222_U46
g13423 not P1_U4008 ; P1_R1222_U47
g13424 not P1_U3051 ; P1_R1222_U48
g13425 not P1_U3055 ; P1_R1222_U49
g13426 not P1_U4009 ; P1_R1222_U50
g13427 not P1_U4010 ; P1_R1222_U51
g13428 not P1_U3056 ; P1_R1222_U52
g13429 not P1_U4011 ; P1_R1222_U53
g13430 not P1_U3063 ; P1_R1222_U54
g13431 not P1_U4014 ; P1_R1222_U55
g13432 not P1_U3073 ; P1_R1222_U56
g13433 not P1_U3501 ; P1_R1222_U57
g13434 not P1_U3071 ; P1_R1222_U58
g13435 not P1_U3067 ; P1_R1222_U59
g13436 nand P1_U3071 P1_U3501 ; P1_R1222_U60
g13437 not P1_U3504 ; P1_R1222_U61
g13438 nand P1_U3082 P1_U3477 ; P1_R1222_U62
g13439 not P1_U3483 ; P1_R1222_U63
g13440 not P1_U3060 ; P1_R1222_U64
g13441 not P1_U3489 ; P1_R1222_U65
g13442 not P1_U3070 ; P1_R1222_U66
g13443 not P1_U3486 ; P1_R1222_U67
g13444 not P1_U3061 ; P1_R1222_U68
g13445 nand P1_U3061 P1_U3486 ; P1_R1222_U69
g13446 not P1_U3492 ; P1_R1222_U70
g13447 not P1_U3078 ; P1_R1222_U71
g13448 not P1_U3495 ; P1_R1222_U72
g13449 not P1_U3077 ; P1_R1222_U73
g13450 not P1_U3498 ; P1_R1222_U74
g13451 not P1_U3072 ; P1_R1222_U75
g13452 not P1_U3507 ; P1_R1222_U76
g13453 not P1_U3080 ; P1_R1222_U77
g13454 nand P1_U3080 P1_U3507 ; P1_R1222_U78
g13455 not P1_U3509 ; P1_R1222_U79
g13456 not P1_U3079 ; P1_R1222_U80
g13457 nand P1_U3079 P1_U3509 ; P1_R1222_U81
g13458 not P1_U4015 ; P1_R1222_U82
g13459 not P1_U4013 ; P1_R1222_U83
g13460 not P1_U3059 ; P1_R1222_U84
g13461 not P1_U4012 ; P1_R1222_U85
g13462 not P1_U3064 ; P1_R1222_U86
g13463 nand P1_U4009 P1_U3055 ; P1_R1222_U87
g13464 not P1_U3052 ; P1_R1222_U88
g13465 not P1_U4007 ; P1_R1222_U89
g13466 nand P1_R1222_U303 P1_R1222_U173 ; P1_R1222_U90
g13467 not P1_U3074 ; P1_R1222_U91
g13468 nand P1_R1222_U78 P1_R1222_U312 ; P1_R1222_U92
g13469 nand P1_R1222_U258 P1_R1222_U257 ; P1_R1222_U93
g13470 nand P1_R1222_U69 P1_R1222_U334 ; P1_R1222_U94
g13471 nand P1_R1222_U454 P1_R1222_U453 ; P1_R1222_U95
g13472 nand P1_R1222_U501 P1_R1222_U500 ; P1_R1222_U96
g13473 nand P1_R1222_U372 P1_R1222_U371 ; P1_R1222_U97
g13474 nand P1_R1222_U377 P1_R1222_U376 ; P1_R1222_U98
g13475 nand P1_R1222_U384 P1_R1222_U383 ; P1_R1222_U99
g13476 nand P1_R1222_U391 P1_R1222_U390 ; P1_R1222_U100
g13477 nand P1_R1222_U396 P1_R1222_U395 ; P1_R1222_U101
g13478 nand P1_R1222_U405 P1_R1222_U404 ; P1_R1222_U102
g13479 nand P1_R1222_U412 P1_R1222_U411 ; P1_R1222_U103
g13480 nand P1_R1222_U419 P1_R1222_U418 ; P1_R1222_U104
g13481 nand P1_R1222_U426 P1_R1222_U425 ; P1_R1222_U105
g13482 nand P1_R1222_U431 P1_R1222_U430 ; P1_R1222_U106
g13483 nand P1_R1222_U438 P1_R1222_U437 ; P1_R1222_U107
g13484 nand P1_R1222_U445 P1_R1222_U444 ; P1_R1222_U108
g13485 nand P1_R1222_U459 P1_R1222_U458 ; P1_R1222_U109
g13486 nand P1_R1222_U464 P1_R1222_U463 ; P1_R1222_U110
g13487 nand P1_R1222_U471 P1_R1222_U470 ; P1_R1222_U111
g13488 nand P1_R1222_U478 P1_R1222_U477 ; P1_R1222_U112
g13489 nand P1_R1222_U485 P1_R1222_U484 ; P1_R1222_U113
g13490 nand P1_R1222_U492 P1_R1222_U491 ; P1_R1222_U114
g13491 nand P1_R1222_U497 P1_R1222_U496 ; P1_R1222_U115
g13492 and P1_U3459 P1_U3066 ; P1_R1222_U116
g13493 and P1_R1222_U186 P1_R1222_U184 ; P1_R1222_U117
g13494 and P1_R1222_U191 P1_R1222_U189 ; P1_R1222_U118
g13495 and P1_R1222_U198 P1_R1222_U197 ; P1_R1222_U119
g13496 and P1_R1222_U379 P1_R1222_U378 P1_R1222_U23 ; P1_R1222_U120
g13497 and P1_R1222_U209 P1_R1222_U6 ; P1_R1222_U121
g13498 and P1_R1222_U217 P1_R1222_U215 ; P1_R1222_U122
g13499 and P1_R1222_U386 P1_R1222_U385 P1_R1222_U35 ; P1_R1222_U123
g13500 and P1_R1222_U223 P1_R1222_U4 ; P1_R1222_U124
g13501 and P1_R1222_U231 P1_R1222_U178 ; P1_R1222_U125
g13502 and P1_R1222_U201 P1_R1222_U7 ; P1_R1222_U126
g13503 and P1_R1222_U236 P1_R1222_U168 ; P1_R1222_U127
g13504 and P1_R1222_U245 P1_R1222_U169 ; P1_R1222_U128
g13505 and P1_R1222_U265 P1_R1222_U264 ; P1_R1222_U129
g13506 and P1_R1222_U10 P1_R1222_U279 ; P1_R1222_U130
g13507 and P1_R1222_U282 P1_R1222_U277 ; P1_R1222_U131
g13508 and P1_R1222_U298 P1_R1222_U295 ; P1_R1222_U132
g13509 and P1_R1222_U365 P1_R1222_U299 ; P1_R1222_U133
g13510 and P1_R1222_U156 P1_R1222_U275 ; P1_R1222_U134
g13511 and P1_R1222_U466 P1_R1222_U465 P1_R1222_U60 ; P1_R1222_U135
g13512 and P1_R1222_U487 P1_R1222_U486 P1_R1222_U169 ; P1_R1222_U136
g13513 and P1_R1222_U340 P1_R1222_U8 ; P1_R1222_U137
g13514 and P1_R1222_U499 P1_R1222_U498 P1_R1222_U168 ; P1_R1222_U138
g13515 and P1_R1222_U347 P1_R1222_U7 ; P1_R1222_U139
g13516 nand P1_R1222_U119 P1_R1222_U199 ; P1_R1222_U140
g13517 nand P1_R1222_U214 P1_R1222_U226 ; P1_R1222_U141
g13518 not P1_U3053 ; P1_R1222_U142
g13519 not P1_U4018 ; P1_R1222_U143
g13520 and P1_R1222_U400 P1_R1222_U399 ; P1_R1222_U144
g13521 nand P1_R1222_U301 P1_R1222_U166 P1_R1222_U361 ; P1_R1222_U145
g13522 and P1_R1222_U407 P1_R1222_U406 ; P1_R1222_U146
g13523 nand P1_R1222_U367 P1_R1222_U366 P1_R1222_U133 ; P1_R1222_U147
g13524 and P1_R1222_U414 P1_R1222_U413 ; P1_R1222_U148
g13525 nand P1_R1222_U362 P1_R1222_U296 P1_R1222_U87 ; P1_R1222_U149
g13526 and P1_R1222_U421 P1_R1222_U420 ; P1_R1222_U150
g13527 nand P1_R1222_U290 P1_R1222_U289 ; P1_R1222_U151
g13528 and P1_R1222_U433 P1_R1222_U432 ; P1_R1222_U152
g13529 nand P1_R1222_U286 P1_R1222_U285 ; P1_R1222_U153
g13530 and P1_R1222_U440 P1_R1222_U439 ; P1_R1222_U154
g13531 nand P1_R1222_U131 P1_R1222_U281 ; P1_R1222_U155
g13532 and P1_R1222_U447 P1_R1222_U446 ; P1_R1222_U156
g13533 and P1_R1222_U452 P1_R1222_U451 ; P1_R1222_U157
g13534 nand P1_R1222_U44 P1_R1222_U324 ; P1_R1222_U158
g13535 nand P1_R1222_U129 P1_R1222_U266 ; P1_R1222_U159
g13536 and P1_R1222_U473 P1_R1222_U472 ; P1_R1222_U160
g13537 nand P1_R1222_U254 P1_R1222_U253 ; P1_R1222_U161
g13538 and P1_R1222_U480 P1_R1222_U479 ; P1_R1222_U162
g13539 nand P1_R1222_U250 P1_R1222_U249 ; P1_R1222_U163
g13540 nand P1_R1222_U240 P1_R1222_U239 ; P1_R1222_U164
g13541 nand P1_R1222_U364 P1_R1222_U363 ; P1_R1222_U165
g13542 nand P1_U3052 P1_R1222_U147 ; P1_R1222_U166
g13543 not P1_R1222_U35 ; P1_R1222_U167
g13544 nand P1_U3480 P1_U3081 ; P1_R1222_U168
g13545 nand P1_U3070 P1_U3489 ; P1_R1222_U169
g13546 nand P1_U3056 P1_U4010 ; P1_R1222_U170
g13547 not P1_R1222_U69 ; P1_R1222_U171
g13548 not P1_R1222_U78 ; P1_R1222_U172
g13549 nand P1_U3063 P1_U4011 ; P1_R1222_U173
g13550 not P1_R1222_U62 ; P1_R1222_U174
g13551 or P1_U3065 P1_U3468 ; P1_R1222_U175
g13552 or P1_U3058 P1_U3465 ; P1_R1222_U176
g13553 or P1_U3462 P1_U3062 ; P1_R1222_U177
g13554 or P1_U3459 P1_U3066 ; P1_R1222_U178
g13555 not P1_R1222_U32 ; P1_R1222_U179
g13556 or P1_U3456 P1_U3076 ; P1_R1222_U180
g13557 not P1_R1222_U43 ; P1_R1222_U181
g13558 not P1_R1222_U44 ; P1_R1222_U182
g13559 nand P1_R1222_U43 P1_R1222_U44 ; P1_R1222_U183
g13560 nand P1_R1222_U116 P1_R1222_U177 ; P1_R1222_U184
g13561 nand P1_R1222_U5 P1_R1222_U183 ; P1_R1222_U185
g13562 nand P1_U3062 P1_U3462 ; P1_R1222_U186
g13563 nand P1_R1222_U117 P1_R1222_U185 ; P1_R1222_U187
g13564 nand P1_R1222_U36 P1_R1222_U35 ; P1_R1222_U188
g13565 nand P1_U3065 P1_R1222_U188 ; P1_R1222_U189
g13566 nand P1_R1222_U4 P1_R1222_U187 ; P1_R1222_U190
g13567 nand P1_U3468 P1_R1222_U167 ; P1_R1222_U191
g13568 not P1_R1222_U42 ; P1_R1222_U192
g13569 or P1_U3068 P1_U3474 ; P1_R1222_U193
g13570 or P1_U3069 P1_U3471 ; P1_R1222_U194
g13571 not P1_R1222_U23 ; P1_R1222_U195
g13572 nand P1_R1222_U24 P1_R1222_U23 ; P1_R1222_U196
g13573 nand P1_U3068 P1_R1222_U196 ; P1_R1222_U197
g13574 nand P1_U3474 P1_R1222_U195 ; P1_R1222_U198
g13575 nand P1_R1222_U6 P1_R1222_U42 ; P1_R1222_U199
g13576 not P1_R1222_U140 ; P1_R1222_U200
g13577 or P1_U3477 P1_U3082 ; P1_R1222_U201
g13578 nand P1_R1222_U201 P1_R1222_U140 ; P1_R1222_U202
g13579 not P1_R1222_U41 ; P1_R1222_U203
g13580 or P1_U3081 P1_U3480 ; P1_R1222_U204
g13581 or P1_U3471 P1_U3069 ; P1_R1222_U205
g13582 nand P1_R1222_U205 P1_R1222_U42 ; P1_R1222_U206
g13583 nand P1_R1222_U120 P1_R1222_U206 ; P1_R1222_U207
g13584 nand P1_R1222_U192 P1_R1222_U23 ; P1_R1222_U208
g13585 nand P1_U3474 P1_U3068 ; P1_R1222_U209
g13586 nand P1_R1222_U121 P1_R1222_U208 ; P1_R1222_U210
g13587 or P1_U3069 P1_U3471 ; P1_R1222_U211
g13588 nand P1_R1222_U182 P1_R1222_U178 ; P1_R1222_U212
g13589 nand P1_U3066 P1_U3459 ; P1_R1222_U213
g13590 not P1_R1222_U46 ; P1_R1222_U214
g13591 nand P1_R1222_U181 P1_R1222_U5 ; P1_R1222_U215
g13592 nand P1_R1222_U46 P1_R1222_U177 ; P1_R1222_U216
g13593 nand P1_U3062 P1_U3462 ; P1_R1222_U217
g13594 not P1_R1222_U45 ; P1_R1222_U218
g13595 or P1_U3465 P1_U3058 ; P1_R1222_U219
g13596 nand P1_R1222_U219 P1_R1222_U45 ; P1_R1222_U220
g13597 nand P1_R1222_U123 P1_R1222_U220 ; P1_R1222_U221
g13598 nand P1_R1222_U218 P1_R1222_U35 ; P1_R1222_U222
g13599 nand P1_U3468 P1_U3065 ; P1_R1222_U223
g13600 nand P1_R1222_U124 P1_R1222_U222 ; P1_R1222_U224
g13601 or P1_U3058 P1_U3465 ; P1_R1222_U225
g13602 nand P1_R1222_U181 P1_R1222_U178 ; P1_R1222_U226
g13603 not P1_R1222_U141 ; P1_R1222_U227
g13604 nand P1_U3062 P1_U3462 ; P1_R1222_U228
g13605 nand P1_R1222_U398 P1_R1222_U397 P1_R1222_U44 P1_R1222_U43 ; P1_R1222_U229
g13606 nand P1_R1222_U44 P1_R1222_U43 ; P1_R1222_U230
g13607 nand P1_U3066 P1_U3459 ; P1_R1222_U231
g13608 nand P1_R1222_U125 P1_R1222_U230 ; P1_R1222_U232
g13609 or P1_U3081 P1_U3480 ; P1_R1222_U233
g13610 or P1_U3060 P1_U3483 ; P1_R1222_U234
g13611 nand P1_R1222_U174 P1_R1222_U7 ; P1_R1222_U235
g13612 nand P1_U3060 P1_U3483 ; P1_R1222_U236
g13613 nand P1_R1222_U127 P1_R1222_U235 ; P1_R1222_U237
g13614 or P1_U3483 P1_U3060 ; P1_R1222_U238
g13615 nand P1_R1222_U126 P1_R1222_U140 ; P1_R1222_U239
g13616 nand P1_R1222_U238 P1_R1222_U237 ; P1_R1222_U240
g13617 not P1_R1222_U164 ; P1_R1222_U241
g13618 or P1_U3078 P1_U3492 ; P1_R1222_U242
g13619 or P1_U3070 P1_U3489 ; P1_R1222_U243
g13620 nand P1_R1222_U171 P1_R1222_U8 ; P1_R1222_U244
g13621 nand P1_U3078 P1_U3492 ; P1_R1222_U245
g13622 nand P1_R1222_U128 P1_R1222_U244 ; P1_R1222_U246
g13623 or P1_U3486 P1_U3061 ; P1_R1222_U247
g13624 or P1_U3492 P1_U3078 ; P1_R1222_U248
g13625 nand P1_R1222_U247 P1_R1222_U164 P1_R1222_U8 ; P1_R1222_U249
g13626 nand P1_R1222_U248 P1_R1222_U246 ; P1_R1222_U250
g13627 not P1_R1222_U163 ; P1_R1222_U251
g13628 or P1_U3495 P1_U3077 ; P1_R1222_U252
g13629 nand P1_R1222_U252 P1_R1222_U163 ; P1_R1222_U253
g13630 nand P1_U3077 P1_U3495 ; P1_R1222_U254
g13631 not P1_R1222_U161 ; P1_R1222_U255
g13632 or P1_U3498 P1_U3072 ; P1_R1222_U256
g13633 nand P1_R1222_U256 P1_R1222_U161 ; P1_R1222_U257
g13634 nand P1_U3072 P1_U3498 ; P1_R1222_U258
g13635 not P1_R1222_U93 ; P1_R1222_U259
g13636 or P1_U3067 P1_U3504 ; P1_R1222_U260
g13637 or P1_U3071 P1_U3501 ; P1_R1222_U261
g13638 not P1_R1222_U60 ; P1_R1222_U262
g13639 nand P1_R1222_U61 P1_R1222_U60 ; P1_R1222_U263
g13640 nand P1_U3067 P1_R1222_U263 ; P1_R1222_U264
g13641 nand P1_U3504 P1_R1222_U262 ; P1_R1222_U265
g13642 nand P1_R1222_U9 P1_R1222_U93 ; P1_R1222_U266
g13643 not P1_R1222_U159 ; P1_R1222_U267
g13644 or P1_U3074 P1_U4015 ; P1_R1222_U268
g13645 or P1_U3079 P1_U3509 ; P1_R1222_U269
g13646 or P1_U3073 P1_U4014 ; P1_R1222_U270
g13647 not P1_R1222_U81 ; P1_R1222_U271
g13648 nand P1_U4015 P1_R1222_U271 ; P1_R1222_U272
g13649 nand P1_R1222_U272 P1_R1222_U91 ; P1_R1222_U273
g13650 nand P1_R1222_U81 P1_R1222_U82 ; P1_R1222_U274
g13651 nand P1_R1222_U274 P1_R1222_U273 ; P1_R1222_U275
g13652 nand P1_R1222_U172 P1_R1222_U10 ; P1_R1222_U276
g13653 nand P1_U3073 P1_U4014 ; P1_R1222_U277
g13654 nand P1_R1222_U275 P1_R1222_U276 ; P1_R1222_U278
g13655 or P1_U3507 P1_U3080 ; P1_R1222_U279
g13656 or P1_U4014 P1_U3073 ; P1_R1222_U280
g13657 nand P1_R1222_U270 P1_R1222_U159 P1_R1222_U130 ; P1_R1222_U281
g13658 nand P1_R1222_U280 P1_R1222_U278 ; P1_R1222_U282
g13659 not P1_R1222_U155 ; P1_R1222_U283
g13660 or P1_U4013 P1_U3059 ; P1_R1222_U284
g13661 nand P1_R1222_U284 P1_R1222_U155 ; P1_R1222_U285
g13662 nand P1_U3059 P1_U4013 ; P1_R1222_U286
g13663 not P1_R1222_U153 ; P1_R1222_U287
g13664 or P1_U4012 P1_U3064 ; P1_R1222_U288
g13665 nand P1_R1222_U288 P1_R1222_U153 ; P1_R1222_U289
g13666 nand P1_U3064 P1_U4012 ; P1_R1222_U290
g13667 not P1_R1222_U151 ; P1_R1222_U291
g13668 or P1_U3056 P1_U4010 ; P1_R1222_U292
g13669 nand P1_R1222_U173 P1_R1222_U170 ; P1_R1222_U293
g13670 not P1_R1222_U87 ; P1_R1222_U294
g13671 or P1_U4011 P1_U3063 ; P1_R1222_U295
g13672 nand P1_R1222_U151 P1_R1222_U295 P1_R1222_U165 ; P1_R1222_U296
g13673 not P1_R1222_U149 ; P1_R1222_U297
g13674 or P1_U4008 P1_U3051 ; P1_R1222_U298
g13675 nand P1_U3051 P1_U4008 ; P1_R1222_U299
g13676 not P1_R1222_U147 ; P1_R1222_U300
g13677 nand P1_U4007 P1_R1222_U147 ; P1_R1222_U301
g13678 not P1_R1222_U145 ; P1_R1222_U302
g13679 nand P1_R1222_U295 P1_R1222_U151 ; P1_R1222_U303
g13680 not P1_R1222_U90 ; P1_R1222_U304
g13681 or P1_U4010 P1_U3056 ; P1_R1222_U305
g13682 nand P1_R1222_U305 P1_R1222_U90 ; P1_R1222_U306
g13683 nand P1_R1222_U306 P1_R1222_U170 P1_R1222_U150 ; P1_R1222_U307
g13684 nand P1_R1222_U304 P1_R1222_U170 ; P1_R1222_U308
g13685 nand P1_U4009 P1_U3055 ; P1_R1222_U309
g13686 nand P1_R1222_U308 P1_R1222_U309 P1_R1222_U165 ; P1_R1222_U310
g13687 or P1_U3056 P1_U4010 ; P1_R1222_U311
g13688 nand P1_R1222_U279 P1_R1222_U159 ; P1_R1222_U312
g13689 not P1_R1222_U92 ; P1_R1222_U313
g13690 nand P1_R1222_U10 P1_R1222_U92 ; P1_R1222_U314
g13691 nand P1_R1222_U134 P1_R1222_U314 ; P1_R1222_U315
g13692 nand P1_R1222_U314 P1_R1222_U275 ; P1_R1222_U316
g13693 nand P1_R1222_U450 P1_R1222_U316 ; P1_R1222_U317
g13694 or P1_U3509 P1_U3079 ; P1_R1222_U318
g13695 nand P1_R1222_U318 P1_R1222_U92 ; P1_R1222_U319
g13696 nand P1_R1222_U319 P1_R1222_U81 P1_R1222_U157 ; P1_R1222_U320
g13697 nand P1_R1222_U313 P1_R1222_U81 ; P1_R1222_U321
g13698 nand P1_U3074 P1_U4015 ; P1_R1222_U322
g13699 nand P1_R1222_U322 P1_R1222_U321 P1_R1222_U10 ; P1_R1222_U323
g13700 or P1_U3456 P1_U3076 ; P1_R1222_U324
g13701 not P1_R1222_U158 ; P1_R1222_U325
g13702 or P1_U3079 P1_U3509 ; P1_R1222_U326
g13703 or P1_U3501 P1_U3071 ; P1_R1222_U327
g13704 nand P1_R1222_U327 P1_R1222_U93 ; P1_R1222_U328
g13705 nand P1_R1222_U135 P1_R1222_U328 ; P1_R1222_U329
g13706 nand P1_R1222_U259 P1_R1222_U60 ; P1_R1222_U330
g13707 nand P1_U3504 P1_U3067 ; P1_R1222_U331
g13708 nand P1_R1222_U331 P1_R1222_U330 P1_R1222_U9 ; P1_R1222_U332
g13709 or P1_U3071 P1_U3501 ; P1_R1222_U333
g13710 nand P1_R1222_U247 P1_R1222_U164 ; P1_R1222_U334
g13711 not P1_R1222_U94 ; P1_R1222_U335
g13712 or P1_U3489 P1_U3070 ; P1_R1222_U336
g13713 nand P1_R1222_U336 P1_R1222_U94 ; P1_R1222_U337
g13714 nand P1_R1222_U136 P1_R1222_U337 ; P1_R1222_U338
g13715 nand P1_R1222_U335 P1_R1222_U169 ; P1_R1222_U339
g13716 nand P1_U3078 P1_U3492 ; P1_R1222_U340
g13717 nand P1_R1222_U137 P1_R1222_U339 ; P1_R1222_U341
g13718 or P1_U3070 P1_U3489 ; P1_R1222_U342
g13719 or P1_U3480 P1_U3081 ; P1_R1222_U343
g13720 nand P1_R1222_U343 P1_R1222_U41 ; P1_R1222_U344
g13721 nand P1_R1222_U138 P1_R1222_U344 ; P1_R1222_U345
g13722 nand P1_R1222_U203 P1_R1222_U168 ; P1_R1222_U346
g13723 nand P1_U3060 P1_U3483 ; P1_R1222_U347
g13724 nand P1_R1222_U139 P1_R1222_U346 ; P1_R1222_U348
g13725 nand P1_R1222_U204 P1_R1222_U168 ; P1_R1222_U349
g13726 nand P1_R1222_U201 P1_R1222_U62 ; P1_R1222_U350
g13727 nand P1_R1222_U211 P1_R1222_U23 ; P1_R1222_U351
g13728 nand P1_R1222_U225 P1_R1222_U35 ; P1_R1222_U352
g13729 nand P1_R1222_U228 P1_R1222_U177 ; P1_R1222_U353
g13730 nand P1_R1222_U311 P1_R1222_U170 ; P1_R1222_U354
g13731 nand P1_R1222_U295 P1_R1222_U173 ; P1_R1222_U355
g13732 nand P1_R1222_U326 P1_R1222_U81 ; P1_R1222_U356
g13733 nand P1_R1222_U279 P1_R1222_U78 ; P1_R1222_U357
g13734 nand P1_R1222_U333 P1_R1222_U60 ; P1_R1222_U358
g13735 nand P1_R1222_U342 P1_R1222_U169 ; P1_R1222_U359
g13736 nand P1_R1222_U247 P1_R1222_U69 ; P1_R1222_U360
g13737 nand P1_U4007 P1_U3052 ; P1_R1222_U361
g13738 nand P1_R1222_U293 P1_R1222_U165 ; P1_R1222_U362
g13739 nand P1_U3055 P1_R1222_U292 ; P1_R1222_U363
g13740 nand P1_U4009 P1_R1222_U292 ; P1_R1222_U364
g13741 nand P1_R1222_U293 P1_R1222_U165 P1_R1222_U298 ; P1_R1222_U365
g13742 nand P1_R1222_U151 P1_R1222_U165 P1_R1222_U132 ; P1_R1222_U366
g13743 nand P1_R1222_U294 P1_R1222_U298 ; P1_R1222_U367
g13744 nand P1_U3081 P1_R1222_U40 ; P1_R1222_U368
g13745 nand P1_U3480 P1_R1222_U39 ; P1_R1222_U369
g13746 nand P1_R1222_U369 P1_R1222_U368 ; P1_R1222_U370
g13747 nand P1_R1222_U349 P1_R1222_U41 ; P1_R1222_U371
g13748 nand P1_R1222_U370 P1_R1222_U203 ; P1_R1222_U372
g13749 nand P1_U3082 P1_R1222_U37 ; P1_R1222_U373
g13750 nand P1_U3477 P1_R1222_U38 ; P1_R1222_U374
g13751 nand P1_R1222_U374 P1_R1222_U373 ; P1_R1222_U375
g13752 nand P1_R1222_U350 P1_R1222_U140 ; P1_R1222_U376
g13753 nand P1_R1222_U200 P1_R1222_U375 ; P1_R1222_U377
g13754 nand P1_U3068 P1_R1222_U24 ; P1_R1222_U378
g13755 nand P1_U3474 P1_R1222_U22 ; P1_R1222_U379
g13756 nand P1_U3069 P1_R1222_U20 ; P1_R1222_U380
g13757 nand P1_U3471 P1_R1222_U21 ; P1_R1222_U381
g13758 nand P1_R1222_U381 P1_R1222_U380 ; P1_R1222_U382
g13759 nand P1_R1222_U351 P1_R1222_U42 ; P1_R1222_U383
g13760 nand P1_R1222_U382 P1_R1222_U192 ; P1_R1222_U384
g13761 nand P1_U3065 P1_R1222_U36 ; P1_R1222_U385
g13762 nand P1_U3468 P1_R1222_U27 ; P1_R1222_U386
g13763 nand P1_U3058 P1_R1222_U25 ; P1_R1222_U387
g13764 nand P1_U3465 P1_R1222_U26 ; P1_R1222_U388
g13765 nand P1_R1222_U388 P1_R1222_U387 ; P1_R1222_U389
g13766 nand P1_R1222_U352 P1_R1222_U45 ; P1_R1222_U390
g13767 nand P1_R1222_U389 P1_R1222_U218 ; P1_R1222_U391
g13768 nand P1_U3062 P1_R1222_U33 ; P1_R1222_U392
g13769 nand P1_U3462 P1_R1222_U34 ; P1_R1222_U393
g13770 nand P1_R1222_U393 P1_R1222_U392 ; P1_R1222_U394
g13771 nand P1_R1222_U353 P1_R1222_U141 ; P1_R1222_U395
g13772 nand P1_R1222_U227 P1_R1222_U394 ; P1_R1222_U396
g13773 nand P1_U3066 P1_R1222_U28 ; P1_R1222_U397
g13774 nand P1_U3459 P1_R1222_U29 ; P1_R1222_U398
g13775 nand P1_U3053 P1_R1222_U143 ; P1_R1222_U399
g13776 nand P1_U4018 P1_R1222_U142 ; P1_R1222_U400
g13777 nand P1_U3053 P1_R1222_U143 ; P1_R1222_U401
g13778 nand P1_U4018 P1_R1222_U142 ; P1_R1222_U402
g13779 nand P1_R1222_U402 P1_R1222_U401 ; P1_R1222_U403
g13780 nand P1_R1222_U144 P1_R1222_U145 ; P1_R1222_U404
g13781 nand P1_R1222_U302 P1_R1222_U403 ; P1_R1222_U405
g13782 nand P1_U3052 P1_R1222_U89 ; P1_R1222_U406
g13783 nand P1_U4007 P1_R1222_U88 ; P1_R1222_U407
g13784 nand P1_U3052 P1_R1222_U89 ; P1_R1222_U408
g13785 nand P1_U4007 P1_R1222_U88 ; P1_R1222_U409
g13786 nand P1_R1222_U409 P1_R1222_U408 ; P1_R1222_U410
g13787 nand P1_R1222_U146 P1_R1222_U147 ; P1_R1222_U411
g13788 nand P1_R1222_U300 P1_R1222_U410 ; P1_R1222_U412
g13789 nand P1_U3051 P1_R1222_U47 ; P1_R1222_U413
g13790 nand P1_U4008 P1_R1222_U48 ; P1_R1222_U414
g13791 nand P1_U3051 P1_R1222_U47 ; P1_R1222_U415
g13792 nand P1_U4008 P1_R1222_U48 ; P1_R1222_U416
g13793 nand P1_R1222_U416 P1_R1222_U415 ; P1_R1222_U417
g13794 nand P1_R1222_U148 P1_R1222_U149 ; P1_R1222_U418
g13795 nand P1_R1222_U297 P1_R1222_U417 ; P1_R1222_U419
g13796 nand P1_U3055 P1_R1222_U50 ; P1_R1222_U420
g13797 nand P1_U4009 P1_R1222_U49 ; P1_R1222_U421
g13798 nand P1_U3056 P1_R1222_U51 ; P1_R1222_U422
g13799 nand P1_U4010 P1_R1222_U52 ; P1_R1222_U423
g13800 nand P1_R1222_U423 P1_R1222_U422 ; P1_R1222_U424
g13801 nand P1_R1222_U354 P1_R1222_U90 ; P1_R1222_U425
g13802 nand P1_R1222_U424 P1_R1222_U304 ; P1_R1222_U426
g13803 nand P1_U3063 P1_R1222_U53 ; P1_R1222_U427
g13804 nand P1_U4011 P1_R1222_U54 ; P1_R1222_U428
g13805 nand P1_R1222_U428 P1_R1222_U427 ; P1_R1222_U429
g13806 nand P1_R1222_U355 P1_R1222_U151 ; P1_R1222_U430
g13807 nand P1_R1222_U291 P1_R1222_U429 ; P1_R1222_U431
g13808 nand P1_U3064 P1_R1222_U85 ; P1_R1222_U432
g13809 nand P1_U4012 P1_R1222_U86 ; P1_R1222_U433
g13810 nand P1_U3064 P1_R1222_U85 ; P1_R1222_U434
g13811 nand P1_U4012 P1_R1222_U86 ; P1_R1222_U435
g13812 nand P1_R1222_U435 P1_R1222_U434 ; P1_R1222_U436
g13813 nand P1_R1222_U152 P1_R1222_U153 ; P1_R1222_U437
g13814 nand P1_R1222_U287 P1_R1222_U436 ; P1_R1222_U438
g13815 nand P1_U3059 P1_R1222_U83 ; P1_R1222_U439
g13816 nand P1_U4013 P1_R1222_U84 ; P1_R1222_U440
g13817 nand P1_U3059 P1_R1222_U83 ; P1_R1222_U441
g13818 nand P1_U4013 P1_R1222_U84 ; P1_R1222_U442
g13819 nand P1_R1222_U442 P1_R1222_U441 ; P1_R1222_U443
g13820 nand P1_R1222_U154 P1_R1222_U155 ; P1_R1222_U444
g13821 nand P1_R1222_U283 P1_R1222_U443 ; P1_R1222_U445
g13822 nand P1_U3073 P1_R1222_U55 ; P1_R1222_U446
g13823 nand P1_U4014 P1_R1222_U56 ; P1_R1222_U447
g13824 nand P1_U3073 P1_R1222_U55 ; P1_R1222_U448
g13825 nand P1_U4014 P1_R1222_U56 ; P1_R1222_U449
g13826 nand P1_R1222_U449 P1_R1222_U448 ; P1_R1222_U450
g13827 nand P1_U3074 P1_R1222_U82 ; P1_R1222_U451
g13828 nand P1_U4015 P1_R1222_U91 ; P1_R1222_U452
g13829 nand P1_R1222_U179 P1_R1222_U158 ; P1_R1222_U453
g13830 nand P1_R1222_U325 P1_R1222_U32 ; P1_R1222_U454
g13831 nand P1_U3079 P1_R1222_U79 ; P1_R1222_U455
g13832 nand P1_U3509 P1_R1222_U80 ; P1_R1222_U456
g13833 nand P1_R1222_U456 P1_R1222_U455 ; P1_R1222_U457
g13834 nand P1_R1222_U356 P1_R1222_U92 ; P1_R1222_U458
g13835 nand P1_R1222_U457 P1_R1222_U313 ; P1_R1222_U459
g13836 nand P1_U3080 P1_R1222_U76 ; P1_R1222_U460
g13837 nand P1_U3507 P1_R1222_U77 ; P1_R1222_U461
g13838 nand P1_R1222_U461 P1_R1222_U460 ; P1_R1222_U462
g13839 nand P1_R1222_U357 P1_R1222_U159 ; P1_R1222_U463
g13840 nand P1_R1222_U267 P1_R1222_U462 ; P1_R1222_U464
g13841 nand P1_U3067 P1_R1222_U61 ; P1_R1222_U465
g13842 nand P1_U3504 P1_R1222_U59 ; P1_R1222_U466
g13843 nand P1_U3071 P1_R1222_U57 ; P1_R1222_U467
g13844 nand P1_U3501 P1_R1222_U58 ; P1_R1222_U468
g13845 nand P1_R1222_U468 P1_R1222_U467 ; P1_R1222_U469
g13846 nand P1_R1222_U358 P1_R1222_U93 ; P1_R1222_U470
g13847 nand P1_R1222_U469 P1_R1222_U259 ; P1_R1222_U471
g13848 nand P1_U3072 P1_R1222_U74 ; P1_R1222_U472
g13849 nand P1_U3498 P1_R1222_U75 ; P1_R1222_U473
g13850 nand P1_U3072 P1_R1222_U74 ; P1_R1222_U474
g13851 nand P1_U3498 P1_R1222_U75 ; P1_R1222_U475
g13852 nand P1_R1222_U475 P1_R1222_U474 ; P1_R1222_U476
g13853 nand P1_R1222_U160 P1_R1222_U161 ; P1_R1222_U477
g13854 nand P1_R1222_U255 P1_R1222_U476 ; P1_R1222_U478
g13855 nand P1_U3077 P1_R1222_U72 ; P1_R1222_U479
g13856 nand P1_U3495 P1_R1222_U73 ; P1_R1222_U480
g13857 nand P1_U3077 P1_R1222_U72 ; P1_R1222_U481
g13858 nand P1_U3495 P1_R1222_U73 ; P1_R1222_U482
g13859 nand P1_R1222_U482 P1_R1222_U481 ; P1_R1222_U483
g13860 nand P1_R1222_U162 P1_R1222_U163 ; P1_R1222_U484
g13861 nand P1_R1222_U251 P1_R1222_U483 ; P1_R1222_U485
g13862 nand P1_U3078 P1_R1222_U70 ; P1_R1222_U486
g13863 nand P1_U3492 P1_R1222_U71 ; P1_R1222_U487
g13864 nand P1_U3070 P1_R1222_U65 ; P1_R1222_U488
g13865 nand P1_U3489 P1_R1222_U66 ; P1_R1222_U489
g13866 nand P1_R1222_U489 P1_R1222_U488 ; P1_R1222_U490
g13867 nand P1_R1222_U359 P1_R1222_U94 ; P1_R1222_U491
g13868 nand P1_R1222_U490 P1_R1222_U335 ; P1_R1222_U492
g13869 nand P1_U3061 P1_R1222_U67 ; P1_R1222_U493
g13870 nand P1_U3486 P1_R1222_U68 ; P1_R1222_U494
g13871 nand P1_R1222_U494 P1_R1222_U493 ; P1_R1222_U495
g13872 nand P1_R1222_U360 P1_R1222_U164 ; P1_R1222_U496
g13873 nand P1_R1222_U241 P1_R1222_U495 ; P1_R1222_U497
g13874 nand P1_U3060 P1_R1222_U63 ; P1_R1222_U498
g13875 nand P1_U3483 P1_R1222_U64 ; P1_R1222_U499
g13876 nand P1_U3075 P1_R1222_U30 ; P1_R1222_U500
g13877 nand P1_U3451 P1_R1222_U31 ; P1_R1222_U501
g13878 not P2_REG3_REG_3__SCAN_IN ; P2_ADD_609_U4
g13879 and P2_ADD_609_U76 P2_ADD_609_U104 ; P2_ADD_609_U5
g13880 not P2_REG3_REG_7__SCAN_IN ; P2_ADD_609_U6
g13881 not P2_REG3_REG_6__SCAN_IN ; P2_ADD_609_U7
g13882 not P2_REG3_REG_5__SCAN_IN ; P2_ADD_609_U8
g13883 not P2_REG3_REG_4__SCAN_IN ; P2_ADD_609_U9
g13884 nand P2_REG3_REG_6__SCAN_IN P2_REG3_REG_4__SCAN_IN P2_REG3_REG_5__SCAN_IN P2_REG3_REG_3__SCAN_IN P2_REG3_REG_7__SCAN_IN ; P2_ADD_609_U10
g13885 not P2_REG3_REG_8__SCAN_IN ; P2_ADD_609_U11
g13886 not P2_REG3_REG_9__SCAN_IN ; P2_ADD_609_U12
g13887 nand P2_ADD_609_U74 P2_ADD_609_U85 ; P2_ADD_609_U13
g13888 not P2_REG3_REG_11__SCAN_IN ; P2_ADD_609_U14
g13889 not P2_REG3_REG_10__SCAN_IN ; P2_ADD_609_U15
g13890 nand P2_ADD_609_U75 P2_ADD_609_U87 ; P2_ADD_609_U16
g13891 not P2_REG3_REG_12__SCAN_IN ; P2_ADD_609_U17
g13892 nand P2_ADD_609_U89 P2_REG3_REG_12__SCAN_IN ; P2_ADD_609_U18
g13893 not P2_REG3_REG_13__SCAN_IN ; P2_ADD_609_U19
g13894 nand P2_ADD_609_U90 P2_REG3_REG_13__SCAN_IN ; P2_ADD_609_U20
g13895 not P2_REG3_REG_14__SCAN_IN ; P2_ADD_609_U21
g13896 nand P2_ADD_609_U91 P2_REG3_REG_14__SCAN_IN ; P2_ADD_609_U22
g13897 not P2_REG3_REG_15__SCAN_IN ; P2_ADD_609_U23
g13898 nand P2_ADD_609_U92 P2_REG3_REG_15__SCAN_IN ; P2_ADD_609_U24
g13899 not P2_REG3_REG_16__SCAN_IN ; P2_ADD_609_U25
g13900 nand P2_ADD_609_U93 P2_REG3_REG_16__SCAN_IN ; P2_ADD_609_U26
g13901 not P2_REG3_REG_17__SCAN_IN ; P2_ADD_609_U27
g13902 nand P2_ADD_609_U94 P2_REG3_REG_17__SCAN_IN ; P2_ADD_609_U28
g13903 not P2_REG3_REG_18__SCAN_IN ; P2_ADD_609_U29
g13904 nand P2_ADD_609_U95 P2_REG3_REG_18__SCAN_IN ; P2_ADD_609_U30
g13905 not P2_REG3_REG_19__SCAN_IN ; P2_ADD_609_U31
g13906 nand P2_ADD_609_U96 P2_REG3_REG_19__SCAN_IN ; P2_ADD_609_U32
g13907 not P2_REG3_REG_20__SCAN_IN ; P2_ADD_609_U33
g13908 nand P2_ADD_609_U97 P2_REG3_REG_20__SCAN_IN ; P2_ADD_609_U34
g13909 not P2_REG3_REG_21__SCAN_IN ; P2_ADD_609_U35
g13910 nand P2_ADD_609_U98 P2_REG3_REG_21__SCAN_IN ; P2_ADD_609_U36
g13911 not P2_REG3_REG_22__SCAN_IN ; P2_ADD_609_U37
g13912 nand P2_ADD_609_U99 P2_REG3_REG_22__SCAN_IN ; P2_ADD_609_U38
g13913 not P2_REG3_REG_23__SCAN_IN ; P2_ADD_609_U39
g13914 nand P2_ADD_609_U100 P2_REG3_REG_23__SCAN_IN ; P2_ADD_609_U40
g13915 not P2_REG3_REG_24__SCAN_IN ; P2_ADD_609_U41
g13916 nand P2_ADD_609_U101 P2_REG3_REG_24__SCAN_IN ; P2_ADD_609_U42
g13917 not P2_REG3_REG_25__SCAN_IN ; P2_ADD_609_U43
g13918 nand P2_ADD_609_U102 P2_REG3_REG_25__SCAN_IN ; P2_ADD_609_U44
g13919 not P2_REG3_REG_26__SCAN_IN ; P2_ADD_609_U45
g13920 nand P2_ADD_609_U103 P2_REG3_REG_26__SCAN_IN ; P2_ADD_609_U46
g13921 not P2_REG3_REG_28__SCAN_IN ; P2_ADD_609_U47
g13922 not P2_REG3_REG_27__SCAN_IN ; P2_ADD_609_U48
g13923 nand P2_ADD_609_U108 P2_ADD_609_U107 ; P2_ADD_609_U49
g13924 nand P2_ADD_609_U110 P2_ADD_609_U109 ; P2_ADD_609_U50
g13925 nand P2_ADD_609_U112 P2_ADD_609_U111 ; P2_ADD_609_U51
g13926 nand P2_ADD_609_U114 P2_ADD_609_U113 ; P2_ADD_609_U52
g13927 nand P2_ADD_609_U116 P2_ADD_609_U115 ; P2_ADD_609_U53
g13928 nand P2_ADD_609_U118 P2_ADD_609_U117 ; P2_ADD_609_U54
g13929 nand P2_ADD_609_U120 P2_ADD_609_U119 ; P2_ADD_609_U55
g13930 nand P2_ADD_609_U122 P2_ADD_609_U121 ; P2_ADD_609_U56
g13931 nand P2_ADD_609_U124 P2_ADD_609_U123 ; P2_ADD_609_U57
g13932 nand P2_ADD_609_U126 P2_ADD_609_U125 ; P2_ADD_609_U58
g13933 nand P2_ADD_609_U128 P2_ADD_609_U127 ; P2_ADD_609_U59
g13934 nand P2_ADD_609_U130 P2_ADD_609_U129 ; P2_ADD_609_U60
g13935 nand P2_ADD_609_U132 P2_ADD_609_U131 ; P2_ADD_609_U61
g13936 nand P2_ADD_609_U134 P2_ADD_609_U133 ; P2_ADD_609_U62
g13937 nand P2_ADD_609_U136 P2_ADD_609_U135 ; P2_ADD_609_U63
g13938 nand P2_ADD_609_U138 P2_ADD_609_U137 ; P2_ADD_609_U64
g13939 nand P2_ADD_609_U140 P2_ADD_609_U139 ; P2_ADD_609_U65
g13940 nand P2_ADD_609_U142 P2_ADD_609_U141 ; P2_ADD_609_U66
g13941 nand P2_ADD_609_U144 P2_ADD_609_U143 ; P2_ADD_609_U67
g13942 nand P2_ADD_609_U146 P2_ADD_609_U145 ; P2_ADD_609_U68
g13943 nand P2_ADD_609_U148 P2_ADD_609_U147 ; P2_ADD_609_U69
g13944 nand P2_ADD_609_U150 P2_ADD_609_U149 ; P2_ADD_609_U70
g13945 nand P2_ADD_609_U152 P2_ADD_609_U151 ; P2_ADD_609_U71
g13946 nand P2_ADD_609_U154 P2_ADD_609_U153 ; P2_ADD_609_U72
g13947 nand P2_ADD_609_U156 P2_ADD_609_U155 ; P2_ADD_609_U73
g13948 and P2_REG3_REG_9__SCAN_IN P2_REG3_REG_8__SCAN_IN ; P2_ADD_609_U74
g13949 and P2_REG3_REG_11__SCAN_IN P2_REG3_REG_10__SCAN_IN ; P2_ADD_609_U75
g13950 and P2_REG3_REG_28__SCAN_IN P2_REG3_REG_27__SCAN_IN ; P2_ADD_609_U76
g13951 nand P2_ADD_609_U85 P2_REG3_REG_8__SCAN_IN ; P2_ADD_609_U77
g13952 nand P2_REG3_REG_6__SCAN_IN P2_REG3_REG_4__SCAN_IN P2_REG3_REG_5__SCAN_IN P2_REG3_REG_3__SCAN_IN ; P2_ADD_609_U78
g13953 nand P2_REG3_REG_4__SCAN_IN P2_REG3_REG_5__SCAN_IN P2_REG3_REG_3__SCAN_IN ; P2_ADD_609_U79
g13954 nand P2_REG3_REG_4__SCAN_IN P2_REG3_REG_3__SCAN_IN ; P2_ADD_609_U80
g13955 nand P2_ADD_609_U104 P2_REG3_REG_27__SCAN_IN ; P2_ADD_609_U81
g13956 nand P2_ADD_609_U87 P2_REG3_REG_10__SCAN_IN ; P2_ADD_609_U82
g13957 not P2_ADD_609_U80 ; P2_ADD_609_U83
g13958 not P2_ADD_609_U78 ; P2_ADD_609_U84
g13959 not P2_ADD_609_U10 ; P2_ADD_609_U85
g13960 not P2_ADD_609_U77 ; P2_ADD_609_U86
g13961 not P2_ADD_609_U13 ; P2_ADD_609_U87
g13962 not P2_ADD_609_U82 ; P2_ADD_609_U88
g13963 not P2_ADD_609_U16 ; P2_ADD_609_U89
g13964 not P2_ADD_609_U18 ; P2_ADD_609_U90
g13965 not P2_ADD_609_U20 ; P2_ADD_609_U91
g13966 not P2_ADD_609_U22 ; P2_ADD_609_U92
g13967 not P2_ADD_609_U24 ; P2_ADD_609_U93
g13968 not P2_ADD_609_U26 ; P2_ADD_609_U94
g13969 not P2_ADD_609_U28 ; P2_ADD_609_U95
g13970 not P2_ADD_609_U30 ; P2_ADD_609_U96
g13971 not P2_ADD_609_U32 ; P2_ADD_609_U97
g13972 not P2_ADD_609_U34 ; P2_ADD_609_U98
g13973 not P2_ADD_609_U36 ; P2_ADD_609_U99
g13974 not P2_ADD_609_U38 ; P2_ADD_609_U100
g13975 not P2_ADD_609_U40 ; P2_ADD_609_U101
g13976 not P2_ADD_609_U42 ; P2_ADD_609_U102
g13977 not P2_ADD_609_U44 ; P2_ADD_609_U103
g13978 not P2_ADD_609_U46 ; P2_ADD_609_U104
g13979 not P2_ADD_609_U81 ; P2_ADD_609_U105
g13980 not P2_ADD_609_U79 ; P2_ADD_609_U106
g13981 nand P2_ADD_609_U77 P2_REG3_REG_9__SCAN_IN ; P2_ADD_609_U107
g13982 nand P2_ADD_609_U86 P2_ADD_609_U12 ; P2_ADD_609_U108
g13983 nand P2_ADD_609_U10 P2_REG3_REG_8__SCAN_IN ; P2_ADD_609_U109
g13984 nand P2_ADD_609_U85 P2_ADD_609_U11 ; P2_ADD_609_U110
g13985 nand P2_ADD_609_U78 P2_REG3_REG_7__SCAN_IN ; P2_ADD_609_U111
g13986 nand P2_ADD_609_U84 P2_ADD_609_U6 ; P2_ADD_609_U112
g13987 nand P2_ADD_609_U79 P2_REG3_REG_6__SCAN_IN ; P2_ADD_609_U113
g13988 nand P2_ADD_609_U106 P2_ADD_609_U7 ; P2_ADD_609_U114
g13989 nand P2_ADD_609_U80 P2_REG3_REG_5__SCAN_IN ; P2_ADD_609_U115
g13990 nand P2_ADD_609_U83 P2_ADD_609_U8 ; P2_ADD_609_U116
g13991 nand P2_ADD_609_U4 P2_REG3_REG_4__SCAN_IN ; P2_ADD_609_U117
g13992 nand P2_ADD_609_U9 P2_REG3_REG_3__SCAN_IN ; P2_ADD_609_U118
g13993 nand P2_ADD_609_U81 P2_REG3_REG_28__SCAN_IN ; P2_ADD_609_U119
g13994 nand P2_ADD_609_U105 P2_ADD_609_U47 ; P2_ADD_609_U120
g13995 nand P2_ADD_609_U46 P2_REG3_REG_27__SCAN_IN ; P2_ADD_609_U121
g13996 nand P2_ADD_609_U104 P2_ADD_609_U48 ; P2_ADD_609_U122
g13997 nand P2_ADD_609_U44 P2_REG3_REG_26__SCAN_IN ; P2_ADD_609_U123
g13998 nand P2_ADD_609_U103 P2_ADD_609_U45 ; P2_ADD_609_U124
g13999 nand P2_ADD_609_U42 P2_REG3_REG_25__SCAN_IN ; P2_ADD_609_U125
g14000 nand P2_ADD_609_U102 P2_ADD_609_U43 ; P2_ADD_609_U126
g14001 nand P2_ADD_609_U40 P2_REG3_REG_24__SCAN_IN ; P2_ADD_609_U127
g14002 nand P2_ADD_609_U101 P2_ADD_609_U41 ; P2_ADD_609_U128
g14003 nand P2_ADD_609_U38 P2_REG3_REG_23__SCAN_IN ; P2_ADD_609_U129
g14004 nand P2_ADD_609_U100 P2_ADD_609_U39 ; P2_ADD_609_U130
g14005 nand P2_ADD_609_U36 P2_REG3_REG_22__SCAN_IN ; P2_ADD_609_U131
g14006 nand P2_ADD_609_U99 P2_ADD_609_U37 ; P2_ADD_609_U132
g14007 nand P2_ADD_609_U34 P2_REG3_REG_21__SCAN_IN ; P2_ADD_609_U133
g14008 nand P2_ADD_609_U98 P2_ADD_609_U35 ; P2_ADD_609_U134
g14009 nand P2_ADD_609_U32 P2_REG3_REG_20__SCAN_IN ; P2_ADD_609_U135
g14010 nand P2_ADD_609_U97 P2_ADD_609_U33 ; P2_ADD_609_U136
g14011 nand P2_ADD_609_U30 P2_REG3_REG_19__SCAN_IN ; P2_ADD_609_U137
g14012 nand P2_ADD_609_U96 P2_ADD_609_U31 ; P2_ADD_609_U138
g14013 nand P2_ADD_609_U28 P2_REG3_REG_18__SCAN_IN ; P2_ADD_609_U139
g14014 nand P2_ADD_609_U95 P2_ADD_609_U29 ; P2_ADD_609_U140
g14015 nand P2_ADD_609_U26 P2_REG3_REG_17__SCAN_IN ; P2_ADD_609_U141
g14016 nand P2_ADD_609_U94 P2_ADD_609_U27 ; P2_ADD_609_U142
g14017 nand P2_ADD_609_U24 P2_REG3_REG_16__SCAN_IN ; P2_ADD_609_U143
g14018 nand P2_ADD_609_U93 P2_ADD_609_U25 ; P2_ADD_609_U144
g14019 nand P2_ADD_609_U22 P2_REG3_REG_15__SCAN_IN ; P2_ADD_609_U145
g14020 nand P2_ADD_609_U92 P2_ADD_609_U23 ; P2_ADD_609_U146
g14021 nand P2_ADD_609_U20 P2_REG3_REG_14__SCAN_IN ; P2_ADD_609_U147
g14022 nand P2_ADD_609_U91 P2_ADD_609_U21 ; P2_ADD_609_U148
g14023 nand P2_ADD_609_U18 P2_REG3_REG_13__SCAN_IN ; P2_ADD_609_U149
g14024 nand P2_ADD_609_U90 P2_ADD_609_U19 ; P2_ADD_609_U150
g14025 nand P2_ADD_609_U16 P2_REG3_REG_12__SCAN_IN ; P2_ADD_609_U151
g14026 nand P2_ADD_609_U89 P2_ADD_609_U17 ; P2_ADD_609_U152
g14027 nand P2_ADD_609_U82 P2_REG3_REG_11__SCAN_IN ; P2_ADD_609_U153
g14028 nand P2_ADD_609_U88 P2_ADD_609_U14 ; P2_ADD_609_U154
g14029 nand P2_ADD_609_U13 P2_REG3_REG_10__SCAN_IN ; P2_ADD_609_U155
g14030 nand P2_ADD_609_U87 P2_ADD_609_U15 ; P2_ADD_609_U156
g14031 and P2_R1340_U179 P2_R1340_U176 P2_R1340_U175 P2_R1340_U173 ; P2_R1340_U6
g14032 not P2_U3456 ; P2_R1340_U7
g14033 not P2_U3459 ; P2_R1340_U8
g14034 not P2_U3462 ; P2_R1340_U9
g14035 not P2_U3182 ; P2_R1340_U10
g14036 not P2_U3181 ; P2_R1340_U11
g14037 not P2_U3180 ; P2_R1340_U12
g14038 not P2_U3179 ; P2_R1340_U13
g14039 not P2_U3178 ; P2_R1340_U14
g14040 not P2_U3177 ; P2_R1340_U15
g14041 not P2_U3465 ; P2_R1340_U16
g14042 not P2_U3468 ; P2_R1340_U17
g14043 not P2_U3471 ; P2_R1340_U18
g14044 not P2_U3474 ; P2_R1340_U19
g14045 not P2_U3477 ; P2_R1340_U20
g14046 not P2_U3480 ; P2_R1340_U21
g14047 not P2_U3176 ; P2_R1340_U22
g14048 not P2_U3175 ; P2_R1340_U23
g14049 not P2_U3174 ; P2_R1340_U24
g14050 not P2_U3173 ; P2_R1340_U25
g14051 not P2_U3172 ; P2_R1340_U26
g14052 not P2_U3171 ; P2_R1340_U27
g14053 not P2_U3483 ; P2_R1340_U28
g14054 not P2_U3486 ; P2_R1340_U29
g14055 not P2_U3489 ; P2_R1340_U30
g14056 not P2_U3492 ; P2_R1340_U31
g14057 not P2_U3495 ; P2_R1340_U32
g14058 not P2_U3498 ; P2_R1340_U33
g14059 not P2_U3170 ; P2_R1340_U34
g14060 not P2_U3169 ; P2_R1340_U35
g14061 not P2_U3168 ; P2_R1340_U36
g14062 not P2_U3167 ; P2_R1340_U37
g14063 not P2_U3501 ; P2_R1340_U38
g14064 not P2_U3504 ; P2_R1340_U39
g14065 not P2_U3166 ; P2_R1340_U40
g14066 not P2_U3165 ; P2_R1340_U41
g14067 not P2_U3506 ; P2_R1340_U42
g14068 not P2_U3976 ; P2_R1340_U43
g14069 not P2_U3164 ; P2_R1340_U44
g14070 not P2_U3163 ; P2_R1340_U45
g14071 not P2_U3975 ; P2_R1340_U46
g14072 not P2_U3974 ; P2_R1340_U47
g14073 not P2_U3162 ; P2_R1340_U48
g14074 not P2_U3161 ; P2_R1340_U49
g14075 not P2_U3973 ; P2_R1340_U50
g14076 not P2_U3972 ; P2_R1340_U51
g14077 not P2_U3160 ; P2_R1340_U52
g14078 not P2_U3159 ; P2_R1340_U53
g14079 not P2_U3971 ; P2_R1340_U54
g14080 not P2_U3970 ; P2_R1340_U55
g14081 not P2_U3158 ; P2_R1340_U56
g14082 not P2_U3157 ; P2_R1340_U57
g14083 not P2_U3969 ; P2_R1340_U58
g14084 not P2_U3968 ; P2_R1340_U59
g14085 not P2_U3156 ; P2_R1340_U60
g14086 not P2_U3155 ; P2_R1340_U61
g14087 not P2_U3979 ; P2_R1340_U62
g14088 not P2_U3153 ; P2_R1340_U63
g14089 not P2_U3977 ; P2_R1340_U64
g14090 and P2_R1340_U99 P2_R1340_U100 P2_R1340_U98 ; P2_R1340_U65
g14091 and P2_R1340_U105 P2_R1340_U104 P2_R1340_U178 ; P2_R1340_U66
g14092 and P2_U3181 P2_R1340_U8 ; P2_R1340_U67
g14093 and P2_R1340_U106 P2_R1340_U103 P2_R1340_U102 P2_R1340_U69 ; P2_R1340_U68
g14094 and P2_R1340_U111 P2_R1340_U107 P2_R1340_U112 ; P2_R1340_U69
g14095 and P2_U3468 P2_R1340_U14 ; P2_R1340_U70
g14096 and P2_R1340_U113 P2_R1340_U110 P2_R1340_U109 P2_R1340_U72 ; P2_R1340_U71
g14097 and P2_R1340_U118 P2_R1340_U114 P2_R1340_U119 ; P2_R1340_U72
g14098 and P2_U3175 P2_R1340_U20 ; P2_R1340_U73
g14099 and P2_R1340_U120 P2_R1340_U117 P2_R1340_U116 P2_R1340_U75 ; P2_R1340_U74
g14100 and P2_R1340_U125 P2_R1340_U121 P2_R1340_U126 ; P2_R1340_U75
g14101 and P2_U3486 P2_R1340_U26 ; P2_R1340_U76
g14102 and P2_R1340_U127 P2_R1340_U124 P2_R1340_U123 P2_R1340_U78 ; P2_R1340_U77
g14103 and P2_R1340_U132 P2_R1340_U128 P2_R1340_U133 ; P2_R1340_U78
g14104 and P2_U3169 P2_R1340_U32 ; P2_R1340_U79
g14105 and P2_R1340_U81 P2_R1340_U131 P2_R1340_U130 ; P2_R1340_U80
g14106 and P2_R1340_U135 P2_R1340_U134 ; P2_R1340_U81
g14107 and P2_R1340_U137 P2_R1340_U138 ; P2_R1340_U82
g14108 and P2_R1340_U140 P2_R1340_U141 ; P2_R1340_U83
g14109 and P2_R1340_U143 P2_R1340_U144 ; P2_R1340_U84
g14110 and P2_R1340_U146 P2_R1340_U147 ; P2_R1340_U85
g14111 and P2_R1340_U149 P2_R1340_U150 ; P2_R1340_U86
g14112 and P2_R1340_U152 P2_R1340_U153 ; P2_R1340_U87
g14113 and P2_R1340_U155 P2_R1340_U156 ; P2_R1340_U88
g14114 and P2_R1340_U158 P2_R1340_U159 ; P2_R1340_U89
g14115 and P2_R1340_U161 P2_R1340_U162 ; P2_R1340_U90
g14116 and P2_R1340_U164 P2_R1340_U165 ; P2_R1340_U91
g14117 and P2_R1340_U170 P2_R1340_U171 ; P2_R1340_U92
g14118 and P2_R1340_U177 P2_R1340_U174 ; P2_R1340_U93
g14119 and P2_U3154 P2_R1340_U177 ; P2_R1340_U94
g14120 not P2_U3978 ; P2_R1340_U95
g14121 not P2_U3183 ; P2_R1340_U96
g14122 not P2_U3184 ; P2_R1340_U97
g14123 nand P2_R1340_U97 P2_R1340_U96 P2_U3448 ; P2_R1340_U98
g14124 nand P2_U3453 P2_R1340_U96 ; P2_R1340_U99
g14125 nand P2_U3456 P2_R1340_U10 ; P2_R1340_U100
g14126 nand P2_R1340_U66 P2_R1340_U65 ; P2_R1340_U101
g14127 nand P2_U3182 P2_R1340_U105 P2_R1340_U104 P2_R1340_U7 ; P2_R1340_U102
g14128 nand P2_R1340_U67 P2_R1340_U105 ; P2_R1340_U103
g14129 nand P2_U3459 P2_R1340_U11 ; P2_R1340_U104
g14130 nand P2_U3462 P2_R1340_U12 ; P2_R1340_U105
g14131 nand P2_U3180 P2_R1340_U9 ; P2_R1340_U106
g14132 nand P2_U3179 P2_R1340_U16 ; P2_R1340_U107
g14133 nand P2_R1340_U101 P2_R1340_U68 ; P2_R1340_U108
g14134 nand P2_U3465 P2_R1340_U112 P2_R1340_U111 P2_R1340_U13 ; P2_R1340_U109
g14135 nand P2_R1340_U70 P2_R1340_U112 ; P2_R1340_U110
g14136 nand P2_U3178 P2_R1340_U17 ; P2_R1340_U111
g14137 nand P2_U3177 P2_R1340_U18 ; P2_R1340_U112
g14138 nand P2_U3471 P2_R1340_U15 ; P2_R1340_U113
g14139 nand P2_U3474 P2_R1340_U22 ; P2_R1340_U114
g14140 nand P2_R1340_U108 P2_R1340_U71 ; P2_R1340_U115
g14141 nand P2_U3176 P2_R1340_U119 P2_R1340_U118 P2_R1340_U19 ; P2_R1340_U116
g14142 nand P2_R1340_U73 P2_R1340_U119 ; P2_R1340_U117
g14143 nand P2_U3477 P2_R1340_U23 ; P2_R1340_U118
g14144 nand P2_U3480 P2_R1340_U24 ; P2_R1340_U119
g14145 nand P2_U3174 P2_R1340_U21 ; P2_R1340_U120
g14146 nand P2_U3173 P2_R1340_U28 ; P2_R1340_U121
g14147 nand P2_R1340_U115 P2_R1340_U74 ; P2_R1340_U122
g14148 nand P2_U3483 P2_R1340_U126 P2_R1340_U125 P2_R1340_U25 ; P2_R1340_U123
g14149 nand P2_R1340_U76 P2_R1340_U126 ; P2_R1340_U124
g14150 nand P2_U3172 P2_R1340_U29 ; P2_R1340_U125
g14151 nand P2_U3171 P2_R1340_U30 ; P2_R1340_U126
g14152 nand P2_U3489 P2_R1340_U27 ; P2_R1340_U127
g14153 nand P2_U3492 P2_R1340_U34 ; P2_R1340_U128
g14154 nand P2_R1340_U122 P2_R1340_U77 ; P2_R1340_U129
g14155 nand P2_U3170 P2_R1340_U133 P2_R1340_U132 P2_R1340_U31 ; P2_R1340_U130
g14156 nand P2_R1340_U79 P2_R1340_U133 ; P2_R1340_U131
g14157 nand P2_U3495 P2_R1340_U35 ; P2_R1340_U132
g14158 nand P2_U3498 P2_R1340_U36 ; P2_R1340_U133
g14159 nand P2_U3168 P2_R1340_U33 ; P2_R1340_U134
g14160 nand P2_U3167 P2_R1340_U38 ; P2_R1340_U135
g14161 nand P2_R1340_U129 P2_R1340_U80 ; P2_R1340_U136
g14162 nand P2_U3501 P2_R1340_U37 ; P2_R1340_U137
g14163 nand P2_U3504 P2_R1340_U40 ; P2_R1340_U138
g14164 nand P2_R1340_U82 P2_R1340_U136 ; P2_R1340_U139
g14165 nand P2_U3166 P2_R1340_U39 ; P2_R1340_U140
g14166 nand P2_U3165 P2_R1340_U42 ; P2_R1340_U141
g14167 nand P2_R1340_U83 P2_R1340_U139 ; P2_R1340_U142
g14168 nand P2_U3506 P2_R1340_U41 ; P2_R1340_U143
g14169 nand P2_U3976 P2_R1340_U44 ; P2_R1340_U144
g14170 nand P2_R1340_U84 P2_R1340_U142 ; P2_R1340_U145
g14171 nand P2_U3164 P2_R1340_U43 ; P2_R1340_U146
g14172 nand P2_U3163 P2_R1340_U46 ; P2_R1340_U147
g14173 nand P2_R1340_U85 P2_R1340_U145 ; P2_R1340_U148
g14174 nand P2_U3975 P2_R1340_U45 ; P2_R1340_U149
g14175 nand P2_U3974 P2_R1340_U48 ; P2_R1340_U150
g14176 nand P2_R1340_U86 P2_R1340_U148 ; P2_R1340_U151
g14177 nand P2_U3162 P2_R1340_U47 ; P2_R1340_U152
g14178 nand P2_U3161 P2_R1340_U50 ; P2_R1340_U153
g14179 nand P2_R1340_U87 P2_R1340_U151 ; P2_R1340_U154
g14180 nand P2_U3973 P2_R1340_U49 ; P2_R1340_U155
g14181 nand P2_U3972 P2_R1340_U52 ; P2_R1340_U156
g14182 nand P2_R1340_U88 P2_R1340_U154 ; P2_R1340_U157
g14183 nand P2_U3160 P2_R1340_U51 ; P2_R1340_U158
g14184 nand P2_U3159 P2_R1340_U54 ; P2_R1340_U159
g14185 nand P2_R1340_U89 P2_R1340_U157 ; P2_R1340_U160
g14186 nand P2_U3971 P2_R1340_U53 ; P2_R1340_U161
g14187 nand P2_U3970 P2_R1340_U56 ; P2_R1340_U162
g14188 nand P2_R1340_U90 P2_R1340_U160 ; P2_R1340_U163
g14189 nand P2_U3158 P2_R1340_U55 ; P2_R1340_U164
g14190 nand P2_U3157 P2_R1340_U58 ; P2_R1340_U165
g14191 nand P2_R1340_U91 P2_R1340_U163 ; P2_R1340_U166
g14192 nand P2_U3969 P2_R1340_U57 ; P2_R1340_U167
g14193 nand P2_U3968 P2_R1340_U60 ; P2_R1340_U168
g14194 nand P2_R1340_U167 P2_R1340_U166 P2_R1340_U168 ; P2_R1340_U169
g14195 nand P2_U3156 P2_R1340_U59 ; P2_R1340_U170
g14196 nand P2_U3155 P2_R1340_U62 ; P2_R1340_U171
g14197 nand P2_R1340_U92 P2_R1340_U169 ; P2_R1340_U172
g14198 nand P2_R1340_U172 P2_R1340_U95 P2_R1340_U93 ; P2_R1340_U173
g14199 nand P2_U3979 P2_R1340_U61 ; P2_R1340_U174
g14200 nand P2_U3977 P2_R1340_U63 ; P2_R1340_U175
g14201 nand P2_R1340_U177 P2_U3154 P2_R1340_U95 ; P2_R1340_U176
g14202 nand P2_U3153 P2_R1340_U64 ; P2_R1340_U177
g14203 nand P2_U3448 P2_U3453 P2_R1340_U97 ; P2_R1340_U178
g14204 nand P2_R1340_U174 P2_R1340_U172 P2_R1340_U94 ; P2_R1340_U179
g14205 and P2_SUB_598_U57 P2_SUB_598_U56 ; P2_SUB_598_U6
g14206 nor P2_IR_REG_25__SCAN_IN P2_IR_REG_26__SCAN_IN P2_IR_REG_27__SCAN_IN ; P2_SUB_598_U7
g14207 nor P2_IR_REG_25__SCAN_IN P2_IR_REG_26__SCAN_IN ; P2_SUB_598_U8
g14208 and P2_SUB_598_U55 P2_SUB_598_U54 P2_SUB_598_U53 P2_SUB_598_U52 ; P2_SUB_598_U9
g14209 nor P2_IR_REG_9__SCAN_IN P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN ; P2_SUB_598_U10
g14210 and P2_SUB_598_U142 P2_SUB_598_U47 ; P2_SUB_598_U11
g14211 and P2_SUB_598_U140 P2_SUB_598_U111 ; P2_SUB_598_U12
g14212 and P2_SUB_598_U139 P2_SUB_598_U43 ; P2_SUB_598_U13
g14213 and P2_SUB_598_U138 P2_SUB_598_U44 ; P2_SUB_598_U14
g14214 and P2_SUB_598_U136 P2_SUB_598_U114 ; P2_SUB_598_U15
g14215 and P2_SUB_598_U135 P2_SUB_598_U96 ; P2_SUB_598_U16
g14216 and P2_SUB_598_U134 P2_SUB_598_U125 ; P2_SUB_598_U17
g14217 and P2_SUB_598_U132 P2_SUB_598_U126 ; P2_SUB_598_U18
g14218 and P2_SUB_598_U131 P2_SUB_598_U91 ; P2_SUB_598_U19
g14219 and P2_SUB_598_U64 P2_SUB_598_U144 ; P2_SUB_598_U20
g14220 and P2_SUB_598_U130 P2_SUB_598_U89 ; P2_SUB_598_U21
g14221 and P2_SUB_598_U124 P2_SUB_598_U116 ; P2_SUB_598_U22
g14222 and P2_SUB_598_U123 P2_SUB_598_U117 ; P2_SUB_598_U23
g14223 and P2_SUB_598_U122 P2_SUB_598_U34 ; P2_SUB_598_U24
g14224 and P2_SUB_598_U109 P2_SUB_598_U101 ; P2_SUB_598_U25
g14225 and P2_SUB_598_U108 P2_SUB_598_U30 ; P2_SUB_598_U26
g14226 and P2_SUB_598_U107 P2_SUB_598_U32 ; P2_SUB_598_U27
g14227 and P2_SUB_598_U105 P2_SUB_598_U103 ; P2_SUB_598_U28
g14228 and P2_SUB_598_U104 P2_SUB_598_U31 ; P2_SUB_598_U29
g14229 or P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_2__SCAN_IN P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN ; P2_SUB_598_U30
g14230 nand P2_SUB_598_U50 P2_SUB_598_U148 ; P2_SUB_598_U31
g14231 nand P2_SUB_598_U51 P2_SUB_598_U148 ; P2_SUB_598_U32
g14232 not P2_IR_REG_7__SCAN_IN ; P2_SUB_598_U33
g14233 or P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_2__SCAN_IN ; P2_SUB_598_U34
g14234 not P2_IR_REG_3__SCAN_IN ; P2_SUB_598_U35
g14235 nand P2_SUB_598_U6 P2_SUB_598_U9 ; P2_SUB_598_U36
g14236 nand P2_SUB_598_U58 P2_SUB_598_U147 ; P2_SUB_598_U37
g14237 nand P2_SUB_598_U118 P2_SUB_598_U80 ; P2_SUB_598_U38
g14238 not P2_IR_REG_25__SCAN_IN ; P2_SUB_598_U39
g14239 nand P2_SUB_598_U62 P2_SUB_598_U9 ; P2_SUB_598_U40
g14240 not P2_IR_REG_23__SCAN_IN ; P2_SUB_598_U41
g14241 not P2_IR_REG_21__SCAN_IN ; P2_SUB_598_U42
g14242 nand P2_SUB_598_U10 P2_SUB_598_U149 ; P2_SUB_598_U43
g14243 nand P2_SUB_598_U69 P2_SUB_598_U112 ; P2_SUB_598_U44
g14244 not P2_IR_REG_16__SCAN_IN ; P2_SUB_598_U45
g14245 not P2_IR_REG_15__SCAN_IN ; P2_SUB_598_U46
g14246 nand P2_SUB_598_U70 P2_SUB_598_U149 ; P2_SUB_598_U47
g14247 not P2_IR_REG_11__SCAN_IN ; P2_SUB_598_U48
g14248 nand P2_SUB_598_U169 P2_SUB_598_U168 ; P2_SUB_598_U49
g14249 nor P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN ; P2_SUB_598_U50
g14250 nor P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_598_U51
g14251 nor P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN P2_IR_REG_13__SCAN_IN P2_IR_REG_14__SCAN_IN ; P2_SUB_598_U52
g14252 nor P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_15__SCAN_IN P2_IR_REG_16__SCAN_IN ; P2_SUB_598_U53
g14253 nor P2_IR_REG_2__SCAN_IN P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN ; P2_SUB_598_U54
g14254 nor P2_IR_REG_6__SCAN_IN P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN P2_IR_REG_9__SCAN_IN ; P2_SUB_598_U55
g14255 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN P2_IR_REG_20__SCAN_IN ; P2_SUB_598_U56
g14256 nor P2_IR_REG_21__SCAN_IN P2_IR_REG_22__SCAN_IN P2_IR_REG_23__SCAN_IN P2_IR_REG_24__SCAN_IN ; P2_SUB_598_U57
g14257 and P2_SUB_598_U7 P2_SUB_598_U82 ; P2_SUB_598_U58
g14258 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN ; P2_SUB_598_U59
g14259 nor P2_IR_REG_19__SCAN_IN P2_IR_REG_20__SCAN_IN ; P2_SUB_598_U60
g14260 nor P2_IR_REG_21__SCAN_IN P2_IR_REG_22__SCAN_IN ; P2_SUB_598_U61
g14261 and P2_SUB_598_U60 P2_SUB_598_U59 P2_SUB_598_U61 ; P2_SUB_598_U62
g14262 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN P2_IR_REG_20__SCAN_IN ; P2_SUB_598_U63
g14263 and P2_SUB_598_U143 P2_SUB_598_U40 ; P2_SUB_598_U64
g14264 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN ; P2_SUB_598_U65
g14265 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN ; P2_SUB_598_U66
g14266 nor P2_IR_REG_13__SCAN_IN P2_IR_REG_14__SCAN_IN P2_IR_REG_15__SCAN_IN ; P2_SUB_598_U67
g14267 and P2_SUB_598_U10 P2_SUB_598_U45 P2_SUB_598_U67 ; P2_SUB_598_U68
g14268 nor P2_IR_REG_13__SCAN_IN P2_IR_REG_14__SCAN_IN ; P2_SUB_598_U69
g14269 nor P2_IR_REG_9__SCAN_IN P2_IR_REG_10__SCAN_IN ; P2_SUB_598_U70
g14270 not P2_IR_REG_9__SCAN_IN ; P2_SUB_598_U71
g14271 and P2_SUB_598_U151 P2_SUB_598_U150 ; P2_SUB_598_U72
g14272 not P2_IR_REG_5__SCAN_IN ; P2_SUB_598_U73
g14273 and P2_SUB_598_U153 P2_SUB_598_U152 ; P2_SUB_598_U74
g14274 not P2_IR_REG_31__SCAN_IN ; P2_SUB_598_U75
g14275 nand P2_SUB_598_U119 P2_SUB_598_U78 ; P2_SUB_598_U76
g14276 and P2_SUB_598_U155 P2_SUB_598_U154 ; P2_SUB_598_U77
g14277 not P2_IR_REG_30__SCAN_IN ; P2_SUB_598_U78
g14278 and P2_SUB_598_U157 P2_SUB_598_U156 ; P2_SUB_598_U79
g14279 not P2_IR_REG_29__SCAN_IN ; P2_SUB_598_U80
g14280 and P2_SUB_598_U159 P2_SUB_598_U158 ; P2_SUB_598_U81
g14281 not P2_IR_REG_28__SCAN_IN ; P2_SUB_598_U82
g14282 nand P2_SUB_598_U6 P2_SUB_598_U7 P2_SUB_598_U9 ; P2_SUB_598_U83
g14283 and P2_SUB_598_U161 P2_SUB_598_U160 ; P2_SUB_598_U84
g14284 not P2_IR_REG_27__SCAN_IN ; P2_SUB_598_U85
g14285 nand P2_SUB_598_U6 P2_SUB_598_U8 P2_SUB_598_U9 ; P2_SUB_598_U86
g14286 and P2_SUB_598_U163 P2_SUB_598_U162 ; P2_SUB_598_U87
g14287 not P2_IR_REG_24__SCAN_IN ; P2_SUB_598_U88
g14288 nand P2_SUB_598_U128 P2_SUB_598_U41 ; P2_SUB_598_U89
g14289 and P2_SUB_598_U165 P2_SUB_598_U164 ; P2_SUB_598_U90
g14290 nand P2_SUB_598_U63 P2_SUB_598_U9 ; P2_SUB_598_U91
g14291 and P2_SUB_598_U167 P2_SUB_598_U166 ; P2_SUB_598_U92
g14292 not P2_IR_REG_1__SCAN_IN ; P2_SUB_598_U93
g14293 not P2_IR_REG_0__SCAN_IN ; P2_SUB_598_U94
g14294 not P2_IR_REG_17__SCAN_IN ; P2_SUB_598_U95
g14295 nand P2_SUB_598_U68 P2_SUB_598_U149 ; P2_SUB_598_U96
g14296 and P2_SUB_598_U171 P2_SUB_598_U170 ; P2_SUB_598_U97
g14297 not P2_IR_REG_13__SCAN_IN ; P2_SUB_598_U98
g14298 and P2_SUB_598_U173 P2_SUB_598_U172 ; P2_SUB_598_U99
g14299 not P2_SUB_598_U34 ; P2_SUB_598_U100
g14300 nand P2_SUB_598_U100 P2_SUB_598_U35 ; P2_SUB_598_U101
g14301 not P2_SUB_598_U32 ; P2_SUB_598_U102
g14302 nand P2_SUB_598_U102 P2_SUB_598_U33 ; P2_SUB_598_U103
g14303 nand P2_SUB_598_U103 P2_IR_REG_8__SCAN_IN ; P2_SUB_598_U104
g14304 nand P2_SUB_598_U32 P2_IR_REG_7__SCAN_IN ; P2_SUB_598_U105
g14305 nand P2_SUB_598_U148 P2_SUB_598_U73 ; P2_SUB_598_U106
g14306 nand P2_SUB_598_U106 P2_IR_REG_6__SCAN_IN ; P2_SUB_598_U107
g14307 nand P2_SUB_598_U101 P2_IR_REG_4__SCAN_IN ; P2_SUB_598_U108
g14308 nand P2_SUB_598_U34 P2_IR_REG_3__SCAN_IN ; P2_SUB_598_U109
g14309 not P2_SUB_598_U47 ; P2_SUB_598_U110
g14310 nand P2_SUB_598_U110 P2_SUB_598_U48 ; P2_SUB_598_U111
g14311 not P2_SUB_598_U43 ; P2_SUB_598_U112
g14312 not P2_SUB_598_U44 ; P2_SUB_598_U113
g14313 nand P2_SUB_598_U113 P2_SUB_598_U46 ; P2_SUB_598_U114
g14314 not P2_SUB_598_U96 ; P2_SUB_598_U115
g14315 nand P2_SUB_598_U147 P2_SUB_598_U39 ; P2_SUB_598_U116
g14316 nand P2_SUB_598_U8 P2_SUB_598_U147 ; P2_SUB_598_U117
g14317 not P2_SUB_598_U37 ; P2_SUB_598_U118
g14318 not P2_SUB_598_U38 ; P2_SUB_598_U119
g14319 not P2_SUB_598_U76 ; P2_SUB_598_U120
g14320 or P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN ; P2_SUB_598_U121
g14321 nand P2_SUB_598_U121 P2_IR_REG_2__SCAN_IN ; P2_SUB_598_U122
g14322 nand P2_SUB_598_U116 P2_IR_REG_26__SCAN_IN ; P2_SUB_598_U123
g14323 nand P2_SUB_598_U36 P2_IR_REG_25__SCAN_IN ; P2_SUB_598_U124
g14324 nand P2_SUB_598_U66 P2_SUB_598_U9 ; P2_SUB_598_U125
g14325 nand P2_SUB_598_U65 P2_SUB_598_U9 ; P2_SUB_598_U126
g14326 not P2_SUB_598_U91 ; P2_SUB_598_U127
g14327 not P2_SUB_598_U40 ; P2_SUB_598_U128
g14328 not P2_SUB_598_U89 ; P2_SUB_598_U129
g14329 nand P2_SUB_598_U40 P2_IR_REG_23__SCAN_IN ; P2_SUB_598_U130
g14330 nand P2_SUB_598_U126 P2_IR_REG_20__SCAN_IN ; P2_SUB_598_U131
g14331 nand P2_SUB_598_U125 P2_IR_REG_19__SCAN_IN ; P2_SUB_598_U132
g14332 nand P2_SUB_598_U9 P2_SUB_598_U95 ; P2_SUB_598_U133
g14333 nand P2_SUB_598_U133 P2_IR_REG_18__SCAN_IN ; P2_SUB_598_U134
g14334 nand P2_SUB_598_U114 P2_IR_REG_16__SCAN_IN ; P2_SUB_598_U135
g14335 nand P2_SUB_598_U44 P2_IR_REG_15__SCAN_IN ; P2_SUB_598_U136
g14336 nand P2_SUB_598_U112 P2_SUB_598_U98 ; P2_SUB_598_U137
g14337 nand P2_SUB_598_U137 P2_IR_REG_14__SCAN_IN ; P2_SUB_598_U138
g14338 nand P2_SUB_598_U111 P2_IR_REG_12__SCAN_IN ; P2_SUB_598_U139
g14339 nand P2_SUB_598_U47 P2_IR_REG_11__SCAN_IN ; P2_SUB_598_U140
g14340 nand P2_SUB_598_U149 P2_SUB_598_U71 ; P2_SUB_598_U141
g14341 nand P2_SUB_598_U141 P2_IR_REG_10__SCAN_IN ; P2_SUB_598_U142
g14342 nand P2_IR_REG_21__SCAN_IN P2_IR_REG_22__SCAN_IN ; P2_SUB_598_U143
g14343 nand P2_SUB_598_U91 P2_IR_REG_22__SCAN_IN ; P2_SUB_598_U144
g14344 not P2_SUB_598_U86 ; P2_SUB_598_U145
g14345 not P2_SUB_598_U83 ; P2_SUB_598_U146
g14346 not P2_SUB_598_U36 ; P2_SUB_598_U147
g14347 not P2_SUB_598_U30 ; P2_SUB_598_U148
g14348 not P2_SUB_598_U31 ; P2_SUB_598_U149
g14349 nand P2_SUB_598_U31 P2_IR_REG_9__SCAN_IN ; P2_SUB_598_U150
g14350 nand P2_SUB_598_U149 P2_SUB_598_U71 ; P2_SUB_598_U151
g14351 nand P2_SUB_598_U30 P2_IR_REG_5__SCAN_IN ; P2_SUB_598_U152
g14352 nand P2_SUB_598_U148 P2_SUB_598_U73 ; P2_SUB_598_U153
g14353 nand P2_SUB_598_U76 P2_IR_REG_31__SCAN_IN ; P2_SUB_598_U154
g14354 nand P2_SUB_598_U120 P2_SUB_598_U75 ; P2_SUB_598_U155
g14355 nand P2_SUB_598_U38 P2_IR_REG_30__SCAN_IN ; P2_SUB_598_U156
g14356 nand P2_SUB_598_U119 P2_SUB_598_U78 ; P2_SUB_598_U157
g14357 nand P2_SUB_598_U37 P2_IR_REG_29__SCAN_IN ; P2_SUB_598_U158
g14358 nand P2_SUB_598_U118 P2_SUB_598_U80 ; P2_SUB_598_U159
g14359 nand P2_SUB_598_U83 P2_IR_REG_28__SCAN_IN ; P2_SUB_598_U160
g14360 nand P2_SUB_598_U146 P2_SUB_598_U82 ; P2_SUB_598_U161
g14361 nand P2_SUB_598_U86 P2_IR_REG_27__SCAN_IN ; P2_SUB_598_U162
g14362 nand P2_SUB_598_U145 P2_SUB_598_U85 ; P2_SUB_598_U163
g14363 nand P2_SUB_598_U89 P2_IR_REG_24__SCAN_IN ; P2_SUB_598_U164
g14364 nand P2_SUB_598_U129 P2_SUB_598_U88 ; P2_SUB_598_U165
g14365 nand P2_SUB_598_U91 P2_IR_REG_21__SCAN_IN ; P2_SUB_598_U166
g14366 nand P2_SUB_598_U127 P2_SUB_598_U42 ; P2_SUB_598_U167
g14367 nand P2_SUB_598_U94 P2_IR_REG_1__SCAN_IN ; P2_SUB_598_U168
g14368 nand P2_SUB_598_U93 P2_IR_REG_0__SCAN_IN ; P2_SUB_598_U169
g14369 nand P2_SUB_598_U96 P2_IR_REG_17__SCAN_IN ; P2_SUB_598_U170
g14370 nand P2_SUB_598_U115 P2_SUB_598_U95 ; P2_SUB_598_U171
g14371 nand P2_SUB_598_U43 P2_IR_REG_13__SCAN_IN ; P2_SUB_598_U172
g14372 nand P2_SUB_598_U112 P2_SUB_598_U98 ; P2_SUB_598_U173
g14373 and P2_U3059 P2_R1299_U7 ; P2_R1299_U6
g14374 not P2_U3056 ; P2_R1299_U7
g14375 and P2_R1312_U129 P2_R1312_U130 ; P2_R1312_U6
g14376 and P2_R1312_U131 P2_R1312_U132 ; P2_R1312_U7
g14377 and P2_R1312_U96 P2_R1312_U134 P2_R1312_U136 P2_R1312_U7 ; P2_R1312_U8
g14378 and P2_R1312_U143 P2_R1312_U144 ; P2_R1312_U9
g14379 and P2_R1312_U146 P2_R1312_U145 ; P2_R1312_U10
g14380 and P2_R1312_U99 P2_R1312_U147 P2_R1312_U100 ; P2_R1312_U11
g14381 and P2_R1312_U101 P2_R1312_U11 ; P2_R1312_U12
g14382 and P2_R1312_U162 P2_R1312_U161 ; P2_R1312_U13
g14383 and P2_R1312_U128 P2_R1312_U127 ; P2_R1312_U14
g14384 and P2_R1312_U85 P2_R1312_U20 ; P2_R1312_U15
g14385 and P2_R1312_U87 P2_R1312_U20 ; P2_R1312_U16
g14386 and P2_R1312_U89 P2_R1312_U20 ; P2_R1312_U17
g14387 and P2_R1312_U90 P2_R1312_U20 ; P2_R1312_U18
g14388 and P2_R1312_U119 P2_R1312_U20 ; P2_R1312_U19
g14389 and P2_R1312_U207 P2_R1312_U206 ; P2_R1312_U20
g14390 nand P2_R1312_U204 P2_R1312_U203 P2_R1312_U14 P2_R1312_U120 ; P2_R1312_U21
g14391 not P2_U3117 ; P2_R1312_U22
g14392 not P2_U3085 ; P2_R1312_U23
g14393 not P2_U3118 ; P2_R1312_U24
g14394 not P2_U3086 ; P2_R1312_U25
g14395 not P2_U3119 ; P2_R1312_U26
g14396 not P2_U3087 ; P2_R1312_U27
g14397 not P2_U3088 ; P2_R1312_U28
g14398 not P2_U3090 ; P2_R1312_U29
g14399 not P2_U3089 ; P2_R1312_U30
g14400 not P2_U3123 ; P2_R1312_U31
g14401 not P2_U3122 ; P2_R1312_U32
g14402 not P2_U3121 ; P2_R1312_U33
g14403 not P2_U3120 ; P2_R1312_U34
g14404 not P2_U3125 ; P2_R1312_U35
g14405 not P2_U3124 ; P2_R1312_U36
g14406 not P2_U3095 ; P2_R1312_U37
g14407 not P2_U3128 ; P2_R1312_U38
g14408 not P2_U3096 ; P2_R1312_U39
g14409 not P2_U3129 ; P2_R1312_U40
g14410 not P2_U3130 ; P2_R1312_U41
g14411 not P2_U3099 ; P2_R1312_U42
g14412 not P2_U3131 ; P2_R1312_U43
g14413 not P2_U3100 ; P2_R1312_U44
g14414 not P2_U3098 ; P2_R1312_U45
g14415 not P2_U3097 ; P2_R1312_U46
g14416 not P2_U3132 ; P2_R1312_U47
g14417 not P2_U3133 ; P2_R1312_U48
g14418 not P2_U3101 ; P2_R1312_U49
g14419 not P2_U3102 ; P2_R1312_U50
g14420 not P2_U3142 ; P2_R1312_U51
g14421 not P2_U3111 ; P2_R1312_U52
g14422 not P2_U3108 ; P2_R1312_U53
g14423 not P2_U3107 ; P2_R1312_U54
g14424 not P2_U3143 ; P2_R1312_U55
g14425 not P2_U3112 ; P2_R1312_U56
g14426 not P2_U3110 ; P2_R1312_U57
g14427 not P2_U3109 ; P2_R1312_U58
g14428 not P2_U3113 ; P2_R1312_U59
g14429 not P2_U3114 ; P2_R1312_U60
g14430 not P2_U3115 ; P2_R1312_U61
g14431 not P2_U3137 ; P2_R1312_U62
g14432 not P2_U3136 ; P2_R1312_U63
g14433 not P2_U3140 ; P2_R1312_U64
g14434 not P2_U3141 ; P2_R1312_U65
g14435 not P2_U3147 ; P2_R1312_U66
g14436 not P2_U3146 ; P2_R1312_U67
g14437 not P2_U3144 ; P2_R1312_U68
g14438 not P2_U3145 ; P2_R1312_U69
g14439 not P2_U3139 ; P2_R1312_U70
g14440 not P2_U3138 ; P2_R1312_U71
g14441 not P2_U3105 ; P2_R1312_U72
g14442 not P2_U3106 ; P2_R1312_U73
g14443 not P2_U3103 ; P2_R1312_U74
g14444 not P2_U3104 ; P2_R1312_U75
g14445 not P2_U3135 ; P2_R1312_U76
g14446 not P2_U3134 ; P2_R1312_U77
g14447 not P2_U3127 ; P2_R1312_U78
g14448 not P2_U3126 ; P2_R1312_U79
g14449 not P2_U3094 ; P2_R1312_U80
g14450 not P2_U3093 ; P2_R1312_U81
g14451 not P2_U3091 ; P2_R1312_U82
g14452 not P2_U3092 ; P2_R1312_U83
g14453 and P2_R1312_U27 P2_U3119 ; P2_R1312_U84
g14454 and P2_R1312_U124 P2_R1312_U82 P2_U3123 P2_R1312_U125 P2_R1312_U123 ; P2_R1312_U85
g14455 and P2_U3122 P2_R1312_U29 ; P2_R1312_U86
g14456 and P2_R1312_U86 P2_R1312_U125 P2_R1312_U123 ; P2_R1312_U87
g14457 and P2_U3121 P2_R1312_U30 ; P2_R1312_U88
g14458 and P2_R1312_U88 P2_R1312_U123 ; P2_R1312_U89
g14459 and P2_U3120 P2_R1312_U28 ; P2_R1312_U90
g14460 and P2_U3128 P2_R1312_U39 ; P2_R1312_U91
g14461 and P2_U3129 P2_R1312_U46 ; P2_R1312_U92
g14462 and P2_R1312_U182 P2_R1312_U181 ; P2_R1312_U93
g14463 and P2_U3099 P2_R1312_U43 ; P2_R1312_U94
g14464 and P2_U3100 P2_R1312_U47 ; P2_R1312_U95
g14465 and P2_R1312_U135 P2_R1312_U133 ; P2_R1312_U96
g14466 and P2_U3111 P2_R1312_U55 ; P2_R1312_U97
g14467 and P2_U3112 P2_R1312_U68 ; P2_R1312_U98
g14468 and P2_R1312_U148 P2_R1312_U142 ; P2_R1312_U99
g14469 and P2_R1312_U9 P2_R1312_U149 ; P2_R1312_U100
g14470 and P2_R1312_U151 P2_R1312_U150 ; P2_R1312_U101
g14471 and P2_R1312_U154 P2_R1312_U155 P2_R1312_U153 ; P2_R1312_U102
g14472 and P2_U3140 P2_R1312_U53 ; P2_R1312_U103
g14473 and P2_U3141 P2_R1312_U58 ; P2_R1312_U104
g14474 and P2_U3147 P2_R1312_U61 ; P2_R1312_U105
g14475 and P2_U3146 P2_R1312_U60 ; P2_R1312_U106
g14476 and P2_R1312_U13 P2_R1312_U108 ; P2_R1312_U107
g14477 and P2_R1312_U167 P2_R1312_U168 ; P2_R1312_U108
g14478 and P2_R1312_U166 P2_R1312_U107 ; P2_R1312_U109
g14479 and P2_U3105 P2_R1312_U62 ; P2_R1312_U110
g14480 and P2_U3106 P2_R1312_U71 ; P2_R1312_U111
g14481 and P2_R1312_U171 P2_R1312_U114 ; P2_R1312_U112
g14482 and P2_R1312_U112 P2_R1312_U172 ; P2_R1312_U113
g14483 and P2_R1312_U174 P2_R1312_U173 ; P2_R1312_U114
g14484 and P2_R1312_U185 P2_R1312_U184 P2_R1312_U138 ; P2_R1312_U115
g14485 and P2_R1312_U117 P2_R1312_U186 ; P2_R1312_U116
g14486 and P2_R1312_U189 P2_R1312_U188 ; P2_R1312_U117
g14487 and P2_R1312_U196 P2_R1312_U194 P2_R1312_U195 ; P2_R1312_U118
g14488 and P2_R1312_U190 P2_R1312_U124 P2_R1312_U118 P2_R1312_U125 P2_R1312_U123 ; P2_R1312_U119
g14489 and P2_R1312_U202 P2_R1312_U201 P2_R1312_U200 P2_R1312_U199 ; P2_R1312_U120
g14490 nand P2_R1312_U198 P2_R1312_U197 ; P2_R1312_U121
g14491 nand P2_U3087 P2_R1312_U26 ; P2_R1312_U122
g14492 nand P2_U3088 P2_R1312_U34 ; P2_R1312_U123
g14493 nand P2_U3090 P2_R1312_U32 ; P2_R1312_U124
g14494 nand P2_U3089 P2_R1312_U33 ; P2_R1312_U125
g14495 nand P2_U3086 P2_R1312_U24 ; P2_R1312_U126
g14496 nand P2_R1312_U209 P2_R1312_U208 P2_R1312_U205 ; P2_R1312_U127
g14497 nand P2_R1312_U20 P2_U3118 P2_R1312_U25 ; P2_R1312_U128
g14498 nand P2_U3130 P2_R1312_U45 ; P2_R1312_U129
g14499 nand P2_U3131 P2_R1312_U42 ; P2_R1312_U130
g14500 nand P2_U3095 P2_R1312_U78 ; P2_R1312_U131
g14501 nand P2_U3096 P2_R1312_U38 ; P2_R1312_U132
g14502 nand P2_R1312_U94 P2_R1312_U129 ; P2_R1312_U133
g14503 nand P2_R1312_U95 P2_R1312_U6 ; P2_R1312_U134
g14504 nand P2_U3098 P2_R1312_U41 ; P2_R1312_U135
g14505 nand P2_U3097 P2_R1312_U40 ; P2_R1312_U136
g14506 nand P2_U3101 P2_R1312_U48 ; P2_R1312_U137
g14507 nand P2_U3125 P2_R1312_U81 ; P2_R1312_U138
g14508 nand P2_U3124 P2_R1312_U83 ; P2_R1312_U139
g14509 nand P2_U3102 P2_R1312_U77 ; P2_R1312_U140
g14510 nand P2_U3142 P2_R1312_U57 ; P2_R1312_U141
g14511 nand P2_R1312_U97 P2_R1312_U141 ; P2_R1312_U142
g14512 nand P2_U3107 P2_R1312_U70 ; P2_R1312_U143
g14513 nand P2_U3108 P2_R1312_U64 ; P2_R1312_U144
g14514 nand P2_U3143 P2_R1312_U52 ; P2_R1312_U145
g14515 nand P2_U3142 P2_R1312_U57 ; P2_R1312_U146
g14516 nand P2_R1312_U98 P2_R1312_U10 ; P2_R1312_U147
g14517 nand P2_U3110 P2_R1312_U51 ; P2_R1312_U148
g14518 nand P2_U3109 P2_R1312_U65 ; P2_R1312_U149
g14519 nand P2_U3113 P2_R1312_U69 ; P2_R1312_U150
g14520 nand P2_U3114 P2_R1312_U67 ; P2_R1312_U151
g14521 nand P2_U3148 P2_U3149 ; P2_R1312_U152
g14522 nand P2_U3116 P2_R1312_U152 ; P2_R1312_U153
g14523 or P2_U3148 P2_U3149 ; P2_R1312_U154
g14524 nand P2_U3115 P2_R1312_U66 ; P2_R1312_U155
g14525 nand P2_R1312_U102 P2_R1312_U12 ; P2_R1312_U156
g14526 nand P2_R1312_U106 P2_R1312_U150 ; P2_R1312_U157
g14527 nand P2_U3144 P2_R1312_U56 ; P2_R1312_U158
g14528 nand P2_U3145 P2_R1312_U59 ; P2_R1312_U159
g14529 nand P2_R1312_U10 P2_R1312_U159 P2_R1312_U158 P2_R1312_U157 ; P2_R1312_U160
g14530 nand P2_U3137 P2_R1312_U72 ; P2_R1312_U161
g14531 nand P2_U3136 P2_R1312_U75 ; P2_R1312_U162
g14532 nand P2_R1312_U103 P2_R1312_U143 ; P2_R1312_U163
g14533 nand P2_R1312_U104 P2_R1312_U9 ; P2_R1312_U164
g14534 nand P2_R1312_U105 P2_R1312_U12 ; P2_R1312_U165
g14535 nand P2_R1312_U11 P2_R1312_U160 ; P2_R1312_U166
g14536 nand P2_U3139 P2_R1312_U54 ; P2_R1312_U167
g14537 nand P2_U3138 P2_R1312_U73 ; P2_R1312_U168
g14538 nand P2_R1312_U165 P2_R1312_U164 P2_R1312_U163 P2_R1312_U156 P2_R1312_U109 ; P2_R1312_U169
g14539 nand P2_U3136 P2_R1312_U75 ; P2_R1312_U170
g14540 nand P2_R1312_U110 P2_R1312_U170 ; P2_R1312_U171
g14541 nand P2_R1312_U111 P2_R1312_U13 ; P2_R1312_U172
g14542 nand P2_U3103 P2_R1312_U76 ; P2_R1312_U173
g14543 nand P2_U3104 P2_R1312_U63 ; P2_R1312_U174
g14544 nand P2_R1312_U169 P2_R1312_U113 ; P2_R1312_U175
g14545 nand P2_U3135 P2_R1312_U74 ; P2_R1312_U176
g14546 nand P2_R1312_U176 P2_R1312_U175 ; P2_R1312_U177
g14547 nand P2_R1312_U177 P2_R1312_U140 ; P2_R1312_U178
g14548 nand P2_U3134 P2_R1312_U50 ; P2_R1312_U179
g14549 nand P2_R1312_U179 P2_R1312_U178 ; P2_R1312_U180
g14550 nand P2_U3132 P2_R1312_U44 ; P2_R1312_U181
g14551 nand P2_U3133 P2_R1312_U49 ; P2_R1312_U182
g14552 nand P2_R1312_U93 P2_R1312_U6 ; P2_R1312_U183
g14553 nand P2_R1312_U91 P2_R1312_U131 ; P2_R1312_U184
g14554 nand P2_R1312_U92 P2_R1312_U7 ; P2_R1312_U185
g14555 nand P2_R1312_U8 P2_R1312_U183 ; P2_R1312_U186
g14556 nand P2_R1312_U180 P2_R1312_U137 P2_R1312_U8 ; P2_R1312_U187
g14557 nand P2_U3127 P2_R1312_U37 ; P2_R1312_U188
g14558 nand P2_U3126 P2_R1312_U80 ; P2_R1312_U189
g14559 nand P2_R1312_U187 P2_R1312_U116 P2_R1312_U115 P2_R1312_U139 ; P2_R1312_U190
g14560 nand P2_U3094 P2_R1312_U79 ; P2_R1312_U191
g14561 nand P2_U3093 P2_R1312_U35 ; P2_R1312_U192
g14562 nand P2_R1312_U192 P2_R1312_U191 ; P2_R1312_U193
g14563 nand P2_R1312_U193 P2_R1312_U138 P2_R1312_U139 ; P2_R1312_U194
g14564 nand P2_U3091 P2_R1312_U31 ; P2_R1312_U195
g14565 nand P2_U3092 P2_R1312_U36 ; P2_R1312_U196
g14566 nand P2_U3118 P2_R1312_U122 ; P2_R1312_U197
g14567 nand P2_R1312_U122 P2_R1312_U25 ; P2_R1312_U198
g14568 nand P2_R1312_U84 P2_R1312_U20 P2_R1312_U126 ; P2_R1312_U199
g14569 nand P2_R1312_U15 P2_R1312_U121 ; P2_R1312_U200
g14570 nand P2_R1312_U16 P2_R1312_U121 ; P2_R1312_U201
g14571 nand P2_R1312_U17 P2_R1312_U121 ; P2_R1312_U202
g14572 nand P2_R1312_U18 P2_R1312_U121 ; P2_R1312_U203
g14573 nand P2_R1312_U19 P2_R1312_U121 ; P2_R1312_U204
g14574 nand P2_U3085 P2_U3117 ; P2_R1312_U205
g14575 nand P2_U3085 P2_R1312_U22 ; P2_R1312_U206
g14576 nand P2_U3117 P2_R1312_U23 ; P2_R1312_U207
g14577 or P2_U3150 P2_U3117 ; P2_R1312_U208
g14578 nand P2_U3150 P2_R1312_U23 ; P2_R1312_U209
g14579 not P2_U3059 ; P2_R1335_U6
g14580 not P2_U3056 ; P2_R1335_U7
g14581 and P2_R1335_U10 P2_R1335_U9 ; P2_R1335_U8
g14582 nand P2_U3056 P2_R1335_U6 ; P2_R1335_U9
g14583 nand P2_U3059 P2_R1335_U7 ; P2_R1335_U10
g14584 and P2_R1209_U95 P2_R1209_U94 ; P2_R1209_U4
g14585 and P2_R1209_U96 P2_R1209_U97 ; P2_R1209_U5
g14586 and P2_R1209_U113 P2_R1209_U112 ; P2_R1209_U6
g14587 and P2_R1209_U155 P2_R1209_U154 ; P2_R1209_U7
g14588 and P2_R1209_U164 P2_R1209_U163 ; P2_R1209_U8
g14589 and P2_R1209_U182 P2_R1209_U181 ; P2_R1209_U9
g14590 and P2_R1209_U218 P2_R1209_U215 ; P2_R1209_U10
g14591 and P2_R1209_U211 P2_R1209_U208 ; P2_R1209_U11
g14592 and P2_R1209_U202 P2_R1209_U199 ; P2_R1209_U12
g14593 and P2_R1209_U196 P2_R1209_U192 ; P2_R1209_U13
g14594 and P2_R1209_U151 P2_R1209_U148 ; P2_R1209_U14
g14595 and P2_R1209_U143 P2_R1209_U140 ; P2_R1209_U15
g14596 and P2_R1209_U129 P2_R1209_U126 ; P2_R1209_U16
g14597 not P2_REG1_REG_6__SCAN_IN ; P2_R1209_U17
g14598 not P2_U3467 ; P2_R1209_U18
g14599 not P2_U3470 ; P2_R1209_U19
g14600 nand P2_U3467 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U20
g14601 not P2_REG1_REG_7__SCAN_IN ; P2_R1209_U21
g14602 not P2_REG1_REG_4__SCAN_IN ; P2_R1209_U22
g14603 not P2_U3461 ; P2_R1209_U23
g14604 not P2_U3464 ; P2_R1209_U24
g14605 not P2_REG1_REG_2__SCAN_IN ; P2_R1209_U25
g14606 not P2_U3455 ; P2_R1209_U26
g14607 not P2_REG1_REG_0__SCAN_IN ; P2_R1209_U27
g14608 not P2_U3446 ; P2_R1209_U28
g14609 nand P2_U3446 P2_REG1_REG_0__SCAN_IN ; P2_R1209_U29
g14610 not P2_REG1_REG_3__SCAN_IN ; P2_R1209_U30
g14611 not P2_U3458 ; P2_R1209_U31
g14612 nand P2_U3461 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U32
g14613 not P2_REG1_REG_5__SCAN_IN ; P2_R1209_U33
g14614 not P2_REG1_REG_8__SCAN_IN ; P2_R1209_U34
g14615 not P2_U3473 ; P2_R1209_U35
g14616 not P2_U3476 ; P2_R1209_U36
g14617 not P2_REG1_REG_9__SCAN_IN ; P2_R1209_U37
g14618 nand P2_R1209_U49 P2_R1209_U121 ; P2_R1209_U38
g14619 nand P2_R1209_U110 P2_R1209_U108 P2_R1209_U109 ; P2_R1209_U39
g14620 nand P2_R1209_U98 P2_R1209_U99 ; P2_R1209_U40
g14621 nand P2_U3452 P2_REG1_REG_1__SCAN_IN ; P2_R1209_U41
g14622 nand P2_R1209_U136 P2_R1209_U134 P2_R1209_U135 ; P2_R1209_U42
g14623 nand P2_R1209_U132 P2_R1209_U131 ; P2_R1209_U43
g14624 not P2_REG1_REG_16__SCAN_IN ; P2_R1209_U44
g14625 not P2_U3497 ; P2_R1209_U45
g14626 not P2_U3500 ; P2_R1209_U46
g14627 nand P2_U3497 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U47
g14628 not P2_REG1_REG_17__SCAN_IN ; P2_R1209_U48
g14629 nand P2_U3473 P2_REG1_REG_8__SCAN_IN ; P2_R1209_U49
g14630 not P2_REG1_REG_10__SCAN_IN ; P2_R1209_U50
g14631 not P2_U3479 ; P2_R1209_U51
g14632 not P2_REG1_REG_12__SCAN_IN ; P2_R1209_U52
g14633 not P2_U3485 ; P2_R1209_U53
g14634 not P2_REG1_REG_11__SCAN_IN ; P2_R1209_U54
g14635 not P2_U3482 ; P2_R1209_U55
g14636 nand P2_U3482 P2_REG1_REG_11__SCAN_IN ; P2_R1209_U56
g14637 not P2_REG1_REG_13__SCAN_IN ; P2_R1209_U57
g14638 not P2_U3488 ; P2_R1209_U58
g14639 not P2_REG1_REG_14__SCAN_IN ; P2_R1209_U59
g14640 not P2_U3491 ; P2_R1209_U60
g14641 not P2_REG1_REG_15__SCAN_IN ; P2_R1209_U61
g14642 not P2_U3494 ; P2_R1209_U62
g14643 not P2_REG1_REG_18__SCAN_IN ; P2_R1209_U63
g14644 not P2_U3503 ; P2_R1209_U64
g14645 nand P2_R1209_U186 P2_R1209_U185 P2_R1209_U187 ; P2_R1209_U65
g14646 nand P2_R1209_U179 P2_R1209_U178 ; P2_R1209_U66
g14647 nand P2_R1209_U56 P2_R1209_U204 ; P2_R1209_U67
g14648 nand P2_R1209_U259 P2_R1209_U258 ; P2_R1209_U68
g14649 nand P2_R1209_U308 P2_R1209_U307 ; P2_R1209_U69
g14650 nand P2_R1209_U231 P2_R1209_U230 ; P2_R1209_U70
g14651 nand P2_R1209_U236 P2_R1209_U235 ; P2_R1209_U71
g14652 nand P2_R1209_U243 P2_R1209_U242 ; P2_R1209_U72
g14653 nand P2_R1209_U250 P2_R1209_U249 ; P2_R1209_U73
g14654 nand P2_R1209_U255 P2_R1209_U254 ; P2_R1209_U74
g14655 nand P2_R1209_U271 P2_R1209_U270 ; P2_R1209_U75
g14656 nand P2_R1209_U278 P2_R1209_U277 ; P2_R1209_U76
g14657 nand P2_R1209_U285 P2_R1209_U284 ; P2_R1209_U77
g14658 nand P2_R1209_U292 P2_R1209_U291 ; P2_R1209_U78
g14659 nand P2_R1209_U299 P2_R1209_U298 ; P2_R1209_U79
g14660 nand P2_R1209_U304 P2_R1209_U303 ; P2_R1209_U80
g14661 nand P2_R1209_U117 P2_R1209_U116 P2_R1209_U118 ; P2_R1209_U81
g14662 nand P2_R1209_U133 P2_R1209_U145 ; P2_R1209_U82
g14663 nand P2_R1209_U41 P2_R1209_U152 ; P2_R1209_U83
g14664 not P2_U3445 ; P2_R1209_U84
g14665 not P2_REG1_REG_19__SCAN_IN ; P2_R1209_U85
g14666 nand P2_R1209_U175 P2_R1209_U174 ; P2_R1209_U86
g14667 nand P2_R1209_U171 P2_R1209_U170 ; P2_R1209_U87
g14668 nand P2_R1209_U161 P2_R1209_U160 ; P2_R1209_U88
g14669 not P2_R1209_U32 ; P2_R1209_U89
g14670 nand P2_U3476 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U90
g14671 nand P2_U3485 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U91
g14672 not P2_R1209_U56 ; P2_R1209_U92
g14673 not P2_R1209_U49 ; P2_R1209_U93
g14674 or P2_U3464 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U94
g14675 or P2_U3461 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U95
g14676 or P2_U3458 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U96
g14677 or P2_U3455 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U97
g14678 not P2_R1209_U29 ; P2_R1209_U98
g14679 or P2_U3452 P2_REG1_REG_1__SCAN_IN ; P2_R1209_U99
g14680 not P2_R1209_U40 ; P2_R1209_U100
g14681 not P2_R1209_U41 ; P2_R1209_U101
g14682 nand P2_R1209_U40 P2_R1209_U41 ; P2_R1209_U102
g14683 nand P2_U3455 P2_R1209_U96 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U103
g14684 nand P2_R1209_U5 P2_R1209_U102 ; P2_R1209_U104
g14685 nand P2_U3458 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U105
g14686 nand P2_R1209_U105 P2_R1209_U103 P2_R1209_U104 ; P2_R1209_U106
g14687 nand P2_R1209_U33 P2_R1209_U32 ; P2_R1209_U107
g14688 nand P2_U3464 P2_R1209_U107 ; P2_R1209_U108
g14689 nand P2_R1209_U4 P2_R1209_U106 ; P2_R1209_U109
g14690 nand P2_R1209_U89 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U110
g14691 not P2_R1209_U39 ; P2_R1209_U111
g14692 or P2_U3470 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U112
g14693 or P2_U3467 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U113
g14694 not P2_R1209_U20 ; P2_R1209_U114
g14695 nand P2_R1209_U21 P2_R1209_U20 ; P2_R1209_U115
g14696 nand P2_U3470 P2_R1209_U115 ; P2_R1209_U116
g14697 nand P2_R1209_U114 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U117
g14698 nand P2_R1209_U6 P2_R1209_U39 ; P2_R1209_U118
g14699 not P2_R1209_U81 ; P2_R1209_U119
g14700 or P2_U3473 P2_REG1_REG_8__SCAN_IN ; P2_R1209_U120
g14701 nand P2_R1209_U120 P2_R1209_U81 ; P2_R1209_U121
g14702 not P2_R1209_U38 ; P2_R1209_U122
g14703 or P2_U3476 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U123
g14704 or P2_U3467 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U124
g14705 nand P2_R1209_U124 P2_R1209_U39 ; P2_R1209_U125
g14706 nand P2_R1209_U238 P2_R1209_U237 P2_R1209_U20 P2_R1209_U125 ; P2_R1209_U126
g14707 nand P2_R1209_U111 P2_R1209_U20 ; P2_R1209_U127
g14708 nand P2_U3470 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U128
g14709 nand P2_R1209_U128 P2_R1209_U6 P2_R1209_U127 ; P2_R1209_U129
g14710 or P2_U3467 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U130
g14711 nand P2_R1209_U101 P2_R1209_U97 ; P2_R1209_U131
g14712 nand P2_U3455 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U132
g14713 not P2_R1209_U43 ; P2_R1209_U133
g14714 nand P2_R1209_U100 P2_R1209_U5 ; P2_R1209_U134
g14715 nand P2_R1209_U43 P2_R1209_U96 ; P2_R1209_U135
g14716 nand P2_U3458 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U136
g14717 not P2_R1209_U42 ; P2_R1209_U137
g14718 or P2_U3461 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U138
g14719 nand P2_R1209_U138 P2_R1209_U42 ; P2_R1209_U139
g14720 nand P2_R1209_U245 P2_R1209_U244 P2_R1209_U32 P2_R1209_U139 ; P2_R1209_U140
g14721 nand P2_R1209_U137 P2_R1209_U32 ; P2_R1209_U141
g14722 nand P2_U3464 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U142
g14723 nand P2_R1209_U142 P2_R1209_U4 P2_R1209_U141 ; P2_R1209_U143
g14724 or P2_U3461 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U144
g14725 nand P2_R1209_U100 P2_R1209_U97 ; P2_R1209_U145
g14726 not P2_R1209_U82 ; P2_R1209_U146
g14727 nand P2_U3458 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U147
g14728 nand P2_R1209_U257 P2_R1209_U256 P2_R1209_U41 P2_R1209_U40 ; P2_R1209_U148
g14729 nand P2_R1209_U41 P2_R1209_U40 ; P2_R1209_U149
g14730 nand P2_U3455 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U150
g14731 nand P2_R1209_U150 P2_R1209_U97 P2_R1209_U149 ; P2_R1209_U151
g14732 or P2_U3452 P2_REG1_REG_1__SCAN_IN ; P2_R1209_U152
g14733 not P2_R1209_U83 ; P2_R1209_U153
g14734 or P2_U3476 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U154
g14735 or P2_U3479 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U155
g14736 nand P2_R1209_U93 P2_R1209_U7 ; P2_R1209_U156
g14737 nand P2_U3479 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U157
g14738 nand P2_R1209_U157 P2_R1209_U90 P2_R1209_U156 ; P2_R1209_U158
g14739 or P2_U3479 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U159
g14740 nand P2_R1209_U120 P2_R1209_U7 P2_R1209_U81 ; P2_R1209_U160
g14741 nand P2_R1209_U159 P2_R1209_U158 ; P2_R1209_U161
g14742 not P2_R1209_U88 ; P2_R1209_U162
g14743 or P2_U3488 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U163
g14744 or P2_U3485 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U164
g14745 nand P2_R1209_U92 P2_R1209_U8 ; P2_R1209_U165
g14746 nand P2_U3488 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U166
g14747 nand P2_R1209_U166 P2_R1209_U91 P2_R1209_U165 ; P2_R1209_U167
g14748 or P2_U3482 P2_REG1_REG_11__SCAN_IN ; P2_R1209_U168
g14749 or P2_U3488 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U169
g14750 nand P2_R1209_U168 P2_R1209_U8 P2_R1209_U88 ; P2_R1209_U170
g14751 nand P2_R1209_U169 P2_R1209_U167 ; P2_R1209_U171
g14752 not P2_R1209_U87 ; P2_R1209_U172
g14753 or P2_U3491 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U173
g14754 nand P2_R1209_U173 P2_R1209_U87 ; P2_R1209_U174
g14755 nand P2_U3491 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U175
g14756 not P2_R1209_U86 ; P2_R1209_U176
g14757 or P2_U3494 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U177
g14758 nand P2_R1209_U177 P2_R1209_U86 ; P2_R1209_U178
g14759 nand P2_U3494 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U179
g14760 not P2_R1209_U66 ; P2_R1209_U180
g14761 or P2_U3500 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U181
g14762 or P2_U3497 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U182
g14763 not P2_R1209_U47 ; P2_R1209_U183
g14764 nand P2_R1209_U48 P2_R1209_U47 ; P2_R1209_U184
g14765 nand P2_U3500 P2_R1209_U184 ; P2_R1209_U185
g14766 nand P2_R1209_U183 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U186
g14767 nand P2_R1209_U9 P2_R1209_U66 ; P2_R1209_U187
g14768 not P2_R1209_U65 ; P2_R1209_U188
g14769 or P2_U3503 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U189
g14770 nand P2_R1209_U189 P2_R1209_U65 ; P2_R1209_U190
g14771 nand P2_U3503 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U191
g14772 nand P2_R1209_U261 P2_R1209_U260 P2_R1209_U191 P2_R1209_U190 ; P2_R1209_U192
g14773 nand P2_U3503 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U193
g14774 nand P2_R1209_U188 P2_R1209_U193 ; P2_R1209_U194
g14775 or P2_U3503 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U195
g14776 nand P2_R1209_U195 P2_R1209_U264 P2_R1209_U194 ; P2_R1209_U196
g14777 or P2_U3497 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U197
g14778 nand P2_R1209_U197 P2_R1209_U66 ; P2_R1209_U198
g14779 nand P2_R1209_U273 P2_R1209_U272 P2_R1209_U47 P2_R1209_U198 ; P2_R1209_U199
g14780 nand P2_R1209_U180 P2_R1209_U47 ; P2_R1209_U200
g14781 nand P2_U3500 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U201
g14782 nand P2_R1209_U201 P2_R1209_U9 P2_R1209_U200 ; P2_R1209_U202
g14783 or P2_U3497 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U203
g14784 nand P2_R1209_U168 P2_R1209_U88 ; P2_R1209_U204
g14785 not P2_R1209_U67 ; P2_R1209_U205
g14786 or P2_U3485 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U206
g14787 nand P2_R1209_U206 P2_R1209_U67 ; P2_R1209_U207
g14788 nand P2_R1209_U294 P2_R1209_U293 P2_R1209_U91 P2_R1209_U207 ; P2_R1209_U208
g14789 nand P2_R1209_U205 P2_R1209_U91 ; P2_R1209_U209
g14790 nand P2_U3488 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U210
g14791 nand P2_R1209_U210 P2_R1209_U8 P2_R1209_U209 ; P2_R1209_U211
g14792 or P2_U3485 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U212
g14793 or P2_U3476 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U213
g14794 nand P2_R1209_U213 P2_R1209_U38 ; P2_R1209_U214
g14795 nand P2_R1209_U306 P2_R1209_U305 P2_R1209_U90 P2_R1209_U214 ; P2_R1209_U215
g14796 nand P2_R1209_U122 P2_R1209_U90 ; P2_R1209_U216
g14797 nand P2_U3479 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U217
g14798 nand P2_R1209_U217 P2_R1209_U7 P2_R1209_U216 ; P2_R1209_U218
g14799 nand P2_R1209_U123 P2_R1209_U90 ; P2_R1209_U219
g14800 nand P2_R1209_U120 P2_R1209_U49 ; P2_R1209_U220
g14801 nand P2_R1209_U130 P2_R1209_U20 ; P2_R1209_U221
g14802 nand P2_R1209_U144 P2_R1209_U32 ; P2_R1209_U222
g14803 nand P2_R1209_U147 P2_R1209_U96 ; P2_R1209_U223
g14804 nand P2_R1209_U203 P2_R1209_U47 ; P2_R1209_U224
g14805 nand P2_R1209_U212 P2_R1209_U91 ; P2_R1209_U225
g14806 nand P2_R1209_U168 P2_R1209_U56 ; P2_R1209_U226
g14807 nand P2_U3476 P2_R1209_U37 ; P2_R1209_U227
g14808 nand P2_R1209_U36 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U228
g14809 nand P2_R1209_U228 P2_R1209_U227 ; P2_R1209_U229
g14810 nand P2_R1209_U219 P2_R1209_U38 ; P2_R1209_U230
g14811 nand P2_R1209_U229 P2_R1209_U122 ; P2_R1209_U231
g14812 nand P2_U3473 P2_R1209_U34 ; P2_R1209_U232
g14813 nand P2_R1209_U35 P2_REG1_REG_8__SCAN_IN ; P2_R1209_U233
g14814 nand P2_R1209_U233 P2_R1209_U232 ; P2_R1209_U234
g14815 nand P2_R1209_U220 P2_R1209_U81 ; P2_R1209_U235
g14816 nand P2_R1209_U119 P2_R1209_U234 ; P2_R1209_U236
g14817 nand P2_U3470 P2_R1209_U21 ; P2_R1209_U237
g14818 nand P2_R1209_U19 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U238
g14819 nand P2_U3467 P2_R1209_U17 ; P2_R1209_U239
g14820 nand P2_R1209_U18 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U240
g14821 nand P2_R1209_U240 P2_R1209_U239 ; P2_R1209_U241
g14822 nand P2_R1209_U221 P2_R1209_U39 ; P2_R1209_U242
g14823 nand P2_R1209_U241 P2_R1209_U111 ; P2_R1209_U243
g14824 nand P2_U3464 P2_R1209_U33 ; P2_R1209_U244
g14825 nand P2_R1209_U24 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U245
g14826 nand P2_U3461 P2_R1209_U22 ; P2_R1209_U246
g14827 nand P2_R1209_U23 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U247
g14828 nand P2_R1209_U247 P2_R1209_U246 ; P2_R1209_U248
g14829 nand P2_R1209_U222 P2_R1209_U42 ; P2_R1209_U249
g14830 nand P2_R1209_U248 P2_R1209_U137 ; P2_R1209_U250
g14831 nand P2_U3458 P2_R1209_U30 ; P2_R1209_U251
g14832 nand P2_R1209_U31 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U252
g14833 nand P2_R1209_U252 P2_R1209_U251 ; P2_R1209_U253
g14834 nand P2_R1209_U223 P2_R1209_U82 ; P2_R1209_U254
g14835 nand P2_R1209_U146 P2_R1209_U253 ; P2_R1209_U255
g14836 nand P2_U3455 P2_R1209_U25 ; P2_R1209_U256
g14837 nand P2_R1209_U26 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U257
g14838 nand P2_R1209_U98 P2_R1209_U83 ; P2_R1209_U258
g14839 nand P2_R1209_U153 P2_R1209_U29 ; P2_R1209_U259
g14840 nand P2_U3445 P2_R1209_U85 ; P2_R1209_U260
g14841 nand P2_R1209_U84 P2_REG1_REG_19__SCAN_IN ; P2_R1209_U261
g14842 nand P2_U3445 P2_R1209_U85 ; P2_R1209_U262
g14843 nand P2_R1209_U84 P2_REG1_REG_19__SCAN_IN ; P2_R1209_U263
g14844 nand P2_R1209_U263 P2_R1209_U262 ; P2_R1209_U264
g14845 nand P2_U3503 P2_R1209_U63 ; P2_R1209_U265
g14846 nand P2_R1209_U64 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U266
g14847 nand P2_U3503 P2_R1209_U63 ; P2_R1209_U267
g14848 nand P2_R1209_U64 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U268
g14849 nand P2_R1209_U268 P2_R1209_U267 ; P2_R1209_U269
g14850 nand P2_R1209_U266 P2_R1209_U265 P2_R1209_U65 ; P2_R1209_U270
g14851 nand P2_R1209_U269 P2_R1209_U188 ; P2_R1209_U271
g14852 nand P2_U3500 P2_R1209_U48 ; P2_R1209_U272
g14853 nand P2_R1209_U46 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U273
g14854 nand P2_U3497 P2_R1209_U44 ; P2_R1209_U274
g14855 nand P2_R1209_U45 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U275
g14856 nand P2_R1209_U275 P2_R1209_U274 ; P2_R1209_U276
g14857 nand P2_R1209_U224 P2_R1209_U66 ; P2_R1209_U277
g14858 nand P2_R1209_U276 P2_R1209_U180 ; P2_R1209_U278
g14859 nand P2_U3494 P2_R1209_U61 ; P2_R1209_U279
g14860 nand P2_R1209_U62 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U280
g14861 nand P2_U3494 P2_R1209_U61 ; P2_R1209_U281
g14862 nand P2_R1209_U62 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U282
g14863 nand P2_R1209_U282 P2_R1209_U281 ; P2_R1209_U283
g14864 nand P2_R1209_U280 P2_R1209_U279 P2_R1209_U86 ; P2_R1209_U284
g14865 nand P2_R1209_U176 P2_R1209_U283 ; P2_R1209_U285
g14866 nand P2_U3491 P2_R1209_U59 ; P2_R1209_U286
g14867 nand P2_R1209_U60 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U287
g14868 nand P2_U3491 P2_R1209_U59 ; P2_R1209_U288
g14869 nand P2_R1209_U60 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U289
g14870 nand P2_R1209_U289 P2_R1209_U288 ; P2_R1209_U290
g14871 nand P2_R1209_U287 P2_R1209_U286 P2_R1209_U87 ; P2_R1209_U291
g14872 nand P2_R1209_U172 P2_R1209_U290 ; P2_R1209_U292
g14873 nand P2_U3488 P2_R1209_U57 ; P2_R1209_U293
g14874 nand P2_R1209_U58 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U294
g14875 nand P2_U3485 P2_R1209_U52 ; P2_R1209_U295
g14876 nand P2_R1209_U53 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U296
g14877 nand P2_R1209_U296 P2_R1209_U295 ; P2_R1209_U297
g14878 nand P2_R1209_U225 P2_R1209_U67 ; P2_R1209_U298
g14879 nand P2_R1209_U297 P2_R1209_U205 ; P2_R1209_U299
g14880 nand P2_U3482 P2_R1209_U54 ; P2_R1209_U300
g14881 nand P2_R1209_U55 P2_REG1_REG_11__SCAN_IN ; P2_R1209_U301
g14882 nand P2_R1209_U301 P2_R1209_U300 ; P2_R1209_U302
g14883 nand P2_R1209_U226 P2_R1209_U88 ; P2_R1209_U303
g14884 nand P2_R1209_U162 P2_R1209_U302 ; P2_R1209_U304
g14885 nand P2_U3479 P2_R1209_U50 ; P2_R1209_U305
g14886 nand P2_R1209_U51 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U306
g14887 nand P2_U3446 P2_R1209_U27 ; P2_R1209_U307
g14888 nand P2_R1209_U28 P2_REG1_REG_0__SCAN_IN ; P2_R1209_U308
g14889 and P2_R1170_U95 P2_R1170_U94 ; P2_R1170_U4
g14890 and P2_R1170_U96 P2_R1170_U97 ; P2_R1170_U5
g14891 and P2_R1170_U113 P2_R1170_U112 ; P2_R1170_U6
g14892 and P2_R1170_U155 P2_R1170_U154 ; P2_R1170_U7
g14893 and P2_R1170_U164 P2_R1170_U163 ; P2_R1170_U8
g14894 and P2_R1170_U182 P2_R1170_U181 ; P2_R1170_U9
g14895 and P2_R1170_U218 P2_R1170_U215 ; P2_R1170_U10
g14896 and P2_R1170_U211 P2_R1170_U208 ; P2_R1170_U11
g14897 and P2_R1170_U202 P2_R1170_U199 ; P2_R1170_U12
g14898 and P2_R1170_U196 P2_R1170_U192 ; P2_R1170_U13
g14899 and P2_R1170_U151 P2_R1170_U148 ; P2_R1170_U14
g14900 and P2_R1170_U143 P2_R1170_U140 ; P2_R1170_U15
g14901 and P2_R1170_U129 P2_R1170_U126 ; P2_R1170_U16
g14902 not P2_REG2_REG_6__SCAN_IN ; P2_R1170_U17
g14903 not P2_U3467 ; P2_R1170_U18
g14904 not P2_U3470 ; P2_R1170_U19
g14905 nand P2_U3467 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U20
g14906 not P2_REG2_REG_7__SCAN_IN ; P2_R1170_U21
g14907 not P2_REG2_REG_4__SCAN_IN ; P2_R1170_U22
g14908 not P2_U3461 ; P2_R1170_U23
g14909 not P2_U3464 ; P2_R1170_U24
g14910 not P2_REG2_REG_2__SCAN_IN ; P2_R1170_U25
g14911 not P2_U3455 ; P2_R1170_U26
g14912 not P2_REG2_REG_0__SCAN_IN ; P2_R1170_U27
g14913 not P2_U3446 ; P2_R1170_U28
g14914 nand P2_U3446 P2_REG2_REG_0__SCAN_IN ; P2_R1170_U29
g14915 not P2_REG2_REG_3__SCAN_IN ; P2_R1170_U30
g14916 not P2_U3458 ; P2_R1170_U31
g14917 nand P2_U3461 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U32
g14918 not P2_REG2_REG_5__SCAN_IN ; P2_R1170_U33
g14919 not P2_REG2_REG_8__SCAN_IN ; P2_R1170_U34
g14920 not P2_U3473 ; P2_R1170_U35
g14921 not P2_U3476 ; P2_R1170_U36
g14922 not P2_REG2_REG_9__SCAN_IN ; P2_R1170_U37
g14923 nand P2_R1170_U49 P2_R1170_U121 ; P2_R1170_U38
g14924 nand P2_R1170_U110 P2_R1170_U108 P2_R1170_U109 ; P2_R1170_U39
g14925 nand P2_R1170_U98 P2_R1170_U99 ; P2_R1170_U40
g14926 nand P2_U3452 P2_REG2_REG_1__SCAN_IN ; P2_R1170_U41
g14927 nand P2_R1170_U136 P2_R1170_U134 P2_R1170_U135 ; P2_R1170_U42
g14928 nand P2_R1170_U132 P2_R1170_U131 ; P2_R1170_U43
g14929 not P2_REG2_REG_16__SCAN_IN ; P2_R1170_U44
g14930 not P2_U3497 ; P2_R1170_U45
g14931 not P2_U3500 ; P2_R1170_U46
g14932 nand P2_U3497 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U47
g14933 not P2_REG2_REG_17__SCAN_IN ; P2_R1170_U48
g14934 nand P2_U3473 P2_REG2_REG_8__SCAN_IN ; P2_R1170_U49
g14935 not P2_REG2_REG_10__SCAN_IN ; P2_R1170_U50
g14936 not P2_U3479 ; P2_R1170_U51
g14937 not P2_REG2_REG_12__SCAN_IN ; P2_R1170_U52
g14938 not P2_U3485 ; P2_R1170_U53
g14939 not P2_REG2_REG_11__SCAN_IN ; P2_R1170_U54
g14940 not P2_U3482 ; P2_R1170_U55
g14941 nand P2_U3482 P2_REG2_REG_11__SCAN_IN ; P2_R1170_U56
g14942 not P2_REG2_REG_13__SCAN_IN ; P2_R1170_U57
g14943 not P2_U3488 ; P2_R1170_U58
g14944 not P2_REG2_REG_14__SCAN_IN ; P2_R1170_U59
g14945 not P2_U3491 ; P2_R1170_U60
g14946 not P2_REG2_REG_15__SCAN_IN ; P2_R1170_U61
g14947 not P2_U3494 ; P2_R1170_U62
g14948 not P2_REG2_REG_18__SCAN_IN ; P2_R1170_U63
g14949 not P2_U3503 ; P2_R1170_U64
g14950 nand P2_R1170_U186 P2_R1170_U185 P2_R1170_U187 ; P2_R1170_U65
g14951 nand P2_R1170_U179 P2_R1170_U178 ; P2_R1170_U66
g14952 nand P2_R1170_U56 P2_R1170_U204 ; P2_R1170_U67
g14953 nand P2_R1170_U259 P2_R1170_U258 ; P2_R1170_U68
g14954 nand P2_R1170_U308 P2_R1170_U307 ; P2_R1170_U69
g14955 nand P2_R1170_U231 P2_R1170_U230 ; P2_R1170_U70
g14956 nand P2_R1170_U236 P2_R1170_U235 ; P2_R1170_U71
g14957 nand P2_R1170_U243 P2_R1170_U242 ; P2_R1170_U72
g14958 nand P2_R1170_U250 P2_R1170_U249 ; P2_R1170_U73
g14959 nand P2_R1170_U255 P2_R1170_U254 ; P2_R1170_U74
g14960 nand P2_R1170_U271 P2_R1170_U270 ; P2_R1170_U75
g14961 nand P2_R1170_U278 P2_R1170_U277 ; P2_R1170_U76
g14962 nand P2_R1170_U285 P2_R1170_U284 ; P2_R1170_U77
g14963 nand P2_R1170_U292 P2_R1170_U291 ; P2_R1170_U78
g14964 nand P2_R1170_U299 P2_R1170_U298 ; P2_R1170_U79
g14965 nand P2_R1170_U304 P2_R1170_U303 ; P2_R1170_U80
g14966 nand P2_R1170_U117 P2_R1170_U116 P2_R1170_U118 ; P2_R1170_U81
g14967 nand P2_R1170_U133 P2_R1170_U145 ; P2_R1170_U82
g14968 nand P2_R1170_U41 P2_R1170_U152 ; P2_R1170_U83
g14969 not P2_U3445 ; P2_R1170_U84
g14970 not P2_REG2_REG_19__SCAN_IN ; P2_R1170_U85
g14971 nand P2_R1170_U175 P2_R1170_U174 ; P2_R1170_U86
g14972 nand P2_R1170_U171 P2_R1170_U170 ; P2_R1170_U87
g14973 nand P2_R1170_U161 P2_R1170_U160 ; P2_R1170_U88
g14974 not P2_R1170_U32 ; P2_R1170_U89
g14975 nand P2_U3476 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U90
g14976 nand P2_U3485 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U91
g14977 not P2_R1170_U56 ; P2_R1170_U92
g14978 not P2_R1170_U49 ; P2_R1170_U93
g14979 or P2_U3464 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U94
g14980 or P2_U3461 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U95
g14981 or P2_U3458 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U96
g14982 or P2_U3455 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U97
g14983 not P2_R1170_U29 ; P2_R1170_U98
g14984 or P2_U3452 P2_REG2_REG_1__SCAN_IN ; P2_R1170_U99
g14985 not P2_R1170_U40 ; P2_R1170_U100
g14986 not P2_R1170_U41 ; P2_R1170_U101
g14987 nand P2_R1170_U40 P2_R1170_U41 ; P2_R1170_U102
g14988 nand P2_U3455 P2_R1170_U96 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U103
g14989 nand P2_R1170_U5 P2_R1170_U102 ; P2_R1170_U104
g14990 nand P2_U3458 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U105
g14991 nand P2_R1170_U105 P2_R1170_U103 P2_R1170_U104 ; P2_R1170_U106
g14992 nand P2_R1170_U33 P2_R1170_U32 ; P2_R1170_U107
g14993 nand P2_U3464 P2_R1170_U107 ; P2_R1170_U108
g14994 nand P2_R1170_U4 P2_R1170_U106 ; P2_R1170_U109
g14995 nand P2_R1170_U89 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U110
g14996 not P2_R1170_U39 ; P2_R1170_U111
g14997 or P2_U3470 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U112
g14998 or P2_U3467 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U113
g14999 not P2_R1170_U20 ; P2_R1170_U114
g15000 nand P2_R1170_U21 P2_R1170_U20 ; P2_R1170_U115
g15001 nand P2_U3470 P2_R1170_U115 ; P2_R1170_U116
g15002 nand P2_R1170_U114 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U117
g15003 nand P2_R1170_U6 P2_R1170_U39 ; P2_R1170_U118
g15004 not P2_R1170_U81 ; P2_R1170_U119
g15005 or P2_U3473 P2_REG2_REG_8__SCAN_IN ; P2_R1170_U120
g15006 nand P2_R1170_U120 P2_R1170_U81 ; P2_R1170_U121
g15007 not P2_R1170_U38 ; P2_R1170_U122
g15008 or P2_U3476 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U123
g15009 or P2_U3467 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U124
g15010 nand P2_R1170_U124 P2_R1170_U39 ; P2_R1170_U125
g15011 nand P2_R1170_U238 P2_R1170_U237 P2_R1170_U20 P2_R1170_U125 ; P2_R1170_U126
g15012 nand P2_R1170_U111 P2_R1170_U20 ; P2_R1170_U127
g15013 nand P2_U3470 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U128
g15014 nand P2_R1170_U128 P2_R1170_U6 P2_R1170_U127 ; P2_R1170_U129
g15015 or P2_U3467 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U130
g15016 nand P2_R1170_U101 P2_R1170_U97 ; P2_R1170_U131
g15017 nand P2_U3455 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U132
g15018 not P2_R1170_U43 ; P2_R1170_U133
g15019 nand P2_R1170_U100 P2_R1170_U5 ; P2_R1170_U134
g15020 nand P2_R1170_U43 P2_R1170_U96 ; P2_R1170_U135
g15021 nand P2_U3458 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U136
g15022 not P2_R1170_U42 ; P2_R1170_U137
g15023 or P2_U3461 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U138
g15024 nand P2_R1170_U138 P2_R1170_U42 ; P2_R1170_U139
g15025 nand P2_R1170_U245 P2_R1170_U244 P2_R1170_U32 P2_R1170_U139 ; P2_R1170_U140
g15026 nand P2_R1170_U137 P2_R1170_U32 ; P2_R1170_U141
g15027 nand P2_U3464 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U142
g15028 nand P2_R1170_U142 P2_R1170_U4 P2_R1170_U141 ; P2_R1170_U143
g15029 or P2_U3461 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U144
g15030 nand P2_R1170_U100 P2_R1170_U97 ; P2_R1170_U145
g15031 not P2_R1170_U82 ; P2_R1170_U146
g15032 nand P2_U3458 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U147
g15033 nand P2_R1170_U257 P2_R1170_U256 P2_R1170_U41 P2_R1170_U40 ; P2_R1170_U148
g15034 nand P2_R1170_U41 P2_R1170_U40 ; P2_R1170_U149
g15035 nand P2_U3455 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U150
g15036 nand P2_R1170_U150 P2_R1170_U97 P2_R1170_U149 ; P2_R1170_U151
g15037 or P2_U3452 P2_REG2_REG_1__SCAN_IN ; P2_R1170_U152
g15038 not P2_R1170_U83 ; P2_R1170_U153
g15039 or P2_U3476 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U154
g15040 or P2_U3479 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U155
g15041 nand P2_R1170_U93 P2_R1170_U7 ; P2_R1170_U156
g15042 nand P2_U3479 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U157
g15043 nand P2_R1170_U157 P2_R1170_U90 P2_R1170_U156 ; P2_R1170_U158
g15044 or P2_U3479 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U159
g15045 nand P2_R1170_U120 P2_R1170_U7 P2_R1170_U81 ; P2_R1170_U160
g15046 nand P2_R1170_U159 P2_R1170_U158 ; P2_R1170_U161
g15047 not P2_R1170_U88 ; P2_R1170_U162
g15048 or P2_U3488 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U163
g15049 or P2_U3485 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U164
g15050 nand P2_R1170_U92 P2_R1170_U8 ; P2_R1170_U165
g15051 nand P2_U3488 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U166
g15052 nand P2_R1170_U166 P2_R1170_U91 P2_R1170_U165 ; P2_R1170_U167
g15053 or P2_U3482 P2_REG2_REG_11__SCAN_IN ; P2_R1170_U168
g15054 or P2_U3488 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U169
g15055 nand P2_R1170_U168 P2_R1170_U8 P2_R1170_U88 ; P2_R1170_U170
g15056 nand P2_R1170_U169 P2_R1170_U167 ; P2_R1170_U171
g15057 not P2_R1170_U87 ; P2_R1170_U172
g15058 or P2_U3491 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U173
g15059 nand P2_R1170_U173 P2_R1170_U87 ; P2_R1170_U174
g15060 nand P2_U3491 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U175
g15061 not P2_R1170_U86 ; P2_R1170_U176
g15062 or P2_U3494 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U177
g15063 nand P2_R1170_U177 P2_R1170_U86 ; P2_R1170_U178
g15064 nand P2_U3494 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U179
g15065 not P2_R1170_U66 ; P2_R1170_U180
g15066 or P2_U3500 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U181
g15067 or P2_U3497 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U182
g15068 not P2_R1170_U47 ; P2_R1170_U183
g15069 nand P2_R1170_U48 P2_R1170_U47 ; P2_R1170_U184
g15070 nand P2_U3500 P2_R1170_U184 ; P2_R1170_U185
g15071 nand P2_R1170_U183 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U186
g15072 nand P2_R1170_U9 P2_R1170_U66 ; P2_R1170_U187
g15073 not P2_R1170_U65 ; P2_R1170_U188
g15074 or P2_U3503 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U189
g15075 nand P2_R1170_U189 P2_R1170_U65 ; P2_R1170_U190
g15076 nand P2_U3503 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U191
g15077 nand P2_R1170_U261 P2_R1170_U260 P2_R1170_U191 P2_R1170_U190 ; P2_R1170_U192
g15078 nand P2_U3503 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U193
g15079 nand P2_R1170_U188 P2_R1170_U193 ; P2_R1170_U194
g15080 or P2_U3503 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U195
g15081 nand P2_R1170_U195 P2_R1170_U264 P2_R1170_U194 ; P2_R1170_U196
g15082 or P2_U3497 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U197
g15083 nand P2_R1170_U197 P2_R1170_U66 ; P2_R1170_U198
g15084 nand P2_R1170_U273 P2_R1170_U272 P2_R1170_U47 P2_R1170_U198 ; P2_R1170_U199
g15085 nand P2_R1170_U180 P2_R1170_U47 ; P2_R1170_U200
g15086 nand P2_U3500 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U201
g15087 nand P2_R1170_U201 P2_R1170_U9 P2_R1170_U200 ; P2_R1170_U202
g15088 or P2_U3497 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U203
g15089 nand P2_R1170_U168 P2_R1170_U88 ; P2_R1170_U204
g15090 not P2_R1170_U67 ; P2_R1170_U205
g15091 or P2_U3485 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U206
g15092 nand P2_R1170_U206 P2_R1170_U67 ; P2_R1170_U207
g15093 nand P2_R1170_U294 P2_R1170_U293 P2_R1170_U91 P2_R1170_U207 ; P2_R1170_U208
g15094 nand P2_R1170_U205 P2_R1170_U91 ; P2_R1170_U209
g15095 nand P2_U3488 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U210
g15096 nand P2_R1170_U210 P2_R1170_U8 P2_R1170_U209 ; P2_R1170_U211
g15097 or P2_U3485 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U212
g15098 or P2_U3476 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U213
g15099 nand P2_R1170_U213 P2_R1170_U38 ; P2_R1170_U214
g15100 nand P2_R1170_U306 P2_R1170_U305 P2_R1170_U90 P2_R1170_U214 ; P2_R1170_U215
g15101 nand P2_R1170_U122 P2_R1170_U90 ; P2_R1170_U216
g15102 nand P2_U3479 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U217
g15103 nand P2_R1170_U217 P2_R1170_U7 P2_R1170_U216 ; P2_R1170_U218
g15104 nand P2_R1170_U123 P2_R1170_U90 ; P2_R1170_U219
g15105 nand P2_R1170_U120 P2_R1170_U49 ; P2_R1170_U220
g15106 nand P2_R1170_U130 P2_R1170_U20 ; P2_R1170_U221
g15107 nand P2_R1170_U144 P2_R1170_U32 ; P2_R1170_U222
g15108 nand P2_R1170_U147 P2_R1170_U96 ; P2_R1170_U223
g15109 nand P2_R1170_U203 P2_R1170_U47 ; P2_R1170_U224
g15110 nand P2_R1170_U212 P2_R1170_U91 ; P2_R1170_U225
g15111 nand P2_R1170_U168 P2_R1170_U56 ; P2_R1170_U226
g15112 nand P2_U3476 P2_R1170_U37 ; P2_R1170_U227
g15113 nand P2_R1170_U36 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U228
g15114 nand P2_R1170_U228 P2_R1170_U227 ; P2_R1170_U229
g15115 nand P2_R1170_U219 P2_R1170_U38 ; P2_R1170_U230
g15116 nand P2_R1170_U229 P2_R1170_U122 ; P2_R1170_U231
g15117 nand P2_U3473 P2_R1170_U34 ; P2_R1170_U232
g15118 nand P2_R1170_U35 P2_REG2_REG_8__SCAN_IN ; P2_R1170_U233
g15119 nand P2_R1170_U233 P2_R1170_U232 ; P2_R1170_U234
g15120 nand P2_R1170_U220 P2_R1170_U81 ; P2_R1170_U235
g15121 nand P2_R1170_U119 P2_R1170_U234 ; P2_R1170_U236
g15122 nand P2_U3470 P2_R1170_U21 ; P2_R1170_U237
g15123 nand P2_R1170_U19 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U238
g15124 nand P2_U3467 P2_R1170_U17 ; P2_R1170_U239
g15125 nand P2_R1170_U18 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U240
g15126 nand P2_R1170_U240 P2_R1170_U239 ; P2_R1170_U241
g15127 nand P2_R1170_U221 P2_R1170_U39 ; P2_R1170_U242
g15128 nand P2_R1170_U241 P2_R1170_U111 ; P2_R1170_U243
g15129 nand P2_U3464 P2_R1170_U33 ; P2_R1170_U244
g15130 nand P2_R1170_U24 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U245
g15131 nand P2_U3461 P2_R1170_U22 ; P2_R1170_U246
g15132 nand P2_R1170_U23 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U247
g15133 nand P2_R1170_U247 P2_R1170_U246 ; P2_R1170_U248
g15134 nand P2_R1170_U222 P2_R1170_U42 ; P2_R1170_U249
g15135 nand P2_R1170_U248 P2_R1170_U137 ; P2_R1170_U250
g15136 nand P2_U3458 P2_R1170_U30 ; P2_R1170_U251
g15137 nand P2_R1170_U31 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U252
g15138 nand P2_R1170_U252 P2_R1170_U251 ; P2_R1170_U253
g15139 nand P2_R1170_U223 P2_R1170_U82 ; P2_R1170_U254
g15140 nand P2_R1170_U146 P2_R1170_U253 ; P2_R1170_U255
g15141 nand P2_U3455 P2_R1170_U25 ; P2_R1170_U256
g15142 nand P2_R1170_U26 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U257
g15143 nand P2_R1170_U98 P2_R1170_U83 ; P2_R1170_U258
g15144 nand P2_R1170_U153 P2_R1170_U29 ; P2_R1170_U259
g15145 nand P2_U3445 P2_R1170_U85 ; P2_R1170_U260
g15146 nand P2_R1170_U84 P2_REG2_REG_19__SCAN_IN ; P2_R1170_U261
g15147 nand P2_U3445 P2_R1170_U85 ; P2_R1170_U262
g15148 nand P2_R1170_U84 P2_REG2_REG_19__SCAN_IN ; P2_R1170_U263
g15149 nand P2_R1170_U263 P2_R1170_U262 ; P2_R1170_U264
g15150 nand P2_U3503 P2_R1170_U63 ; P2_R1170_U265
g15151 nand P2_R1170_U64 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U266
g15152 nand P2_U3503 P2_R1170_U63 ; P2_R1170_U267
g15153 nand P2_R1170_U64 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U268
g15154 nand P2_R1170_U268 P2_R1170_U267 ; P2_R1170_U269
g15155 nand P2_R1170_U266 P2_R1170_U265 P2_R1170_U65 ; P2_R1170_U270
g15156 nand P2_R1170_U269 P2_R1170_U188 ; P2_R1170_U271
g15157 nand P2_U3500 P2_R1170_U48 ; P2_R1170_U272
g15158 nand P2_R1170_U46 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U273
g15159 nand P2_U3497 P2_R1170_U44 ; P2_R1170_U274
g15160 nand P2_R1170_U45 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U275
g15161 nand P2_R1170_U275 P2_R1170_U274 ; P2_R1170_U276
g15162 nand P2_R1170_U224 P2_R1170_U66 ; P2_R1170_U277
g15163 nand P2_R1170_U276 P2_R1170_U180 ; P2_R1170_U278
g15164 nand P2_U3494 P2_R1170_U61 ; P2_R1170_U279
g15165 nand P2_R1170_U62 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U280
g15166 nand P2_U3494 P2_R1170_U61 ; P2_R1170_U281
g15167 nand P2_R1170_U62 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U282
g15168 nand P2_R1170_U282 P2_R1170_U281 ; P2_R1170_U283
g15169 nand P2_R1170_U280 P2_R1170_U279 P2_R1170_U86 ; P2_R1170_U284
g15170 nand P2_R1170_U176 P2_R1170_U283 ; P2_R1170_U285
g15171 nand P2_U3491 P2_R1170_U59 ; P2_R1170_U286
g15172 nand P2_R1170_U60 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U287
g15173 nand P2_U3491 P2_R1170_U59 ; P2_R1170_U288
g15174 nand P2_R1170_U60 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U289
g15175 nand P2_R1170_U289 P2_R1170_U288 ; P2_R1170_U290
g15176 nand P2_R1170_U287 P2_R1170_U286 P2_R1170_U87 ; P2_R1170_U291
g15177 nand P2_R1170_U172 P2_R1170_U290 ; P2_R1170_U292
g15178 nand P2_U3488 P2_R1170_U57 ; P2_R1170_U293
g15179 nand P2_R1170_U58 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U294
g15180 nand P2_U3485 P2_R1170_U52 ; P2_R1170_U295
g15181 nand P2_R1170_U53 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U296
g15182 nand P2_R1170_U296 P2_R1170_U295 ; P2_R1170_U297
g15183 nand P2_R1170_U225 P2_R1170_U67 ; P2_R1170_U298
g15184 nand P2_R1170_U297 P2_R1170_U205 ; P2_R1170_U299
g15185 nand P2_U3482 P2_R1170_U54 ; P2_R1170_U300
g15186 nand P2_R1170_U55 P2_REG2_REG_11__SCAN_IN ; P2_R1170_U301
g15187 nand P2_R1170_U301 P2_R1170_U300 ; P2_R1170_U302
g15188 nand P2_R1170_U226 P2_R1170_U88 ; P2_R1170_U303
g15189 nand P2_R1170_U162 P2_R1170_U302 ; P2_R1170_U304
g15190 nand P2_U3479 P2_R1170_U50 ; P2_R1170_U305
g15191 nand P2_R1170_U51 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U306
g15192 nand P2_U3446 P2_R1170_U27 ; P2_R1170_U307
g15193 nand P2_R1170_U28 P2_REG2_REG_0__SCAN_IN ; P2_R1170_U308
g15194 and P2_R1275_U135 P2_R1275_U35 ; P2_R1275_U6
g15195 and P2_R1275_U133 P2_R1275_U36 ; P2_R1275_U7
g15196 and P2_R1275_U132 P2_R1275_U37 ; P2_R1275_U8
g15197 and P2_R1275_U131 P2_R1275_U38 ; P2_R1275_U9
g15198 and P2_R1275_U129 P2_R1275_U39 ; P2_R1275_U10
g15199 and P2_R1275_U128 P2_R1275_U40 ; P2_R1275_U11
g15200 and P2_R1275_U127 P2_R1275_U41 ; P2_R1275_U12
g15201 and P2_R1275_U125 P2_R1275_U42 ; P2_R1275_U13
g15202 and P2_R1275_U123 P2_R1275_U43 ; P2_R1275_U14
g15203 and P2_R1275_U121 P2_R1275_U44 ; P2_R1275_U15
g15204 and P2_R1275_U119 P2_R1275_U45 ; P2_R1275_U16
g15205 and P2_R1275_U117 P2_R1275_U46 ; P2_R1275_U17
g15206 and P2_R1275_U115 P2_R1275_U25 ; P2_R1275_U18
g15207 and P2_R1275_U113 P2_R1275_U67 ; P2_R1275_U19
g15208 and P2_R1275_U98 P2_R1275_U26 ; P2_R1275_U20
g15209 and P2_R1275_U97 P2_R1275_U27 ; P2_R1275_U21
g15210 and P2_R1275_U96 P2_R1275_U28 ; P2_R1275_U22
g15211 and P2_R1275_U94 P2_R1275_U29 ; P2_R1275_U23
g15212 and P2_R1275_U93 P2_R1275_U30 ; P2_R1275_U24
g15213 or P2_U3453 P2_U3448 P2_U3456 ; P2_R1275_U25
g15214 nand P2_R1275_U87 P2_R1275_U34 ; P2_R1275_U26
g15215 nand P2_R1275_U88 P2_R1275_U33 ; P2_R1275_U27
g15216 nand P2_R1275_U56 P2_R1275_U89 ; P2_R1275_U28
g15217 nand P2_R1275_U90 P2_R1275_U32 ; P2_R1275_U29
g15218 nand P2_R1275_U91 P2_R1275_U31 ; P2_R1275_U30
g15219 not P2_U3474 ; P2_R1275_U31
g15220 not P2_U3471 ; P2_R1275_U32
g15221 not P2_U3462 ; P2_R1275_U33
g15222 not P2_U3459 ; P2_R1275_U34
g15223 nand P2_R1275_U57 P2_R1275_U92 ; P2_R1275_U35
g15224 nand P2_R1275_U99 P2_R1275_U54 ; P2_R1275_U36
g15225 nand P2_R1275_U100 P2_R1275_U53 ; P2_R1275_U37
g15226 nand P2_R1275_U58 P2_R1275_U101 ; P2_R1275_U38
g15227 nand P2_R1275_U102 P2_R1275_U52 ; P2_R1275_U39
g15228 nand P2_R1275_U103 P2_R1275_U51 ; P2_R1275_U40
g15229 nand P2_R1275_U59 P2_R1275_U104 ; P2_R1275_U41
g15230 nand P2_R1275_U60 P2_R1275_U105 ; P2_R1275_U42
g15231 nand P2_R1275_U61 P2_R1275_U106 ; P2_R1275_U43
g15232 nand P2_R1275_U107 P2_R1275_U75 P2_R1275_U50 ; P2_R1275_U44
g15233 nand P2_R1275_U108 P2_R1275_U73 P2_R1275_U49 ; P2_R1275_U45
g15234 nand P2_R1275_U109 P2_R1275_U71 P2_R1275_U48 ; P2_R1275_U46
g15235 not P2_U3978 ; P2_R1275_U47
g15236 not P2_U3968 ; P2_R1275_U48
g15237 not P2_U3970 ; P2_R1275_U49
g15238 not P2_U3972 ; P2_R1275_U50
g15239 not P2_U3498 ; P2_R1275_U51
g15240 not P2_U3495 ; P2_R1275_U52
g15241 not P2_U3486 ; P2_R1275_U53
g15242 not P2_U3483 ; P2_R1275_U54
g15243 nand P2_R1275_U153 P2_R1275_U152 ; P2_R1275_U55
g15244 nor P2_U3465 P2_U3468 ; P2_R1275_U56
g15245 nor P2_U3480 P2_U3477 ; P2_R1275_U57
g15246 nor P2_U3489 P2_U3492 ; P2_R1275_U58
g15247 nor P2_U3501 P2_U3504 ; P2_R1275_U59
g15248 nor P2_U3506 P2_U3976 ; P2_R1275_U60
g15249 nor P2_U3975 P2_U3974 ; P2_R1275_U61
g15250 not P2_U3477 ; P2_R1275_U62
g15251 and P2_R1275_U137 P2_R1275_U136 ; P2_R1275_U63
g15252 not P2_U3465 ; P2_R1275_U64
g15253 and P2_R1275_U139 P2_R1275_U138 ; P2_R1275_U65
g15254 not P2_U3977 ; P2_R1275_U66
g15255 nand P2_R1275_U110 P2_R1275_U69 P2_R1275_U47 ; P2_R1275_U67
g15256 and P2_R1275_U141 P2_R1275_U140 ; P2_R1275_U68
g15257 not P2_U3979 ; P2_R1275_U69
g15258 and P2_R1275_U143 P2_R1275_U142 ; P2_R1275_U70
g15259 not P2_U3969 ; P2_R1275_U71
g15260 and P2_R1275_U145 P2_R1275_U144 ; P2_R1275_U72
g15261 not P2_U3971 ; P2_R1275_U73
g15262 and P2_R1275_U147 P2_R1275_U146 ; P2_R1275_U74
g15263 not P2_U3973 ; P2_R1275_U75
g15264 and P2_R1275_U149 P2_R1275_U148 ; P2_R1275_U76
g15265 not P2_U3975 ; P2_R1275_U77
g15266 and P2_R1275_U151 P2_R1275_U150 ; P2_R1275_U78
g15267 not P2_U3453 ; P2_R1275_U79
g15268 not P2_U3448 ; P2_R1275_U80
g15269 not P2_U3506 ; P2_R1275_U81
g15270 and P2_R1275_U155 P2_R1275_U154 ; P2_R1275_U82
g15271 not P2_U3501 ; P2_R1275_U83
g15272 and P2_R1275_U157 P2_R1275_U156 ; P2_R1275_U84
g15273 not P2_U3489 ; P2_R1275_U85
g15274 and P2_R1275_U159 P2_R1275_U158 ; P2_R1275_U86
g15275 not P2_R1275_U25 ; P2_R1275_U87
g15276 not P2_R1275_U26 ; P2_R1275_U88
g15277 not P2_R1275_U27 ; P2_R1275_U89
g15278 not P2_R1275_U28 ; P2_R1275_U90
g15279 not P2_R1275_U29 ; P2_R1275_U91
g15280 not P2_R1275_U30 ; P2_R1275_U92
g15281 nand P2_U3474 P2_R1275_U29 ; P2_R1275_U93
g15282 nand P2_U3471 P2_R1275_U28 ; P2_R1275_U94
g15283 nand P2_R1275_U89 P2_R1275_U64 ; P2_R1275_U95
g15284 nand P2_U3468 P2_R1275_U95 ; P2_R1275_U96
g15285 nand P2_U3462 P2_R1275_U26 ; P2_R1275_U97
g15286 nand P2_U3459 P2_R1275_U25 ; P2_R1275_U98
g15287 not P2_R1275_U35 ; P2_R1275_U99
g15288 not P2_R1275_U36 ; P2_R1275_U100
g15289 not P2_R1275_U37 ; P2_R1275_U101
g15290 not P2_R1275_U38 ; P2_R1275_U102
g15291 not P2_R1275_U39 ; P2_R1275_U103
g15292 not P2_R1275_U40 ; P2_R1275_U104
g15293 not P2_R1275_U41 ; P2_R1275_U105
g15294 not P2_R1275_U42 ; P2_R1275_U106
g15295 not P2_R1275_U43 ; P2_R1275_U107
g15296 not P2_R1275_U44 ; P2_R1275_U108
g15297 not P2_R1275_U45 ; P2_R1275_U109
g15298 not P2_R1275_U46 ; P2_R1275_U110
g15299 not P2_R1275_U67 ; P2_R1275_U111
g15300 nand P2_R1275_U110 P2_R1275_U69 ; P2_R1275_U112
g15301 nand P2_U3978 P2_R1275_U112 ; P2_R1275_U113
g15302 or P2_U3453 P2_U3448 ; P2_R1275_U114
g15303 nand P2_U3456 P2_R1275_U114 ; P2_R1275_U115
g15304 nand P2_R1275_U109 P2_R1275_U71 ; P2_R1275_U116
g15305 nand P2_U3968 P2_R1275_U116 ; P2_R1275_U117
g15306 nand P2_R1275_U108 P2_R1275_U73 ; P2_R1275_U118
g15307 nand P2_U3970 P2_R1275_U118 ; P2_R1275_U119
g15308 nand P2_R1275_U107 P2_R1275_U75 ; P2_R1275_U120
g15309 nand P2_U3972 P2_R1275_U120 ; P2_R1275_U121
g15310 nand P2_R1275_U106 P2_R1275_U77 ; P2_R1275_U122
g15311 nand P2_U3974 P2_R1275_U122 ; P2_R1275_U123
g15312 nand P2_R1275_U105 P2_R1275_U81 ; P2_R1275_U124
g15313 nand P2_U3976 P2_R1275_U124 ; P2_R1275_U125
g15314 nand P2_R1275_U104 P2_R1275_U83 ; P2_R1275_U126
g15315 nand P2_U3504 P2_R1275_U126 ; P2_R1275_U127
g15316 nand P2_U3498 P2_R1275_U39 ; P2_R1275_U128
g15317 nand P2_U3495 P2_R1275_U38 ; P2_R1275_U129
g15318 nand P2_R1275_U101 P2_R1275_U85 ; P2_R1275_U130
g15319 nand P2_U3492 P2_R1275_U130 ; P2_R1275_U131
g15320 nand P2_U3486 P2_R1275_U36 ; P2_R1275_U132
g15321 nand P2_U3483 P2_R1275_U35 ; P2_R1275_U133
g15322 nand P2_R1275_U92 P2_R1275_U62 ; P2_R1275_U134
g15323 nand P2_U3480 P2_R1275_U134 ; P2_R1275_U135
g15324 nand P2_U3477 P2_R1275_U30 ; P2_R1275_U136
g15325 nand P2_R1275_U92 P2_R1275_U62 ; P2_R1275_U137
g15326 nand P2_U3465 P2_R1275_U27 ; P2_R1275_U138
g15327 nand P2_R1275_U89 P2_R1275_U64 ; P2_R1275_U139
g15328 nand P2_U3977 P2_R1275_U67 ; P2_R1275_U140
g15329 nand P2_R1275_U111 P2_R1275_U66 ; P2_R1275_U141
g15330 nand P2_U3979 P2_R1275_U46 ; P2_R1275_U142
g15331 nand P2_R1275_U110 P2_R1275_U69 ; P2_R1275_U143
g15332 nand P2_U3969 P2_R1275_U45 ; P2_R1275_U144
g15333 nand P2_R1275_U109 P2_R1275_U71 ; P2_R1275_U145
g15334 nand P2_U3971 P2_R1275_U44 ; P2_R1275_U146
g15335 nand P2_R1275_U108 P2_R1275_U73 ; P2_R1275_U147
g15336 nand P2_U3973 P2_R1275_U43 ; P2_R1275_U148
g15337 nand P2_R1275_U107 P2_R1275_U75 ; P2_R1275_U149
g15338 nand P2_U3975 P2_R1275_U42 ; P2_R1275_U150
g15339 nand P2_R1275_U106 P2_R1275_U77 ; P2_R1275_U151
g15340 nand P2_U3453 P2_R1275_U80 ; P2_R1275_U152
g15341 nand P2_U3448 P2_R1275_U79 ; P2_R1275_U153
g15342 nand P2_U3506 P2_R1275_U41 ; P2_R1275_U154
g15343 nand P2_R1275_U105 P2_R1275_U81 ; P2_R1275_U155
g15344 nand P2_U3501 P2_R1275_U40 ; P2_R1275_U156
g15345 nand P2_R1275_U104 P2_R1275_U83 ; P2_R1275_U157
g15346 nand P2_U3489 P2_R1275_U37 ; P2_R1275_U158
g15347 nand P2_R1275_U101 P2_R1275_U85 ; P2_R1275_U159
g15348 and P2_LT_719_U115 P2_LT_719_U116 ; P2_LT_719_U6
g15349 and P2_LT_719_U122 P2_LT_719_U121 P2_LT_719_U120 P2_LT_719_U118 ; P2_LT_719_U7
g15350 and P2_LT_719_U75 P2_LT_719_U7 ; P2_LT_719_U8
g15351 and P2_LT_719_U8 P2_LT_719_U126 ; P2_LT_719_U9
g15352 and P2_LT_719_U111 P2_LT_719_U112 P2_LT_719_U109 ; P2_LT_719_U10
g15353 and P2_LT_719_U186 P2_LT_719_U185 P2_LT_719_U105 P2_LT_719_U106 ; P2_LT_719_U11
g15354 not P2_U3979 ; P2_LT_719_U12
g15355 not P2_U3592 ; P2_LT_719_U13
g15356 not P2_U3599 ; P2_LT_719_U14
g15357 not P2_U3600 ; P2_LT_719_U15
g15358 not P2_U3974 ; P2_LT_719_U16
g15359 not P2_U3606 ; P2_LT_719_U17
g15360 not P2_U3605 ; P2_LT_719_U18
g15361 not P2_U3498 ; P2_LT_719_U19
g15362 not P2_U3495 ; P2_LT_719_U20
g15363 not P2_U3492 ; P2_LT_719_U21
g15364 not P2_U3611 ; P2_LT_719_U22
g15365 not P2_U3480 ; P2_LT_719_U23
g15366 not P2_U3477 ; P2_LT_719_U24
g15367 not P2_U3471 ; P2_LT_719_U25
g15368 not P2_U3474 ; P2_LT_719_U26
g15369 not P2_U3468 ; P2_LT_719_U27
g15370 not P2_U3465 ; P2_LT_719_U28
g15371 not P2_U3462 ; P2_LT_719_U29
g15372 not P2_U3459 ; P2_LT_719_U30
g15373 not P2_U3604 ; P2_LT_719_U31
g15374 not P2_U3456 ; P2_LT_719_U32
g15375 not P2_U3453 ; P2_LT_719_U33
g15376 not P2_U3612 ; P2_LT_719_U34
g15377 not P2_U3593 ; P2_LT_719_U35
g15378 not P2_U3590 ; P2_LT_719_U36
g15379 not P2_U3589 ; P2_LT_719_U37
g15380 not P2_U3588 ; P2_LT_719_U38
g15381 not P2_U3587 ; P2_LT_719_U39
g15382 not P2_U3586 ; P2_LT_719_U40
g15383 not P2_U3585 ; P2_LT_719_U41
g15384 not P2_U3584 ; P2_LT_719_U42
g15385 not P2_U3614 ; P2_LT_719_U43
g15386 not P2_U3613 ; P2_LT_719_U44
g15387 not P2_U3486 ; P2_LT_719_U45
g15388 not P2_U3483 ; P2_LT_719_U46
g15389 not P2_U3489 ; P2_LT_719_U47
g15390 not P2_U3610 ; P2_LT_719_U48
g15391 not P2_U3609 ; P2_LT_719_U49
g15392 not P2_U3608 ; P2_LT_719_U50
g15393 not P2_U3607 ; P2_LT_719_U51
g15394 not P2_U3975 ; P2_LT_719_U52
g15395 not P2_U3504 ; P2_LT_719_U53
g15396 not P2_U3501 ; P2_LT_719_U54
g15397 not P2_U3506 ; P2_LT_719_U55
g15398 not P2_U3976 ; P2_LT_719_U56
g15399 not P2_U3603 ; P2_LT_719_U57
g15400 not P2_U3602 ; P2_LT_719_U58
g15401 not P2_U3601 ; P2_LT_719_U59
g15402 not P2_U3973 ; P2_LT_719_U60
g15403 not P2_U3972 ; P2_LT_719_U61
g15404 nand P2_LT_719_U179 P2_LT_719_U178 ; P2_LT_719_U62
g15405 not P2_U3598 ; P2_LT_719_U63
g15406 not P2_U3970 ; P2_LT_719_U64
g15407 not P2_U3591 ; P2_LT_719_U65
g15408 not P2_U3969 ; P2_LT_719_U66
g15409 not P2_U3968 ; P2_LT_719_U67
g15410 not P2_U3978 ; P2_LT_719_U68
g15411 not P2_U3594 ; P2_LT_719_U69
g15412 not P2_U3596 ; P2_LT_719_U70
g15413 not P2_U3597 ; P2_LT_719_U71
g15414 not P2_U3977 ; P2_LT_719_U72
g15415 not P2_U3595 ; P2_LT_719_U73
g15416 and P2_U3448 P2_LT_719_U107 ; P2_LT_719_U74
g15417 and P2_LT_719_U124 P2_LT_719_U123 P2_LT_719_U125 ; P2_LT_719_U75
g15418 and P2_LT_719_U128 P2_LT_719_U129 ; P2_LT_719_U76
g15419 and P2_LT_719_U76 P2_LT_719_U127 ; P2_LT_719_U77
g15420 and P2_U3593 P2_LT_719_U32 ; P2_LT_719_U78
g15421 and P2_U3590 P2_LT_719_U30 ; P2_LT_719_U79
g15422 and P2_LT_719_U124 P2_LT_719_U123 ; P2_LT_719_U80
g15423 and P2_LT_719_U140 P2_LT_719_U141 ; P2_LT_719_U81
g15424 and P2_LT_719_U120 P2_LT_719_U118 ; P2_LT_719_U82
g15425 and P2_LT_719_U146 P2_LT_719_U84 ; P2_LT_719_U83
g15426 and P2_LT_719_U148 P2_LT_719_U147 ; P2_LT_719_U84
g15427 and P2_LT_719_U145 P2_LT_719_U83 ; P2_LT_719_U85
g15428 and P2_U3483 P2_LT_719_U44 ; P2_LT_719_U86
g15429 and P2_LT_719_U151 P2_LT_719_U88 ; P2_LT_719_U87
g15430 and P2_LT_719_U152 P2_LT_719_U150 ; P2_LT_719_U88
g15431 and P2_LT_719_U155 P2_LT_719_U132 ; P2_LT_719_U89
g15432 and P2_LT_719_U153 P2_LT_719_U117 ; P2_LT_719_U90
g15433 and P2_LT_719_U6 P2_LT_719_U92 ; P2_LT_719_U91
g15434 and P2_LT_719_U161 P2_LT_719_U162 ; P2_LT_719_U92
g15435 and P2_U3504 P2_LT_719_U17 ; P2_LT_719_U93
g15436 and P2_U3501 P2_LT_719_U51 ; P2_LT_719_U94
g15437 and P2_LT_719_U164 P2_LT_719_U166 ; P2_LT_719_U95
g15438 and P2_LT_719_U168 P2_LT_719_U167 P2_LT_719_U169 P2_LT_719_U95 ; P2_LT_719_U96
g15439 and P2_U3603 P2_LT_719_U56 ; P2_LT_719_U97
g15440 and P2_LT_719_U171 P2_LT_719_U172 P2_LT_719_U173 ; P2_LT_719_U98
g15441 and P2_LT_719_U176 P2_LT_719_U165 ; P2_LT_719_U99
g15442 and P2_LT_719_U174 P2_LT_719_U113 ; P2_LT_719_U100
g15443 and P2_LT_719_U10 P2_LT_719_U184 ; P2_LT_719_U101
g15444 and P2_U3594 P2_LT_719_U12 ; P2_LT_719_U102
g15445 and P2_LT_719_U104 P2_LT_719_U109 ; P2_LT_719_U103
g15446 and P2_U3595 P2_LT_719_U67 ; P2_LT_719_U104
g15447 and P2_LT_719_U189 P2_LT_719_U188 ; P2_LT_719_U105
g15448 and P2_LT_719_U191 P2_LT_719_U192 P2_LT_719_U190 ; P2_LT_719_U106
g15449 not P2_U3615 ; P2_LT_719_U107
g15450 nand P2_LT_719_U194 P2_LT_719_U193 ; P2_LT_719_U108
g15451 nand P2_U3591 P2_LT_719_U72 ; P2_LT_719_U109
g15452 nand P2_U3979 P2_LT_719_U69 ; P2_LT_719_U110
g15453 nand P2_U3969 P2_LT_719_U70 ; P2_LT_719_U111
g15454 nand P2_U3968 P2_LT_719_U73 ; P2_LT_719_U112
g15455 nand P2_U3599 P2_LT_719_U61 ; P2_LT_719_U113
g15456 nand P2_U3498 P2_LT_719_U50 ; P2_LT_719_U114
g15457 nand P2_U3605 P2_LT_719_U55 ; P2_LT_719_U115
g15458 nand P2_U3606 P2_LT_719_U53 ; P2_LT_719_U116
g15459 nand P2_U3495 P2_LT_719_U49 ; P2_LT_719_U117
g15460 nand P2_U3480 P2_LT_719_U43 ; P2_LT_719_U118
g15461 nand P2_U3604 P2_LT_719_U33 ; P2_LT_719_U119
g15462 nand P2_U3477 P2_LT_719_U42 ; P2_LT_719_U120
g15463 nand P2_U3471 P2_LT_719_U40 ; P2_LT_719_U121
g15464 nand P2_U3474 P2_LT_719_U41 ; P2_LT_719_U122
g15465 nand P2_U3468 P2_LT_719_U39 ; P2_LT_719_U123
g15466 nand P2_U3465 P2_LT_719_U38 ; P2_LT_719_U124
g15467 nand P2_U3462 P2_LT_719_U37 ; P2_LT_719_U125
g15468 nand P2_U3459 P2_LT_719_U36 ; P2_LT_719_U126
g15469 nand P2_LT_719_U74 P2_LT_719_U119 ; P2_LT_719_U127
g15470 nand P2_U3456 P2_LT_719_U35 ; P2_LT_719_U128
g15471 nand P2_U3453 P2_LT_719_U31 ; P2_LT_719_U129
g15472 nand P2_LT_719_U77 P2_LT_719_U9 ; P2_LT_719_U130
g15473 nand P2_U3612 P2_LT_719_U45 ; P2_LT_719_U131
g15474 nand P2_U3611 P2_LT_719_U47 ; P2_LT_719_U132
g15475 nand P2_U3585 P2_LT_719_U26 ; P2_LT_719_U133
g15476 nand P2_U3584 P2_LT_719_U24 ; P2_LT_719_U134
g15477 nand P2_LT_719_U134 P2_LT_719_U133 ; P2_LT_719_U135
g15478 nand P2_U3589 P2_LT_719_U29 ; P2_LT_719_U136
g15479 nand P2_U3588 P2_LT_719_U28 ; P2_LT_719_U137
g15480 nand P2_LT_719_U137 P2_LT_719_U136 ; P2_LT_719_U138
g15481 nand P2_LT_719_U80 P2_LT_719_U138 ; P2_LT_719_U139
g15482 nand P2_U3587 P2_LT_719_U27 ; P2_LT_719_U140
g15483 nand P2_U3586 P2_LT_719_U25 ; P2_LT_719_U141
g15484 nand P2_LT_719_U81 P2_LT_719_U139 ; P2_LT_719_U142
g15485 nand P2_LT_719_U78 P2_LT_719_U9 ; P2_LT_719_U143
g15486 nand P2_LT_719_U79 P2_LT_719_U8 ; P2_LT_719_U144
g15487 nand P2_LT_719_U7 P2_LT_719_U142 ; P2_LT_719_U145
g15488 nand P2_LT_719_U82 P2_LT_719_U135 ; P2_LT_719_U146
g15489 nand P2_U3614 P2_LT_719_U23 ; P2_LT_719_U147
g15490 nand P2_U3613 P2_LT_719_U46 ; P2_LT_719_U148
g15491 nand P2_LT_719_U144 P2_LT_719_U143 P2_LT_719_U131 P2_LT_719_U130 P2_LT_719_U85 ; P2_LT_719_U149
g15492 nand P2_U3486 P2_LT_719_U34 ; P2_LT_719_U150
g15493 nand P2_LT_719_U86 P2_LT_719_U131 ; P2_LT_719_U151
g15494 nand P2_U3489 P2_LT_719_U22 ; P2_LT_719_U152
g15495 nand P2_U3492 P2_LT_719_U48 ; P2_LT_719_U153
g15496 nand P2_LT_719_U149 P2_LT_719_U87 ; P2_LT_719_U154
g15497 nand P2_U3610 P2_LT_719_U21 ; P2_LT_719_U155
g15498 nand P2_LT_719_U89 P2_LT_719_U154 ; P2_LT_719_U156
g15499 nand P2_LT_719_U90 P2_LT_719_U156 ; P2_LT_719_U157
g15500 nand P2_U3609 P2_LT_719_U20 ; P2_LT_719_U158
g15501 nand P2_LT_719_U158 P2_LT_719_U157 ; P2_LT_719_U159
g15502 nand P2_LT_719_U159 P2_LT_719_U114 ; P2_LT_719_U160
g15503 nand P2_U3608 P2_LT_719_U19 ; P2_LT_719_U161
g15504 nand P2_U3607 P2_LT_719_U54 ; P2_LT_719_U162
g15505 nand P2_LT_719_U160 P2_LT_719_U91 ; P2_LT_719_U163
g15506 nand P2_U3975 P2_LT_719_U58 ; P2_LT_719_U164
g15507 nand P2_U3974 P2_LT_719_U59 ; P2_LT_719_U165
g15508 nand P2_LT_719_U93 P2_LT_719_U115 ; P2_LT_719_U166
g15509 nand P2_LT_719_U94 P2_LT_719_U6 ; P2_LT_719_U167
g15510 nand P2_U3506 P2_LT_719_U18 ; P2_LT_719_U168
g15511 nand P2_U3976 P2_LT_719_U57 ; P2_LT_719_U169
g15512 nand P2_LT_719_U163 P2_LT_719_U96 ; P2_LT_719_U170
g15513 nand P2_LT_719_U97 P2_LT_719_U164 ; P2_LT_719_U171
g15514 nand P2_U3602 P2_LT_719_U52 ; P2_LT_719_U172
g15515 nand P2_U3601 P2_LT_719_U16 ; P2_LT_719_U173
g15516 nand P2_U3600 P2_LT_719_U60 ; P2_LT_719_U174
g15517 nand P2_LT_719_U170 P2_LT_719_U98 ; P2_LT_719_U175
g15518 nand P2_U3973 P2_LT_719_U15 ; P2_LT_719_U176
g15519 nand P2_LT_719_U99 P2_LT_719_U175 ; P2_LT_719_U177
g15520 nand P2_LT_719_U100 P2_LT_719_U177 ; P2_LT_719_U178
g15521 nand P2_U3972 P2_LT_719_U14 ; P2_LT_719_U179
g15522 not P2_LT_719_U62 ; P2_LT_719_U180
g15523 nand P2_U3598 P2_LT_719_U180 ; P2_LT_719_U181
g15524 nand P2_U3971 P2_LT_719_U181 ; P2_LT_719_U182
g15525 nand P2_LT_719_U62 P2_LT_719_U63 ; P2_LT_719_U183
g15526 nand P2_U3970 P2_LT_719_U71 ; P2_LT_719_U184
g15527 nand P2_LT_719_U182 P2_LT_719_U183 P2_LT_719_U108 P2_LT_719_U101 ; P2_LT_719_U185
g15528 nand P2_LT_719_U109 P2_U3592 P2_LT_719_U68 ; P2_LT_719_U186
g15529 nand P2_U3978 P2_LT_719_U13 ; P2_LT_719_U187
g15530 nand P2_LT_719_U109 P2_LT_719_U102 P2_LT_719_U187 ; P2_LT_719_U188
g15531 nand P2_U3596 P2_LT_719_U10 P2_LT_719_U108 P2_LT_719_U66 ; P2_LT_719_U189
g15532 nand P2_U3597 P2_LT_719_U10 P2_LT_719_U108 P2_LT_719_U64 ; P2_LT_719_U190
g15533 nand P2_U3977 P2_LT_719_U65 ; P2_LT_719_U191
g15534 nand P2_LT_719_U108 P2_LT_719_U103 ; P2_LT_719_U192
g15535 nand P2_U3592 P2_LT_719_U110 ; P2_LT_719_U193
g15536 nand P2_LT_719_U110 P2_LT_719_U68 ; P2_LT_719_U194
g15537 and P2_R1179_U205 P2_R1179_U204 ; P2_R1179_U6
g15538 and P2_R1179_U244 P2_R1179_U243 ; P2_R1179_U7
g15539 and P2_R1179_U261 P2_R1179_U260 ; P2_R1179_U8
g15540 and P2_R1179_U285 P2_R1179_U284 ; P2_R1179_U9
g15541 and P2_R1179_U384 P2_R1179_U383 ; P2_R1179_U10
g15542 nand P2_R1179_U340 P2_R1179_U343 ; P2_R1179_U11
g15543 nand P2_R1179_U329 P2_R1179_U332 ; P2_R1179_U12
g15544 nand P2_R1179_U318 P2_R1179_U321 ; P2_R1179_U13
g15545 nand P2_R1179_U310 P2_R1179_U312 ; P2_R1179_U14
g15546 nand P2_R1179_U349 P2_R1179_U177 P2_R1179_U156 ; P2_R1179_U15
g15547 nand P2_R1179_U238 P2_R1179_U240 ; P2_R1179_U16
g15548 nand P2_R1179_U230 P2_R1179_U233 ; P2_R1179_U17
g15549 nand P2_R1179_U222 P2_R1179_U224 ; P2_R1179_U18
g15550 nand P2_R1179_U166 P2_R1179_U346 ; P2_R1179_U19
g15551 not P2_U3471 ; P2_R1179_U20
g15552 not P2_U3465 ; P2_R1179_U21
g15553 not P2_U3456 ; P2_R1179_U22
g15554 not P2_U3448 ; P2_R1179_U23
g15555 not P2_U3078 ; P2_R1179_U24
g15556 not P2_U3459 ; P2_R1179_U25
g15557 not P2_U3068 ; P2_R1179_U26
g15558 nand P2_U3068 P2_R1179_U22 ; P2_R1179_U27
g15559 not P2_U3064 ; P2_R1179_U28
g15560 not P2_U3468 ; P2_R1179_U29
g15561 not P2_U3462 ; P2_R1179_U30
g15562 not P2_U3071 ; P2_R1179_U31
g15563 not P2_U3067 ; P2_R1179_U32
g15564 not P2_U3060 ; P2_R1179_U33
g15565 nand P2_U3060 P2_R1179_U30 ; P2_R1179_U34
g15566 not P2_U3474 ; P2_R1179_U35
g15567 not P2_U3070 ; P2_R1179_U36
g15568 nand P2_U3070 P2_R1179_U20 ; P2_R1179_U37
g15569 not P2_U3084 ; P2_R1179_U38
g15570 not P2_U3477 ; P2_R1179_U39
g15571 not P2_U3083 ; P2_R1179_U40
g15572 nand P2_R1179_U211 P2_R1179_U210 ; P2_R1179_U41
g15573 nand P2_R1179_U34 P2_R1179_U226 ; P2_R1179_U42
g15574 nand P2_R1179_U195 P2_R1179_U179 P2_R1179_U347 ; P2_R1179_U43
g15575 not P2_U3970 ; P2_R1179_U44
g15576 not P2_U3974 ; P2_R1179_U45
g15577 not P2_U3495 ; P2_R1179_U46
g15578 not P2_U3480 ; P2_R1179_U47
g15579 not P2_U3483 ; P2_R1179_U48
g15580 not P2_U3063 ; P2_R1179_U49
g15581 not P2_U3062 ; P2_R1179_U50
g15582 nand P2_U3083 P2_R1179_U39 ; P2_R1179_U51
g15583 not P2_U3486 ; P2_R1179_U52
g15584 not P2_U3072 ; P2_R1179_U53
g15585 not P2_U3489 ; P2_R1179_U54
g15586 not P2_U3080 ; P2_R1179_U55
g15587 not P2_U3498 ; P2_R1179_U56
g15588 not P2_U3492 ; P2_R1179_U57
g15589 not P2_U3073 ; P2_R1179_U58
g15590 not P2_U3074 ; P2_R1179_U59
g15591 not P2_U3079 ; P2_R1179_U60
g15592 nand P2_U3079 P2_R1179_U57 ; P2_R1179_U61
g15593 not P2_U3501 ; P2_R1179_U62
g15594 not P2_U3069 ; P2_R1179_U63
g15595 not P2_U3082 ; P2_R1179_U64
g15596 not P2_U3506 ; P2_R1179_U65
g15597 not P2_U3081 ; P2_R1179_U66
g15598 not P2_U3976 ; P2_R1179_U67
g15599 not P2_U3076 ; P2_R1179_U68
g15600 not P2_U3973 ; P2_R1179_U69
g15601 not P2_U3975 ; P2_R1179_U70
g15602 not P2_U3066 ; P2_R1179_U71
g15603 not P2_U3061 ; P2_R1179_U72
g15604 not P2_U3075 ; P2_R1179_U73
g15605 nand P2_U3075 P2_R1179_U70 ; P2_R1179_U74
g15606 not P2_U3972 ; P2_R1179_U75
g15607 not P2_U3065 ; P2_R1179_U76
g15608 not P2_U3971 ; P2_R1179_U77
g15609 not P2_U3058 ; P2_R1179_U78
g15610 not P2_U3969 ; P2_R1179_U79
g15611 not P2_U3057 ; P2_R1179_U80
g15612 nand P2_U3057 P2_R1179_U44 ; P2_R1179_U81
g15613 not P2_U3053 ; P2_R1179_U82
g15614 not P2_U3968 ; P2_R1179_U83
g15615 not P2_U3054 ; P2_R1179_U84
g15616 nand P2_R1179_U299 P2_R1179_U298 ; P2_R1179_U85
g15617 nand P2_R1179_U74 P2_R1179_U314 ; P2_R1179_U86
g15618 nand P2_R1179_U61 P2_R1179_U325 ; P2_R1179_U87
g15619 nand P2_R1179_U51 P2_R1179_U336 ; P2_R1179_U88
g15620 not P2_U3077 ; P2_R1179_U89
g15621 nand P2_R1179_U394 P2_R1179_U393 ; P2_R1179_U90
g15622 nand P2_R1179_U408 P2_R1179_U407 ; P2_R1179_U91
g15623 nand P2_R1179_U413 P2_R1179_U412 ; P2_R1179_U92
g15624 nand P2_R1179_U429 P2_R1179_U428 ; P2_R1179_U93
g15625 nand P2_R1179_U434 P2_R1179_U433 ; P2_R1179_U94
g15626 nand P2_R1179_U439 P2_R1179_U438 ; P2_R1179_U95
g15627 nand P2_R1179_U444 P2_R1179_U443 ; P2_R1179_U96
g15628 nand P2_R1179_U449 P2_R1179_U448 ; P2_R1179_U97
g15629 nand P2_R1179_U465 P2_R1179_U464 ; P2_R1179_U98
g15630 nand P2_R1179_U470 P2_R1179_U469 ; P2_R1179_U99
g15631 nand P2_R1179_U353 P2_R1179_U352 ; P2_R1179_U100
g15632 nand P2_R1179_U362 P2_R1179_U361 ; P2_R1179_U101
g15633 nand P2_R1179_U369 P2_R1179_U368 ; P2_R1179_U102
g15634 nand P2_R1179_U373 P2_R1179_U372 ; P2_R1179_U103
g15635 nand P2_R1179_U382 P2_R1179_U381 ; P2_R1179_U104
g15636 nand P2_R1179_U403 P2_R1179_U402 ; P2_R1179_U105
g15637 nand P2_R1179_U420 P2_R1179_U419 ; P2_R1179_U106
g15638 nand P2_R1179_U424 P2_R1179_U423 ; P2_R1179_U107
g15639 nand P2_R1179_U456 P2_R1179_U455 ; P2_R1179_U108
g15640 nand P2_R1179_U460 P2_R1179_U459 ; P2_R1179_U109
g15641 nand P2_R1179_U477 P2_R1179_U476 ; P2_R1179_U110
g15642 and P2_R1179_U197 P2_R1179_U187 ; P2_R1179_U111
g15643 and P2_R1179_U200 P2_R1179_U201 ; P2_R1179_U112
g15644 and P2_R1179_U208 P2_R1179_U203 P2_R1179_U188 ; P2_R1179_U113
g15645 and P2_R1179_U213 P2_R1179_U189 ; P2_R1179_U114
g15646 and P2_R1179_U216 P2_R1179_U217 ; P2_R1179_U115
g15647 and P2_R1179_U355 P2_R1179_U354 P2_R1179_U37 ; P2_R1179_U116
g15648 and P2_R1179_U358 P2_R1179_U189 ; P2_R1179_U117
g15649 and P2_R1179_U232 P2_R1179_U6 ; P2_R1179_U118
g15650 and P2_R1179_U365 P2_R1179_U188 ; P2_R1179_U119
g15651 and P2_R1179_U375 P2_R1179_U374 P2_R1179_U27 ; P2_R1179_U120
g15652 and P2_R1179_U378 P2_R1179_U187 ; P2_R1179_U121
g15653 and P2_R1179_U242 P2_R1179_U219 P2_R1179_U183 ; P2_R1179_U122
g15654 and P2_R1179_U264 P2_R1179_U184 P2_R1179_U259 ; P2_R1179_U123
g15655 and P2_R1179_U288 P2_R1179_U185 P2_R1179_U283 ; P2_R1179_U124
g15656 and P2_R1179_U301 P2_R1179_U186 ; P2_R1179_U125
g15657 and P2_R1179_U304 P2_R1179_U305 ; P2_R1179_U126
g15658 and P2_R1179_U304 P2_R1179_U305 ; P2_R1179_U127
g15659 and P2_R1179_U10 P2_R1179_U308 ; P2_R1179_U128
g15660 nand P2_R1179_U391 P2_R1179_U390 ; P2_R1179_U129
g15661 and P2_R1179_U396 P2_R1179_U395 P2_R1179_U81 ; P2_R1179_U130
g15662 and P2_R1179_U399 P2_R1179_U186 ; P2_R1179_U131
g15663 nand P2_R1179_U405 P2_R1179_U404 ; P2_R1179_U132
g15664 nand P2_R1179_U410 P2_R1179_U409 ; P2_R1179_U133
g15665 and P2_R1179_U320 P2_R1179_U9 ; P2_R1179_U134
g15666 and P2_R1179_U416 P2_R1179_U185 ; P2_R1179_U135
g15667 nand P2_R1179_U426 P2_R1179_U425 ; P2_R1179_U136
g15668 nand P2_R1179_U431 P2_R1179_U430 ; P2_R1179_U137
g15669 nand P2_R1179_U436 P2_R1179_U435 ; P2_R1179_U138
g15670 nand P2_R1179_U441 P2_R1179_U440 ; P2_R1179_U139
g15671 nand P2_R1179_U446 P2_R1179_U445 ; P2_R1179_U140
g15672 and P2_R1179_U331 P2_R1179_U8 ; P2_R1179_U141
g15673 and P2_R1179_U452 P2_R1179_U184 ; P2_R1179_U142
g15674 nand P2_R1179_U462 P2_R1179_U461 ; P2_R1179_U143
g15675 nand P2_R1179_U467 P2_R1179_U466 ; P2_R1179_U144
g15676 and P2_R1179_U342 P2_R1179_U7 ; P2_R1179_U145
g15677 and P2_R1179_U473 P2_R1179_U183 ; P2_R1179_U146
g15678 and P2_R1179_U351 P2_R1179_U350 ; P2_R1179_U147
g15679 nand P2_R1179_U115 P2_R1179_U214 ; P2_R1179_U148
g15680 and P2_R1179_U360 P2_R1179_U359 ; P2_R1179_U149
g15681 and P2_R1179_U367 P2_R1179_U366 ; P2_R1179_U150
g15682 and P2_R1179_U371 P2_R1179_U370 ; P2_R1179_U151
g15683 nand P2_R1179_U112 P2_R1179_U198 ; P2_R1179_U152
g15684 and P2_R1179_U380 P2_R1179_U379 ; P2_R1179_U153
g15685 not P2_U3979 ; P2_R1179_U154
g15686 not P2_U3055 ; P2_R1179_U155
g15687 and P2_R1179_U389 P2_R1179_U388 ; P2_R1179_U156
g15688 nand P2_R1179_U126 P2_R1179_U302 ; P2_R1179_U157
g15689 and P2_R1179_U401 P2_R1179_U400 ; P2_R1179_U158
g15690 nand P2_R1179_U295 P2_R1179_U294 ; P2_R1179_U159
g15691 nand P2_R1179_U291 P2_R1179_U290 ; P2_R1179_U160
g15692 and P2_R1179_U418 P2_R1179_U417 ; P2_R1179_U161
g15693 and P2_R1179_U422 P2_R1179_U421 ; P2_R1179_U162
g15694 nand P2_R1179_U281 P2_R1179_U280 ; P2_R1179_U163
g15695 nand P2_R1179_U277 P2_R1179_U276 ; P2_R1179_U164
g15696 not P2_U3453 ; P2_R1179_U165
g15697 nand P2_U3448 P2_R1179_U89 ; P2_R1179_U166
g15698 nand P2_R1179_U273 P2_R1179_U178 P2_R1179_U348 ; P2_R1179_U167
g15699 not P2_U3504 ; P2_R1179_U168
g15700 nand P2_R1179_U271 P2_R1179_U270 ; P2_R1179_U169
g15701 nand P2_R1179_U267 P2_R1179_U266 ; P2_R1179_U170
g15702 and P2_R1179_U454 P2_R1179_U453 ; P2_R1179_U171
g15703 and P2_R1179_U458 P2_R1179_U457 ; P2_R1179_U172
g15704 nand P2_R1179_U257 P2_R1179_U256 ; P2_R1179_U173
g15705 nand P2_R1179_U253 P2_R1179_U252 ; P2_R1179_U174
g15706 nand P2_R1179_U249 P2_R1179_U248 ; P2_R1179_U175
g15707 and P2_R1179_U475 P2_R1179_U474 ; P2_R1179_U176
g15708 nand P2_R1179_U307 P2_R1179_U157 P2_R1179_U387 ; P2_R1179_U177
g15709 nand P2_R1179_U169 P2_R1179_U168 ; P2_R1179_U178
g15710 nand P2_R1179_U166 P2_R1179_U165 ; P2_R1179_U179
g15711 not P2_R1179_U81 ; P2_R1179_U180
g15712 not P2_R1179_U27 ; P2_R1179_U181
g15713 not P2_R1179_U37 ; P2_R1179_U182
g15714 nand P2_U3480 P2_R1179_U50 ; P2_R1179_U183
g15715 nand P2_U3495 P2_R1179_U59 ; P2_R1179_U184
g15716 nand P2_U3974 P2_R1179_U72 ; P2_R1179_U185
g15717 nand P2_U3970 P2_R1179_U80 ; P2_R1179_U186
g15718 nand P2_U3456 P2_R1179_U26 ; P2_R1179_U187
g15719 nand P2_U3465 P2_R1179_U32 ; P2_R1179_U188
g15720 nand P2_U3471 P2_R1179_U36 ; P2_R1179_U189
g15721 not P2_R1179_U61 ; P2_R1179_U190
g15722 not P2_R1179_U74 ; P2_R1179_U191
g15723 not P2_R1179_U34 ; P2_R1179_U192
g15724 not P2_R1179_U51 ; P2_R1179_U193
g15725 not P2_R1179_U166 ; P2_R1179_U194
g15726 nand P2_U3078 P2_R1179_U166 ; P2_R1179_U195
g15727 not P2_R1179_U43 ; P2_R1179_U196
g15728 nand P2_U3459 P2_R1179_U28 ; P2_R1179_U197
g15729 nand P2_R1179_U111 P2_R1179_U43 ; P2_R1179_U198
g15730 nand P2_R1179_U28 P2_R1179_U27 ; P2_R1179_U199
g15731 nand P2_R1179_U199 P2_R1179_U25 ; P2_R1179_U200
g15732 nand P2_U3064 P2_R1179_U181 ; P2_R1179_U201
g15733 not P2_R1179_U152 ; P2_R1179_U202
g15734 nand P2_U3468 P2_R1179_U31 ; P2_R1179_U203
g15735 nand P2_U3071 P2_R1179_U29 ; P2_R1179_U204
g15736 nand P2_U3067 P2_R1179_U21 ; P2_R1179_U205
g15737 nand P2_R1179_U192 P2_R1179_U188 ; P2_R1179_U206
g15738 nand P2_R1179_U6 P2_R1179_U206 ; P2_R1179_U207
g15739 nand P2_U3462 P2_R1179_U33 ; P2_R1179_U208
g15740 nand P2_U3468 P2_R1179_U31 ; P2_R1179_U209
g15741 nand P2_R1179_U152 P2_R1179_U113 ; P2_R1179_U210
g15742 nand P2_R1179_U209 P2_R1179_U207 ; P2_R1179_U211
g15743 not P2_R1179_U41 ; P2_R1179_U212
g15744 nand P2_U3474 P2_R1179_U38 ; P2_R1179_U213
g15745 nand P2_R1179_U114 P2_R1179_U41 ; P2_R1179_U214
g15746 nand P2_R1179_U38 P2_R1179_U37 ; P2_R1179_U215
g15747 nand P2_R1179_U215 P2_R1179_U35 ; P2_R1179_U216
g15748 nand P2_U3084 P2_R1179_U182 ; P2_R1179_U217
g15749 not P2_R1179_U148 ; P2_R1179_U218
g15750 nand P2_U3477 P2_R1179_U40 ; P2_R1179_U219
g15751 nand P2_R1179_U219 P2_R1179_U51 ; P2_R1179_U220
g15752 nand P2_R1179_U212 P2_R1179_U37 ; P2_R1179_U221
g15753 nand P2_R1179_U117 P2_R1179_U221 ; P2_R1179_U222
g15754 nand P2_R1179_U41 P2_R1179_U189 ; P2_R1179_U223
g15755 nand P2_R1179_U116 P2_R1179_U223 ; P2_R1179_U224
g15756 nand P2_R1179_U37 P2_R1179_U189 ; P2_R1179_U225
g15757 nand P2_R1179_U208 P2_R1179_U152 ; P2_R1179_U226
g15758 not P2_R1179_U42 ; P2_R1179_U227
g15759 nand P2_U3067 P2_R1179_U21 ; P2_R1179_U228
g15760 nand P2_R1179_U227 P2_R1179_U228 ; P2_R1179_U229
g15761 nand P2_R1179_U119 P2_R1179_U229 ; P2_R1179_U230
g15762 nand P2_R1179_U42 P2_R1179_U188 ; P2_R1179_U231
g15763 nand P2_U3468 P2_R1179_U31 ; P2_R1179_U232
g15764 nand P2_R1179_U118 P2_R1179_U231 ; P2_R1179_U233
g15765 nand P2_U3067 P2_R1179_U21 ; P2_R1179_U234
g15766 nand P2_R1179_U188 P2_R1179_U234 ; P2_R1179_U235
g15767 nand P2_R1179_U208 P2_R1179_U34 ; P2_R1179_U236
g15768 nand P2_R1179_U196 P2_R1179_U27 ; P2_R1179_U237
g15769 nand P2_R1179_U121 P2_R1179_U237 ; P2_R1179_U238
g15770 nand P2_R1179_U43 P2_R1179_U187 ; P2_R1179_U239
g15771 nand P2_R1179_U120 P2_R1179_U239 ; P2_R1179_U240
g15772 nand P2_R1179_U27 P2_R1179_U187 ; P2_R1179_U241
g15773 nand P2_U3483 P2_R1179_U49 ; P2_R1179_U242
g15774 nand P2_U3063 P2_R1179_U48 ; P2_R1179_U243
g15775 nand P2_U3062 P2_R1179_U47 ; P2_R1179_U244
g15776 nand P2_R1179_U193 P2_R1179_U183 ; P2_R1179_U245
g15777 nand P2_R1179_U7 P2_R1179_U245 ; P2_R1179_U246
g15778 nand P2_U3483 P2_R1179_U49 ; P2_R1179_U247
g15779 nand P2_R1179_U148 P2_R1179_U122 ; P2_R1179_U248
g15780 nand P2_R1179_U247 P2_R1179_U246 ; P2_R1179_U249
g15781 not P2_R1179_U175 ; P2_R1179_U250
g15782 nand P2_U3486 P2_R1179_U53 ; P2_R1179_U251
g15783 nand P2_R1179_U251 P2_R1179_U175 ; P2_R1179_U252
g15784 nand P2_U3072 P2_R1179_U52 ; P2_R1179_U253
g15785 not P2_R1179_U174 ; P2_R1179_U254
g15786 nand P2_U3489 P2_R1179_U55 ; P2_R1179_U255
g15787 nand P2_R1179_U255 P2_R1179_U174 ; P2_R1179_U256
g15788 nand P2_U3080 P2_R1179_U54 ; P2_R1179_U257
g15789 not P2_R1179_U173 ; P2_R1179_U258
g15790 nand P2_U3498 P2_R1179_U58 ; P2_R1179_U259
g15791 nand P2_U3073 P2_R1179_U56 ; P2_R1179_U260
g15792 nand P2_U3074 P2_R1179_U46 ; P2_R1179_U261
g15793 nand P2_R1179_U190 P2_R1179_U184 ; P2_R1179_U262
g15794 nand P2_R1179_U8 P2_R1179_U262 ; P2_R1179_U263
g15795 nand P2_U3492 P2_R1179_U60 ; P2_R1179_U264
g15796 nand P2_U3498 P2_R1179_U58 ; P2_R1179_U265
g15797 nand P2_R1179_U173 P2_R1179_U123 ; P2_R1179_U266
g15798 nand P2_R1179_U265 P2_R1179_U263 ; P2_R1179_U267
g15799 not P2_R1179_U170 ; P2_R1179_U268
g15800 nand P2_U3501 P2_R1179_U63 ; P2_R1179_U269
g15801 nand P2_R1179_U269 P2_R1179_U170 ; P2_R1179_U270
g15802 nand P2_U3069 P2_R1179_U62 ; P2_R1179_U271
g15803 not P2_R1179_U169 ; P2_R1179_U272
g15804 nand P2_U3082 P2_R1179_U169 ; P2_R1179_U273
g15805 not P2_R1179_U167 ; P2_R1179_U274
g15806 nand P2_U3506 P2_R1179_U66 ; P2_R1179_U275
g15807 nand P2_R1179_U275 P2_R1179_U167 ; P2_R1179_U276
g15808 nand P2_U3081 P2_R1179_U65 ; P2_R1179_U277
g15809 not P2_R1179_U164 ; P2_R1179_U278
g15810 nand P2_U3976 P2_R1179_U68 ; P2_R1179_U279
g15811 nand P2_R1179_U279 P2_R1179_U164 ; P2_R1179_U280
g15812 nand P2_U3076 P2_R1179_U67 ; P2_R1179_U281
g15813 not P2_R1179_U163 ; P2_R1179_U282
g15814 nand P2_U3973 P2_R1179_U71 ; P2_R1179_U283
g15815 nand P2_U3066 P2_R1179_U69 ; P2_R1179_U284
g15816 nand P2_U3061 P2_R1179_U45 ; P2_R1179_U285
g15817 nand P2_R1179_U191 P2_R1179_U185 ; P2_R1179_U286
g15818 nand P2_R1179_U9 P2_R1179_U286 ; P2_R1179_U287
g15819 nand P2_U3975 P2_R1179_U73 ; P2_R1179_U288
g15820 nand P2_U3973 P2_R1179_U71 ; P2_R1179_U289
g15821 nand P2_R1179_U163 P2_R1179_U124 ; P2_R1179_U290
g15822 nand P2_R1179_U289 P2_R1179_U287 ; P2_R1179_U291
g15823 not P2_R1179_U160 ; P2_R1179_U292
g15824 nand P2_U3972 P2_R1179_U76 ; P2_R1179_U293
g15825 nand P2_R1179_U293 P2_R1179_U160 ; P2_R1179_U294
g15826 nand P2_U3065 P2_R1179_U75 ; P2_R1179_U295
g15827 not P2_R1179_U159 ; P2_R1179_U296
g15828 nand P2_U3971 P2_R1179_U78 ; P2_R1179_U297
g15829 nand P2_R1179_U297 P2_R1179_U159 ; P2_R1179_U298
g15830 nand P2_U3058 P2_R1179_U77 ; P2_R1179_U299
g15831 not P2_R1179_U85 ; P2_R1179_U300
g15832 nand P2_U3969 P2_R1179_U82 ; P2_R1179_U301
g15833 nand P2_R1179_U125 P2_R1179_U85 ; P2_R1179_U302
g15834 nand P2_R1179_U82 P2_R1179_U81 ; P2_R1179_U303
g15835 nand P2_R1179_U303 P2_R1179_U79 ; P2_R1179_U304
g15836 nand P2_U3053 P2_R1179_U180 ; P2_R1179_U305
g15837 not P2_R1179_U157 ; P2_R1179_U306
g15838 nand P2_U3968 P2_R1179_U84 ; P2_R1179_U307
g15839 nand P2_U3054 P2_R1179_U83 ; P2_R1179_U308
g15840 nand P2_R1179_U300 P2_R1179_U81 ; P2_R1179_U309
g15841 nand P2_R1179_U131 P2_R1179_U309 ; P2_R1179_U310
g15842 nand P2_R1179_U85 P2_R1179_U186 ; P2_R1179_U311
g15843 nand P2_R1179_U130 P2_R1179_U311 ; P2_R1179_U312
g15844 nand P2_R1179_U81 P2_R1179_U186 ; P2_R1179_U313
g15845 nand P2_R1179_U288 P2_R1179_U163 ; P2_R1179_U314
g15846 not P2_R1179_U86 ; P2_R1179_U315
g15847 nand P2_U3061 P2_R1179_U45 ; P2_R1179_U316
g15848 nand P2_R1179_U315 P2_R1179_U316 ; P2_R1179_U317
g15849 nand P2_R1179_U135 P2_R1179_U317 ; P2_R1179_U318
g15850 nand P2_R1179_U86 P2_R1179_U185 ; P2_R1179_U319
g15851 nand P2_U3973 P2_R1179_U71 ; P2_R1179_U320
g15852 nand P2_R1179_U134 P2_R1179_U319 ; P2_R1179_U321
g15853 nand P2_U3061 P2_R1179_U45 ; P2_R1179_U322
g15854 nand P2_R1179_U185 P2_R1179_U322 ; P2_R1179_U323
g15855 nand P2_R1179_U288 P2_R1179_U74 ; P2_R1179_U324
g15856 nand P2_R1179_U264 P2_R1179_U173 ; P2_R1179_U325
g15857 not P2_R1179_U87 ; P2_R1179_U326
g15858 nand P2_U3074 P2_R1179_U46 ; P2_R1179_U327
g15859 nand P2_R1179_U326 P2_R1179_U327 ; P2_R1179_U328
g15860 nand P2_R1179_U142 P2_R1179_U328 ; P2_R1179_U329
g15861 nand P2_R1179_U87 P2_R1179_U184 ; P2_R1179_U330
g15862 nand P2_U3498 P2_R1179_U58 ; P2_R1179_U331
g15863 nand P2_R1179_U141 P2_R1179_U330 ; P2_R1179_U332
g15864 nand P2_U3074 P2_R1179_U46 ; P2_R1179_U333
g15865 nand P2_R1179_U184 P2_R1179_U333 ; P2_R1179_U334
g15866 nand P2_R1179_U264 P2_R1179_U61 ; P2_R1179_U335
g15867 nand P2_R1179_U219 P2_R1179_U148 ; P2_R1179_U336
g15868 not P2_R1179_U88 ; P2_R1179_U337
g15869 nand P2_U3062 P2_R1179_U47 ; P2_R1179_U338
g15870 nand P2_R1179_U337 P2_R1179_U338 ; P2_R1179_U339
g15871 nand P2_R1179_U146 P2_R1179_U339 ; P2_R1179_U340
g15872 nand P2_R1179_U88 P2_R1179_U183 ; P2_R1179_U341
g15873 nand P2_U3483 P2_R1179_U49 ; P2_R1179_U342
g15874 nand P2_R1179_U145 P2_R1179_U341 ; P2_R1179_U343
g15875 nand P2_U3062 P2_R1179_U47 ; P2_R1179_U344
g15876 nand P2_R1179_U183 P2_R1179_U344 ; P2_R1179_U345
g15877 nand P2_U3077 P2_R1179_U23 ; P2_R1179_U346
g15878 nand P2_U3078 P2_R1179_U165 ; P2_R1179_U347
g15879 nand P2_U3082 P2_R1179_U168 ; P2_R1179_U348
g15880 nand P2_R1179_U127 P2_R1179_U302 P2_R1179_U128 ; P2_R1179_U349
g15881 nand P2_U3477 P2_R1179_U40 ; P2_R1179_U350
g15882 nand P2_U3083 P2_R1179_U39 ; P2_R1179_U351
g15883 nand P2_R1179_U220 P2_R1179_U148 ; P2_R1179_U352
g15884 nand P2_R1179_U218 P2_R1179_U147 ; P2_R1179_U353
g15885 nand P2_U3474 P2_R1179_U38 ; P2_R1179_U354
g15886 nand P2_U3084 P2_R1179_U35 ; P2_R1179_U355
g15887 nand P2_U3474 P2_R1179_U38 ; P2_R1179_U356
g15888 nand P2_U3084 P2_R1179_U35 ; P2_R1179_U357
g15889 nand P2_R1179_U357 P2_R1179_U356 ; P2_R1179_U358
g15890 nand P2_U3471 P2_R1179_U36 ; P2_R1179_U359
g15891 nand P2_U3070 P2_R1179_U20 ; P2_R1179_U360
g15892 nand P2_R1179_U225 P2_R1179_U41 ; P2_R1179_U361
g15893 nand P2_R1179_U149 P2_R1179_U212 ; P2_R1179_U362
g15894 nand P2_U3468 P2_R1179_U31 ; P2_R1179_U363
g15895 nand P2_U3071 P2_R1179_U29 ; P2_R1179_U364
g15896 nand P2_R1179_U364 P2_R1179_U363 ; P2_R1179_U365
g15897 nand P2_U3465 P2_R1179_U32 ; P2_R1179_U366
g15898 nand P2_U3067 P2_R1179_U21 ; P2_R1179_U367
g15899 nand P2_R1179_U235 P2_R1179_U42 ; P2_R1179_U368
g15900 nand P2_R1179_U150 P2_R1179_U227 ; P2_R1179_U369
g15901 nand P2_U3462 P2_R1179_U33 ; P2_R1179_U370
g15902 nand P2_U3060 P2_R1179_U30 ; P2_R1179_U371
g15903 nand P2_R1179_U236 P2_R1179_U152 ; P2_R1179_U372
g15904 nand P2_R1179_U202 P2_R1179_U151 ; P2_R1179_U373
g15905 nand P2_U3459 P2_R1179_U28 ; P2_R1179_U374
g15906 nand P2_U3064 P2_R1179_U25 ; P2_R1179_U375
g15907 nand P2_U3459 P2_R1179_U28 ; P2_R1179_U376
g15908 nand P2_U3064 P2_R1179_U25 ; P2_R1179_U377
g15909 nand P2_R1179_U377 P2_R1179_U376 ; P2_R1179_U378
g15910 nand P2_U3456 P2_R1179_U26 ; P2_R1179_U379
g15911 nand P2_U3068 P2_R1179_U22 ; P2_R1179_U380
g15912 nand P2_R1179_U241 P2_R1179_U43 ; P2_R1179_U381
g15913 nand P2_R1179_U153 P2_R1179_U196 ; P2_R1179_U382
g15914 nand P2_U3979 P2_R1179_U155 ; P2_R1179_U383
g15915 nand P2_U3055 P2_R1179_U154 ; P2_R1179_U384
g15916 nand P2_U3979 P2_R1179_U155 ; P2_R1179_U385
g15917 nand P2_U3055 P2_R1179_U154 ; P2_R1179_U386
g15918 nand P2_R1179_U386 P2_R1179_U385 ; P2_R1179_U387
g15919 nand P2_U3968 P2_R1179_U10 P2_R1179_U84 ; P2_R1179_U388
g15920 nand P2_R1179_U387 P2_R1179_U83 P2_U3054 ; P2_R1179_U389
g15921 nand P2_U3968 P2_R1179_U84 ; P2_R1179_U390
g15922 nand P2_U3054 P2_R1179_U83 ; P2_R1179_U391
g15923 not P2_R1179_U129 ; P2_R1179_U392
g15924 nand P2_R1179_U306 P2_R1179_U392 ; P2_R1179_U393
g15925 nand P2_R1179_U129 P2_R1179_U157 ; P2_R1179_U394
g15926 nand P2_U3969 P2_R1179_U82 ; P2_R1179_U395
g15927 nand P2_U3053 P2_R1179_U79 ; P2_R1179_U396
g15928 nand P2_U3969 P2_R1179_U82 ; P2_R1179_U397
g15929 nand P2_U3053 P2_R1179_U79 ; P2_R1179_U398
g15930 nand P2_R1179_U398 P2_R1179_U397 ; P2_R1179_U399
g15931 nand P2_U3970 P2_R1179_U80 ; P2_R1179_U400
g15932 nand P2_U3057 P2_R1179_U44 ; P2_R1179_U401
g15933 nand P2_R1179_U313 P2_R1179_U85 ; P2_R1179_U402
g15934 nand P2_R1179_U158 P2_R1179_U300 ; P2_R1179_U403
g15935 nand P2_U3971 P2_R1179_U78 ; P2_R1179_U404
g15936 nand P2_U3058 P2_R1179_U77 ; P2_R1179_U405
g15937 not P2_R1179_U132 ; P2_R1179_U406
g15938 nand P2_R1179_U296 P2_R1179_U406 ; P2_R1179_U407
g15939 nand P2_R1179_U132 P2_R1179_U159 ; P2_R1179_U408
g15940 nand P2_U3972 P2_R1179_U76 ; P2_R1179_U409
g15941 nand P2_U3065 P2_R1179_U75 ; P2_R1179_U410
g15942 not P2_R1179_U133 ; P2_R1179_U411
g15943 nand P2_R1179_U292 P2_R1179_U411 ; P2_R1179_U412
g15944 nand P2_R1179_U133 P2_R1179_U160 ; P2_R1179_U413
g15945 nand P2_U3973 P2_R1179_U71 ; P2_R1179_U414
g15946 nand P2_U3066 P2_R1179_U69 ; P2_R1179_U415
g15947 nand P2_R1179_U415 P2_R1179_U414 ; P2_R1179_U416
g15948 nand P2_U3974 P2_R1179_U72 ; P2_R1179_U417
g15949 nand P2_U3061 P2_R1179_U45 ; P2_R1179_U418
g15950 nand P2_R1179_U323 P2_R1179_U86 ; P2_R1179_U419
g15951 nand P2_R1179_U161 P2_R1179_U315 ; P2_R1179_U420
g15952 nand P2_U3975 P2_R1179_U73 ; P2_R1179_U421
g15953 nand P2_U3075 P2_R1179_U70 ; P2_R1179_U422
g15954 nand P2_R1179_U324 P2_R1179_U163 ; P2_R1179_U423
g15955 nand P2_R1179_U282 P2_R1179_U162 ; P2_R1179_U424
g15956 nand P2_U3976 P2_R1179_U68 ; P2_R1179_U425
g15957 nand P2_U3076 P2_R1179_U67 ; P2_R1179_U426
g15958 not P2_R1179_U136 ; P2_R1179_U427
g15959 nand P2_R1179_U278 P2_R1179_U427 ; P2_R1179_U428
g15960 nand P2_R1179_U136 P2_R1179_U164 ; P2_R1179_U429
g15961 nand P2_U3453 P2_R1179_U24 ; P2_R1179_U430
g15962 nand P2_U3078 P2_R1179_U165 ; P2_R1179_U431
g15963 not P2_R1179_U137 ; P2_R1179_U432
g15964 nand P2_R1179_U194 P2_R1179_U432 ; P2_R1179_U433
g15965 nand P2_R1179_U137 P2_R1179_U166 ; P2_R1179_U434
g15966 nand P2_U3506 P2_R1179_U66 ; P2_R1179_U435
g15967 nand P2_U3081 P2_R1179_U65 ; P2_R1179_U436
g15968 not P2_R1179_U138 ; P2_R1179_U437
g15969 nand P2_R1179_U274 P2_R1179_U437 ; P2_R1179_U438
g15970 nand P2_R1179_U138 P2_R1179_U167 ; P2_R1179_U439
g15971 nand P2_U3504 P2_R1179_U64 ; P2_R1179_U440
g15972 nand P2_U3082 P2_R1179_U168 ; P2_R1179_U441
g15973 not P2_R1179_U139 ; P2_R1179_U442
g15974 nand P2_R1179_U272 P2_R1179_U442 ; P2_R1179_U443
g15975 nand P2_R1179_U139 P2_R1179_U169 ; P2_R1179_U444
g15976 nand P2_U3501 P2_R1179_U63 ; P2_R1179_U445
g15977 nand P2_U3069 P2_R1179_U62 ; P2_R1179_U446
g15978 not P2_R1179_U140 ; P2_R1179_U447
g15979 nand P2_R1179_U268 P2_R1179_U447 ; P2_R1179_U448
g15980 nand P2_R1179_U140 P2_R1179_U170 ; P2_R1179_U449
g15981 nand P2_U3498 P2_R1179_U58 ; P2_R1179_U450
g15982 nand P2_U3073 P2_R1179_U56 ; P2_R1179_U451
g15983 nand P2_R1179_U451 P2_R1179_U450 ; P2_R1179_U452
g15984 nand P2_U3495 P2_R1179_U59 ; P2_R1179_U453
g15985 nand P2_U3074 P2_R1179_U46 ; P2_R1179_U454
g15986 nand P2_R1179_U334 P2_R1179_U87 ; P2_R1179_U455
g15987 nand P2_R1179_U171 P2_R1179_U326 ; P2_R1179_U456
g15988 nand P2_U3492 P2_R1179_U60 ; P2_R1179_U457
g15989 nand P2_U3079 P2_R1179_U57 ; P2_R1179_U458
g15990 nand P2_R1179_U335 P2_R1179_U173 ; P2_R1179_U459
g15991 nand P2_R1179_U258 P2_R1179_U172 ; P2_R1179_U460
g15992 nand P2_U3489 P2_R1179_U55 ; P2_R1179_U461
g15993 nand P2_U3080 P2_R1179_U54 ; P2_R1179_U462
g15994 not P2_R1179_U143 ; P2_R1179_U463
g15995 nand P2_R1179_U254 P2_R1179_U463 ; P2_R1179_U464
g15996 nand P2_R1179_U143 P2_R1179_U174 ; P2_R1179_U465
g15997 nand P2_U3486 P2_R1179_U53 ; P2_R1179_U466
g15998 nand P2_U3072 P2_R1179_U52 ; P2_R1179_U467
g15999 not P2_R1179_U144 ; P2_R1179_U468
g16000 nand P2_R1179_U250 P2_R1179_U468 ; P2_R1179_U469
g16001 nand P2_R1179_U144 P2_R1179_U175 ; P2_R1179_U470
g16002 nand P2_U3483 P2_R1179_U49 ; P2_R1179_U471
g16003 nand P2_U3063 P2_R1179_U48 ; P2_R1179_U472
g16004 nand P2_R1179_U472 P2_R1179_U471 ; P2_R1179_U473
g16005 nand P2_U3480 P2_R1179_U50 ; P2_R1179_U474
g16006 nand P2_U3062 P2_R1179_U47 ; P2_R1179_U475
g16007 nand P2_R1179_U345 P2_R1179_U88 ; P2_R1179_U476
g16008 nand P2_R1179_U176 P2_R1179_U337 ; P2_R1179_U477
g16009 and P2_R1215_U179 P2_R1215_U178 ; P2_R1215_U4
g16010 and P2_R1215_U197 P2_R1215_U196 ; P2_R1215_U5
g16011 and P2_R1215_U237 P2_R1215_U236 ; P2_R1215_U6
g16012 and P2_R1215_U246 P2_R1215_U245 ; P2_R1215_U7
g16013 and P2_R1215_U264 P2_R1215_U263 ; P2_R1215_U8
g16014 and P2_R1215_U272 P2_R1215_U271 ; P2_R1215_U9
g16015 and P2_R1215_U351 P2_R1215_U348 ; P2_R1215_U10
g16016 and P2_R1215_U344 P2_R1215_U341 ; P2_R1215_U11
g16017 and P2_R1215_U335 P2_R1215_U332 ; P2_R1215_U12
g16018 and P2_R1215_U326 P2_R1215_U323 ; P2_R1215_U13
g16019 and P2_R1215_U320 P2_R1215_U318 ; P2_R1215_U14
g16020 and P2_R1215_U313 P2_R1215_U310 ; P2_R1215_U15
g16021 and P2_R1215_U235 P2_R1215_U232 ; P2_R1215_U16
g16022 and P2_R1215_U227 P2_R1215_U224 ; P2_R1215_U17
g16023 and P2_R1215_U213 P2_R1215_U210 ; P2_R1215_U18
g16024 not P2_U3468 ; P2_R1215_U19
g16025 not P2_U3071 ; P2_R1215_U20
g16026 not P2_U3070 ; P2_R1215_U21
g16027 nand P2_U3071 P2_U3468 ; P2_R1215_U22
g16028 not P2_U3471 ; P2_R1215_U23
g16029 not P2_U3462 ; P2_R1215_U24
g16030 not P2_U3060 ; P2_R1215_U25
g16031 not P2_U3067 ; P2_R1215_U26
g16032 not P2_U3456 ; P2_R1215_U27
g16033 not P2_U3068 ; P2_R1215_U28
g16034 not P2_U3448 ; P2_R1215_U29
g16035 not P2_U3077 ; P2_R1215_U30
g16036 nand P2_U3077 P2_U3448 ; P2_R1215_U31
g16037 not P2_U3459 ; P2_R1215_U32
g16038 not P2_U3064 ; P2_R1215_U33
g16039 nand P2_U3060 P2_U3462 ; P2_R1215_U34
g16040 not P2_U3465 ; P2_R1215_U35
g16041 not P2_U3474 ; P2_R1215_U36
g16042 not P2_U3084 ; P2_R1215_U37
g16043 not P2_U3083 ; P2_R1215_U38
g16044 not P2_U3477 ; P2_R1215_U39
g16045 nand P2_R1215_U61 P2_R1215_U205 ; P2_R1215_U40
g16046 nand P2_R1215_U117 P2_R1215_U193 ; P2_R1215_U41
g16047 nand P2_R1215_U182 P2_R1215_U183 ; P2_R1215_U42
g16048 nand P2_U3453 P2_U3078 ; P2_R1215_U43
g16049 nand P2_R1215_U122 P2_R1215_U219 ; P2_R1215_U44
g16050 nand P2_R1215_U216 P2_R1215_U215 ; P2_R1215_U45
g16051 not P2_U3969 ; P2_R1215_U46
g16052 not P2_U3053 ; P2_R1215_U47
g16053 not P2_U3057 ; P2_R1215_U48
g16054 not P2_U3970 ; P2_R1215_U49
g16055 not P2_U3971 ; P2_R1215_U50
g16056 not P2_U3058 ; P2_R1215_U51
g16057 not P2_U3972 ; P2_R1215_U52
g16058 not P2_U3065 ; P2_R1215_U53
g16059 not P2_U3975 ; P2_R1215_U54
g16060 not P2_U3075 ; P2_R1215_U55
g16061 not P2_U3498 ; P2_R1215_U56
g16062 not P2_U3073 ; P2_R1215_U57
g16063 not P2_U3069 ; P2_R1215_U58
g16064 nand P2_U3073 P2_U3498 ; P2_R1215_U59
g16065 not P2_U3501 ; P2_R1215_U60
g16066 nand P2_U3084 P2_U3474 ; P2_R1215_U61
g16067 not P2_U3480 ; P2_R1215_U62
g16068 not P2_U3062 ; P2_R1215_U63
g16069 not P2_U3486 ; P2_R1215_U64
g16070 not P2_U3072 ; P2_R1215_U65
g16071 not P2_U3483 ; P2_R1215_U66
g16072 not P2_U3063 ; P2_R1215_U67
g16073 nand P2_U3063 P2_U3483 ; P2_R1215_U68
g16074 not P2_U3489 ; P2_R1215_U69
g16075 not P2_U3080 ; P2_R1215_U70
g16076 not P2_U3492 ; P2_R1215_U71
g16077 not P2_U3079 ; P2_R1215_U72
g16078 not P2_U3495 ; P2_R1215_U73
g16079 not P2_U3074 ; P2_R1215_U74
g16080 not P2_U3504 ; P2_R1215_U75
g16081 not P2_U3082 ; P2_R1215_U76
g16082 nand P2_U3082 P2_U3504 ; P2_R1215_U77
g16083 not P2_U3506 ; P2_R1215_U78
g16084 not P2_U3081 ; P2_R1215_U79
g16085 nand P2_U3081 P2_U3506 ; P2_R1215_U80
g16086 not P2_U3976 ; P2_R1215_U81
g16087 not P2_U3974 ; P2_R1215_U82
g16088 not P2_U3061 ; P2_R1215_U83
g16089 not P2_U3973 ; P2_R1215_U84
g16090 not P2_U3066 ; P2_R1215_U85
g16091 nand P2_U3970 P2_U3057 ; P2_R1215_U86
g16092 not P2_U3054 ; P2_R1215_U87
g16093 not P2_U3968 ; P2_R1215_U88
g16094 nand P2_R1215_U306 P2_R1215_U176 ; P2_R1215_U89
g16095 not P2_U3076 ; P2_R1215_U90
g16096 nand P2_R1215_U77 P2_R1215_U315 ; P2_R1215_U91
g16097 nand P2_R1215_U261 P2_R1215_U260 ; P2_R1215_U92
g16098 nand P2_R1215_U68 P2_R1215_U337 ; P2_R1215_U93
g16099 nand P2_R1215_U457 P2_R1215_U456 ; P2_R1215_U94
g16100 nand P2_R1215_U504 P2_R1215_U503 ; P2_R1215_U95
g16101 nand P2_R1215_U375 P2_R1215_U374 ; P2_R1215_U96
g16102 nand P2_R1215_U380 P2_R1215_U379 ; P2_R1215_U97
g16103 nand P2_R1215_U387 P2_R1215_U386 ; P2_R1215_U98
g16104 nand P2_R1215_U394 P2_R1215_U393 ; P2_R1215_U99
g16105 nand P2_R1215_U399 P2_R1215_U398 ; P2_R1215_U100
g16106 nand P2_R1215_U408 P2_R1215_U407 ; P2_R1215_U101
g16107 nand P2_R1215_U415 P2_R1215_U414 ; P2_R1215_U102
g16108 nand P2_R1215_U422 P2_R1215_U421 ; P2_R1215_U103
g16109 nand P2_R1215_U429 P2_R1215_U428 ; P2_R1215_U104
g16110 nand P2_R1215_U434 P2_R1215_U433 ; P2_R1215_U105
g16111 nand P2_R1215_U441 P2_R1215_U440 ; P2_R1215_U106
g16112 nand P2_R1215_U448 P2_R1215_U447 ; P2_R1215_U107
g16113 nand P2_R1215_U462 P2_R1215_U461 ; P2_R1215_U108
g16114 nand P2_R1215_U467 P2_R1215_U466 ; P2_R1215_U109
g16115 nand P2_R1215_U474 P2_R1215_U473 ; P2_R1215_U110
g16116 nand P2_R1215_U481 P2_R1215_U480 ; P2_R1215_U111
g16117 nand P2_R1215_U488 P2_R1215_U487 ; P2_R1215_U112
g16118 nand P2_R1215_U495 P2_R1215_U494 ; P2_R1215_U113
g16119 nand P2_R1215_U500 P2_R1215_U499 ; P2_R1215_U114
g16120 and P2_R1215_U189 P2_R1215_U187 ; P2_R1215_U115
g16121 and P2_R1215_U4 P2_R1215_U180 ; P2_R1215_U116
g16122 and P2_R1215_U194 P2_R1215_U192 ; P2_R1215_U117
g16123 and P2_R1215_U201 P2_R1215_U200 ; P2_R1215_U118
g16124 and P2_R1215_U382 P2_R1215_U381 P2_R1215_U22 ; P2_R1215_U119
g16125 and P2_R1215_U212 P2_R1215_U5 ; P2_R1215_U120
g16126 and P2_R1215_U181 P2_R1215_U180 ; P2_R1215_U121
g16127 and P2_R1215_U220 P2_R1215_U218 ; P2_R1215_U122
g16128 and P2_R1215_U389 P2_R1215_U388 P2_R1215_U34 ; P2_R1215_U123
g16129 and P2_R1215_U226 P2_R1215_U4 ; P2_R1215_U124
g16130 and P2_R1215_U234 P2_R1215_U181 ; P2_R1215_U125
g16131 and P2_R1215_U204 P2_R1215_U6 ; P2_R1215_U126
g16132 and P2_R1215_U239 P2_R1215_U171 ; P2_R1215_U127
g16133 and P2_R1215_U250 P2_R1215_U7 ; P2_R1215_U128
g16134 and P2_R1215_U248 P2_R1215_U172 ; P2_R1215_U129
g16135 and P2_R1215_U268 P2_R1215_U267 ; P2_R1215_U130
g16136 and P2_R1215_U9 P2_R1215_U282 P2_R1215_U273 ; P2_R1215_U131
g16137 and P2_R1215_U285 P2_R1215_U280 ; P2_R1215_U132
g16138 and P2_R1215_U301 P2_R1215_U298 ; P2_R1215_U133
g16139 and P2_R1215_U368 P2_R1215_U302 ; P2_R1215_U134
g16140 and P2_R1215_U424 P2_R1215_U423 P2_R1215_U173 ; P2_R1215_U135
g16141 and P2_R1215_U160 P2_R1215_U278 ; P2_R1215_U136
g16142 and P2_R1215_U455 P2_R1215_U454 P2_R1215_U80 ; P2_R1215_U137
g16143 and P2_R1215_U325 P2_R1215_U9 ; P2_R1215_U138
g16144 and P2_R1215_U469 P2_R1215_U468 P2_R1215_U59 ; P2_R1215_U139
g16145 and P2_R1215_U334 P2_R1215_U8 ; P2_R1215_U140
g16146 and P2_R1215_U490 P2_R1215_U489 P2_R1215_U172 ; P2_R1215_U141
g16147 and P2_R1215_U343 P2_R1215_U7 ; P2_R1215_U142
g16148 and P2_R1215_U502 P2_R1215_U501 P2_R1215_U171 ; P2_R1215_U143
g16149 and P2_R1215_U350 P2_R1215_U6 ; P2_R1215_U144
g16150 nand P2_R1215_U118 P2_R1215_U202 ; P2_R1215_U145
g16151 nand P2_R1215_U217 P2_R1215_U229 ; P2_R1215_U146
g16152 not P2_U3055 ; P2_R1215_U147
g16153 not P2_U3979 ; P2_R1215_U148
g16154 and P2_R1215_U403 P2_R1215_U402 ; P2_R1215_U149
g16155 nand P2_R1215_U304 P2_R1215_U169 P2_R1215_U364 ; P2_R1215_U150
g16156 and P2_R1215_U410 P2_R1215_U409 ; P2_R1215_U151
g16157 nand P2_R1215_U370 P2_R1215_U369 P2_R1215_U134 ; P2_R1215_U152
g16158 and P2_R1215_U417 P2_R1215_U416 ; P2_R1215_U153
g16159 nand P2_R1215_U365 P2_R1215_U299 P2_R1215_U86 ; P2_R1215_U154
g16160 nand P2_R1215_U293 P2_R1215_U292 ; P2_R1215_U155
g16161 and P2_R1215_U436 P2_R1215_U435 ; P2_R1215_U156
g16162 nand P2_R1215_U289 P2_R1215_U288 ; P2_R1215_U157
g16163 and P2_R1215_U443 P2_R1215_U442 ; P2_R1215_U158
g16164 nand P2_R1215_U132 P2_R1215_U284 ; P2_R1215_U159
g16165 and P2_R1215_U450 P2_R1215_U449 ; P2_R1215_U160
g16166 nand P2_R1215_U43 P2_R1215_U327 ; P2_R1215_U161
g16167 nand P2_R1215_U130 P2_R1215_U269 ; P2_R1215_U162
g16168 and P2_R1215_U476 P2_R1215_U475 ; P2_R1215_U163
g16169 nand P2_R1215_U257 P2_R1215_U256 ; P2_R1215_U164
g16170 and P2_R1215_U483 P2_R1215_U482 ; P2_R1215_U165
g16171 nand P2_R1215_U253 P2_R1215_U252 ; P2_R1215_U166
g16172 nand P2_R1215_U243 P2_R1215_U242 ; P2_R1215_U167
g16173 nand P2_R1215_U367 P2_R1215_U366 ; P2_R1215_U168
g16174 nand P2_U3054 P2_R1215_U152 ; P2_R1215_U169
g16175 not P2_R1215_U34 ; P2_R1215_U170
g16176 nand P2_U3477 P2_U3083 ; P2_R1215_U171
g16177 nand P2_U3072 P2_U3486 ; P2_R1215_U172
g16178 nand P2_U3058 P2_U3971 ; P2_R1215_U173
g16179 not P2_R1215_U68 ; P2_R1215_U174
g16180 not P2_R1215_U77 ; P2_R1215_U175
g16181 nand P2_U3065 P2_U3972 ; P2_R1215_U176
g16182 not P2_R1215_U61 ; P2_R1215_U177
g16183 or P2_U3067 P2_U3465 ; P2_R1215_U178
g16184 or P2_U3060 P2_U3462 ; P2_R1215_U179
g16185 or P2_U3459 P2_U3064 ; P2_R1215_U180
g16186 or P2_U3456 P2_U3068 ; P2_R1215_U181
g16187 not P2_R1215_U31 ; P2_R1215_U182
g16188 or P2_U3453 P2_U3078 ; P2_R1215_U183
g16189 not P2_R1215_U42 ; P2_R1215_U184
g16190 not P2_R1215_U43 ; P2_R1215_U185
g16191 nand P2_R1215_U42 P2_R1215_U43 ; P2_R1215_U186
g16192 nand P2_U3068 P2_U3456 ; P2_R1215_U187
g16193 nand P2_R1215_U186 P2_R1215_U181 ; P2_R1215_U188
g16194 nand P2_U3064 P2_U3459 ; P2_R1215_U189
g16195 nand P2_R1215_U115 P2_R1215_U188 ; P2_R1215_U190
g16196 nand P2_R1215_U35 P2_R1215_U34 ; P2_R1215_U191
g16197 nand P2_U3067 P2_R1215_U191 ; P2_R1215_U192
g16198 nand P2_R1215_U116 P2_R1215_U190 ; P2_R1215_U193
g16199 nand P2_U3465 P2_R1215_U170 ; P2_R1215_U194
g16200 not P2_R1215_U41 ; P2_R1215_U195
g16201 or P2_U3070 P2_U3471 ; P2_R1215_U196
g16202 or P2_U3071 P2_U3468 ; P2_R1215_U197
g16203 not P2_R1215_U22 ; P2_R1215_U198
g16204 nand P2_R1215_U23 P2_R1215_U22 ; P2_R1215_U199
g16205 nand P2_U3070 P2_R1215_U199 ; P2_R1215_U200
g16206 nand P2_U3471 P2_R1215_U198 ; P2_R1215_U201
g16207 nand P2_R1215_U5 P2_R1215_U41 ; P2_R1215_U202
g16208 not P2_R1215_U145 ; P2_R1215_U203
g16209 or P2_U3474 P2_U3084 ; P2_R1215_U204
g16210 nand P2_R1215_U204 P2_R1215_U145 ; P2_R1215_U205
g16211 not P2_R1215_U40 ; P2_R1215_U206
g16212 or P2_U3083 P2_U3477 ; P2_R1215_U207
g16213 or P2_U3468 P2_U3071 ; P2_R1215_U208
g16214 nand P2_R1215_U208 P2_R1215_U41 ; P2_R1215_U209
g16215 nand P2_R1215_U119 P2_R1215_U209 ; P2_R1215_U210
g16216 nand P2_R1215_U195 P2_R1215_U22 ; P2_R1215_U211
g16217 nand P2_U3471 P2_U3070 ; P2_R1215_U212
g16218 nand P2_R1215_U120 P2_R1215_U211 ; P2_R1215_U213
g16219 or P2_U3071 P2_U3468 ; P2_R1215_U214
g16220 nand P2_R1215_U185 P2_R1215_U181 ; P2_R1215_U215
g16221 nand P2_U3068 P2_U3456 ; P2_R1215_U216
g16222 not P2_R1215_U45 ; P2_R1215_U217
g16223 nand P2_R1215_U121 P2_R1215_U184 ; P2_R1215_U218
g16224 nand P2_R1215_U45 P2_R1215_U180 ; P2_R1215_U219
g16225 nand P2_U3064 P2_U3459 ; P2_R1215_U220
g16226 not P2_R1215_U44 ; P2_R1215_U221
g16227 or P2_U3462 P2_U3060 ; P2_R1215_U222
g16228 nand P2_R1215_U222 P2_R1215_U44 ; P2_R1215_U223
g16229 nand P2_R1215_U123 P2_R1215_U223 ; P2_R1215_U224
g16230 nand P2_R1215_U221 P2_R1215_U34 ; P2_R1215_U225
g16231 nand P2_U3465 P2_U3067 ; P2_R1215_U226
g16232 nand P2_R1215_U124 P2_R1215_U225 ; P2_R1215_U227
g16233 or P2_U3060 P2_U3462 ; P2_R1215_U228
g16234 nand P2_R1215_U184 P2_R1215_U181 ; P2_R1215_U229
g16235 not P2_R1215_U146 ; P2_R1215_U230
g16236 nand P2_U3064 P2_U3459 ; P2_R1215_U231
g16237 nand P2_R1215_U401 P2_R1215_U400 P2_R1215_U43 P2_R1215_U42 ; P2_R1215_U232
g16238 nand P2_R1215_U43 P2_R1215_U42 ; P2_R1215_U233
g16239 nand P2_U3068 P2_U3456 ; P2_R1215_U234
g16240 nand P2_R1215_U125 P2_R1215_U233 ; P2_R1215_U235
g16241 or P2_U3083 P2_U3477 ; P2_R1215_U236
g16242 or P2_U3062 P2_U3480 ; P2_R1215_U237
g16243 nand P2_R1215_U177 P2_R1215_U6 ; P2_R1215_U238
g16244 nand P2_U3062 P2_U3480 ; P2_R1215_U239
g16245 nand P2_R1215_U127 P2_R1215_U238 ; P2_R1215_U240
g16246 or P2_U3480 P2_U3062 ; P2_R1215_U241
g16247 nand P2_R1215_U126 P2_R1215_U145 ; P2_R1215_U242
g16248 nand P2_R1215_U241 P2_R1215_U240 ; P2_R1215_U243
g16249 not P2_R1215_U167 ; P2_R1215_U244
g16250 or P2_U3080 P2_U3489 ; P2_R1215_U245
g16251 or P2_U3072 P2_U3486 ; P2_R1215_U246
g16252 nand P2_R1215_U174 P2_R1215_U7 ; P2_R1215_U247
g16253 nand P2_U3080 P2_U3489 ; P2_R1215_U248
g16254 nand P2_R1215_U129 P2_R1215_U247 ; P2_R1215_U249
g16255 or P2_U3483 P2_U3063 ; P2_R1215_U250
g16256 or P2_U3489 P2_U3080 ; P2_R1215_U251
g16257 nand P2_R1215_U128 P2_R1215_U167 ; P2_R1215_U252
g16258 nand P2_R1215_U251 P2_R1215_U249 ; P2_R1215_U253
g16259 not P2_R1215_U166 ; P2_R1215_U254
g16260 or P2_U3492 P2_U3079 ; P2_R1215_U255
g16261 nand P2_R1215_U255 P2_R1215_U166 ; P2_R1215_U256
g16262 nand P2_U3079 P2_U3492 ; P2_R1215_U257
g16263 not P2_R1215_U164 ; P2_R1215_U258
g16264 or P2_U3495 P2_U3074 ; P2_R1215_U259
g16265 nand P2_R1215_U259 P2_R1215_U164 ; P2_R1215_U260
g16266 nand P2_U3074 P2_U3495 ; P2_R1215_U261
g16267 not P2_R1215_U92 ; P2_R1215_U262
g16268 or P2_U3069 P2_U3501 ; P2_R1215_U263
g16269 or P2_U3073 P2_U3498 ; P2_R1215_U264
g16270 not P2_R1215_U59 ; P2_R1215_U265
g16271 nand P2_R1215_U60 P2_R1215_U59 ; P2_R1215_U266
g16272 nand P2_U3069 P2_R1215_U266 ; P2_R1215_U267
g16273 nand P2_U3501 P2_R1215_U265 ; P2_R1215_U268
g16274 nand P2_R1215_U8 P2_R1215_U92 ; P2_R1215_U269
g16275 not P2_R1215_U162 ; P2_R1215_U270
g16276 or P2_U3076 P2_U3976 ; P2_R1215_U271
g16277 or P2_U3081 P2_U3506 ; P2_R1215_U272
g16278 or P2_U3075 P2_U3975 ; P2_R1215_U273
g16279 not P2_R1215_U80 ; P2_R1215_U274
g16280 nand P2_U3976 P2_R1215_U274 ; P2_R1215_U275
g16281 nand P2_R1215_U275 P2_R1215_U90 ; P2_R1215_U276
g16282 nand P2_R1215_U80 P2_R1215_U81 ; P2_R1215_U277
g16283 nand P2_R1215_U277 P2_R1215_U276 ; P2_R1215_U278
g16284 nand P2_R1215_U175 P2_R1215_U9 ; P2_R1215_U279
g16285 nand P2_U3075 P2_U3975 ; P2_R1215_U280
g16286 nand P2_R1215_U278 P2_R1215_U279 ; P2_R1215_U281
g16287 or P2_U3504 P2_U3082 ; P2_R1215_U282
g16288 or P2_U3975 P2_U3075 ; P2_R1215_U283
g16289 nand P2_R1215_U162 P2_R1215_U131 ; P2_R1215_U284
g16290 nand P2_R1215_U283 P2_R1215_U281 ; P2_R1215_U285
g16291 not P2_R1215_U159 ; P2_R1215_U286
g16292 or P2_U3974 P2_U3061 ; P2_R1215_U287
g16293 nand P2_R1215_U287 P2_R1215_U159 ; P2_R1215_U288
g16294 nand P2_U3061 P2_U3974 ; P2_R1215_U289
g16295 not P2_R1215_U157 ; P2_R1215_U290
g16296 or P2_U3973 P2_U3066 ; P2_R1215_U291
g16297 nand P2_R1215_U291 P2_R1215_U157 ; P2_R1215_U292
g16298 nand P2_U3066 P2_U3973 ; P2_R1215_U293
g16299 not P2_R1215_U155 ; P2_R1215_U294
g16300 or P2_U3058 P2_U3971 ; P2_R1215_U295
g16301 nand P2_R1215_U176 P2_R1215_U173 ; P2_R1215_U296
g16302 not P2_R1215_U86 ; P2_R1215_U297
g16303 or P2_U3972 P2_U3065 ; P2_R1215_U298
g16304 nand P2_R1215_U155 P2_R1215_U298 P2_R1215_U168 ; P2_R1215_U299
g16305 not P2_R1215_U154 ; P2_R1215_U300
g16306 or P2_U3969 P2_U3053 ; P2_R1215_U301
g16307 nand P2_U3053 P2_U3969 ; P2_R1215_U302
g16308 not P2_R1215_U152 ; P2_R1215_U303
g16309 nand P2_U3968 P2_R1215_U152 ; P2_R1215_U304
g16310 not P2_R1215_U150 ; P2_R1215_U305
g16311 nand P2_R1215_U298 P2_R1215_U155 ; P2_R1215_U306
g16312 not P2_R1215_U89 ; P2_R1215_U307
g16313 or P2_U3971 P2_U3058 ; P2_R1215_U308
g16314 nand P2_R1215_U308 P2_R1215_U89 ; P2_R1215_U309
g16315 nand P2_R1215_U135 P2_R1215_U309 ; P2_R1215_U310
g16316 nand P2_R1215_U307 P2_R1215_U173 ; P2_R1215_U311
g16317 nand P2_U3970 P2_U3057 ; P2_R1215_U312
g16318 nand P2_R1215_U311 P2_R1215_U312 P2_R1215_U168 ; P2_R1215_U313
g16319 or P2_U3058 P2_U3971 ; P2_R1215_U314
g16320 nand P2_R1215_U282 P2_R1215_U162 ; P2_R1215_U315
g16321 not P2_R1215_U91 ; P2_R1215_U316
g16322 nand P2_R1215_U9 P2_R1215_U91 ; P2_R1215_U317
g16323 nand P2_R1215_U136 P2_R1215_U317 ; P2_R1215_U318
g16324 nand P2_R1215_U317 P2_R1215_U278 ; P2_R1215_U319
g16325 nand P2_R1215_U453 P2_R1215_U319 ; P2_R1215_U320
g16326 or P2_U3506 P2_U3081 ; P2_R1215_U321
g16327 nand P2_R1215_U321 P2_R1215_U91 ; P2_R1215_U322
g16328 nand P2_R1215_U137 P2_R1215_U322 ; P2_R1215_U323
g16329 nand P2_R1215_U316 P2_R1215_U80 ; P2_R1215_U324
g16330 nand P2_U3076 P2_U3976 ; P2_R1215_U325
g16331 nand P2_R1215_U138 P2_R1215_U324 ; P2_R1215_U326
g16332 or P2_U3453 P2_U3078 ; P2_R1215_U327
g16333 not P2_R1215_U161 ; P2_R1215_U328
g16334 or P2_U3081 P2_U3506 ; P2_R1215_U329
g16335 or P2_U3498 P2_U3073 ; P2_R1215_U330
g16336 nand P2_R1215_U330 P2_R1215_U92 ; P2_R1215_U331
g16337 nand P2_R1215_U139 P2_R1215_U331 ; P2_R1215_U332
g16338 nand P2_R1215_U262 P2_R1215_U59 ; P2_R1215_U333
g16339 nand P2_U3501 P2_U3069 ; P2_R1215_U334
g16340 nand P2_R1215_U140 P2_R1215_U333 ; P2_R1215_U335
g16341 or P2_U3073 P2_U3498 ; P2_R1215_U336
g16342 nand P2_R1215_U250 P2_R1215_U167 ; P2_R1215_U337
g16343 not P2_R1215_U93 ; P2_R1215_U338
g16344 or P2_U3486 P2_U3072 ; P2_R1215_U339
g16345 nand P2_R1215_U339 P2_R1215_U93 ; P2_R1215_U340
g16346 nand P2_R1215_U141 P2_R1215_U340 ; P2_R1215_U341
g16347 nand P2_R1215_U338 P2_R1215_U172 ; P2_R1215_U342
g16348 nand P2_U3080 P2_U3489 ; P2_R1215_U343
g16349 nand P2_R1215_U142 P2_R1215_U342 ; P2_R1215_U344
g16350 or P2_U3072 P2_U3486 ; P2_R1215_U345
g16351 or P2_U3477 P2_U3083 ; P2_R1215_U346
g16352 nand P2_R1215_U346 P2_R1215_U40 ; P2_R1215_U347
g16353 nand P2_R1215_U143 P2_R1215_U347 ; P2_R1215_U348
g16354 nand P2_R1215_U206 P2_R1215_U171 ; P2_R1215_U349
g16355 nand P2_U3062 P2_U3480 ; P2_R1215_U350
g16356 nand P2_R1215_U144 P2_R1215_U349 ; P2_R1215_U351
g16357 nand P2_R1215_U207 P2_R1215_U171 ; P2_R1215_U352
g16358 nand P2_R1215_U204 P2_R1215_U61 ; P2_R1215_U353
g16359 nand P2_R1215_U214 P2_R1215_U22 ; P2_R1215_U354
g16360 nand P2_R1215_U228 P2_R1215_U34 ; P2_R1215_U355
g16361 nand P2_R1215_U231 P2_R1215_U180 ; P2_R1215_U356
g16362 nand P2_R1215_U314 P2_R1215_U173 ; P2_R1215_U357
g16363 nand P2_R1215_U298 P2_R1215_U176 ; P2_R1215_U358
g16364 nand P2_R1215_U329 P2_R1215_U80 ; P2_R1215_U359
g16365 nand P2_R1215_U282 P2_R1215_U77 ; P2_R1215_U360
g16366 nand P2_R1215_U336 P2_R1215_U59 ; P2_R1215_U361
g16367 nand P2_R1215_U345 P2_R1215_U172 ; P2_R1215_U362
g16368 nand P2_R1215_U250 P2_R1215_U68 ; P2_R1215_U363
g16369 nand P2_U3968 P2_U3054 ; P2_R1215_U364
g16370 nand P2_R1215_U296 P2_R1215_U168 ; P2_R1215_U365
g16371 nand P2_U3057 P2_R1215_U295 ; P2_R1215_U366
g16372 nand P2_U3970 P2_R1215_U295 ; P2_R1215_U367
g16373 nand P2_R1215_U296 P2_R1215_U168 P2_R1215_U301 ; P2_R1215_U368
g16374 nand P2_R1215_U155 P2_R1215_U168 P2_R1215_U133 ; P2_R1215_U369
g16375 nand P2_R1215_U297 P2_R1215_U301 ; P2_R1215_U370
g16376 nand P2_U3083 P2_R1215_U39 ; P2_R1215_U371
g16377 nand P2_U3477 P2_R1215_U38 ; P2_R1215_U372
g16378 nand P2_R1215_U372 P2_R1215_U371 ; P2_R1215_U373
g16379 nand P2_R1215_U352 P2_R1215_U40 ; P2_R1215_U374
g16380 nand P2_R1215_U373 P2_R1215_U206 ; P2_R1215_U375
g16381 nand P2_U3084 P2_R1215_U36 ; P2_R1215_U376
g16382 nand P2_U3474 P2_R1215_U37 ; P2_R1215_U377
g16383 nand P2_R1215_U377 P2_R1215_U376 ; P2_R1215_U378
g16384 nand P2_R1215_U353 P2_R1215_U145 ; P2_R1215_U379
g16385 nand P2_R1215_U203 P2_R1215_U378 ; P2_R1215_U380
g16386 nand P2_U3070 P2_R1215_U23 ; P2_R1215_U381
g16387 nand P2_U3471 P2_R1215_U21 ; P2_R1215_U382
g16388 nand P2_U3071 P2_R1215_U19 ; P2_R1215_U383
g16389 nand P2_U3468 P2_R1215_U20 ; P2_R1215_U384
g16390 nand P2_R1215_U384 P2_R1215_U383 ; P2_R1215_U385
g16391 nand P2_R1215_U354 P2_R1215_U41 ; P2_R1215_U386
g16392 nand P2_R1215_U385 P2_R1215_U195 ; P2_R1215_U387
g16393 nand P2_U3067 P2_R1215_U35 ; P2_R1215_U388
g16394 nand P2_U3465 P2_R1215_U26 ; P2_R1215_U389
g16395 nand P2_U3060 P2_R1215_U24 ; P2_R1215_U390
g16396 nand P2_U3462 P2_R1215_U25 ; P2_R1215_U391
g16397 nand P2_R1215_U391 P2_R1215_U390 ; P2_R1215_U392
g16398 nand P2_R1215_U355 P2_R1215_U44 ; P2_R1215_U393
g16399 nand P2_R1215_U392 P2_R1215_U221 ; P2_R1215_U394
g16400 nand P2_U3064 P2_R1215_U32 ; P2_R1215_U395
g16401 nand P2_U3459 P2_R1215_U33 ; P2_R1215_U396
g16402 nand P2_R1215_U396 P2_R1215_U395 ; P2_R1215_U397
g16403 nand P2_R1215_U356 P2_R1215_U146 ; P2_R1215_U398
g16404 nand P2_R1215_U230 P2_R1215_U397 ; P2_R1215_U399
g16405 nand P2_U3068 P2_R1215_U27 ; P2_R1215_U400
g16406 nand P2_U3456 P2_R1215_U28 ; P2_R1215_U401
g16407 nand P2_U3055 P2_R1215_U148 ; P2_R1215_U402
g16408 nand P2_U3979 P2_R1215_U147 ; P2_R1215_U403
g16409 nand P2_U3055 P2_R1215_U148 ; P2_R1215_U404
g16410 nand P2_U3979 P2_R1215_U147 ; P2_R1215_U405
g16411 nand P2_R1215_U405 P2_R1215_U404 ; P2_R1215_U406
g16412 nand P2_R1215_U149 P2_R1215_U150 ; P2_R1215_U407
g16413 nand P2_R1215_U305 P2_R1215_U406 ; P2_R1215_U408
g16414 nand P2_U3054 P2_R1215_U88 ; P2_R1215_U409
g16415 nand P2_U3968 P2_R1215_U87 ; P2_R1215_U410
g16416 nand P2_U3054 P2_R1215_U88 ; P2_R1215_U411
g16417 nand P2_U3968 P2_R1215_U87 ; P2_R1215_U412
g16418 nand P2_R1215_U412 P2_R1215_U411 ; P2_R1215_U413
g16419 nand P2_R1215_U151 P2_R1215_U152 ; P2_R1215_U414
g16420 nand P2_R1215_U303 P2_R1215_U413 ; P2_R1215_U415
g16421 nand P2_U3053 P2_R1215_U46 ; P2_R1215_U416
g16422 nand P2_U3969 P2_R1215_U47 ; P2_R1215_U417
g16423 nand P2_U3053 P2_R1215_U46 ; P2_R1215_U418
g16424 nand P2_U3969 P2_R1215_U47 ; P2_R1215_U419
g16425 nand P2_R1215_U419 P2_R1215_U418 ; P2_R1215_U420
g16426 nand P2_R1215_U153 P2_R1215_U154 ; P2_R1215_U421
g16427 nand P2_R1215_U300 P2_R1215_U420 ; P2_R1215_U422
g16428 nand P2_U3057 P2_R1215_U49 ; P2_R1215_U423
g16429 nand P2_U3970 P2_R1215_U48 ; P2_R1215_U424
g16430 nand P2_U3058 P2_R1215_U50 ; P2_R1215_U425
g16431 nand P2_U3971 P2_R1215_U51 ; P2_R1215_U426
g16432 nand P2_R1215_U426 P2_R1215_U425 ; P2_R1215_U427
g16433 nand P2_R1215_U357 P2_R1215_U89 ; P2_R1215_U428
g16434 nand P2_R1215_U427 P2_R1215_U307 ; P2_R1215_U429
g16435 nand P2_U3065 P2_R1215_U52 ; P2_R1215_U430
g16436 nand P2_U3972 P2_R1215_U53 ; P2_R1215_U431
g16437 nand P2_R1215_U431 P2_R1215_U430 ; P2_R1215_U432
g16438 nand P2_R1215_U358 P2_R1215_U155 ; P2_R1215_U433
g16439 nand P2_R1215_U294 P2_R1215_U432 ; P2_R1215_U434
g16440 nand P2_U3066 P2_R1215_U84 ; P2_R1215_U435
g16441 nand P2_U3973 P2_R1215_U85 ; P2_R1215_U436
g16442 nand P2_U3066 P2_R1215_U84 ; P2_R1215_U437
g16443 nand P2_U3973 P2_R1215_U85 ; P2_R1215_U438
g16444 nand P2_R1215_U438 P2_R1215_U437 ; P2_R1215_U439
g16445 nand P2_R1215_U156 P2_R1215_U157 ; P2_R1215_U440
g16446 nand P2_R1215_U290 P2_R1215_U439 ; P2_R1215_U441
g16447 nand P2_U3061 P2_R1215_U82 ; P2_R1215_U442
g16448 nand P2_U3974 P2_R1215_U83 ; P2_R1215_U443
g16449 nand P2_U3061 P2_R1215_U82 ; P2_R1215_U444
g16450 nand P2_U3974 P2_R1215_U83 ; P2_R1215_U445
g16451 nand P2_R1215_U445 P2_R1215_U444 ; P2_R1215_U446
g16452 nand P2_R1215_U158 P2_R1215_U159 ; P2_R1215_U447
g16453 nand P2_R1215_U286 P2_R1215_U446 ; P2_R1215_U448
g16454 nand P2_U3075 P2_R1215_U54 ; P2_R1215_U449
g16455 nand P2_U3975 P2_R1215_U55 ; P2_R1215_U450
g16456 nand P2_U3075 P2_R1215_U54 ; P2_R1215_U451
g16457 nand P2_U3975 P2_R1215_U55 ; P2_R1215_U452
g16458 nand P2_R1215_U452 P2_R1215_U451 ; P2_R1215_U453
g16459 nand P2_U3076 P2_R1215_U81 ; P2_R1215_U454
g16460 nand P2_U3976 P2_R1215_U90 ; P2_R1215_U455
g16461 nand P2_R1215_U182 P2_R1215_U161 ; P2_R1215_U456
g16462 nand P2_R1215_U328 P2_R1215_U31 ; P2_R1215_U457
g16463 nand P2_U3081 P2_R1215_U78 ; P2_R1215_U458
g16464 nand P2_U3506 P2_R1215_U79 ; P2_R1215_U459
g16465 nand P2_R1215_U459 P2_R1215_U458 ; P2_R1215_U460
g16466 nand P2_R1215_U359 P2_R1215_U91 ; P2_R1215_U461
g16467 nand P2_R1215_U460 P2_R1215_U316 ; P2_R1215_U462
g16468 nand P2_U3082 P2_R1215_U75 ; P2_R1215_U463
g16469 nand P2_U3504 P2_R1215_U76 ; P2_R1215_U464
g16470 nand P2_R1215_U464 P2_R1215_U463 ; P2_R1215_U465
g16471 nand P2_R1215_U360 P2_R1215_U162 ; P2_R1215_U466
g16472 nand P2_R1215_U270 P2_R1215_U465 ; P2_R1215_U467
g16473 nand P2_U3069 P2_R1215_U60 ; P2_R1215_U468
g16474 nand P2_U3501 P2_R1215_U58 ; P2_R1215_U469
g16475 nand P2_U3073 P2_R1215_U56 ; P2_R1215_U470
g16476 nand P2_U3498 P2_R1215_U57 ; P2_R1215_U471
g16477 nand P2_R1215_U471 P2_R1215_U470 ; P2_R1215_U472
g16478 nand P2_R1215_U361 P2_R1215_U92 ; P2_R1215_U473
g16479 nand P2_R1215_U472 P2_R1215_U262 ; P2_R1215_U474
g16480 nand P2_U3074 P2_R1215_U73 ; P2_R1215_U475
g16481 nand P2_U3495 P2_R1215_U74 ; P2_R1215_U476
g16482 nand P2_U3074 P2_R1215_U73 ; P2_R1215_U477
g16483 nand P2_U3495 P2_R1215_U74 ; P2_R1215_U478
g16484 nand P2_R1215_U478 P2_R1215_U477 ; P2_R1215_U479
g16485 nand P2_R1215_U163 P2_R1215_U164 ; P2_R1215_U480
g16486 nand P2_R1215_U258 P2_R1215_U479 ; P2_R1215_U481
g16487 nand P2_U3079 P2_R1215_U71 ; P2_R1215_U482
g16488 nand P2_U3492 P2_R1215_U72 ; P2_R1215_U483
g16489 nand P2_U3079 P2_R1215_U71 ; P2_R1215_U484
g16490 nand P2_U3492 P2_R1215_U72 ; P2_R1215_U485
g16491 nand P2_R1215_U485 P2_R1215_U484 ; P2_R1215_U486
g16492 nand P2_R1215_U165 P2_R1215_U166 ; P2_R1215_U487
g16493 nand P2_R1215_U254 P2_R1215_U486 ; P2_R1215_U488
g16494 nand P2_U3080 P2_R1215_U69 ; P2_R1215_U489
g16495 nand P2_U3489 P2_R1215_U70 ; P2_R1215_U490
g16496 nand P2_U3072 P2_R1215_U64 ; P2_R1215_U491
g16497 nand P2_U3486 P2_R1215_U65 ; P2_R1215_U492
g16498 nand P2_R1215_U492 P2_R1215_U491 ; P2_R1215_U493
g16499 nand P2_R1215_U362 P2_R1215_U93 ; P2_R1215_U494
g16500 nand P2_R1215_U493 P2_R1215_U338 ; P2_R1215_U495
g16501 nand P2_U3063 P2_R1215_U66 ; P2_R1215_U496
g16502 nand P2_U3483 P2_R1215_U67 ; P2_R1215_U497
g16503 nand P2_R1215_U497 P2_R1215_U496 ; P2_R1215_U498
g16504 nand P2_R1215_U363 P2_R1215_U167 ; P2_R1215_U499
g16505 nand P2_R1215_U244 P2_R1215_U498 ; P2_R1215_U500
g16506 nand P2_U3062 P2_R1215_U62 ; P2_R1215_U501
g16507 nand P2_U3480 P2_R1215_U63 ; P2_R1215_U502
g16508 nand P2_U3077 P2_R1215_U29 ; P2_R1215_U503
g16509 nand P2_U3448 P2_R1215_U30 ; P2_R1215_U504
g16510 and P2_R1164_U179 P2_R1164_U178 ; P2_R1164_U4
g16511 and P2_R1164_U197 P2_R1164_U196 ; P2_R1164_U5
g16512 and P2_R1164_U237 P2_R1164_U236 ; P2_R1164_U6
g16513 and P2_R1164_U246 P2_R1164_U245 ; P2_R1164_U7
g16514 and P2_R1164_U264 P2_R1164_U263 ; P2_R1164_U8
g16515 and P2_R1164_U272 P2_R1164_U271 ; P2_R1164_U9
g16516 and P2_R1164_U351 P2_R1164_U348 ; P2_R1164_U10
g16517 and P2_R1164_U344 P2_R1164_U341 ; P2_R1164_U11
g16518 and P2_R1164_U335 P2_R1164_U332 ; P2_R1164_U12
g16519 and P2_R1164_U326 P2_R1164_U323 ; P2_R1164_U13
g16520 and P2_R1164_U320 P2_R1164_U318 ; P2_R1164_U14
g16521 and P2_R1164_U313 P2_R1164_U310 ; P2_R1164_U15
g16522 and P2_R1164_U235 P2_R1164_U232 ; P2_R1164_U16
g16523 and P2_R1164_U227 P2_R1164_U224 ; P2_R1164_U17
g16524 and P2_R1164_U213 P2_R1164_U210 ; P2_R1164_U18
g16525 not P2_U3468 ; P2_R1164_U19
g16526 not P2_U3071 ; P2_R1164_U20
g16527 not P2_U3070 ; P2_R1164_U21
g16528 nand P2_U3071 P2_U3468 ; P2_R1164_U22
g16529 not P2_U3471 ; P2_R1164_U23
g16530 not P2_U3462 ; P2_R1164_U24
g16531 not P2_U3060 ; P2_R1164_U25
g16532 not P2_U3067 ; P2_R1164_U26
g16533 not P2_U3456 ; P2_R1164_U27
g16534 not P2_U3068 ; P2_R1164_U28
g16535 not P2_U3448 ; P2_R1164_U29
g16536 not P2_U3077 ; P2_R1164_U30
g16537 nand P2_U3077 P2_U3448 ; P2_R1164_U31
g16538 not P2_U3459 ; P2_R1164_U32
g16539 not P2_U3064 ; P2_R1164_U33
g16540 nand P2_U3060 P2_U3462 ; P2_R1164_U34
g16541 not P2_U3465 ; P2_R1164_U35
g16542 not P2_U3474 ; P2_R1164_U36
g16543 not P2_U3084 ; P2_R1164_U37
g16544 not P2_U3083 ; P2_R1164_U38
g16545 not P2_U3477 ; P2_R1164_U39
g16546 nand P2_R1164_U63 P2_R1164_U205 ; P2_R1164_U40
g16547 nand P2_R1164_U117 P2_R1164_U193 ; P2_R1164_U41
g16548 nand P2_R1164_U182 P2_R1164_U183 ; P2_R1164_U42
g16549 nand P2_U3453 P2_U3078 ; P2_R1164_U43
g16550 nand P2_R1164_U122 P2_R1164_U219 ; P2_R1164_U44
g16551 nand P2_R1164_U216 P2_R1164_U215 ; P2_R1164_U45
g16552 not P2_U3969 ; P2_R1164_U46
g16553 not P2_U3053 ; P2_R1164_U47
g16554 not P2_U3057 ; P2_R1164_U48
g16555 not P2_U3970 ; P2_R1164_U49
g16556 not P2_U3971 ; P2_R1164_U50
g16557 not P2_U3058 ; P2_R1164_U51
g16558 not P2_U3972 ; P2_R1164_U52
g16559 not P2_U3065 ; P2_R1164_U53
g16560 not P2_U3975 ; P2_R1164_U54
g16561 not P2_U3075 ; P2_R1164_U55
g16562 not P2_U3498 ; P2_R1164_U56
g16563 not P2_U3073 ; P2_R1164_U57
g16564 not P2_U3069 ; P2_R1164_U58
g16565 nand P2_U3073 P2_U3498 ; P2_R1164_U59
g16566 not P2_U3501 ; P2_R1164_U60
g16567 not P2_U3480 ; P2_R1164_U61
g16568 not P2_U3062 ; P2_R1164_U62
g16569 nand P2_U3084 P2_U3474 ; P2_R1164_U63
g16570 not P2_U3486 ; P2_R1164_U64
g16571 not P2_U3072 ; P2_R1164_U65
g16572 not P2_U3483 ; P2_R1164_U66
g16573 not P2_U3063 ; P2_R1164_U67
g16574 nand P2_U3063 P2_U3483 ; P2_R1164_U68
g16575 not P2_U3489 ; P2_R1164_U69
g16576 not P2_U3080 ; P2_R1164_U70
g16577 not P2_U3492 ; P2_R1164_U71
g16578 not P2_U3079 ; P2_R1164_U72
g16579 not P2_U3495 ; P2_R1164_U73
g16580 not P2_U3074 ; P2_R1164_U74
g16581 not P2_U3504 ; P2_R1164_U75
g16582 not P2_U3082 ; P2_R1164_U76
g16583 nand P2_U3082 P2_U3504 ; P2_R1164_U77
g16584 not P2_U3506 ; P2_R1164_U78
g16585 not P2_U3081 ; P2_R1164_U79
g16586 nand P2_U3081 P2_U3506 ; P2_R1164_U80
g16587 not P2_U3976 ; P2_R1164_U81
g16588 not P2_U3974 ; P2_R1164_U82
g16589 not P2_U3061 ; P2_R1164_U83
g16590 not P2_U3973 ; P2_R1164_U84
g16591 not P2_U3066 ; P2_R1164_U85
g16592 nand P2_U3970 P2_U3057 ; P2_R1164_U86
g16593 not P2_U3054 ; P2_R1164_U87
g16594 not P2_U3968 ; P2_R1164_U88
g16595 nand P2_R1164_U306 P2_R1164_U176 ; P2_R1164_U89
g16596 not P2_U3076 ; P2_R1164_U90
g16597 nand P2_R1164_U77 P2_R1164_U315 ; P2_R1164_U91
g16598 nand P2_R1164_U261 P2_R1164_U260 ; P2_R1164_U92
g16599 nand P2_R1164_U68 P2_R1164_U337 ; P2_R1164_U93
g16600 nand P2_R1164_U457 P2_R1164_U456 ; P2_R1164_U94
g16601 nand P2_R1164_U504 P2_R1164_U503 ; P2_R1164_U95
g16602 nand P2_R1164_U375 P2_R1164_U374 ; P2_R1164_U96
g16603 nand P2_R1164_U380 P2_R1164_U379 ; P2_R1164_U97
g16604 nand P2_R1164_U387 P2_R1164_U386 ; P2_R1164_U98
g16605 nand P2_R1164_U394 P2_R1164_U393 ; P2_R1164_U99
g16606 nand P2_R1164_U399 P2_R1164_U398 ; P2_R1164_U100
g16607 nand P2_R1164_U408 P2_R1164_U407 ; P2_R1164_U101
g16608 nand P2_R1164_U415 P2_R1164_U414 ; P2_R1164_U102
g16609 nand P2_R1164_U422 P2_R1164_U421 ; P2_R1164_U103
g16610 nand P2_R1164_U429 P2_R1164_U428 ; P2_R1164_U104
g16611 nand P2_R1164_U434 P2_R1164_U433 ; P2_R1164_U105
g16612 nand P2_R1164_U441 P2_R1164_U440 ; P2_R1164_U106
g16613 nand P2_R1164_U448 P2_R1164_U447 ; P2_R1164_U107
g16614 nand P2_R1164_U462 P2_R1164_U461 ; P2_R1164_U108
g16615 nand P2_R1164_U467 P2_R1164_U466 ; P2_R1164_U109
g16616 nand P2_R1164_U474 P2_R1164_U473 ; P2_R1164_U110
g16617 nand P2_R1164_U481 P2_R1164_U480 ; P2_R1164_U111
g16618 nand P2_R1164_U488 P2_R1164_U487 ; P2_R1164_U112
g16619 nand P2_R1164_U495 P2_R1164_U494 ; P2_R1164_U113
g16620 nand P2_R1164_U500 P2_R1164_U499 ; P2_R1164_U114
g16621 and P2_R1164_U189 P2_R1164_U187 ; P2_R1164_U115
g16622 and P2_R1164_U4 P2_R1164_U180 ; P2_R1164_U116
g16623 and P2_R1164_U194 P2_R1164_U192 ; P2_R1164_U117
g16624 and P2_R1164_U201 P2_R1164_U200 ; P2_R1164_U118
g16625 and P2_R1164_U382 P2_R1164_U381 P2_R1164_U22 ; P2_R1164_U119
g16626 and P2_R1164_U212 P2_R1164_U5 ; P2_R1164_U120
g16627 and P2_R1164_U181 P2_R1164_U180 ; P2_R1164_U121
g16628 and P2_R1164_U220 P2_R1164_U218 ; P2_R1164_U122
g16629 and P2_R1164_U389 P2_R1164_U388 P2_R1164_U34 ; P2_R1164_U123
g16630 and P2_R1164_U226 P2_R1164_U4 ; P2_R1164_U124
g16631 and P2_R1164_U234 P2_R1164_U181 ; P2_R1164_U125
g16632 and P2_R1164_U204 P2_R1164_U6 ; P2_R1164_U126
g16633 and P2_R1164_U243 P2_R1164_U239 ; P2_R1164_U127
g16634 and P2_R1164_U250 P2_R1164_U7 ; P2_R1164_U128
g16635 and P2_R1164_U248 P2_R1164_U172 ; P2_R1164_U129
g16636 and P2_R1164_U268 P2_R1164_U267 ; P2_R1164_U130
g16637 and P2_R1164_U9 P2_R1164_U282 P2_R1164_U273 ; P2_R1164_U131
g16638 and P2_R1164_U285 P2_R1164_U280 ; P2_R1164_U132
g16639 and P2_R1164_U301 P2_R1164_U298 ; P2_R1164_U133
g16640 and P2_R1164_U368 P2_R1164_U302 ; P2_R1164_U134
g16641 and P2_R1164_U424 P2_R1164_U423 P2_R1164_U173 ; P2_R1164_U135
g16642 and P2_R1164_U160 P2_R1164_U278 ; P2_R1164_U136
g16643 and P2_R1164_U455 P2_R1164_U454 P2_R1164_U80 ; P2_R1164_U137
g16644 and P2_R1164_U325 P2_R1164_U9 ; P2_R1164_U138
g16645 and P2_R1164_U469 P2_R1164_U468 P2_R1164_U59 ; P2_R1164_U139
g16646 and P2_R1164_U334 P2_R1164_U8 ; P2_R1164_U140
g16647 and P2_R1164_U490 P2_R1164_U489 P2_R1164_U172 ; P2_R1164_U141
g16648 and P2_R1164_U343 P2_R1164_U7 ; P2_R1164_U142
g16649 and P2_R1164_U502 P2_R1164_U501 P2_R1164_U171 ; P2_R1164_U143
g16650 and P2_R1164_U350 P2_R1164_U6 ; P2_R1164_U144
g16651 nand P2_R1164_U118 P2_R1164_U202 ; P2_R1164_U145
g16652 nand P2_R1164_U217 P2_R1164_U229 ; P2_R1164_U146
g16653 not P2_U3055 ; P2_R1164_U147
g16654 not P2_U3979 ; P2_R1164_U148
g16655 and P2_R1164_U403 P2_R1164_U402 ; P2_R1164_U149
g16656 nand P2_R1164_U304 P2_R1164_U169 P2_R1164_U364 ; P2_R1164_U150
g16657 and P2_R1164_U410 P2_R1164_U409 ; P2_R1164_U151
g16658 nand P2_R1164_U370 P2_R1164_U369 P2_R1164_U134 ; P2_R1164_U152
g16659 and P2_R1164_U417 P2_R1164_U416 ; P2_R1164_U153
g16660 nand P2_R1164_U365 P2_R1164_U299 P2_R1164_U86 ; P2_R1164_U154
g16661 nand P2_R1164_U293 P2_R1164_U292 ; P2_R1164_U155
g16662 and P2_R1164_U436 P2_R1164_U435 ; P2_R1164_U156
g16663 nand P2_R1164_U289 P2_R1164_U288 ; P2_R1164_U157
g16664 and P2_R1164_U443 P2_R1164_U442 ; P2_R1164_U158
g16665 nand P2_R1164_U132 P2_R1164_U284 ; P2_R1164_U159
g16666 and P2_R1164_U450 P2_R1164_U449 ; P2_R1164_U160
g16667 nand P2_R1164_U43 P2_R1164_U327 ; P2_R1164_U161
g16668 nand P2_R1164_U130 P2_R1164_U269 ; P2_R1164_U162
g16669 and P2_R1164_U476 P2_R1164_U475 ; P2_R1164_U163
g16670 nand P2_R1164_U257 P2_R1164_U256 ; P2_R1164_U164
g16671 and P2_R1164_U483 P2_R1164_U482 ; P2_R1164_U165
g16672 nand P2_R1164_U253 P2_R1164_U252 ; P2_R1164_U166
g16673 nand P2_R1164_U127 P2_R1164_U242 ; P2_R1164_U167
g16674 nand P2_R1164_U367 P2_R1164_U366 ; P2_R1164_U168
g16675 nand P2_U3054 P2_R1164_U152 ; P2_R1164_U169
g16676 not P2_R1164_U34 ; P2_R1164_U170
g16677 nand P2_U3477 P2_U3083 ; P2_R1164_U171
g16678 nand P2_U3072 P2_U3486 ; P2_R1164_U172
g16679 nand P2_U3058 P2_U3971 ; P2_R1164_U173
g16680 not P2_R1164_U68 ; P2_R1164_U174
g16681 not P2_R1164_U77 ; P2_R1164_U175
g16682 nand P2_U3065 P2_U3972 ; P2_R1164_U176
g16683 not P2_R1164_U63 ; P2_R1164_U177
g16684 or P2_U3067 P2_U3465 ; P2_R1164_U178
g16685 or P2_U3060 P2_U3462 ; P2_R1164_U179
g16686 or P2_U3459 P2_U3064 ; P2_R1164_U180
g16687 or P2_U3456 P2_U3068 ; P2_R1164_U181
g16688 not P2_R1164_U31 ; P2_R1164_U182
g16689 or P2_U3453 P2_U3078 ; P2_R1164_U183
g16690 not P2_R1164_U42 ; P2_R1164_U184
g16691 not P2_R1164_U43 ; P2_R1164_U185
g16692 nand P2_R1164_U42 P2_R1164_U43 ; P2_R1164_U186
g16693 nand P2_U3068 P2_U3456 ; P2_R1164_U187
g16694 nand P2_R1164_U186 P2_R1164_U181 ; P2_R1164_U188
g16695 nand P2_U3064 P2_U3459 ; P2_R1164_U189
g16696 nand P2_R1164_U115 P2_R1164_U188 ; P2_R1164_U190
g16697 nand P2_R1164_U35 P2_R1164_U34 ; P2_R1164_U191
g16698 nand P2_U3067 P2_R1164_U191 ; P2_R1164_U192
g16699 nand P2_R1164_U116 P2_R1164_U190 ; P2_R1164_U193
g16700 nand P2_U3465 P2_R1164_U170 ; P2_R1164_U194
g16701 not P2_R1164_U41 ; P2_R1164_U195
g16702 or P2_U3070 P2_U3471 ; P2_R1164_U196
g16703 or P2_U3071 P2_U3468 ; P2_R1164_U197
g16704 not P2_R1164_U22 ; P2_R1164_U198
g16705 nand P2_R1164_U23 P2_R1164_U22 ; P2_R1164_U199
g16706 nand P2_U3070 P2_R1164_U199 ; P2_R1164_U200
g16707 nand P2_U3471 P2_R1164_U198 ; P2_R1164_U201
g16708 nand P2_R1164_U5 P2_R1164_U41 ; P2_R1164_U202
g16709 not P2_R1164_U145 ; P2_R1164_U203
g16710 or P2_U3474 P2_U3084 ; P2_R1164_U204
g16711 nand P2_R1164_U204 P2_R1164_U145 ; P2_R1164_U205
g16712 not P2_R1164_U40 ; P2_R1164_U206
g16713 or P2_U3083 P2_U3477 ; P2_R1164_U207
g16714 or P2_U3468 P2_U3071 ; P2_R1164_U208
g16715 nand P2_R1164_U208 P2_R1164_U41 ; P2_R1164_U209
g16716 nand P2_R1164_U119 P2_R1164_U209 ; P2_R1164_U210
g16717 nand P2_R1164_U195 P2_R1164_U22 ; P2_R1164_U211
g16718 nand P2_U3471 P2_U3070 ; P2_R1164_U212
g16719 nand P2_R1164_U120 P2_R1164_U211 ; P2_R1164_U213
g16720 or P2_U3071 P2_U3468 ; P2_R1164_U214
g16721 nand P2_R1164_U185 P2_R1164_U181 ; P2_R1164_U215
g16722 nand P2_U3068 P2_U3456 ; P2_R1164_U216
g16723 not P2_R1164_U45 ; P2_R1164_U217
g16724 nand P2_R1164_U121 P2_R1164_U184 ; P2_R1164_U218
g16725 nand P2_R1164_U45 P2_R1164_U180 ; P2_R1164_U219
g16726 nand P2_U3064 P2_U3459 ; P2_R1164_U220
g16727 not P2_R1164_U44 ; P2_R1164_U221
g16728 or P2_U3462 P2_U3060 ; P2_R1164_U222
g16729 nand P2_R1164_U222 P2_R1164_U44 ; P2_R1164_U223
g16730 nand P2_R1164_U123 P2_R1164_U223 ; P2_R1164_U224
g16731 nand P2_R1164_U221 P2_R1164_U34 ; P2_R1164_U225
g16732 nand P2_U3465 P2_U3067 ; P2_R1164_U226
g16733 nand P2_R1164_U124 P2_R1164_U225 ; P2_R1164_U227
g16734 or P2_U3060 P2_U3462 ; P2_R1164_U228
g16735 nand P2_R1164_U184 P2_R1164_U181 ; P2_R1164_U229
g16736 not P2_R1164_U146 ; P2_R1164_U230
g16737 nand P2_U3064 P2_U3459 ; P2_R1164_U231
g16738 nand P2_R1164_U401 P2_R1164_U400 P2_R1164_U43 P2_R1164_U42 ; P2_R1164_U232
g16739 nand P2_R1164_U43 P2_R1164_U42 ; P2_R1164_U233
g16740 nand P2_U3068 P2_U3456 ; P2_R1164_U234
g16741 nand P2_R1164_U125 P2_R1164_U233 ; P2_R1164_U235
g16742 or P2_U3083 P2_U3477 ; P2_R1164_U236
g16743 or P2_U3062 P2_U3480 ; P2_R1164_U237
g16744 nand P2_R1164_U177 P2_R1164_U6 ; P2_R1164_U238
g16745 nand P2_U3062 P2_U3480 ; P2_R1164_U239
g16746 nand P2_R1164_U171 P2_R1164_U238 ; P2_R1164_U240
g16747 or P2_U3480 P2_U3062 ; P2_R1164_U241
g16748 nand P2_R1164_U126 P2_R1164_U145 ; P2_R1164_U242
g16749 nand P2_R1164_U241 P2_R1164_U240 ; P2_R1164_U243
g16750 not P2_R1164_U167 ; P2_R1164_U244
g16751 or P2_U3080 P2_U3489 ; P2_R1164_U245
g16752 or P2_U3072 P2_U3486 ; P2_R1164_U246
g16753 nand P2_R1164_U174 P2_R1164_U7 ; P2_R1164_U247
g16754 nand P2_U3080 P2_U3489 ; P2_R1164_U248
g16755 nand P2_R1164_U129 P2_R1164_U247 ; P2_R1164_U249
g16756 or P2_U3483 P2_U3063 ; P2_R1164_U250
g16757 or P2_U3489 P2_U3080 ; P2_R1164_U251
g16758 nand P2_R1164_U128 P2_R1164_U167 ; P2_R1164_U252
g16759 nand P2_R1164_U251 P2_R1164_U249 ; P2_R1164_U253
g16760 not P2_R1164_U166 ; P2_R1164_U254
g16761 or P2_U3492 P2_U3079 ; P2_R1164_U255
g16762 nand P2_R1164_U255 P2_R1164_U166 ; P2_R1164_U256
g16763 nand P2_U3079 P2_U3492 ; P2_R1164_U257
g16764 not P2_R1164_U164 ; P2_R1164_U258
g16765 or P2_U3495 P2_U3074 ; P2_R1164_U259
g16766 nand P2_R1164_U259 P2_R1164_U164 ; P2_R1164_U260
g16767 nand P2_U3074 P2_U3495 ; P2_R1164_U261
g16768 not P2_R1164_U92 ; P2_R1164_U262
g16769 or P2_U3069 P2_U3501 ; P2_R1164_U263
g16770 or P2_U3073 P2_U3498 ; P2_R1164_U264
g16771 not P2_R1164_U59 ; P2_R1164_U265
g16772 nand P2_R1164_U60 P2_R1164_U59 ; P2_R1164_U266
g16773 nand P2_U3069 P2_R1164_U266 ; P2_R1164_U267
g16774 nand P2_U3501 P2_R1164_U265 ; P2_R1164_U268
g16775 nand P2_R1164_U8 P2_R1164_U92 ; P2_R1164_U269
g16776 not P2_R1164_U162 ; P2_R1164_U270
g16777 or P2_U3076 P2_U3976 ; P2_R1164_U271
g16778 or P2_U3081 P2_U3506 ; P2_R1164_U272
g16779 or P2_U3075 P2_U3975 ; P2_R1164_U273
g16780 not P2_R1164_U80 ; P2_R1164_U274
g16781 nand P2_U3976 P2_R1164_U274 ; P2_R1164_U275
g16782 nand P2_R1164_U275 P2_R1164_U90 ; P2_R1164_U276
g16783 nand P2_R1164_U80 P2_R1164_U81 ; P2_R1164_U277
g16784 nand P2_R1164_U277 P2_R1164_U276 ; P2_R1164_U278
g16785 nand P2_R1164_U175 P2_R1164_U9 ; P2_R1164_U279
g16786 nand P2_U3075 P2_U3975 ; P2_R1164_U280
g16787 nand P2_R1164_U278 P2_R1164_U279 ; P2_R1164_U281
g16788 or P2_U3504 P2_U3082 ; P2_R1164_U282
g16789 or P2_U3975 P2_U3075 ; P2_R1164_U283
g16790 nand P2_R1164_U162 P2_R1164_U131 ; P2_R1164_U284
g16791 nand P2_R1164_U283 P2_R1164_U281 ; P2_R1164_U285
g16792 not P2_R1164_U159 ; P2_R1164_U286
g16793 or P2_U3974 P2_U3061 ; P2_R1164_U287
g16794 nand P2_R1164_U287 P2_R1164_U159 ; P2_R1164_U288
g16795 nand P2_U3061 P2_U3974 ; P2_R1164_U289
g16796 not P2_R1164_U157 ; P2_R1164_U290
g16797 or P2_U3973 P2_U3066 ; P2_R1164_U291
g16798 nand P2_R1164_U291 P2_R1164_U157 ; P2_R1164_U292
g16799 nand P2_U3066 P2_U3973 ; P2_R1164_U293
g16800 not P2_R1164_U155 ; P2_R1164_U294
g16801 or P2_U3058 P2_U3971 ; P2_R1164_U295
g16802 nand P2_R1164_U176 P2_R1164_U173 ; P2_R1164_U296
g16803 not P2_R1164_U86 ; P2_R1164_U297
g16804 or P2_U3972 P2_U3065 ; P2_R1164_U298
g16805 nand P2_R1164_U155 P2_R1164_U298 P2_R1164_U168 ; P2_R1164_U299
g16806 not P2_R1164_U154 ; P2_R1164_U300
g16807 or P2_U3969 P2_U3053 ; P2_R1164_U301
g16808 nand P2_U3053 P2_U3969 ; P2_R1164_U302
g16809 not P2_R1164_U152 ; P2_R1164_U303
g16810 nand P2_U3968 P2_R1164_U152 ; P2_R1164_U304
g16811 not P2_R1164_U150 ; P2_R1164_U305
g16812 nand P2_R1164_U298 P2_R1164_U155 ; P2_R1164_U306
g16813 not P2_R1164_U89 ; P2_R1164_U307
g16814 or P2_U3971 P2_U3058 ; P2_R1164_U308
g16815 nand P2_R1164_U308 P2_R1164_U89 ; P2_R1164_U309
g16816 nand P2_R1164_U135 P2_R1164_U309 ; P2_R1164_U310
g16817 nand P2_R1164_U307 P2_R1164_U173 ; P2_R1164_U311
g16818 nand P2_U3970 P2_U3057 ; P2_R1164_U312
g16819 nand P2_R1164_U311 P2_R1164_U312 P2_R1164_U168 ; P2_R1164_U313
g16820 or P2_U3058 P2_U3971 ; P2_R1164_U314
g16821 nand P2_R1164_U282 P2_R1164_U162 ; P2_R1164_U315
g16822 not P2_R1164_U91 ; P2_R1164_U316
g16823 nand P2_R1164_U9 P2_R1164_U91 ; P2_R1164_U317
g16824 nand P2_R1164_U136 P2_R1164_U317 ; P2_R1164_U318
g16825 nand P2_R1164_U317 P2_R1164_U278 ; P2_R1164_U319
g16826 nand P2_R1164_U453 P2_R1164_U319 ; P2_R1164_U320
g16827 or P2_U3506 P2_U3081 ; P2_R1164_U321
g16828 nand P2_R1164_U321 P2_R1164_U91 ; P2_R1164_U322
g16829 nand P2_R1164_U137 P2_R1164_U322 ; P2_R1164_U323
g16830 nand P2_R1164_U316 P2_R1164_U80 ; P2_R1164_U324
g16831 nand P2_U3076 P2_U3976 ; P2_R1164_U325
g16832 nand P2_R1164_U138 P2_R1164_U324 ; P2_R1164_U326
g16833 or P2_U3453 P2_U3078 ; P2_R1164_U327
g16834 not P2_R1164_U161 ; P2_R1164_U328
g16835 or P2_U3081 P2_U3506 ; P2_R1164_U329
g16836 or P2_U3498 P2_U3073 ; P2_R1164_U330
g16837 nand P2_R1164_U330 P2_R1164_U92 ; P2_R1164_U331
g16838 nand P2_R1164_U139 P2_R1164_U331 ; P2_R1164_U332
g16839 nand P2_R1164_U262 P2_R1164_U59 ; P2_R1164_U333
g16840 nand P2_U3501 P2_U3069 ; P2_R1164_U334
g16841 nand P2_R1164_U140 P2_R1164_U333 ; P2_R1164_U335
g16842 or P2_U3073 P2_U3498 ; P2_R1164_U336
g16843 nand P2_R1164_U250 P2_R1164_U167 ; P2_R1164_U337
g16844 not P2_R1164_U93 ; P2_R1164_U338
g16845 or P2_U3486 P2_U3072 ; P2_R1164_U339
g16846 nand P2_R1164_U339 P2_R1164_U93 ; P2_R1164_U340
g16847 nand P2_R1164_U141 P2_R1164_U340 ; P2_R1164_U341
g16848 nand P2_R1164_U338 P2_R1164_U172 ; P2_R1164_U342
g16849 nand P2_U3080 P2_U3489 ; P2_R1164_U343
g16850 nand P2_R1164_U142 P2_R1164_U342 ; P2_R1164_U344
g16851 or P2_U3072 P2_U3486 ; P2_R1164_U345
g16852 or P2_U3477 P2_U3083 ; P2_R1164_U346
g16853 nand P2_R1164_U346 P2_R1164_U40 ; P2_R1164_U347
g16854 nand P2_R1164_U143 P2_R1164_U347 ; P2_R1164_U348
g16855 nand P2_R1164_U206 P2_R1164_U171 ; P2_R1164_U349
g16856 nand P2_U3062 P2_U3480 ; P2_R1164_U350
g16857 nand P2_R1164_U144 P2_R1164_U349 ; P2_R1164_U351
g16858 nand P2_R1164_U207 P2_R1164_U171 ; P2_R1164_U352
g16859 nand P2_R1164_U204 P2_R1164_U63 ; P2_R1164_U353
g16860 nand P2_R1164_U214 P2_R1164_U22 ; P2_R1164_U354
g16861 nand P2_R1164_U228 P2_R1164_U34 ; P2_R1164_U355
g16862 nand P2_R1164_U231 P2_R1164_U180 ; P2_R1164_U356
g16863 nand P2_R1164_U314 P2_R1164_U173 ; P2_R1164_U357
g16864 nand P2_R1164_U298 P2_R1164_U176 ; P2_R1164_U358
g16865 nand P2_R1164_U329 P2_R1164_U80 ; P2_R1164_U359
g16866 nand P2_R1164_U282 P2_R1164_U77 ; P2_R1164_U360
g16867 nand P2_R1164_U336 P2_R1164_U59 ; P2_R1164_U361
g16868 nand P2_R1164_U345 P2_R1164_U172 ; P2_R1164_U362
g16869 nand P2_R1164_U250 P2_R1164_U68 ; P2_R1164_U363
g16870 nand P2_U3968 P2_U3054 ; P2_R1164_U364
g16871 nand P2_R1164_U296 P2_R1164_U168 ; P2_R1164_U365
g16872 nand P2_U3057 P2_R1164_U295 ; P2_R1164_U366
g16873 nand P2_U3970 P2_R1164_U295 ; P2_R1164_U367
g16874 nand P2_R1164_U296 P2_R1164_U168 P2_R1164_U301 ; P2_R1164_U368
g16875 nand P2_R1164_U155 P2_R1164_U168 P2_R1164_U133 ; P2_R1164_U369
g16876 nand P2_R1164_U297 P2_R1164_U301 ; P2_R1164_U370
g16877 nand P2_U3083 P2_R1164_U39 ; P2_R1164_U371
g16878 nand P2_U3477 P2_R1164_U38 ; P2_R1164_U372
g16879 nand P2_R1164_U372 P2_R1164_U371 ; P2_R1164_U373
g16880 nand P2_R1164_U352 P2_R1164_U40 ; P2_R1164_U374
g16881 nand P2_R1164_U373 P2_R1164_U206 ; P2_R1164_U375
g16882 nand P2_U3084 P2_R1164_U36 ; P2_R1164_U376
g16883 nand P2_U3474 P2_R1164_U37 ; P2_R1164_U377
g16884 nand P2_R1164_U377 P2_R1164_U376 ; P2_R1164_U378
g16885 nand P2_R1164_U353 P2_R1164_U145 ; P2_R1164_U379
g16886 nand P2_R1164_U203 P2_R1164_U378 ; P2_R1164_U380
g16887 nand P2_U3070 P2_R1164_U23 ; P2_R1164_U381
g16888 nand P2_U3471 P2_R1164_U21 ; P2_R1164_U382
g16889 nand P2_U3071 P2_R1164_U19 ; P2_R1164_U383
g16890 nand P2_U3468 P2_R1164_U20 ; P2_R1164_U384
g16891 nand P2_R1164_U384 P2_R1164_U383 ; P2_R1164_U385
g16892 nand P2_R1164_U354 P2_R1164_U41 ; P2_R1164_U386
g16893 nand P2_R1164_U385 P2_R1164_U195 ; P2_R1164_U387
g16894 nand P2_U3067 P2_R1164_U35 ; P2_R1164_U388
g16895 nand P2_U3465 P2_R1164_U26 ; P2_R1164_U389
g16896 nand P2_U3060 P2_R1164_U24 ; P2_R1164_U390
g16897 nand P2_U3462 P2_R1164_U25 ; P2_R1164_U391
g16898 nand P2_R1164_U391 P2_R1164_U390 ; P2_R1164_U392
g16899 nand P2_R1164_U355 P2_R1164_U44 ; P2_R1164_U393
g16900 nand P2_R1164_U392 P2_R1164_U221 ; P2_R1164_U394
g16901 nand P2_U3064 P2_R1164_U32 ; P2_R1164_U395
g16902 nand P2_U3459 P2_R1164_U33 ; P2_R1164_U396
g16903 nand P2_R1164_U396 P2_R1164_U395 ; P2_R1164_U397
g16904 nand P2_R1164_U356 P2_R1164_U146 ; P2_R1164_U398
g16905 nand P2_R1164_U230 P2_R1164_U397 ; P2_R1164_U399
g16906 nand P2_U3068 P2_R1164_U27 ; P2_R1164_U400
g16907 nand P2_U3456 P2_R1164_U28 ; P2_R1164_U401
g16908 nand P2_U3055 P2_R1164_U148 ; P2_R1164_U402
g16909 nand P2_U3979 P2_R1164_U147 ; P2_R1164_U403
g16910 nand P2_U3055 P2_R1164_U148 ; P2_R1164_U404
g16911 nand P2_U3979 P2_R1164_U147 ; P2_R1164_U405
g16912 nand P2_R1164_U405 P2_R1164_U404 ; P2_R1164_U406
g16913 nand P2_R1164_U149 P2_R1164_U150 ; P2_R1164_U407
g16914 nand P2_R1164_U305 P2_R1164_U406 ; P2_R1164_U408
g16915 nand P2_U3054 P2_R1164_U88 ; P2_R1164_U409
g16916 nand P2_U3968 P2_R1164_U87 ; P2_R1164_U410
g16917 nand P2_U3054 P2_R1164_U88 ; P2_R1164_U411
g16918 nand P2_U3968 P2_R1164_U87 ; P2_R1164_U412
g16919 nand P2_R1164_U412 P2_R1164_U411 ; P2_R1164_U413
g16920 nand P2_R1164_U151 P2_R1164_U152 ; P2_R1164_U414
g16921 nand P2_R1164_U303 P2_R1164_U413 ; P2_R1164_U415
g16922 nand P2_U3053 P2_R1164_U46 ; P2_R1164_U416
g16923 nand P2_U3969 P2_R1164_U47 ; P2_R1164_U417
g16924 nand P2_U3053 P2_R1164_U46 ; P2_R1164_U418
g16925 nand P2_U3969 P2_R1164_U47 ; P2_R1164_U419
g16926 nand P2_R1164_U419 P2_R1164_U418 ; P2_R1164_U420
g16927 nand P2_R1164_U153 P2_R1164_U154 ; P2_R1164_U421
g16928 nand P2_R1164_U300 P2_R1164_U420 ; P2_R1164_U422
g16929 nand P2_U3057 P2_R1164_U49 ; P2_R1164_U423
g16930 nand P2_U3970 P2_R1164_U48 ; P2_R1164_U424
g16931 nand P2_U3058 P2_R1164_U50 ; P2_R1164_U425
g16932 nand P2_U3971 P2_R1164_U51 ; P2_R1164_U426
g16933 nand P2_R1164_U426 P2_R1164_U425 ; P2_R1164_U427
g16934 nand P2_R1164_U357 P2_R1164_U89 ; P2_R1164_U428
g16935 nand P2_R1164_U427 P2_R1164_U307 ; P2_R1164_U429
g16936 nand P2_U3065 P2_R1164_U52 ; P2_R1164_U430
g16937 nand P2_U3972 P2_R1164_U53 ; P2_R1164_U431
g16938 nand P2_R1164_U431 P2_R1164_U430 ; P2_R1164_U432
g16939 nand P2_R1164_U358 P2_R1164_U155 ; P2_R1164_U433
g16940 nand P2_R1164_U294 P2_R1164_U432 ; P2_R1164_U434
g16941 nand P2_U3066 P2_R1164_U84 ; P2_R1164_U435
g16942 nand P2_U3973 P2_R1164_U85 ; P2_R1164_U436
g16943 nand P2_U3066 P2_R1164_U84 ; P2_R1164_U437
g16944 nand P2_U3973 P2_R1164_U85 ; P2_R1164_U438
g16945 nand P2_R1164_U438 P2_R1164_U437 ; P2_R1164_U439
g16946 nand P2_R1164_U156 P2_R1164_U157 ; P2_R1164_U440
g16947 nand P2_R1164_U290 P2_R1164_U439 ; P2_R1164_U441
g16948 nand P2_U3061 P2_R1164_U82 ; P2_R1164_U442
g16949 nand P2_U3974 P2_R1164_U83 ; P2_R1164_U443
g16950 nand P2_U3061 P2_R1164_U82 ; P2_R1164_U444
g16951 nand P2_U3974 P2_R1164_U83 ; P2_R1164_U445
g16952 nand P2_R1164_U445 P2_R1164_U444 ; P2_R1164_U446
g16953 nand P2_R1164_U158 P2_R1164_U159 ; P2_R1164_U447
g16954 nand P2_R1164_U286 P2_R1164_U446 ; P2_R1164_U448
g16955 nand P2_U3075 P2_R1164_U54 ; P2_R1164_U449
g16956 nand P2_U3975 P2_R1164_U55 ; P2_R1164_U450
g16957 nand P2_U3075 P2_R1164_U54 ; P2_R1164_U451
g16958 nand P2_U3975 P2_R1164_U55 ; P2_R1164_U452
g16959 nand P2_R1164_U452 P2_R1164_U451 ; P2_R1164_U453
g16960 nand P2_U3076 P2_R1164_U81 ; P2_R1164_U454
g16961 nand P2_U3976 P2_R1164_U90 ; P2_R1164_U455
g16962 nand P2_R1164_U182 P2_R1164_U161 ; P2_R1164_U456
g16963 nand P2_R1164_U328 P2_R1164_U31 ; P2_R1164_U457
g16964 nand P2_U3081 P2_R1164_U78 ; P2_R1164_U458
g16965 nand P2_U3506 P2_R1164_U79 ; P2_R1164_U459
g16966 nand P2_R1164_U459 P2_R1164_U458 ; P2_R1164_U460
g16967 nand P2_R1164_U359 P2_R1164_U91 ; P2_R1164_U461
g16968 nand P2_R1164_U460 P2_R1164_U316 ; P2_R1164_U462
g16969 nand P2_U3082 P2_R1164_U75 ; P2_R1164_U463
g16970 nand P2_U3504 P2_R1164_U76 ; P2_R1164_U464
g16971 nand P2_R1164_U464 P2_R1164_U463 ; P2_R1164_U465
g16972 nand P2_R1164_U360 P2_R1164_U162 ; P2_R1164_U466
g16973 nand P2_R1164_U270 P2_R1164_U465 ; P2_R1164_U467
g16974 nand P2_U3069 P2_R1164_U60 ; P2_R1164_U468
g16975 nand P2_U3501 P2_R1164_U58 ; P2_R1164_U469
g16976 nand P2_U3073 P2_R1164_U56 ; P2_R1164_U470
g16977 nand P2_U3498 P2_R1164_U57 ; P2_R1164_U471
g16978 nand P2_R1164_U471 P2_R1164_U470 ; P2_R1164_U472
g16979 nand P2_R1164_U361 P2_R1164_U92 ; P2_R1164_U473
g16980 nand P2_R1164_U472 P2_R1164_U262 ; P2_R1164_U474
g16981 nand P2_U3074 P2_R1164_U73 ; P2_R1164_U475
g16982 nand P2_U3495 P2_R1164_U74 ; P2_R1164_U476
g16983 nand P2_U3074 P2_R1164_U73 ; P2_R1164_U477
g16984 nand P2_U3495 P2_R1164_U74 ; P2_R1164_U478
g16985 nand P2_R1164_U478 P2_R1164_U477 ; P2_R1164_U479
g16986 nand P2_R1164_U163 P2_R1164_U164 ; P2_R1164_U480
g16987 nand P2_R1164_U258 P2_R1164_U479 ; P2_R1164_U481
g16988 nand P2_U3079 P2_R1164_U71 ; P2_R1164_U482
g16989 nand P2_U3492 P2_R1164_U72 ; P2_R1164_U483
g16990 nand P2_U3079 P2_R1164_U71 ; P2_R1164_U484
g16991 nand P2_U3492 P2_R1164_U72 ; P2_R1164_U485
g16992 nand P2_R1164_U485 P2_R1164_U484 ; P2_R1164_U486
g16993 nand P2_R1164_U165 P2_R1164_U166 ; P2_R1164_U487
g16994 nand P2_R1164_U254 P2_R1164_U486 ; P2_R1164_U488
g16995 nand P2_U3080 P2_R1164_U69 ; P2_R1164_U489
g16996 nand P2_U3489 P2_R1164_U70 ; P2_R1164_U490
g16997 nand P2_U3072 P2_R1164_U64 ; P2_R1164_U491
g16998 nand P2_U3486 P2_R1164_U65 ; P2_R1164_U492
g16999 nand P2_R1164_U492 P2_R1164_U491 ; P2_R1164_U493
g17000 nand P2_R1164_U362 P2_R1164_U93 ; P2_R1164_U494
g17001 nand P2_R1164_U493 P2_R1164_U338 ; P2_R1164_U495
g17002 nand P2_U3063 P2_R1164_U66 ; P2_R1164_U496
g17003 nand P2_U3483 P2_R1164_U67 ; P2_R1164_U497
g17004 nand P2_R1164_U497 P2_R1164_U496 ; P2_R1164_U498
g17005 nand P2_R1164_U363 P2_R1164_U167 ; P2_R1164_U499
g17006 nand P2_R1164_U244 P2_R1164_U498 ; P2_R1164_U500
g17007 nand P2_U3062 P2_R1164_U61 ; P2_R1164_U501
g17008 nand P2_U3480 P2_R1164_U62 ; P2_R1164_U502
g17009 nand P2_U3077 P2_R1164_U29 ; P2_R1164_U503
g17010 nand P2_U3448 P2_R1164_U30 ; P2_R1164_U504
g17011 and P2_R1233_U179 P2_R1233_U178 ; P2_R1233_U4
g17012 and P2_R1233_U197 P2_R1233_U196 ; P2_R1233_U5
g17013 and P2_R1233_U237 P2_R1233_U236 ; P2_R1233_U6
g17014 and P2_R1233_U246 P2_R1233_U245 ; P2_R1233_U7
g17015 and P2_R1233_U264 P2_R1233_U263 ; P2_R1233_U8
g17016 and P2_R1233_U272 P2_R1233_U271 ; P2_R1233_U9
g17017 and P2_R1233_U351 P2_R1233_U348 ; P2_R1233_U10
g17018 and P2_R1233_U344 P2_R1233_U341 ; P2_R1233_U11
g17019 and P2_R1233_U335 P2_R1233_U332 ; P2_R1233_U12
g17020 and P2_R1233_U326 P2_R1233_U323 ; P2_R1233_U13
g17021 and P2_R1233_U320 P2_R1233_U318 ; P2_R1233_U14
g17022 and P2_R1233_U313 P2_R1233_U310 ; P2_R1233_U15
g17023 and P2_R1233_U235 P2_R1233_U232 ; P2_R1233_U16
g17024 and P2_R1233_U227 P2_R1233_U224 ; P2_R1233_U17
g17025 and P2_R1233_U213 P2_R1233_U210 ; P2_R1233_U18
g17026 not P2_U3468 ; P2_R1233_U19
g17027 not P2_U3071 ; P2_R1233_U20
g17028 not P2_U3070 ; P2_R1233_U21
g17029 nand P2_U3071 P2_U3468 ; P2_R1233_U22
g17030 not P2_U3471 ; P2_R1233_U23
g17031 not P2_U3462 ; P2_R1233_U24
g17032 not P2_U3060 ; P2_R1233_U25
g17033 not P2_U3067 ; P2_R1233_U26
g17034 not P2_U3456 ; P2_R1233_U27
g17035 not P2_U3068 ; P2_R1233_U28
g17036 not P2_U3448 ; P2_R1233_U29
g17037 not P2_U3077 ; P2_R1233_U30
g17038 nand P2_U3077 P2_U3448 ; P2_R1233_U31
g17039 not P2_U3459 ; P2_R1233_U32
g17040 not P2_U3064 ; P2_R1233_U33
g17041 nand P2_U3060 P2_U3462 ; P2_R1233_U34
g17042 not P2_U3465 ; P2_R1233_U35
g17043 not P2_U3474 ; P2_R1233_U36
g17044 not P2_U3084 ; P2_R1233_U37
g17045 not P2_U3083 ; P2_R1233_U38
g17046 not P2_U3477 ; P2_R1233_U39
g17047 nand P2_R1233_U63 P2_R1233_U205 ; P2_R1233_U40
g17048 nand P2_R1233_U117 P2_R1233_U193 ; P2_R1233_U41
g17049 nand P2_R1233_U182 P2_R1233_U183 ; P2_R1233_U42
g17050 nand P2_U3453 P2_U3078 ; P2_R1233_U43
g17051 nand P2_R1233_U122 P2_R1233_U219 ; P2_R1233_U44
g17052 nand P2_R1233_U216 P2_R1233_U215 ; P2_R1233_U45
g17053 not P2_U3969 ; P2_R1233_U46
g17054 not P2_U3053 ; P2_R1233_U47
g17055 not P2_U3057 ; P2_R1233_U48
g17056 not P2_U3970 ; P2_R1233_U49
g17057 not P2_U3971 ; P2_R1233_U50
g17058 not P2_U3058 ; P2_R1233_U51
g17059 not P2_U3972 ; P2_R1233_U52
g17060 not P2_U3065 ; P2_R1233_U53
g17061 not P2_U3975 ; P2_R1233_U54
g17062 not P2_U3075 ; P2_R1233_U55
g17063 not P2_U3498 ; P2_R1233_U56
g17064 not P2_U3073 ; P2_R1233_U57
g17065 not P2_U3069 ; P2_R1233_U58
g17066 nand P2_U3073 P2_U3498 ; P2_R1233_U59
g17067 not P2_U3501 ; P2_R1233_U60
g17068 not P2_U3480 ; P2_R1233_U61
g17069 not P2_U3062 ; P2_R1233_U62
g17070 nand P2_U3084 P2_U3474 ; P2_R1233_U63
g17071 not P2_U3486 ; P2_R1233_U64
g17072 not P2_U3072 ; P2_R1233_U65
g17073 not P2_U3483 ; P2_R1233_U66
g17074 not P2_U3063 ; P2_R1233_U67
g17075 nand P2_U3063 P2_U3483 ; P2_R1233_U68
g17076 not P2_U3489 ; P2_R1233_U69
g17077 not P2_U3080 ; P2_R1233_U70
g17078 not P2_U3492 ; P2_R1233_U71
g17079 not P2_U3079 ; P2_R1233_U72
g17080 not P2_U3495 ; P2_R1233_U73
g17081 not P2_U3074 ; P2_R1233_U74
g17082 not P2_U3504 ; P2_R1233_U75
g17083 not P2_U3082 ; P2_R1233_U76
g17084 nand P2_U3082 P2_U3504 ; P2_R1233_U77
g17085 not P2_U3506 ; P2_R1233_U78
g17086 not P2_U3081 ; P2_R1233_U79
g17087 nand P2_U3081 P2_U3506 ; P2_R1233_U80
g17088 not P2_U3976 ; P2_R1233_U81
g17089 not P2_U3974 ; P2_R1233_U82
g17090 not P2_U3061 ; P2_R1233_U83
g17091 not P2_U3973 ; P2_R1233_U84
g17092 not P2_U3066 ; P2_R1233_U85
g17093 nand P2_U3970 P2_U3057 ; P2_R1233_U86
g17094 not P2_U3054 ; P2_R1233_U87
g17095 not P2_U3968 ; P2_R1233_U88
g17096 nand P2_R1233_U306 P2_R1233_U176 ; P2_R1233_U89
g17097 not P2_U3076 ; P2_R1233_U90
g17098 nand P2_R1233_U77 P2_R1233_U315 ; P2_R1233_U91
g17099 nand P2_R1233_U261 P2_R1233_U260 ; P2_R1233_U92
g17100 nand P2_R1233_U68 P2_R1233_U337 ; P2_R1233_U93
g17101 nand P2_R1233_U457 P2_R1233_U456 ; P2_R1233_U94
g17102 nand P2_R1233_U504 P2_R1233_U503 ; P2_R1233_U95
g17103 nand P2_R1233_U375 P2_R1233_U374 ; P2_R1233_U96
g17104 nand P2_R1233_U380 P2_R1233_U379 ; P2_R1233_U97
g17105 nand P2_R1233_U387 P2_R1233_U386 ; P2_R1233_U98
g17106 nand P2_R1233_U394 P2_R1233_U393 ; P2_R1233_U99
g17107 nand P2_R1233_U399 P2_R1233_U398 ; P2_R1233_U100
g17108 nand P2_R1233_U408 P2_R1233_U407 ; P2_R1233_U101
g17109 nand P2_R1233_U415 P2_R1233_U414 ; P2_R1233_U102
g17110 nand P2_R1233_U422 P2_R1233_U421 ; P2_R1233_U103
g17111 nand P2_R1233_U429 P2_R1233_U428 ; P2_R1233_U104
g17112 nand P2_R1233_U434 P2_R1233_U433 ; P2_R1233_U105
g17113 nand P2_R1233_U441 P2_R1233_U440 ; P2_R1233_U106
g17114 nand P2_R1233_U448 P2_R1233_U447 ; P2_R1233_U107
g17115 nand P2_R1233_U462 P2_R1233_U461 ; P2_R1233_U108
g17116 nand P2_R1233_U467 P2_R1233_U466 ; P2_R1233_U109
g17117 nand P2_R1233_U474 P2_R1233_U473 ; P2_R1233_U110
g17118 nand P2_R1233_U481 P2_R1233_U480 ; P2_R1233_U111
g17119 nand P2_R1233_U488 P2_R1233_U487 ; P2_R1233_U112
g17120 nand P2_R1233_U495 P2_R1233_U494 ; P2_R1233_U113
g17121 nand P2_R1233_U500 P2_R1233_U499 ; P2_R1233_U114
g17122 and P2_R1233_U189 P2_R1233_U187 ; P2_R1233_U115
g17123 and P2_R1233_U4 P2_R1233_U180 ; P2_R1233_U116
g17124 and P2_R1233_U194 P2_R1233_U192 ; P2_R1233_U117
g17125 and P2_R1233_U201 P2_R1233_U200 ; P2_R1233_U118
g17126 and P2_R1233_U382 P2_R1233_U381 P2_R1233_U22 ; P2_R1233_U119
g17127 and P2_R1233_U212 P2_R1233_U5 ; P2_R1233_U120
g17128 and P2_R1233_U181 P2_R1233_U180 ; P2_R1233_U121
g17129 and P2_R1233_U220 P2_R1233_U218 ; P2_R1233_U122
g17130 and P2_R1233_U389 P2_R1233_U388 P2_R1233_U34 ; P2_R1233_U123
g17131 and P2_R1233_U226 P2_R1233_U4 ; P2_R1233_U124
g17132 and P2_R1233_U234 P2_R1233_U181 ; P2_R1233_U125
g17133 and P2_R1233_U204 P2_R1233_U6 ; P2_R1233_U126
g17134 and P2_R1233_U243 P2_R1233_U239 ; P2_R1233_U127
g17135 and P2_R1233_U250 P2_R1233_U7 ; P2_R1233_U128
g17136 and P2_R1233_U248 P2_R1233_U172 ; P2_R1233_U129
g17137 and P2_R1233_U268 P2_R1233_U267 ; P2_R1233_U130
g17138 and P2_R1233_U9 P2_R1233_U282 P2_R1233_U273 ; P2_R1233_U131
g17139 and P2_R1233_U285 P2_R1233_U280 ; P2_R1233_U132
g17140 and P2_R1233_U301 P2_R1233_U298 ; P2_R1233_U133
g17141 and P2_R1233_U368 P2_R1233_U302 ; P2_R1233_U134
g17142 and P2_R1233_U424 P2_R1233_U423 P2_R1233_U173 ; P2_R1233_U135
g17143 and P2_R1233_U160 P2_R1233_U278 ; P2_R1233_U136
g17144 and P2_R1233_U455 P2_R1233_U454 P2_R1233_U80 ; P2_R1233_U137
g17145 and P2_R1233_U325 P2_R1233_U9 ; P2_R1233_U138
g17146 and P2_R1233_U469 P2_R1233_U468 P2_R1233_U59 ; P2_R1233_U139
g17147 and P2_R1233_U334 P2_R1233_U8 ; P2_R1233_U140
g17148 and P2_R1233_U490 P2_R1233_U489 P2_R1233_U172 ; P2_R1233_U141
g17149 and P2_R1233_U343 P2_R1233_U7 ; P2_R1233_U142
g17150 and P2_R1233_U502 P2_R1233_U501 P2_R1233_U171 ; P2_R1233_U143
g17151 and P2_R1233_U350 P2_R1233_U6 ; P2_R1233_U144
g17152 nand P2_R1233_U118 P2_R1233_U202 ; P2_R1233_U145
g17153 nand P2_R1233_U217 P2_R1233_U229 ; P2_R1233_U146
g17154 not P2_U3055 ; P2_R1233_U147
g17155 not P2_U3979 ; P2_R1233_U148
g17156 and P2_R1233_U403 P2_R1233_U402 ; P2_R1233_U149
g17157 nand P2_R1233_U304 P2_R1233_U169 P2_R1233_U364 ; P2_R1233_U150
g17158 and P2_R1233_U410 P2_R1233_U409 ; P2_R1233_U151
g17159 nand P2_R1233_U370 P2_R1233_U369 P2_R1233_U134 ; P2_R1233_U152
g17160 and P2_R1233_U417 P2_R1233_U416 ; P2_R1233_U153
g17161 nand P2_R1233_U365 P2_R1233_U299 P2_R1233_U86 ; P2_R1233_U154
g17162 nand P2_R1233_U293 P2_R1233_U292 ; P2_R1233_U155
g17163 and P2_R1233_U436 P2_R1233_U435 ; P2_R1233_U156
g17164 nand P2_R1233_U289 P2_R1233_U288 ; P2_R1233_U157
g17165 and P2_R1233_U443 P2_R1233_U442 ; P2_R1233_U158
g17166 nand P2_R1233_U132 P2_R1233_U284 ; P2_R1233_U159
g17167 and P2_R1233_U450 P2_R1233_U449 ; P2_R1233_U160
g17168 nand P2_R1233_U43 P2_R1233_U327 ; P2_R1233_U161
g17169 nand P2_R1233_U130 P2_R1233_U269 ; P2_R1233_U162
g17170 and P2_R1233_U476 P2_R1233_U475 ; P2_R1233_U163
g17171 nand P2_R1233_U257 P2_R1233_U256 ; P2_R1233_U164
g17172 and P2_R1233_U483 P2_R1233_U482 ; P2_R1233_U165
g17173 nand P2_R1233_U253 P2_R1233_U252 ; P2_R1233_U166
g17174 nand P2_R1233_U127 P2_R1233_U242 ; P2_R1233_U167
g17175 nand P2_R1233_U367 P2_R1233_U366 ; P2_R1233_U168
g17176 nand P2_U3054 P2_R1233_U152 ; P2_R1233_U169
g17177 not P2_R1233_U34 ; P2_R1233_U170
g17178 nand P2_U3477 P2_U3083 ; P2_R1233_U171
g17179 nand P2_U3072 P2_U3486 ; P2_R1233_U172
g17180 nand P2_U3058 P2_U3971 ; P2_R1233_U173
g17181 not P2_R1233_U68 ; P2_R1233_U174
g17182 not P2_R1233_U77 ; P2_R1233_U175
g17183 nand P2_U3065 P2_U3972 ; P2_R1233_U176
g17184 not P2_R1233_U63 ; P2_R1233_U177
g17185 or P2_U3067 P2_U3465 ; P2_R1233_U178
g17186 or P2_U3060 P2_U3462 ; P2_R1233_U179
g17187 or P2_U3459 P2_U3064 ; P2_R1233_U180
g17188 or P2_U3456 P2_U3068 ; P2_R1233_U181
g17189 not P2_R1233_U31 ; P2_R1233_U182
g17190 or P2_U3453 P2_U3078 ; P2_R1233_U183
g17191 not P2_R1233_U42 ; P2_R1233_U184
g17192 not P2_R1233_U43 ; P2_R1233_U185
g17193 nand P2_R1233_U42 P2_R1233_U43 ; P2_R1233_U186
g17194 nand P2_U3068 P2_U3456 ; P2_R1233_U187
g17195 nand P2_R1233_U186 P2_R1233_U181 ; P2_R1233_U188
g17196 nand P2_U3064 P2_U3459 ; P2_R1233_U189
g17197 nand P2_R1233_U115 P2_R1233_U188 ; P2_R1233_U190
g17198 nand P2_R1233_U35 P2_R1233_U34 ; P2_R1233_U191
g17199 nand P2_U3067 P2_R1233_U191 ; P2_R1233_U192
g17200 nand P2_R1233_U116 P2_R1233_U190 ; P2_R1233_U193
g17201 nand P2_U3465 P2_R1233_U170 ; P2_R1233_U194
g17202 not P2_R1233_U41 ; P2_R1233_U195
g17203 or P2_U3070 P2_U3471 ; P2_R1233_U196
g17204 or P2_U3071 P2_U3468 ; P2_R1233_U197
g17205 not P2_R1233_U22 ; P2_R1233_U198
g17206 nand P2_R1233_U23 P2_R1233_U22 ; P2_R1233_U199
g17207 nand P2_U3070 P2_R1233_U199 ; P2_R1233_U200
g17208 nand P2_U3471 P2_R1233_U198 ; P2_R1233_U201
g17209 nand P2_R1233_U5 P2_R1233_U41 ; P2_R1233_U202
g17210 not P2_R1233_U145 ; P2_R1233_U203
g17211 or P2_U3474 P2_U3084 ; P2_R1233_U204
g17212 nand P2_R1233_U204 P2_R1233_U145 ; P2_R1233_U205
g17213 not P2_R1233_U40 ; P2_R1233_U206
g17214 or P2_U3083 P2_U3477 ; P2_R1233_U207
g17215 or P2_U3468 P2_U3071 ; P2_R1233_U208
g17216 nand P2_R1233_U208 P2_R1233_U41 ; P2_R1233_U209
g17217 nand P2_R1233_U119 P2_R1233_U209 ; P2_R1233_U210
g17218 nand P2_R1233_U195 P2_R1233_U22 ; P2_R1233_U211
g17219 nand P2_U3471 P2_U3070 ; P2_R1233_U212
g17220 nand P2_R1233_U120 P2_R1233_U211 ; P2_R1233_U213
g17221 or P2_U3071 P2_U3468 ; P2_R1233_U214
g17222 nand P2_R1233_U185 P2_R1233_U181 ; P2_R1233_U215
g17223 nand P2_U3068 P2_U3456 ; P2_R1233_U216
g17224 not P2_R1233_U45 ; P2_R1233_U217
g17225 nand P2_R1233_U121 P2_R1233_U184 ; P2_R1233_U218
g17226 nand P2_R1233_U45 P2_R1233_U180 ; P2_R1233_U219
g17227 nand P2_U3064 P2_U3459 ; P2_R1233_U220
g17228 not P2_R1233_U44 ; P2_R1233_U221
g17229 or P2_U3462 P2_U3060 ; P2_R1233_U222
g17230 nand P2_R1233_U222 P2_R1233_U44 ; P2_R1233_U223
g17231 nand P2_R1233_U123 P2_R1233_U223 ; P2_R1233_U224
g17232 nand P2_R1233_U221 P2_R1233_U34 ; P2_R1233_U225
g17233 nand P2_U3465 P2_U3067 ; P2_R1233_U226
g17234 nand P2_R1233_U124 P2_R1233_U225 ; P2_R1233_U227
g17235 or P2_U3060 P2_U3462 ; P2_R1233_U228
g17236 nand P2_R1233_U184 P2_R1233_U181 ; P2_R1233_U229
g17237 not P2_R1233_U146 ; P2_R1233_U230
g17238 nand P2_U3064 P2_U3459 ; P2_R1233_U231
g17239 nand P2_R1233_U401 P2_R1233_U400 P2_R1233_U43 P2_R1233_U42 ; P2_R1233_U232
g17240 nand P2_R1233_U43 P2_R1233_U42 ; P2_R1233_U233
g17241 nand P2_U3068 P2_U3456 ; P2_R1233_U234
g17242 nand P2_R1233_U125 P2_R1233_U233 ; P2_R1233_U235
g17243 or P2_U3083 P2_U3477 ; P2_R1233_U236
g17244 or P2_U3062 P2_U3480 ; P2_R1233_U237
g17245 nand P2_R1233_U177 P2_R1233_U6 ; P2_R1233_U238
g17246 nand P2_U3062 P2_U3480 ; P2_R1233_U239
g17247 nand P2_R1233_U171 P2_R1233_U238 ; P2_R1233_U240
g17248 or P2_U3480 P2_U3062 ; P2_R1233_U241
g17249 nand P2_R1233_U126 P2_R1233_U145 ; P2_R1233_U242
g17250 nand P2_R1233_U241 P2_R1233_U240 ; P2_R1233_U243
g17251 not P2_R1233_U167 ; P2_R1233_U244
g17252 or P2_U3080 P2_U3489 ; P2_R1233_U245
g17253 or P2_U3072 P2_U3486 ; P2_R1233_U246
g17254 nand P2_R1233_U174 P2_R1233_U7 ; P2_R1233_U247
g17255 nand P2_U3080 P2_U3489 ; P2_R1233_U248
g17256 nand P2_R1233_U129 P2_R1233_U247 ; P2_R1233_U249
g17257 or P2_U3483 P2_U3063 ; P2_R1233_U250
g17258 or P2_U3489 P2_U3080 ; P2_R1233_U251
g17259 nand P2_R1233_U128 P2_R1233_U167 ; P2_R1233_U252
g17260 nand P2_R1233_U251 P2_R1233_U249 ; P2_R1233_U253
g17261 not P2_R1233_U166 ; P2_R1233_U254
g17262 or P2_U3492 P2_U3079 ; P2_R1233_U255
g17263 nand P2_R1233_U255 P2_R1233_U166 ; P2_R1233_U256
g17264 nand P2_U3079 P2_U3492 ; P2_R1233_U257
g17265 not P2_R1233_U164 ; P2_R1233_U258
g17266 or P2_U3495 P2_U3074 ; P2_R1233_U259
g17267 nand P2_R1233_U259 P2_R1233_U164 ; P2_R1233_U260
g17268 nand P2_U3074 P2_U3495 ; P2_R1233_U261
g17269 not P2_R1233_U92 ; P2_R1233_U262
g17270 or P2_U3069 P2_U3501 ; P2_R1233_U263
g17271 or P2_U3073 P2_U3498 ; P2_R1233_U264
g17272 not P2_R1233_U59 ; P2_R1233_U265
g17273 nand P2_R1233_U60 P2_R1233_U59 ; P2_R1233_U266
g17274 nand P2_U3069 P2_R1233_U266 ; P2_R1233_U267
g17275 nand P2_U3501 P2_R1233_U265 ; P2_R1233_U268
g17276 nand P2_R1233_U8 P2_R1233_U92 ; P2_R1233_U269
g17277 not P2_R1233_U162 ; P2_R1233_U270
g17278 or P2_U3076 P2_U3976 ; P2_R1233_U271
g17279 or P2_U3081 P2_U3506 ; P2_R1233_U272
g17280 or P2_U3075 P2_U3975 ; P2_R1233_U273
g17281 not P2_R1233_U80 ; P2_R1233_U274
g17282 nand P2_U3976 P2_R1233_U274 ; P2_R1233_U275
g17283 nand P2_R1233_U275 P2_R1233_U90 ; P2_R1233_U276
g17284 nand P2_R1233_U80 P2_R1233_U81 ; P2_R1233_U277
g17285 nand P2_R1233_U277 P2_R1233_U276 ; P2_R1233_U278
g17286 nand P2_R1233_U175 P2_R1233_U9 ; P2_R1233_U279
g17287 nand P2_U3075 P2_U3975 ; P2_R1233_U280
g17288 nand P2_R1233_U278 P2_R1233_U279 ; P2_R1233_U281
g17289 or P2_U3504 P2_U3082 ; P2_R1233_U282
g17290 or P2_U3975 P2_U3075 ; P2_R1233_U283
g17291 nand P2_R1233_U162 P2_R1233_U131 ; P2_R1233_U284
g17292 nand P2_R1233_U283 P2_R1233_U281 ; P2_R1233_U285
g17293 not P2_R1233_U159 ; P2_R1233_U286
g17294 or P2_U3974 P2_U3061 ; P2_R1233_U287
g17295 nand P2_R1233_U287 P2_R1233_U159 ; P2_R1233_U288
g17296 nand P2_U3061 P2_U3974 ; P2_R1233_U289
g17297 not P2_R1233_U157 ; P2_R1233_U290
g17298 or P2_U3973 P2_U3066 ; P2_R1233_U291
g17299 nand P2_R1233_U291 P2_R1233_U157 ; P2_R1233_U292
g17300 nand P2_U3066 P2_U3973 ; P2_R1233_U293
g17301 not P2_R1233_U155 ; P2_R1233_U294
g17302 or P2_U3058 P2_U3971 ; P2_R1233_U295
g17303 nand P2_R1233_U176 P2_R1233_U173 ; P2_R1233_U296
g17304 not P2_R1233_U86 ; P2_R1233_U297
g17305 or P2_U3972 P2_U3065 ; P2_R1233_U298
g17306 nand P2_R1233_U155 P2_R1233_U298 P2_R1233_U168 ; P2_R1233_U299
g17307 not P2_R1233_U154 ; P2_R1233_U300
g17308 or P2_U3969 P2_U3053 ; P2_R1233_U301
g17309 nand P2_U3053 P2_U3969 ; P2_R1233_U302
g17310 not P2_R1233_U152 ; P2_R1233_U303
g17311 nand P2_U3968 P2_R1233_U152 ; P2_R1233_U304
g17312 not P2_R1233_U150 ; P2_R1233_U305
g17313 nand P2_R1233_U298 P2_R1233_U155 ; P2_R1233_U306
g17314 not P2_R1233_U89 ; P2_R1233_U307
g17315 or P2_U3971 P2_U3058 ; P2_R1233_U308
g17316 nand P2_R1233_U308 P2_R1233_U89 ; P2_R1233_U309
g17317 nand P2_R1233_U135 P2_R1233_U309 ; P2_R1233_U310
g17318 nand P2_R1233_U307 P2_R1233_U173 ; P2_R1233_U311
g17319 nand P2_U3970 P2_U3057 ; P2_R1233_U312
g17320 nand P2_R1233_U311 P2_R1233_U312 P2_R1233_U168 ; P2_R1233_U313
g17321 or P2_U3058 P2_U3971 ; P2_R1233_U314
g17322 nand P2_R1233_U282 P2_R1233_U162 ; P2_R1233_U315
g17323 not P2_R1233_U91 ; P2_R1233_U316
g17324 nand P2_R1233_U9 P2_R1233_U91 ; P2_R1233_U317
g17325 nand P2_R1233_U136 P2_R1233_U317 ; P2_R1233_U318
g17326 nand P2_R1233_U317 P2_R1233_U278 ; P2_R1233_U319
g17327 nand P2_R1233_U453 P2_R1233_U319 ; P2_R1233_U320
g17328 or P2_U3506 P2_U3081 ; P2_R1233_U321
g17329 nand P2_R1233_U321 P2_R1233_U91 ; P2_R1233_U322
g17330 nand P2_R1233_U137 P2_R1233_U322 ; P2_R1233_U323
g17331 nand P2_R1233_U316 P2_R1233_U80 ; P2_R1233_U324
g17332 nand P2_U3076 P2_U3976 ; P2_R1233_U325
g17333 nand P2_R1233_U138 P2_R1233_U324 ; P2_R1233_U326
g17334 or P2_U3453 P2_U3078 ; P2_R1233_U327
g17335 not P2_R1233_U161 ; P2_R1233_U328
g17336 or P2_U3081 P2_U3506 ; P2_R1233_U329
g17337 or P2_U3498 P2_U3073 ; P2_R1233_U330
g17338 nand P2_R1233_U330 P2_R1233_U92 ; P2_R1233_U331
g17339 nand P2_R1233_U139 P2_R1233_U331 ; P2_R1233_U332
g17340 nand P2_R1233_U262 P2_R1233_U59 ; P2_R1233_U333
g17341 nand P2_U3501 P2_U3069 ; P2_R1233_U334
g17342 nand P2_R1233_U140 P2_R1233_U333 ; P2_R1233_U335
g17343 or P2_U3073 P2_U3498 ; P2_R1233_U336
g17344 nand P2_R1233_U250 P2_R1233_U167 ; P2_R1233_U337
g17345 not P2_R1233_U93 ; P2_R1233_U338
g17346 or P2_U3486 P2_U3072 ; P2_R1233_U339
g17347 nand P2_R1233_U339 P2_R1233_U93 ; P2_R1233_U340
g17348 nand P2_R1233_U141 P2_R1233_U340 ; P2_R1233_U341
g17349 nand P2_R1233_U338 P2_R1233_U172 ; P2_R1233_U342
g17350 nand P2_U3080 P2_U3489 ; P2_R1233_U343
g17351 nand P2_R1233_U142 P2_R1233_U342 ; P2_R1233_U344
g17352 or P2_U3072 P2_U3486 ; P2_R1233_U345
g17353 or P2_U3477 P2_U3083 ; P2_R1233_U346
g17354 nand P2_R1233_U346 P2_R1233_U40 ; P2_R1233_U347
g17355 nand P2_R1233_U143 P2_R1233_U347 ; P2_R1233_U348
g17356 nand P2_R1233_U206 P2_R1233_U171 ; P2_R1233_U349
g17357 nand P2_U3062 P2_U3480 ; P2_R1233_U350
g17358 nand P2_R1233_U144 P2_R1233_U349 ; P2_R1233_U351
g17359 nand P2_R1233_U207 P2_R1233_U171 ; P2_R1233_U352
g17360 nand P2_R1233_U204 P2_R1233_U63 ; P2_R1233_U353
g17361 nand P2_R1233_U214 P2_R1233_U22 ; P2_R1233_U354
g17362 nand P2_R1233_U228 P2_R1233_U34 ; P2_R1233_U355
g17363 nand P2_R1233_U231 P2_R1233_U180 ; P2_R1233_U356
g17364 nand P2_R1233_U314 P2_R1233_U173 ; P2_R1233_U357
g17365 nand P2_R1233_U298 P2_R1233_U176 ; P2_R1233_U358
g17366 nand P2_R1233_U329 P2_R1233_U80 ; P2_R1233_U359
g17367 nand P2_R1233_U282 P2_R1233_U77 ; P2_R1233_U360
g17368 nand P2_R1233_U336 P2_R1233_U59 ; P2_R1233_U361
g17369 nand P2_R1233_U345 P2_R1233_U172 ; P2_R1233_U362
g17370 nand P2_R1233_U250 P2_R1233_U68 ; P2_R1233_U363
g17371 nand P2_U3968 P2_U3054 ; P2_R1233_U364
g17372 nand P2_R1233_U296 P2_R1233_U168 ; P2_R1233_U365
g17373 nand P2_U3057 P2_R1233_U295 ; P2_R1233_U366
g17374 nand P2_U3970 P2_R1233_U295 ; P2_R1233_U367
g17375 nand P2_R1233_U296 P2_R1233_U168 P2_R1233_U301 ; P2_R1233_U368
g17376 nand P2_R1233_U155 P2_R1233_U168 P2_R1233_U133 ; P2_R1233_U369
g17377 nand P2_R1233_U297 P2_R1233_U301 ; P2_R1233_U370
g17378 nand P2_U3083 P2_R1233_U39 ; P2_R1233_U371
g17379 nand P2_U3477 P2_R1233_U38 ; P2_R1233_U372
g17380 nand P2_R1233_U372 P2_R1233_U371 ; P2_R1233_U373
g17381 nand P2_R1233_U352 P2_R1233_U40 ; P2_R1233_U374
g17382 nand P2_R1233_U373 P2_R1233_U206 ; P2_R1233_U375
g17383 nand P2_U3084 P2_R1233_U36 ; P2_R1233_U376
g17384 nand P2_U3474 P2_R1233_U37 ; P2_R1233_U377
g17385 nand P2_R1233_U377 P2_R1233_U376 ; P2_R1233_U378
g17386 nand P2_R1233_U353 P2_R1233_U145 ; P2_R1233_U379
g17387 nand P2_R1233_U203 P2_R1233_U378 ; P2_R1233_U380
g17388 nand P2_U3070 P2_R1233_U23 ; P2_R1233_U381
g17389 nand P2_U3471 P2_R1233_U21 ; P2_R1233_U382
g17390 nand P2_U3071 P2_R1233_U19 ; P2_R1233_U383
g17391 nand P2_U3468 P2_R1233_U20 ; P2_R1233_U384
g17392 nand P2_R1233_U384 P2_R1233_U383 ; P2_R1233_U385
g17393 nand P2_R1233_U354 P2_R1233_U41 ; P2_R1233_U386
g17394 nand P2_R1233_U385 P2_R1233_U195 ; P2_R1233_U387
g17395 nand P2_U3067 P2_R1233_U35 ; P2_R1233_U388
g17396 nand P2_U3465 P2_R1233_U26 ; P2_R1233_U389
g17397 nand P2_U3060 P2_R1233_U24 ; P2_R1233_U390
g17398 nand P2_U3462 P2_R1233_U25 ; P2_R1233_U391
g17399 nand P2_R1233_U391 P2_R1233_U390 ; P2_R1233_U392
g17400 nand P2_R1233_U355 P2_R1233_U44 ; P2_R1233_U393
g17401 nand P2_R1233_U392 P2_R1233_U221 ; P2_R1233_U394
g17402 nand P2_U3064 P2_R1233_U32 ; P2_R1233_U395
g17403 nand P2_U3459 P2_R1233_U33 ; P2_R1233_U396
g17404 nand P2_R1233_U396 P2_R1233_U395 ; P2_R1233_U397
g17405 nand P2_R1233_U356 P2_R1233_U146 ; P2_R1233_U398
g17406 nand P2_R1233_U230 P2_R1233_U397 ; P2_R1233_U399
g17407 nand P2_U3068 P2_R1233_U27 ; P2_R1233_U400
g17408 nand P2_U3456 P2_R1233_U28 ; P2_R1233_U401
g17409 nand P2_U3055 P2_R1233_U148 ; P2_R1233_U402
g17410 nand P2_U3979 P2_R1233_U147 ; P2_R1233_U403
g17411 nand P2_U3055 P2_R1233_U148 ; P2_R1233_U404
g17412 nand P2_U3979 P2_R1233_U147 ; P2_R1233_U405
g17413 nand P2_R1233_U405 P2_R1233_U404 ; P2_R1233_U406
g17414 nand P2_R1233_U149 P2_R1233_U150 ; P2_R1233_U407
g17415 nand P2_R1233_U305 P2_R1233_U406 ; P2_R1233_U408
g17416 nand P2_U3054 P2_R1233_U88 ; P2_R1233_U409
g17417 nand P2_U3968 P2_R1233_U87 ; P2_R1233_U410
g17418 nand P2_U3054 P2_R1233_U88 ; P2_R1233_U411
g17419 nand P2_U3968 P2_R1233_U87 ; P2_R1233_U412
g17420 nand P2_R1233_U412 P2_R1233_U411 ; P2_R1233_U413
g17421 nand P2_R1233_U151 P2_R1233_U152 ; P2_R1233_U414
g17422 nand P2_R1233_U303 P2_R1233_U413 ; P2_R1233_U415
g17423 nand P2_U3053 P2_R1233_U46 ; P2_R1233_U416
g17424 nand P2_U3969 P2_R1233_U47 ; P2_R1233_U417
g17425 nand P2_U3053 P2_R1233_U46 ; P2_R1233_U418
g17426 nand P2_U3969 P2_R1233_U47 ; P2_R1233_U419
g17427 nand P2_R1233_U419 P2_R1233_U418 ; P2_R1233_U420
g17428 nand P2_R1233_U153 P2_R1233_U154 ; P2_R1233_U421
g17429 nand P2_R1233_U300 P2_R1233_U420 ; P2_R1233_U422
g17430 nand P2_U3057 P2_R1233_U49 ; P2_R1233_U423
g17431 nand P2_U3970 P2_R1233_U48 ; P2_R1233_U424
g17432 nand P2_U3058 P2_R1233_U50 ; P2_R1233_U425
g17433 nand P2_U3971 P2_R1233_U51 ; P2_R1233_U426
g17434 nand P2_R1233_U426 P2_R1233_U425 ; P2_R1233_U427
g17435 nand P2_R1233_U357 P2_R1233_U89 ; P2_R1233_U428
g17436 nand P2_R1233_U427 P2_R1233_U307 ; P2_R1233_U429
g17437 nand P2_U3065 P2_R1233_U52 ; P2_R1233_U430
g17438 nand P2_U3972 P2_R1233_U53 ; P2_R1233_U431
g17439 nand P2_R1233_U431 P2_R1233_U430 ; P2_R1233_U432
g17440 nand P2_R1233_U358 P2_R1233_U155 ; P2_R1233_U433
g17441 nand P2_R1233_U294 P2_R1233_U432 ; P2_R1233_U434
g17442 nand P2_U3066 P2_R1233_U84 ; P2_R1233_U435
g17443 nand P2_U3973 P2_R1233_U85 ; P2_R1233_U436
g17444 nand P2_U3066 P2_R1233_U84 ; P2_R1233_U437
g17445 nand P2_U3973 P2_R1233_U85 ; P2_R1233_U438
g17446 nand P2_R1233_U438 P2_R1233_U437 ; P2_R1233_U439
g17447 nand P2_R1233_U156 P2_R1233_U157 ; P2_R1233_U440
g17448 nand P2_R1233_U290 P2_R1233_U439 ; P2_R1233_U441
g17449 nand P2_U3061 P2_R1233_U82 ; P2_R1233_U442
g17450 nand P2_U3974 P2_R1233_U83 ; P2_R1233_U443
g17451 nand P2_U3061 P2_R1233_U82 ; P2_R1233_U444
g17452 nand P2_U3974 P2_R1233_U83 ; P2_R1233_U445
g17453 nand P2_R1233_U445 P2_R1233_U444 ; P2_R1233_U446
g17454 nand P2_R1233_U158 P2_R1233_U159 ; P2_R1233_U447
g17455 nand P2_R1233_U286 P2_R1233_U446 ; P2_R1233_U448
g17456 nand P2_U3075 P2_R1233_U54 ; P2_R1233_U449
g17457 nand P2_U3975 P2_R1233_U55 ; P2_R1233_U450
g17458 nand P2_U3075 P2_R1233_U54 ; P2_R1233_U451
g17459 nand P2_U3975 P2_R1233_U55 ; P2_R1233_U452
g17460 nand P2_R1233_U452 P2_R1233_U451 ; P2_R1233_U453
g17461 nand P2_U3076 P2_R1233_U81 ; P2_R1233_U454
g17462 nand P2_U3976 P2_R1233_U90 ; P2_R1233_U455
g17463 nand P2_R1233_U182 P2_R1233_U161 ; P2_R1233_U456
g17464 nand P2_R1233_U328 P2_R1233_U31 ; P2_R1233_U457
g17465 nand P2_U3081 P2_R1233_U78 ; P2_R1233_U458
g17466 nand P2_U3506 P2_R1233_U79 ; P2_R1233_U459
g17467 nand P2_R1233_U459 P2_R1233_U458 ; P2_R1233_U460
g17468 nand P2_R1233_U359 P2_R1233_U91 ; P2_R1233_U461
g17469 nand P2_R1233_U460 P2_R1233_U316 ; P2_R1233_U462
g17470 nand P2_U3082 P2_R1233_U75 ; P2_R1233_U463
g17471 nand P2_U3504 P2_R1233_U76 ; P2_R1233_U464
g17472 nand P2_R1233_U464 P2_R1233_U463 ; P2_R1233_U465
g17473 nand P2_R1233_U360 P2_R1233_U162 ; P2_R1233_U466
g17474 nand P2_R1233_U270 P2_R1233_U465 ; P2_R1233_U467
g17475 nand P2_U3069 P2_R1233_U60 ; P2_R1233_U468
g17476 nand P2_U3501 P2_R1233_U58 ; P2_R1233_U469
g17477 nand P2_U3073 P2_R1233_U56 ; P2_R1233_U470
g17478 nand P2_U3498 P2_R1233_U57 ; P2_R1233_U471
g17479 nand P2_R1233_U471 P2_R1233_U470 ; P2_R1233_U472
g17480 nand P2_R1233_U361 P2_R1233_U92 ; P2_R1233_U473
g17481 nand P2_R1233_U472 P2_R1233_U262 ; P2_R1233_U474
g17482 nand P2_U3074 P2_R1233_U73 ; P2_R1233_U475
g17483 nand P2_U3495 P2_R1233_U74 ; P2_R1233_U476
g17484 nand P2_U3074 P2_R1233_U73 ; P2_R1233_U477
g17485 nand P2_U3495 P2_R1233_U74 ; P2_R1233_U478
g17486 nand P2_R1233_U478 P2_R1233_U477 ; P2_R1233_U479
g17487 nand P2_R1233_U163 P2_R1233_U164 ; P2_R1233_U480
g17488 nand P2_R1233_U258 P2_R1233_U479 ; P2_R1233_U481
g17489 nand P2_U3079 P2_R1233_U71 ; P2_R1233_U482
g17490 nand P2_U3492 P2_R1233_U72 ; P2_R1233_U483
g17491 nand P2_U3079 P2_R1233_U71 ; P2_R1233_U484
g17492 nand P2_U3492 P2_R1233_U72 ; P2_R1233_U485
g17493 nand P2_R1233_U485 P2_R1233_U484 ; P2_R1233_U486
g17494 nand P2_R1233_U165 P2_R1233_U166 ; P2_R1233_U487
g17495 nand P2_R1233_U254 P2_R1233_U486 ; P2_R1233_U488
g17496 nand P2_U3080 P2_R1233_U69 ; P2_R1233_U489
g17497 nand P2_U3489 P2_R1233_U70 ; P2_R1233_U490
g17498 nand P2_U3072 P2_R1233_U64 ; P2_R1233_U491
g17499 nand P2_U3486 P2_R1233_U65 ; P2_R1233_U492
g17500 nand P2_R1233_U492 P2_R1233_U491 ; P2_R1233_U493
g17501 nand P2_R1233_U362 P2_R1233_U93 ; P2_R1233_U494
g17502 nand P2_R1233_U493 P2_R1233_U338 ; P2_R1233_U495
g17503 nand P2_U3063 P2_R1233_U66 ; P2_R1233_U496
g17504 nand P2_U3483 P2_R1233_U67 ; P2_R1233_U497
g17505 nand P2_R1233_U497 P2_R1233_U496 ; P2_R1233_U498
g17506 nand P2_R1233_U363 P2_R1233_U167 ; P2_R1233_U499
g17507 nand P2_R1233_U244 P2_R1233_U498 ; P2_R1233_U500
g17508 nand P2_U3062 P2_R1233_U61 ; P2_R1233_U501
g17509 nand P2_U3480 P2_R1233_U62 ; P2_R1233_U502
g17510 nand P2_U3077 P2_R1233_U29 ; P2_R1233_U503
g17511 nand P2_U3448 P2_R1233_U30 ; P2_R1233_U504
g17512 and P2_R1176_U211 P2_R1176_U210 ; P2_R1176_U4
g17513 and P2_R1176_U224 P2_R1176_U223 ; P2_R1176_U5
g17514 and P2_R1176_U256 P2_R1176_U255 ; P2_R1176_U6
g17515 and P2_R1176_U274 P2_R1176_U273 ; P2_R1176_U7
g17516 and P2_R1176_U286 P2_R1176_U285 ; P2_R1176_U8
g17517 and P2_R1176_U344 P2_R1176_U341 ; P2_R1176_U9
g17518 and P2_R1176_U335 P2_R1176_U332 ; P2_R1176_U10
g17519 and P2_R1176_U328 P2_R1176_U325 ; P2_R1176_U11
g17520 and P2_R1176_U319 P2_R1176_U316 ; P2_R1176_U12
g17521 and P2_R1176_U247 P2_R1176_U244 ; P2_R1176_U13
g17522 and P2_R1176_U240 P2_R1176_U237 ; P2_R1176_U14
g17523 not P2_U3214 ; P2_R1176_U15
g17524 not P2_U3207 ; P2_R1176_U16
g17525 nand P2_U3207 P2_R1176_U56 ; P2_R1176_U17
g17526 not P2_U3206 ; P2_R1176_U18
g17527 not P2_U3211 ; P2_R1176_U19
g17528 nand P2_U3211 P2_R1176_U58 ; P2_R1176_U20
g17529 not P2_U3210 ; P2_R1176_U21
g17530 not P2_U3213 ; P2_R1176_U22
g17531 not P2_U3212 ; P2_R1176_U23
g17532 not P2_U3209 ; P2_R1176_U24
g17533 not P2_U3208 ; P2_R1176_U25
g17534 not P2_U3205 ; P2_R1176_U26
g17535 not P2_U3204 ; P2_R1176_U27
g17536 nand P2_R1176_U221 P2_R1176_U220 ; P2_R1176_U28
g17537 nand P2_R1176_U208 P2_R1176_U207 ; P2_R1176_U29
g17538 not P2_U3186 ; P2_R1176_U30
g17539 not P2_U3187 ; P2_R1176_U31
g17540 not P2_U3188 ; P2_R1176_U32
g17541 not P2_U3189 ; P2_R1176_U33
g17542 not P2_U3197 ; P2_R1176_U34
g17543 nand P2_U3197 P2_R1176_U69 ; P2_R1176_U35
g17544 not P2_U3196 ; P2_R1176_U36
g17545 not P2_U3203 ; P2_R1176_U37
g17546 not P2_U3201 ; P2_R1176_U38
g17547 not P2_U3202 ; P2_R1176_U39
g17548 nand P2_U3202 P2_R1176_U72 ; P2_R1176_U40
g17549 not P2_U3200 ; P2_R1176_U41
g17550 not P2_U3199 ; P2_R1176_U42
g17551 not P2_U3198 ; P2_R1176_U43
g17552 not P2_U3195 ; P2_R1176_U44
g17553 not P2_U3193 ; P2_R1176_U45
g17554 not P2_U3194 ; P2_R1176_U46
g17555 nand P2_U3194 P2_R1176_U78 ; P2_R1176_U47
g17556 not P2_U3192 ; P2_R1176_U48
g17557 not P2_U3191 ; P2_R1176_U49
g17558 not P2_U3190 ; P2_R1176_U50
g17559 nand P2_U3187 P2_R1176_U67 ; P2_R1176_U51
g17560 nand P2_R1176_U47 P2_R1176_U321 ; P2_R1176_U52
g17561 nand P2_R1176_U271 P2_R1176_U270 ; P2_R1176_U53
g17562 nand P2_R1176_U40 P2_R1176_U337 ; P2_R1176_U54
g17563 nand P2_R1176_U366 P2_R1176_U365 ; P2_R1176_U55
g17564 nand P2_R1176_U395 P2_R1176_U394 ; P2_R1176_U56
g17565 nand P2_R1176_U392 P2_R1176_U391 ; P2_R1176_U57
g17566 nand P2_R1176_U386 P2_R1176_U385 ; P2_R1176_U58
g17567 nand P2_R1176_U383 P2_R1176_U382 ; P2_R1176_U59
g17568 nand P2_R1176_U377 P2_R1176_U376 ; P2_R1176_U60
g17569 nand P2_R1176_U380 P2_R1176_U379 ; P2_R1176_U61
g17570 nand P2_R1176_U374 P2_R1176_U373 ; P2_R1176_U62
g17571 nand P2_R1176_U389 P2_R1176_U388 ; P2_R1176_U63
g17572 nand P2_R1176_U398 P2_R1176_U397 ; P2_R1176_U64
g17573 nand P2_R1176_U438 P2_R1176_U437 ; P2_R1176_U65
g17574 nand P2_R1176_U483 P2_R1176_U482 ; P2_R1176_U66
g17575 nand P2_R1176_U486 P2_R1176_U485 ; P2_R1176_U67
g17576 nand P2_R1176_U489 P2_R1176_U488 ; P2_R1176_U68
g17577 nand P2_R1176_U462 P2_R1176_U461 ; P2_R1176_U69
g17578 nand P2_R1176_U459 P2_R1176_U458 ; P2_R1176_U70
g17579 nand P2_R1176_U441 P2_R1176_U440 ; P2_R1176_U71
g17580 nand P2_R1176_U450 P2_R1176_U449 ; P2_R1176_U72
g17581 nand P2_R1176_U444 P2_R1176_U443 ; P2_R1176_U73
g17582 nand P2_R1176_U447 P2_R1176_U446 ; P2_R1176_U74
g17583 nand P2_R1176_U453 P2_R1176_U452 ; P2_R1176_U75
g17584 nand P2_R1176_U456 P2_R1176_U455 ; P2_R1176_U76
g17585 nand P2_R1176_U465 P2_R1176_U464 ; P2_R1176_U77
g17586 nand P2_R1176_U474 P2_R1176_U473 ; P2_R1176_U78
g17587 nand P2_R1176_U468 P2_R1176_U467 ; P2_R1176_U79
g17588 nand P2_R1176_U471 P2_R1176_U470 ; P2_R1176_U80
g17589 nand P2_R1176_U477 P2_R1176_U476 ; P2_R1176_U81
g17590 nand P2_R1176_U480 P2_R1176_U479 ; P2_R1176_U82
g17591 nand P2_R1176_U495 P2_R1176_U494 ; P2_R1176_U83
g17592 nand P2_R1176_U602 P2_R1176_U601 ; P2_R1176_U84
g17593 nand P2_R1176_U401 P2_R1176_U400 ; P2_R1176_U85
g17594 nand P2_R1176_U408 P2_R1176_U407 ; P2_R1176_U86
g17595 nand P2_R1176_U415 P2_R1176_U414 ; P2_R1176_U87
g17596 nand P2_R1176_U422 P2_R1176_U421 ; P2_R1176_U88
g17597 nand P2_R1176_U429 P2_R1176_U428 ; P2_R1176_U89
g17598 nand P2_R1176_U436 P2_R1176_U435 ; P2_R1176_U90
g17599 nand P2_R1176_U498 P2_R1176_U497 ; P2_R1176_U91
g17600 nand P2_R1176_U505 P2_R1176_U504 ; P2_R1176_U92
g17601 nand P2_R1176_U512 P2_R1176_U511 ; P2_R1176_U93
g17602 nand P2_R1176_U517 P2_R1176_U516 ; P2_R1176_U94
g17603 nand P2_R1176_U524 P2_R1176_U523 ; P2_R1176_U95
g17604 nand P2_R1176_U531 P2_R1176_U530 ; P2_R1176_U96
g17605 nand P2_R1176_U538 P2_R1176_U537 ; P2_R1176_U97
g17606 nand P2_R1176_U545 P2_R1176_U544 ; P2_R1176_U98
g17607 nand P2_R1176_U550 P2_R1176_U549 ; P2_R1176_U99
g17608 nand P2_R1176_U557 P2_R1176_U556 ; P2_R1176_U100
g17609 nand P2_R1176_U564 P2_R1176_U563 ; P2_R1176_U101
g17610 nand P2_R1176_U571 P2_R1176_U570 ; P2_R1176_U102
g17611 nand P2_R1176_U578 P2_R1176_U577 ; P2_R1176_U103
g17612 nand P2_R1176_U585 P2_R1176_U584 ; P2_R1176_U104
g17613 nand P2_R1176_U590 P2_R1176_U589 ; P2_R1176_U105
g17614 nand P2_R1176_U597 P2_R1176_U596 ; P2_R1176_U106
g17615 and P2_R1176_U214 P2_R1176_U213 ; P2_R1176_U107
g17616 and P2_R1176_U228 P2_R1176_U227 ; P2_R1176_U108
g17617 and P2_R1176_U410 P2_R1176_U409 P2_R1176_U17 ; P2_R1176_U109
g17618 and P2_R1176_U239 P2_R1176_U5 ; P2_R1176_U110
g17619 and P2_R1176_U431 P2_R1176_U430 P2_R1176_U20 ; P2_R1176_U111
g17620 and P2_R1176_U246 P2_R1176_U4 ; P2_R1176_U112
g17621 and P2_R1176_U260 P2_R1176_U6 ; P2_R1176_U113
g17622 and P2_R1176_U258 P2_R1176_U196 ; P2_R1176_U114
g17623 and P2_R1176_U278 P2_R1176_U277 ; P2_R1176_U115
g17624 and P2_R1176_U290 P2_R1176_U8 ; P2_R1176_U116
g17625 and P2_R1176_U288 P2_R1176_U197 ; P2_R1176_U117
g17626 and P2_R1176_U306 P2_R1176_U192 ; P2_R1176_U118
g17627 and P2_R1176_U364 P2_R1176_U51 ; P2_R1176_U119
g17628 and P2_R1176_U311 P2_R1176_U306 ; P2_R1176_U120
g17629 and P2_R1176_U361 P2_R1176_U310 ; P2_R1176_U121
g17630 nand P2_R1176_U492 P2_R1176_U491 ; P2_R1176_U122
g17631 and P2_R1176_U357 P2_R1176_U51 ; P2_R1176_U123
g17632 and P2_R1176_U507 P2_R1176_U506 P2_R1176_U198 ; P2_R1176_U124
g17633 and P2_R1176_U201 P2_R1176_U198 ; P2_R1176_U125
g17634 and P2_R1176_U318 P2_R1176_U192 ; P2_R1176_U126
g17635 and P2_R1176_U533 P2_R1176_U532 P2_R1176_U197 ; P2_R1176_U127
g17636 and P2_R1176_U327 P2_R1176_U8 ; P2_R1176_U128
g17637 and P2_R1176_U559 P2_R1176_U558 P2_R1176_U35 ; P2_R1176_U129
g17638 and P2_R1176_U334 P2_R1176_U7 ; P2_R1176_U130
g17639 and P2_R1176_U580 P2_R1176_U579 P2_R1176_U196 ; P2_R1176_U131
g17640 and P2_R1176_U343 P2_R1176_U6 ; P2_R1176_U132
g17641 nand P2_R1176_U599 P2_R1176_U598 ; P2_R1176_U133
g17642 not P2_U3477 ; P2_R1176_U134
g17643 and P2_R1176_U369 P2_R1176_U368 ; P2_R1176_U135
g17644 not P2_U3462 ; P2_R1176_U136
g17645 not P2_U3448 ; P2_R1176_U137
g17646 not P2_U3453 ; P2_R1176_U138
g17647 not P2_U3459 ; P2_R1176_U139
g17648 not P2_U3456 ; P2_R1176_U140
g17649 not P2_U3465 ; P2_R1176_U141
g17650 not P2_U3471 ; P2_R1176_U142
g17651 not P2_U3468 ; P2_R1176_U143
g17652 not P2_U3474 ; P2_R1176_U144
g17653 nand P2_R1176_U233 P2_R1176_U232 ; P2_R1176_U145
g17654 and P2_R1176_U403 P2_R1176_U402 ; P2_R1176_U146
g17655 nand P2_R1176_U108 P2_R1176_U229 ; P2_R1176_U147
g17656 and P2_R1176_U417 P2_R1176_U416 ; P2_R1176_U148
g17657 nand P2_R1176_U217 P2_R1176_U194 P2_R1176_U355 ; P2_R1176_U149
g17658 and P2_R1176_U424 P2_R1176_U423 ; P2_R1176_U150
g17659 nand P2_R1176_U107 P2_R1176_U215 ; P2_R1176_U151
g17660 not P2_U3969 ; P2_R1176_U152
g17661 not P2_U3480 ; P2_R1176_U153
g17662 not P2_U3489 ; P2_R1176_U154
g17663 not P2_U3486 ; P2_R1176_U155
g17664 not P2_U3483 ; P2_R1176_U156
g17665 not P2_U3492 ; P2_R1176_U157
g17666 not P2_U3495 ; P2_R1176_U158
g17667 not P2_U3501 ; P2_R1176_U159
g17668 not P2_U3498 ; P2_R1176_U160
g17669 not P2_U3504 ; P2_R1176_U161
g17670 not P2_U3975 ; P2_R1176_U162
g17671 not P2_U3976 ; P2_R1176_U163
g17672 not P2_U3506 ; P2_R1176_U164
g17673 not P2_U3974 ; P2_R1176_U165
g17674 not P2_U3973 ; P2_R1176_U166
g17675 not P2_U3971 ; P2_R1176_U167
g17676 not P2_U3970 ; P2_R1176_U168
g17677 not P2_U3972 ; P2_R1176_U169
g17678 not P2_U3185 ; P2_R1176_U170
g17679 not P2_U3968 ; P2_R1176_U171
g17680 and P2_R1176_U500 P2_R1176_U499 ; P2_R1176_U172
g17681 nand P2_R1176_U123 P2_R1176_U307 ; P2_R1176_U173
g17682 nand P2_R1176_U201 P2_R1176_U312 ; P2_R1176_U174
g17683 nand P2_R1176_U301 P2_R1176_U300 ; P2_R1176_U175
g17684 and P2_R1176_U519 P2_R1176_U518 ; P2_R1176_U176
g17685 nand P2_R1176_U297 P2_R1176_U296 ; P2_R1176_U177
g17686 and P2_R1176_U526 P2_R1176_U525 ; P2_R1176_U178
g17687 nand P2_R1176_U293 P2_R1176_U292 ; P2_R1176_U179
g17688 and P2_R1176_U540 P2_R1176_U539 ; P2_R1176_U180
g17689 nand P2_R1176_U204 P2_R1176_U203 ; P2_R1176_U181
g17690 nand P2_R1176_U283 P2_R1176_U282 ; P2_R1176_U182
g17691 and P2_R1176_U552 P2_R1176_U551 ; P2_R1176_U183
g17692 nand P2_R1176_U115 P2_R1176_U279 ; P2_R1176_U184
g17693 and P2_R1176_U566 P2_R1176_U565 ; P2_R1176_U185
g17694 nand P2_R1176_U267 P2_R1176_U266 ; P2_R1176_U186
g17695 and P2_R1176_U573 P2_R1176_U572 ; P2_R1176_U187
g17696 nand P2_R1176_U263 P2_R1176_U262 ; P2_R1176_U188
g17697 nand P2_R1176_U253 P2_R1176_U252 ; P2_R1176_U189
g17698 and P2_R1176_U592 P2_R1176_U591 ; P2_R1176_U190
g17699 nand P2_R1176_U249 P2_R1176_U193 P2_R1176_U360 ; P2_R1176_U191
g17700 nand P2_R1176_U359 P2_R1176_U358 ; P2_R1176_U192
g17701 nand P2_R1176_U55 P2_R1176_U145 ; P2_R1176_U193
g17702 nand P2_R1176_U62 P2_R1176_U151 ; P2_R1176_U194
g17703 not P2_R1176_U20 ; P2_R1176_U195
g17704 nand P2_U3201 P2_R1176_U74 ; P2_R1176_U196
g17705 nand P2_U3193 P2_R1176_U80 ; P2_R1176_U197
g17706 nand P2_U3188 P2_R1176_U66 ; P2_R1176_U198
g17707 not P2_R1176_U40 ; P2_R1176_U199
g17708 not P2_R1176_U47 ; P2_R1176_U200
g17709 nand P2_U3189 P2_R1176_U68 ; P2_R1176_U201
g17710 nand P2_R1176_U378 P2_R1176_U15 ; P2_R1176_U202
g17711 nand P2_U3213 P2_R1176_U202 ; P2_R1176_U203
g17712 nand P2_U3214 P2_R1176_U60 ; P2_R1176_U204
g17713 not P2_R1176_U181 ; P2_R1176_U205
g17714 nand P2_R1176_U381 P2_R1176_U23 ; P2_R1176_U206
g17715 nand P2_R1176_U206 P2_R1176_U181 ; P2_R1176_U207
g17716 nand P2_U3212 P2_R1176_U61 ; P2_R1176_U208
g17717 not P2_R1176_U29 ; P2_R1176_U209
g17718 nand P2_R1176_U384 P2_R1176_U21 ; P2_R1176_U210
g17719 nand P2_R1176_U387 P2_R1176_U19 ; P2_R1176_U211
g17720 nand P2_R1176_U21 P2_R1176_U20 ; P2_R1176_U212
g17721 nand P2_R1176_U59 P2_R1176_U212 ; P2_R1176_U213
g17722 nand P2_U3210 P2_R1176_U195 ; P2_R1176_U214
g17723 nand P2_R1176_U4 P2_R1176_U29 ; P2_R1176_U215
g17724 not P2_R1176_U151 ; P2_R1176_U216
g17725 nand P2_U3209 P2_R1176_U151 ; P2_R1176_U217
g17726 not P2_R1176_U149 ; P2_R1176_U218
g17727 nand P2_R1176_U390 P2_R1176_U25 ; P2_R1176_U219
g17728 nand P2_R1176_U219 P2_R1176_U149 ; P2_R1176_U220
g17729 nand P2_U3208 P2_R1176_U63 ; P2_R1176_U221
g17730 not P2_R1176_U28 ; P2_R1176_U222
g17731 nand P2_R1176_U393 P2_R1176_U18 ; P2_R1176_U223
g17732 nand P2_R1176_U396 P2_R1176_U16 ; P2_R1176_U224
g17733 not P2_R1176_U17 ; P2_R1176_U225
g17734 nand P2_R1176_U18 P2_R1176_U17 ; P2_R1176_U226
g17735 nand P2_R1176_U57 P2_R1176_U226 ; P2_R1176_U227
g17736 nand P2_U3206 P2_R1176_U225 ; P2_R1176_U228
g17737 nand P2_R1176_U5 P2_R1176_U28 ; P2_R1176_U229
g17738 not P2_R1176_U147 ; P2_R1176_U230
g17739 nand P2_R1176_U399 P2_R1176_U26 ; P2_R1176_U231
g17740 nand P2_R1176_U231 P2_R1176_U147 ; P2_R1176_U232
g17741 nand P2_U3205 P2_R1176_U64 ; P2_R1176_U233
g17742 not P2_R1176_U145 ; P2_R1176_U234
g17743 nand P2_R1176_U396 P2_R1176_U16 ; P2_R1176_U235
g17744 nand P2_R1176_U235 P2_R1176_U28 ; P2_R1176_U236
g17745 nand P2_R1176_U109 P2_R1176_U236 ; P2_R1176_U237
g17746 nand P2_R1176_U222 P2_R1176_U17 ; P2_R1176_U238
g17747 nand P2_U3206 P2_R1176_U57 ; P2_R1176_U239
g17748 nand P2_R1176_U110 P2_R1176_U238 ; P2_R1176_U240
g17749 nand P2_R1176_U396 P2_R1176_U16 ; P2_R1176_U241
g17750 nand P2_R1176_U387 P2_R1176_U19 ; P2_R1176_U242
g17751 nand P2_R1176_U242 P2_R1176_U29 ; P2_R1176_U243
g17752 nand P2_R1176_U111 P2_R1176_U243 ; P2_R1176_U244
g17753 nand P2_R1176_U209 P2_R1176_U20 ; P2_R1176_U245
g17754 nand P2_U3210 P2_R1176_U59 ; P2_R1176_U246
g17755 nand P2_R1176_U112 P2_R1176_U245 ; P2_R1176_U247
g17756 nand P2_R1176_U387 P2_R1176_U19 ; P2_R1176_U248
g17757 nand P2_U3204 P2_R1176_U145 ; P2_R1176_U249
g17758 not P2_R1176_U191 ; P2_R1176_U250
g17759 nand P2_R1176_U442 P2_R1176_U37 ; P2_R1176_U251
g17760 nand P2_R1176_U251 P2_R1176_U191 ; P2_R1176_U252
g17761 nand P2_U3203 P2_R1176_U71 ; P2_R1176_U253
g17762 not P2_R1176_U189 ; P2_R1176_U254
g17763 nand P2_R1176_U445 P2_R1176_U41 ; P2_R1176_U255
g17764 nand P2_R1176_U448 P2_R1176_U38 ; P2_R1176_U256
g17765 nand P2_R1176_U199 P2_R1176_U6 ; P2_R1176_U257
g17766 nand P2_U3200 P2_R1176_U73 ; P2_R1176_U258
g17767 nand P2_R1176_U114 P2_R1176_U257 ; P2_R1176_U259
g17768 nand P2_R1176_U451 P2_R1176_U39 ; P2_R1176_U260
g17769 nand P2_R1176_U445 P2_R1176_U41 ; P2_R1176_U261
g17770 nand P2_R1176_U113 P2_R1176_U189 ; P2_R1176_U262
g17771 nand P2_R1176_U261 P2_R1176_U259 ; P2_R1176_U263
g17772 not P2_R1176_U188 ; P2_R1176_U264
g17773 nand P2_R1176_U454 P2_R1176_U42 ; P2_R1176_U265
g17774 nand P2_R1176_U265 P2_R1176_U188 ; P2_R1176_U266
g17775 nand P2_U3199 P2_R1176_U75 ; P2_R1176_U267
g17776 not P2_R1176_U186 ; P2_R1176_U268
g17777 nand P2_R1176_U457 P2_R1176_U43 ; P2_R1176_U269
g17778 nand P2_R1176_U269 P2_R1176_U186 ; P2_R1176_U270
g17779 nand P2_U3198 P2_R1176_U76 ; P2_R1176_U271
g17780 not P2_R1176_U53 ; P2_R1176_U272
g17781 nand P2_R1176_U460 P2_R1176_U36 ; P2_R1176_U273
g17782 nand P2_R1176_U463 P2_R1176_U34 ; P2_R1176_U274
g17783 not P2_R1176_U35 ; P2_R1176_U275
g17784 nand P2_R1176_U36 P2_R1176_U35 ; P2_R1176_U276
g17785 nand P2_R1176_U70 P2_R1176_U276 ; P2_R1176_U277
g17786 nand P2_U3196 P2_R1176_U275 ; P2_R1176_U278
g17787 nand P2_R1176_U7 P2_R1176_U53 ; P2_R1176_U279
g17788 not P2_R1176_U184 ; P2_R1176_U280
g17789 nand P2_R1176_U466 P2_R1176_U44 ; P2_R1176_U281
g17790 nand P2_R1176_U281 P2_R1176_U184 ; P2_R1176_U282
g17791 nand P2_U3195 P2_R1176_U77 ; P2_R1176_U283
g17792 not P2_R1176_U182 ; P2_R1176_U284
g17793 nand P2_R1176_U469 P2_R1176_U48 ; P2_R1176_U285
g17794 nand P2_R1176_U472 P2_R1176_U45 ; P2_R1176_U286
g17795 nand P2_R1176_U200 P2_R1176_U8 ; P2_R1176_U287
g17796 nand P2_U3192 P2_R1176_U79 ; P2_R1176_U288
g17797 nand P2_R1176_U117 P2_R1176_U287 ; P2_R1176_U289
g17798 nand P2_R1176_U475 P2_R1176_U46 ; P2_R1176_U290
g17799 nand P2_R1176_U469 P2_R1176_U48 ; P2_R1176_U291
g17800 nand P2_R1176_U116 P2_R1176_U182 ; P2_R1176_U292
g17801 nand P2_R1176_U291 P2_R1176_U289 ; P2_R1176_U293
g17802 not P2_R1176_U179 ; P2_R1176_U294
g17803 nand P2_R1176_U478 P2_R1176_U49 ; P2_R1176_U295
g17804 nand P2_R1176_U295 P2_R1176_U179 ; P2_R1176_U296
g17805 nand P2_U3191 P2_R1176_U81 ; P2_R1176_U297
g17806 not P2_R1176_U177 ; P2_R1176_U298
g17807 nand P2_R1176_U481 P2_R1176_U50 ; P2_R1176_U299
g17808 nand P2_R1176_U299 P2_R1176_U177 ; P2_R1176_U300
g17809 nand P2_U3190 P2_R1176_U82 ; P2_R1176_U301
g17810 not P2_R1176_U175 ; P2_R1176_U302
g17811 nand P2_R1176_U484 P2_R1176_U32 ; P2_R1176_U303
g17812 nand P2_R1176_U201 P2_R1176_U198 ; P2_R1176_U304
g17813 not P2_R1176_U51 ; P2_R1176_U305
g17814 nand P2_R1176_U490 P2_R1176_U33 ; P2_R1176_U306
g17815 nand P2_R1176_U118 P2_R1176_U175 ; P2_R1176_U307
g17816 not P2_R1176_U173 ; P2_R1176_U308
g17817 nand P2_R1176_U439 P2_R1176_U30 ; P2_R1176_U309
g17818 nand P2_U3186 P2_R1176_U65 ; P2_R1176_U310
g17819 nand P2_R1176_U439 P2_R1176_U30 ; P2_R1176_U311
g17820 nand P2_R1176_U306 P2_R1176_U175 ; P2_R1176_U312
g17821 not P2_R1176_U174 ; P2_R1176_U313
g17822 nand P2_R1176_U484 P2_R1176_U32 ; P2_R1176_U314
g17823 nand P2_R1176_U314 P2_R1176_U174 ; P2_R1176_U315
g17824 nand P2_R1176_U124 P2_R1176_U315 ; P2_R1176_U316
g17825 nand P2_R1176_U125 P2_R1176_U312 ; P2_R1176_U317
g17826 nand P2_U3187 P2_R1176_U67 ; P2_R1176_U318
g17827 nand P2_R1176_U126 P2_R1176_U317 ; P2_R1176_U319
g17828 nand P2_R1176_U484 P2_R1176_U32 ; P2_R1176_U320
g17829 nand P2_R1176_U290 P2_R1176_U182 ; P2_R1176_U321
g17830 not P2_R1176_U52 ; P2_R1176_U322
g17831 nand P2_R1176_U472 P2_R1176_U45 ; P2_R1176_U323
g17832 nand P2_R1176_U323 P2_R1176_U52 ; P2_R1176_U324
g17833 nand P2_R1176_U127 P2_R1176_U324 ; P2_R1176_U325
g17834 nand P2_R1176_U322 P2_R1176_U197 ; P2_R1176_U326
g17835 nand P2_U3192 P2_R1176_U79 ; P2_R1176_U327
g17836 nand P2_R1176_U128 P2_R1176_U326 ; P2_R1176_U328
g17837 nand P2_R1176_U472 P2_R1176_U45 ; P2_R1176_U329
g17838 nand P2_R1176_U463 P2_R1176_U34 ; P2_R1176_U330
g17839 nand P2_R1176_U330 P2_R1176_U53 ; P2_R1176_U331
g17840 nand P2_R1176_U129 P2_R1176_U331 ; P2_R1176_U332
g17841 nand P2_R1176_U272 P2_R1176_U35 ; P2_R1176_U333
g17842 nand P2_U3196 P2_R1176_U70 ; P2_R1176_U334
g17843 nand P2_R1176_U130 P2_R1176_U333 ; P2_R1176_U335
g17844 nand P2_R1176_U463 P2_R1176_U34 ; P2_R1176_U336
g17845 nand P2_R1176_U260 P2_R1176_U189 ; P2_R1176_U337
g17846 not P2_R1176_U54 ; P2_R1176_U338
g17847 nand P2_R1176_U448 P2_R1176_U38 ; P2_R1176_U339
g17848 nand P2_R1176_U339 P2_R1176_U54 ; P2_R1176_U340
g17849 nand P2_R1176_U131 P2_R1176_U340 ; P2_R1176_U341
g17850 nand P2_R1176_U338 P2_R1176_U196 ; P2_R1176_U342
g17851 nand P2_U3200 P2_R1176_U73 ; P2_R1176_U343
g17852 nand P2_R1176_U132 P2_R1176_U342 ; P2_R1176_U344
g17853 nand P2_R1176_U448 P2_R1176_U38 ; P2_R1176_U345
g17854 nand P2_R1176_U241 P2_R1176_U17 ; P2_R1176_U346
g17855 nand P2_R1176_U248 P2_R1176_U20 ; P2_R1176_U347
g17856 nand P2_R1176_U320 P2_R1176_U198 ; P2_R1176_U348
g17857 nand P2_R1176_U306 P2_R1176_U201 ; P2_R1176_U349
g17858 nand P2_R1176_U329 P2_R1176_U197 ; P2_R1176_U350
g17859 nand P2_R1176_U290 P2_R1176_U47 ; P2_R1176_U351
g17860 nand P2_R1176_U336 P2_R1176_U35 ; P2_R1176_U352
g17861 nand P2_R1176_U345 P2_R1176_U196 ; P2_R1176_U353
g17862 nand P2_R1176_U260 P2_R1176_U40 ; P2_R1176_U354
g17863 nand P2_U3209 P2_R1176_U62 ; P2_R1176_U355
g17864 nand P2_R1176_U357 P2_R1176_U307 P2_R1176_U119 ; P2_R1176_U356
g17865 nand P2_R1176_U304 P2_R1176_U192 ; P2_R1176_U357
g17866 nand P2_R1176_U67 P2_R1176_U303 ; P2_R1176_U358
g17867 nand P2_U3187 P2_R1176_U303 ; P2_R1176_U359
g17868 nand P2_U3204 P2_R1176_U55 ; P2_R1176_U360
g17869 nand P2_R1176_U304 P2_R1176_U192 P2_R1176_U311 ; P2_R1176_U361
g17870 nand P2_R1176_U175 P2_R1176_U192 P2_R1176_U120 ; P2_R1176_U362
g17871 nand P2_R1176_U305 P2_R1176_U311 ; P2_R1176_U363
g17872 nand P2_U3186 P2_R1176_U65 ; P2_R1176_U364
g17873 nand P2_U3214 P2_R1176_U134 ; P2_R1176_U365
g17874 nand P2_U3477 P2_R1176_U15 ; P2_R1176_U366
g17875 not P2_R1176_U55 ; P2_R1176_U367
g17876 nand P2_R1176_U367 P2_U3204 ; P2_R1176_U368
g17877 nand P2_R1176_U55 P2_R1176_U27 ; P2_R1176_U369
g17878 nand P2_R1176_U367 P2_U3204 ; P2_R1176_U370
g17879 nand P2_R1176_U55 P2_R1176_U27 ; P2_R1176_U371
g17880 nand P2_R1176_U371 P2_R1176_U370 ; P2_R1176_U372
g17881 nand P2_U3214 P2_R1176_U136 ; P2_R1176_U373
g17882 nand P2_U3462 P2_R1176_U15 ; P2_R1176_U374
g17883 not P2_R1176_U62 ; P2_R1176_U375
g17884 nand P2_U3214 P2_R1176_U137 ; P2_R1176_U376
g17885 nand P2_U3448 P2_R1176_U15 ; P2_R1176_U377
g17886 not P2_R1176_U60 ; P2_R1176_U378
g17887 nand P2_U3214 P2_R1176_U138 ; P2_R1176_U379
g17888 nand P2_U3453 P2_R1176_U15 ; P2_R1176_U380
g17889 not P2_R1176_U61 ; P2_R1176_U381
g17890 nand P2_U3214 P2_R1176_U139 ; P2_R1176_U382
g17891 nand P2_U3459 P2_R1176_U15 ; P2_R1176_U383
g17892 not P2_R1176_U59 ; P2_R1176_U384
g17893 nand P2_U3214 P2_R1176_U140 ; P2_R1176_U385
g17894 nand P2_U3456 P2_R1176_U15 ; P2_R1176_U386
g17895 not P2_R1176_U58 ; P2_R1176_U387
g17896 nand P2_U3214 P2_R1176_U141 ; P2_R1176_U388
g17897 nand P2_U3465 P2_R1176_U15 ; P2_R1176_U389
g17898 not P2_R1176_U63 ; P2_R1176_U390
g17899 nand P2_U3214 P2_R1176_U142 ; P2_R1176_U391
g17900 nand P2_U3471 P2_R1176_U15 ; P2_R1176_U392
g17901 not P2_R1176_U57 ; P2_R1176_U393
g17902 nand P2_U3214 P2_R1176_U143 ; P2_R1176_U394
g17903 nand P2_U3468 P2_R1176_U15 ; P2_R1176_U395
g17904 not P2_R1176_U56 ; P2_R1176_U396
g17905 nand P2_U3214 P2_R1176_U144 ; P2_R1176_U397
g17906 nand P2_U3474 P2_R1176_U15 ; P2_R1176_U398
g17907 not P2_R1176_U64 ; P2_R1176_U399
g17908 nand P2_R1176_U135 P2_R1176_U145 ; P2_R1176_U400
g17909 nand P2_R1176_U234 P2_R1176_U372 ; P2_R1176_U401
g17910 nand P2_R1176_U399 P2_U3205 ; P2_R1176_U402
g17911 nand P2_R1176_U64 P2_R1176_U26 ; P2_R1176_U403
g17912 nand P2_R1176_U399 P2_U3205 ; P2_R1176_U404
g17913 nand P2_R1176_U64 P2_R1176_U26 ; P2_R1176_U405
g17914 nand P2_R1176_U405 P2_R1176_U404 ; P2_R1176_U406
g17915 nand P2_R1176_U146 P2_R1176_U147 ; P2_R1176_U407
g17916 nand P2_R1176_U230 P2_R1176_U406 ; P2_R1176_U408
g17917 nand P2_R1176_U393 P2_U3206 ; P2_R1176_U409
g17918 nand P2_R1176_U57 P2_R1176_U18 ; P2_R1176_U410
g17919 nand P2_R1176_U396 P2_U3207 ; P2_R1176_U411
g17920 nand P2_R1176_U56 P2_R1176_U16 ; P2_R1176_U412
g17921 nand P2_R1176_U412 P2_R1176_U411 ; P2_R1176_U413
g17922 nand P2_R1176_U346 P2_R1176_U28 ; P2_R1176_U414
g17923 nand P2_R1176_U413 P2_R1176_U222 ; P2_R1176_U415
g17924 nand P2_R1176_U390 P2_U3208 ; P2_R1176_U416
g17925 nand P2_R1176_U63 P2_R1176_U25 ; P2_R1176_U417
g17926 nand P2_R1176_U390 P2_U3208 ; P2_R1176_U418
g17927 nand P2_R1176_U63 P2_R1176_U25 ; P2_R1176_U419
g17928 nand P2_R1176_U419 P2_R1176_U418 ; P2_R1176_U420
g17929 nand P2_R1176_U148 P2_R1176_U149 ; P2_R1176_U421
g17930 nand P2_R1176_U218 P2_R1176_U420 ; P2_R1176_U422
g17931 nand P2_R1176_U375 P2_U3209 ; P2_R1176_U423
g17932 nand P2_R1176_U62 P2_R1176_U24 ; P2_R1176_U424
g17933 nand P2_R1176_U375 P2_U3209 ; P2_R1176_U425
g17934 nand P2_R1176_U62 P2_R1176_U24 ; P2_R1176_U426
g17935 nand P2_R1176_U426 P2_R1176_U425 ; P2_R1176_U427
g17936 nand P2_R1176_U150 P2_R1176_U151 ; P2_R1176_U428
g17937 nand P2_R1176_U216 P2_R1176_U427 ; P2_R1176_U429
g17938 nand P2_R1176_U384 P2_U3210 ; P2_R1176_U430
g17939 nand P2_R1176_U59 P2_R1176_U21 ; P2_R1176_U431
g17940 nand P2_R1176_U387 P2_U3211 ; P2_R1176_U432
g17941 nand P2_R1176_U58 P2_R1176_U19 ; P2_R1176_U433
g17942 nand P2_R1176_U433 P2_R1176_U432 ; P2_R1176_U434
g17943 nand P2_R1176_U347 P2_R1176_U29 ; P2_R1176_U435
g17944 nand P2_R1176_U434 P2_R1176_U209 ; P2_R1176_U436
g17945 nand P2_U3214 P2_R1176_U152 ; P2_R1176_U437
g17946 nand P2_U3969 P2_R1176_U15 ; P2_R1176_U438
g17947 not P2_R1176_U65 ; P2_R1176_U439
g17948 nand P2_U3214 P2_R1176_U153 ; P2_R1176_U440
g17949 nand P2_U3480 P2_R1176_U15 ; P2_R1176_U441
g17950 not P2_R1176_U71 ; P2_R1176_U442
g17951 nand P2_U3214 P2_R1176_U154 ; P2_R1176_U443
g17952 nand P2_U3489 P2_R1176_U15 ; P2_R1176_U444
g17953 not P2_R1176_U73 ; P2_R1176_U445
g17954 nand P2_U3214 P2_R1176_U155 ; P2_R1176_U446
g17955 nand P2_U3486 P2_R1176_U15 ; P2_R1176_U447
g17956 not P2_R1176_U74 ; P2_R1176_U448
g17957 nand P2_U3214 P2_R1176_U156 ; P2_R1176_U449
g17958 nand P2_U3483 P2_R1176_U15 ; P2_R1176_U450
g17959 not P2_R1176_U72 ; P2_R1176_U451
g17960 nand P2_U3214 P2_R1176_U157 ; P2_R1176_U452
g17961 nand P2_U3492 P2_R1176_U15 ; P2_R1176_U453
g17962 not P2_R1176_U75 ; P2_R1176_U454
g17963 nand P2_U3214 P2_R1176_U158 ; P2_R1176_U455
g17964 nand P2_U3495 P2_R1176_U15 ; P2_R1176_U456
g17965 not P2_R1176_U76 ; P2_R1176_U457
g17966 nand P2_U3214 P2_R1176_U159 ; P2_R1176_U458
g17967 nand P2_U3501 P2_R1176_U15 ; P2_R1176_U459
g17968 not P2_R1176_U70 ; P2_R1176_U460
g17969 nand P2_U3214 P2_R1176_U160 ; P2_R1176_U461
g17970 nand P2_U3498 P2_R1176_U15 ; P2_R1176_U462
g17971 not P2_R1176_U69 ; P2_R1176_U463
g17972 nand P2_U3214 P2_R1176_U161 ; P2_R1176_U464
g17973 nand P2_U3504 P2_R1176_U15 ; P2_R1176_U465
g17974 not P2_R1176_U77 ; P2_R1176_U466
g17975 nand P2_U3214 P2_R1176_U162 ; P2_R1176_U467
g17976 nand P2_U3975 P2_R1176_U15 ; P2_R1176_U468
g17977 not P2_R1176_U79 ; P2_R1176_U469
g17978 nand P2_U3214 P2_R1176_U163 ; P2_R1176_U470
g17979 nand P2_U3976 P2_R1176_U15 ; P2_R1176_U471
g17980 not P2_R1176_U80 ; P2_R1176_U472
g17981 nand P2_U3214 P2_R1176_U164 ; P2_R1176_U473
g17982 nand P2_U3506 P2_R1176_U15 ; P2_R1176_U474
g17983 not P2_R1176_U78 ; P2_R1176_U475
g17984 nand P2_U3214 P2_R1176_U165 ; P2_R1176_U476
g17985 nand P2_U3974 P2_R1176_U15 ; P2_R1176_U477
g17986 not P2_R1176_U81 ; P2_R1176_U478
g17987 nand P2_U3214 P2_R1176_U166 ; P2_R1176_U479
g17988 nand P2_U3973 P2_R1176_U15 ; P2_R1176_U480
g17989 not P2_R1176_U82 ; P2_R1176_U481
g17990 nand P2_U3214 P2_R1176_U167 ; P2_R1176_U482
g17991 nand P2_U3971 P2_R1176_U15 ; P2_R1176_U483
g17992 not P2_R1176_U66 ; P2_R1176_U484
g17993 nand P2_U3214 P2_R1176_U168 ; P2_R1176_U485
g17994 nand P2_U3970 P2_R1176_U15 ; P2_R1176_U486
g17995 not P2_R1176_U67 ; P2_R1176_U487
g17996 nand P2_U3214 P2_R1176_U169 ; P2_R1176_U488
g17997 nand P2_U3972 P2_R1176_U15 ; P2_R1176_U489
g17998 not P2_R1176_U68 ; P2_R1176_U490
g17999 nand P2_U3214 P2_R1176_U170 ; P2_R1176_U491
g18000 nand P2_U3185 P2_R1176_U15 ; P2_R1176_U492
g18001 not P2_R1176_U122 ; P2_R1176_U493
g18002 nand P2_U3968 P2_R1176_U493 ; P2_R1176_U494
g18003 nand P2_R1176_U122 P2_R1176_U171 ; P2_R1176_U495
g18004 not P2_R1176_U83 ; P2_R1176_U496
g18005 nand P2_R1176_U356 P2_R1176_U309 P2_R1176_U496 ; P2_R1176_U497
g18006 nand P2_R1176_U363 P2_R1176_U362 P2_R1176_U121 P2_R1176_U83 ; P2_R1176_U498
g18007 nand P2_R1176_U439 P2_U3186 ; P2_R1176_U499
g18008 nand P2_R1176_U65 P2_R1176_U30 ; P2_R1176_U500
g18009 nand P2_R1176_U439 P2_U3186 ; P2_R1176_U501
g18010 nand P2_R1176_U65 P2_R1176_U30 ; P2_R1176_U502
g18011 nand P2_R1176_U502 P2_R1176_U501 ; P2_R1176_U503
g18012 nand P2_R1176_U172 P2_R1176_U173 ; P2_R1176_U504
g18013 nand P2_R1176_U308 P2_R1176_U503 ; P2_R1176_U505
g18014 nand P2_R1176_U487 P2_U3187 ; P2_R1176_U506
g18015 nand P2_R1176_U67 P2_R1176_U31 ; P2_R1176_U507
g18016 nand P2_R1176_U484 P2_U3188 ; P2_R1176_U508
g18017 nand P2_R1176_U66 P2_R1176_U32 ; P2_R1176_U509
g18018 nand P2_R1176_U509 P2_R1176_U508 ; P2_R1176_U510
g18019 nand P2_R1176_U348 P2_R1176_U174 ; P2_R1176_U511
g18020 nand P2_R1176_U313 P2_R1176_U510 ; P2_R1176_U512
g18021 nand P2_R1176_U490 P2_U3189 ; P2_R1176_U513
g18022 nand P2_R1176_U68 P2_R1176_U33 ; P2_R1176_U514
g18023 nand P2_R1176_U514 P2_R1176_U513 ; P2_R1176_U515
g18024 nand P2_R1176_U349 P2_R1176_U175 ; P2_R1176_U516
g18025 nand P2_R1176_U302 P2_R1176_U515 ; P2_R1176_U517
g18026 nand P2_R1176_U481 P2_U3190 ; P2_R1176_U518
g18027 nand P2_R1176_U82 P2_R1176_U50 ; P2_R1176_U519
g18028 nand P2_R1176_U481 P2_U3190 ; P2_R1176_U520
g18029 nand P2_R1176_U82 P2_R1176_U50 ; P2_R1176_U521
g18030 nand P2_R1176_U521 P2_R1176_U520 ; P2_R1176_U522
g18031 nand P2_R1176_U176 P2_R1176_U177 ; P2_R1176_U523
g18032 nand P2_R1176_U298 P2_R1176_U522 ; P2_R1176_U524
g18033 nand P2_R1176_U478 P2_U3191 ; P2_R1176_U525
g18034 nand P2_R1176_U81 P2_R1176_U49 ; P2_R1176_U526
g18035 nand P2_R1176_U478 P2_U3191 ; P2_R1176_U527
g18036 nand P2_R1176_U81 P2_R1176_U49 ; P2_R1176_U528
g18037 nand P2_R1176_U528 P2_R1176_U527 ; P2_R1176_U529
g18038 nand P2_R1176_U178 P2_R1176_U179 ; P2_R1176_U530
g18039 nand P2_R1176_U294 P2_R1176_U529 ; P2_R1176_U531
g18040 nand P2_R1176_U469 P2_U3192 ; P2_R1176_U532
g18041 nand P2_R1176_U79 P2_R1176_U48 ; P2_R1176_U533
g18042 nand P2_R1176_U472 P2_U3193 ; P2_R1176_U534
g18043 nand P2_R1176_U80 P2_R1176_U45 ; P2_R1176_U535
g18044 nand P2_R1176_U535 P2_R1176_U534 ; P2_R1176_U536
g18045 nand P2_R1176_U350 P2_R1176_U52 ; P2_R1176_U537
g18046 nand P2_R1176_U536 P2_R1176_U322 ; P2_R1176_U538
g18047 nand P2_R1176_U381 P2_U3212 ; P2_R1176_U539
g18048 nand P2_R1176_U61 P2_R1176_U23 ; P2_R1176_U540
g18049 nand P2_R1176_U381 P2_U3212 ; P2_R1176_U541
g18050 nand P2_R1176_U61 P2_R1176_U23 ; P2_R1176_U542
g18051 nand P2_R1176_U542 P2_R1176_U541 ; P2_R1176_U543
g18052 nand P2_R1176_U180 P2_R1176_U181 ; P2_R1176_U544
g18053 nand P2_R1176_U205 P2_R1176_U543 ; P2_R1176_U545
g18054 nand P2_R1176_U475 P2_U3194 ; P2_R1176_U546
g18055 nand P2_R1176_U78 P2_R1176_U46 ; P2_R1176_U547
g18056 nand P2_R1176_U547 P2_R1176_U546 ; P2_R1176_U548
g18057 nand P2_R1176_U351 P2_R1176_U182 ; P2_R1176_U549
g18058 nand P2_R1176_U284 P2_R1176_U548 ; P2_R1176_U550
g18059 nand P2_R1176_U466 P2_U3195 ; P2_R1176_U551
g18060 nand P2_R1176_U77 P2_R1176_U44 ; P2_R1176_U552
g18061 nand P2_R1176_U466 P2_U3195 ; P2_R1176_U553
g18062 nand P2_R1176_U77 P2_R1176_U44 ; P2_R1176_U554
g18063 nand P2_R1176_U554 P2_R1176_U553 ; P2_R1176_U555
g18064 nand P2_R1176_U183 P2_R1176_U184 ; P2_R1176_U556
g18065 nand P2_R1176_U280 P2_R1176_U555 ; P2_R1176_U557
g18066 nand P2_R1176_U460 P2_U3196 ; P2_R1176_U558
g18067 nand P2_R1176_U70 P2_R1176_U36 ; P2_R1176_U559
g18068 nand P2_R1176_U463 P2_U3197 ; P2_R1176_U560
g18069 nand P2_R1176_U69 P2_R1176_U34 ; P2_R1176_U561
g18070 nand P2_R1176_U561 P2_R1176_U560 ; P2_R1176_U562
g18071 nand P2_R1176_U352 P2_R1176_U53 ; P2_R1176_U563
g18072 nand P2_R1176_U562 P2_R1176_U272 ; P2_R1176_U564
g18073 nand P2_R1176_U457 P2_U3198 ; P2_R1176_U565
g18074 nand P2_R1176_U76 P2_R1176_U43 ; P2_R1176_U566
g18075 nand P2_R1176_U457 P2_U3198 ; P2_R1176_U567
g18076 nand P2_R1176_U76 P2_R1176_U43 ; P2_R1176_U568
g18077 nand P2_R1176_U568 P2_R1176_U567 ; P2_R1176_U569
g18078 nand P2_R1176_U185 P2_R1176_U186 ; P2_R1176_U570
g18079 nand P2_R1176_U268 P2_R1176_U569 ; P2_R1176_U571
g18080 nand P2_R1176_U454 P2_U3199 ; P2_R1176_U572
g18081 nand P2_R1176_U75 P2_R1176_U42 ; P2_R1176_U573
g18082 nand P2_R1176_U454 P2_U3199 ; P2_R1176_U574
g18083 nand P2_R1176_U75 P2_R1176_U42 ; P2_R1176_U575
g18084 nand P2_R1176_U575 P2_R1176_U574 ; P2_R1176_U576
g18085 nand P2_R1176_U187 P2_R1176_U188 ; P2_R1176_U577
g18086 nand P2_R1176_U264 P2_R1176_U576 ; P2_R1176_U578
g18087 nand P2_R1176_U445 P2_U3200 ; P2_R1176_U579
g18088 nand P2_R1176_U73 P2_R1176_U41 ; P2_R1176_U580
g18089 nand P2_R1176_U448 P2_U3201 ; P2_R1176_U581
g18090 nand P2_R1176_U74 P2_R1176_U38 ; P2_R1176_U582
g18091 nand P2_R1176_U582 P2_R1176_U581 ; P2_R1176_U583
g18092 nand P2_R1176_U353 P2_R1176_U54 ; P2_R1176_U584
g18093 nand P2_R1176_U583 P2_R1176_U338 ; P2_R1176_U585
g18094 nand P2_R1176_U451 P2_U3202 ; P2_R1176_U586
g18095 nand P2_R1176_U72 P2_R1176_U39 ; P2_R1176_U587
g18096 nand P2_R1176_U587 P2_R1176_U586 ; P2_R1176_U588
g18097 nand P2_R1176_U354 P2_R1176_U189 ; P2_R1176_U589
g18098 nand P2_R1176_U254 P2_R1176_U588 ; P2_R1176_U590
g18099 nand P2_R1176_U442 P2_U3203 ; P2_R1176_U591
g18100 nand P2_R1176_U71 P2_R1176_U37 ; P2_R1176_U592
g18101 nand P2_R1176_U442 P2_U3203 ; P2_R1176_U593
g18102 nand P2_R1176_U71 P2_R1176_U37 ; P2_R1176_U594
g18103 nand P2_R1176_U594 P2_R1176_U593 ; P2_R1176_U595
g18104 nand P2_R1176_U190 P2_R1176_U191 ; P2_R1176_U596
g18105 nand P2_R1176_U250 P2_R1176_U595 ; P2_R1176_U597
g18106 nand P2_U3213 P2_R1176_U15 ; P2_R1176_U598
g18107 nand P2_U3214 P2_R1176_U22 ; P2_R1176_U599
g18108 not P2_R1176_U133 ; P2_R1176_U600
g18109 nand P2_R1176_U60 P2_R1176_U600 ; P2_R1176_U601
g18110 nand P2_R1176_U133 P2_R1176_U378 ; P2_R1176_U602
g18111 and P2_R1131_U179 P2_R1131_U178 ; P2_R1131_U4
g18112 and P2_R1131_U197 P2_R1131_U196 ; P2_R1131_U5
g18113 and P2_R1131_U237 P2_R1131_U236 ; P2_R1131_U6
g18114 and P2_R1131_U246 P2_R1131_U245 ; P2_R1131_U7
g18115 and P2_R1131_U264 P2_R1131_U263 ; P2_R1131_U8
g18116 and P2_R1131_U272 P2_R1131_U271 ; P2_R1131_U9
g18117 and P2_R1131_U351 P2_R1131_U348 ; P2_R1131_U10
g18118 and P2_R1131_U344 P2_R1131_U341 ; P2_R1131_U11
g18119 and P2_R1131_U335 P2_R1131_U332 ; P2_R1131_U12
g18120 and P2_R1131_U326 P2_R1131_U323 ; P2_R1131_U13
g18121 and P2_R1131_U320 P2_R1131_U318 ; P2_R1131_U14
g18122 and P2_R1131_U313 P2_R1131_U310 ; P2_R1131_U15
g18123 and P2_R1131_U235 P2_R1131_U232 ; P2_R1131_U16
g18124 and P2_R1131_U227 P2_R1131_U224 ; P2_R1131_U17
g18125 and P2_R1131_U213 P2_R1131_U210 ; P2_R1131_U18
g18126 not P2_U3468 ; P2_R1131_U19
g18127 not P2_U3071 ; P2_R1131_U20
g18128 not P2_U3070 ; P2_R1131_U21
g18129 nand P2_U3071 P2_U3468 ; P2_R1131_U22
g18130 not P2_U3471 ; P2_R1131_U23
g18131 not P2_U3462 ; P2_R1131_U24
g18132 not P2_U3060 ; P2_R1131_U25
g18133 not P2_U3067 ; P2_R1131_U26
g18134 not P2_U3456 ; P2_R1131_U27
g18135 not P2_U3068 ; P2_R1131_U28
g18136 not P2_U3448 ; P2_R1131_U29
g18137 not P2_U3077 ; P2_R1131_U30
g18138 nand P2_U3077 P2_U3448 ; P2_R1131_U31
g18139 not P2_U3459 ; P2_R1131_U32
g18140 not P2_U3064 ; P2_R1131_U33
g18141 nand P2_U3060 P2_U3462 ; P2_R1131_U34
g18142 not P2_U3465 ; P2_R1131_U35
g18143 not P2_U3474 ; P2_R1131_U36
g18144 not P2_U3084 ; P2_R1131_U37
g18145 not P2_U3083 ; P2_R1131_U38
g18146 not P2_U3477 ; P2_R1131_U39
g18147 nand P2_R1131_U61 P2_R1131_U205 ; P2_R1131_U40
g18148 nand P2_R1131_U117 P2_R1131_U193 ; P2_R1131_U41
g18149 nand P2_R1131_U182 P2_R1131_U183 ; P2_R1131_U42
g18150 nand P2_U3453 P2_U3078 ; P2_R1131_U43
g18151 nand P2_R1131_U122 P2_R1131_U219 ; P2_R1131_U44
g18152 nand P2_R1131_U216 P2_R1131_U215 ; P2_R1131_U45
g18153 not P2_U3969 ; P2_R1131_U46
g18154 not P2_U3053 ; P2_R1131_U47
g18155 not P2_U3057 ; P2_R1131_U48
g18156 not P2_U3970 ; P2_R1131_U49
g18157 not P2_U3971 ; P2_R1131_U50
g18158 not P2_U3058 ; P2_R1131_U51
g18159 not P2_U3972 ; P2_R1131_U52
g18160 not P2_U3065 ; P2_R1131_U53
g18161 not P2_U3975 ; P2_R1131_U54
g18162 not P2_U3075 ; P2_R1131_U55
g18163 not P2_U3498 ; P2_R1131_U56
g18164 not P2_U3073 ; P2_R1131_U57
g18165 not P2_U3069 ; P2_R1131_U58
g18166 nand P2_U3073 P2_U3498 ; P2_R1131_U59
g18167 not P2_U3501 ; P2_R1131_U60
g18168 nand P2_U3084 P2_U3474 ; P2_R1131_U61
g18169 not P2_U3480 ; P2_R1131_U62
g18170 not P2_U3062 ; P2_R1131_U63
g18171 not P2_U3486 ; P2_R1131_U64
g18172 not P2_U3072 ; P2_R1131_U65
g18173 not P2_U3483 ; P2_R1131_U66
g18174 not P2_U3063 ; P2_R1131_U67
g18175 nand P2_U3063 P2_U3483 ; P2_R1131_U68
g18176 not P2_U3489 ; P2_R1131_U69
g18177 not P2_U3080 ; P2_R1131_U70
g18178 not P2_U3492 ; P2_R1131_U71
g18179 not P2_U3079 ; P2_R1131_U72
g18180 not P2_U3495 ; P2_R1131_U73
g18181 not P2_U3074 ; P2_R1131_U74
g18182 not P2_U3504 ; P2_R1131_U75
g18183 not P2_U3082 ; P2_R1131_U76
g18184 nand P2_U3082 P2_U3504 ; P2_R1131_U77
g18185 not P2_U3506 ; P2_R1131_U78
g18186 not P2_U3081 ; P2_R1131_U79
g18187 nand P2_U3081 P2_U3506 ; P2_R1131_U80
g18188 not P2_U3976 ; P2_R1131_U81
g18189 not P2_U3974 ; P2_R1131_U82
g18190 not P2_U3061 ; P2_R1131_U83
g18191 not P2_U3973 ; P2_R1131_U84
g18192 not P2_U3066 ; P2_R1131_U85
g18193 nand P2_U3970 P2_U3057 ; P2_R1131_U86
g18194 not P2_U3054 ; P2_R1131_U87
g18195 not P2_U3968 ; P2_R1131_U88
g18196 nand P2_R1131_U306 P2_R1131_U176 ; P2_R1131_U89
g18197 not P2_U3076 ; P2_R1131_U90
g18198 nand P2_R1131_U77 P2_R1131_U315 ; P2_R1131_U91
g18199 nand P2_R1131_U261 P2_R1131_U260 ; P2_R1131_U92
g18200 nand P2_R1131_U68 P2_R1131_U337 ; P2_R1131_U93
g18201 nand P2_R1131_U457 P2_R1131_U456 ; P2_R1131_U94
g18202 nand P2_R1131_U504 P2_R1131_U503 ; P2_R1131_U95
g18203 nand P2_R1131_U375 P2_R1131_U374 ; P2_R1131_U96
g18204 nand P2_R1131_U380 P2_R1131_U379 ; P2_R1131_U97
g18205 nand P2_R1131_U387 P2_R1131_U386 ; P2_R1131_U98
g18206 nand P2_R1131_U394 P2_R1131_U393 ; P2_R1131_U99
g18207 nand P2_R1131_U399 P2_R1131_U398 ; P2_R1131_U100
g18208 nand P2_R1131_U408 P2_R1131_U407 ; P2_R1131_U101
g18209 nand P2_R1131_U415 P2_R1131_U414 ; P2_R1131_U102
g18210 nand P2_R1131_U422 P2_R1131_U421 ; P2_R1131_U103
g18211 nand P2_R1131_U429 P2_R1131_U428 ; P2_R1131_U104
g18212 nand P2_R1131_U434 P2_R1131_U433 ; P2_R1131_U105
g18213 nand P2_R1131_U441 P2_R1131_U440 ; P2_R1131_U106
g18214 nand P2_R1131_U448 P2_R1131_U447 ; P2_R1131_U107
g18215 nand P2_R1131_U462 P2_R1131_U461 ; P2_R1131_U108
g18216 nand P2_R1131_U467 P2_R1131_U466 ; P2_R1131_U109
g18217 nand P2_R1131_U474 P2_R1131_U473 ; P2_R1131_U110
g18218 nand P2_R1131_U481 P2_R1131_U480 ; P2_R1131_U111
g18219 nand P2_R1131_U488 P2_R1131_U487 ; P2_R1131_U112
g18220 nand P2_R1131_U495 P2_R1131_U494 ; P2_R1131_U113
g18221 nand P2_R1131_U500 P2_R1131_U499 ; P2_R1131_U114
g18222 and P2_R1131_U189 P2_R1131_U187 ; P2_R1131_U115
g18223 and P2_R1131_U4 P2_R1131_U180 ; P2_R1131_U116
g18224 and P2_R1131_U194 P2_R1131_U192 ; P2_R1131_U117
g18225 and P2_R1131_U201 P2_R1131_U200 ; P2_R1131_U118
g18226 and P2_R1131_U382 P2_R1131_U381 P2_R1131_U22 ; P2_R1131_U119
g18227 and P2_R1131_U212 P2_R1131_U5 ; P2_R1131_U120
g18228 and P2_R1131_U181 P2_R1131_U180 ; P2_R1131_U121
g18229 and P2_R1131_U220 P2_R1131_U218 ; P2_R1131_U122
g18230 and P2_R1131_U389 P2_R1131_U388 P2_R1131_U34 ; P2_R1131_U123
g18231 and P2_R1131_U226 P2_R1131_U4 ; P2_R1131_U124
g18232 and P2_R1131_U234 P2_R1131_U181 ; P2_R1131_U125
g18233 and P2_R1131_U204 P2_R1131_U6 ; P2_R1131_U126
g18234 and P2_R1131_U239 P2_R1131_U171 ; P2_R1131_U127
g18235 and P2_R1131_U250 P2_R1131_U7 ; P2_R1131_U128
g18236 and P2_R1131_U248 P2_R1131_U172 ; P2_R1131_U129
g18237 and P2_R1131_U268 P2_R1131_U267 ; P2_R1131_U130
g18238 and P2_R1131_U9 P2_R1131_U282 P2_R1131_U273 ; P2_R1131_U131
g18239 and P2_R1131_U285 P2_R1131_U280 ; P2_R1131_U132
g18240 and P2_R1131_U301 P2_R1131_U298 ; P2_R1131_U133
g18241 and P2_R1131_U368 P2_R1131_U302 ; P2_R1131_U134
g18242 and P2_R1131_U424 P2_R1131_U423 P2_R1131_U173 ; P2_R1131_U135
g18243 and P2_R1131_U160 P2_R1131_U278 ; P2_R1131_U136
g18244 and P2_R1131_U455 P2_R1131_U454 P2_R1131_U80 ; P2_R1131_U137
g18245 and P2_R1131_U325 P2_R1131_U9 ; P2_R1131_U138
g18246 and P2_R1131_U469 P2_R1131_U468 P2_R1131_U59 ; P2_R1131_U139
g18247 and P2_R1131_U334 P2_R1131_U8 ; P2_R1131_U140
g18248 and P2_R1131_U490 P2_R1131_U489 P2_R1131_U172 ; P2_R1131_U141
g18249 and P2_R1131_U343 P2_R1131_U7 ; P2_R1131_U142
g18250 and P2_R1131_U502 P2_R1131_U501 P2_R1131_U171 ; P2_R1131_U143
g18251 and P2_R1131_U350 P2_R1131_U6 ; P2_R1131_U144
g18252 nand P2_R1131_U118 P2_R1131_U202 ; P2_R1131_U145
g18253 nand P2_R1131_U217 P2_R1131_U229 ; P2_R1131_U146
g18254 not P2_U3055 ; P2_R1131_U147
g18255 not P2_U3979 ; P2_R1131_U148
g18256 and P2_R1131_U403 P2_R1131_U402 ; P2_R1131_U149
g18257 nand P2_R1131_U304 P2_R1131_U169 P2_R1131_U364 ; P2_R1131_U150
g18258 and P2_R1131_U410 P2_R1131_U409 ; P2_R1131_U151
g18259 nand P2_R1131_U370 P2_R1131_U369 P2_R1131_U134 ; P2_R1131_U152
g18260 and P2_R1131_U417 P2_R1131_U416 ; P2_R1131_U153
g18261 nand P2_R1131_U365 P2_R1131_U299 P2_R1131_U86 ; P2_R1131_U154
g18262 nand P2_R1131_U293 P2_R1131_U292 ; P2_R1131_U155
g18263 and P2_R1131_U436 P2_R1131_U435 ; P2_R1131_U156
g18264 nand P2_R1131_U289 P2_R1131_U288 ; P2_R1131_U157
g18265 and P2_R1131_U443 P2_R1131_U442 ; P2_R1131_U158
g18266 nand P2_R1131_U132 P2_R1131_U284 ; P2_R1131_U159
g18267 and P2_R1131_U450 P2_R1131_U449 ; P2_R1131_U160
g18268 nand P2_R1131_U43 P2_R1131_U327 ; P2_R1131_U161
g18269 nand P2_R1131_U130 P2_R1131_U269 ; P2_R1131_U162
g18270 and P2_R1131_U476 P2_R1131_U475 ; P2_R1131_U163
g18271 nand P2_R1131_U257 P2_R1131_U256 ; P2_R1131_U164
g18272 and P2_R1131_U483 P2_R1131_U482 ; P2_R1131_U165
g18273 nand P2_R1131_U253 P2_R1131_U252 ; P2_R1131_U166
g18274 nand P2_R1131_U243 P2_R1131_U242 ; P2_R1131_U167
g18275 nand P2_R1131_U367 P2_R1131_U366 ; P2_R1131_U168
g18276 nand P2_U3054 P2_R1131_U152 ; P2_R1131_U169
g18277 not P2_R1131_U34 ; P2_R1131_U170
g18278 nand P2_U3477 P2_U3083 ; P2_R1131_U171
g18279 nand P2_U3072 P2_U3486 ; P2_R1131_U172
g18280 nand P2_U3058 P2_U3971 ; P2_R1131_U173
g18281 not P2_R1131_U68 ; P2_R1131_U174
g18282 not P2_R1131_U77 ; P2_R1131_U175
g18283 nand P2_U3065 P2_U3972 ; P2_R1131_U176
g18284 not P2_R1131_U61 ; P2_R1131_U177
g18285 or P2_U3067 P2_U3465 ; P2_R1131_U178
g18286 or P2_U3060 P2_U3462 ; P2_R1131_U179
g18287 or P2_U3459 P2_U3064 ; P2_R1131_U180
g18288 or P2_U3456 P2_U3068 ; P2_R1131_U181
g18289 not P2_R1131_U31 ; P2_R1131_U182
g18290 or P2_U3453 P2_U3078 ; P2_R1131_U183
g18291 not P2_R1131_U42 ; P2_R1131_U184
g18292 not P2_R1131_U43 ; P2_R1131_U185
g18293 nand P2_R1131_U42 P2_R1131_U43 ; P2_R1131_U186
g18294 nand P2_U3068 P2_U3456 ; P2_R1131_U187
g18295 nand P2_R1131_U186 P2_R1131_U181 ; P2_R1131_U188
g18296 nand P2_U3064 P2_U3459 ; P2_R1131_U189
g18297 nand P2_R1131_U115 P2_R1131_U188 ; P2_R1131_U190
g18298 nand P2_R1131_U35 P2_R1131_U34 ; P2_R1131_U191
g18299 nand P2_U3067 P2_R1131_U191 ; P2_R1131_U192
g18300 nand P2_R1131_U116 P2_R1131_U190 ; P2_R1131_U193
g18301 nand P2_U3465 P2_R1131_U170 ; P2_R1131_U194
g18302 not P2_R1131_U41 ; P2_R1131_U195
g18303 or P2_U3070 P2_U3471 ; P2_R1131_U196
g18304 or P2_U3071 P2_U3468 ; P2_R1131_U197
g18305 not P2_R1131_U22 ; P2_R1131_U198
g18306 nand P2_R1131_U23 P2_R1131_U22 ; P2_R1131_U199
g18307 nand P2_U3070 P2_R1131_U199 ; P2_R1131_U200
g18308 nand P2_U3471 P2_R1131_U198 ; P2_R1131_U201
g18309 nand P2_R1131_U5 P2_R1131_U41 ; P2_R1131_U202
g18310 not P2_R1131_U145 ; P2_R1131_U203
g18311 or P2_U3474 P2_U3084 ; P2_R1131_U204
g18312 nand P2_R1131_U204 P2_R1131_U145 ; P2_R1131_U205
g18313 not P2_R1131_U40 ; P2_R1131_U206
g18314 or P2_U3083 P2_U3477 ; P2_R1131_U207
g18315 or P2_U3468 P2_U3071 ; P2_R1131_U208
g18316 nand P2_R1131_U208 P2_R1131_U41 ; P2_R1131_U209
g18317 nand P2_R1131_U119 P2_R1131_U209 ; P2_R1131_U210
g18318 nand P2_R1131_U195 P2_R1131_U22 ; P2_R1131_U211
g18319 nand P2_U3471 P2_U3070 ; P2_R1131_U212
g18320 nand P2_R1131_U120 P2_R1131_U211 ; P2_R1131_U213
g18321 or P2_U3071 P2_U3468 ; P2_R1131_U214
g18322 nand P2_R1131_U185 P2_R1131_U181 ; P2_R1131_U215
g18323 nand P2_U3068 P2_U3456 ; P2_R1131_U216
g18324 not P2_R1131_U45 ; P2_R1131_U217
g18325 nand P2_R1131_U121 P2_R1131_U184 ; P2_R1131_U218
g18326 nand P2_R1131_U45 P2_R1131_U180 ; P2_R1131_U219
g18327 nand P2_U3064 P2_U3459 ; P2_R1131_U220
g18328 not P2_R1131_U44 ; P2_R1131_U221
g18329 or P2_U3462 P2_U3060 ; P2_R1131_U222
g18330 nand P2_R1131_U222 P2_R1131_U44 ; P2_R1131_U223
g18331 nand P2_R1131_U123 P2_R1131_U223 ; P2_R1131_U224
g18332 nand P2_R1131_U221 P2_R1131_U34 ; P2_R1131_U225
g18333 nand P2_U3465 P2_U3067 ; P2_R1131_U226
g18334 nand P2_R1131_U124 P2_R1131_U225 ; P2_R1131_U227
g18335 or P2_U3060 P2_U3462 ; P2_R1131_U228
g18336 nand P2_R1131_U184 P2_R1131_U181 ; P2_R1131_U229
g18337 not P2_R1131_U146 ; P2_R1131_U230
g18338 nand P2_U3064 P2_U3459 ; P2_R1131_U231
g18339 nand P2_R1131_U401 P2_R1131_U400 P2_R1131_U43 P2_R1131_U42 ; P2_R1131_U232
g18340 nand P2_R1131_U43 P2_R1131_U42 ; P2_R1131_U233
g18341 nand P2_U3068 P2_U3456 ; P2_R1131_U234
g18342 nand P2_R1131_U125 P2_R1131_U233 ; P2_R1131_U235
g18343 or P2_U3083 P2_U3477 ; P2_R1131_U236
g18344 or P2_U3062 P2_U3480 ; P2_R1131_U237
g18345 nand P2_R1131_U177 P2_R1131_U6 ; P2_R1131_U238
g18346 nand P2_U3062 P2_U3480 ; P2_R1131_U239
g18347 nand P2_R1131_U127 P2_R1131_U238 ; P2_R1131_U240
g18348 or P2_U3480 P2_U3062 ; P2_R1131_U241
g18349 nand P2_R1131_U126 P2_R1131_U145 ; P2_R1131_U242
g18350 nand P2_R1131_U241 P2_R1131_U240 ; P2_R1131_U243
g18351 not P2_R1131_U167 ; P2_R1131_U244
g18352 or P2_U3080 P2_U3489 ; P2_R1131_U245
g18353 or P2_U3072 P2_U3486 ; P2_R1131_U246
g18354 nand P2_R1131_U174 P2_R1131_U7 ; P2_R1131_U247
g18355 nand P2_U3080 P2_U3489 ; P2_R1131_U248
g18356 nand P2_R1131_U129 P2_R1131_U247 ; P2_R1131_U249
g18357 or P2_U3483 P2_U3063 ; P2_R1131_U250
g18358 or P2_U3489 P2_U3080 ; P2_R1131_U251
g18359 nand P2_R1131_U128 P2_R1131_U167 ; P2_R1131_U252
g18360 nand P2_R1131_U251 P2_R1131_U249 ; P2_R1131_U253
g18361 not P2_R1131_U166 ; P2_R1131_U254
g18362 or P2_U3492 P2_U3079 ; P2_R1131_U255
g18363 nand P2_R1131_U255 P2_R1131_U166 ; P2_R1131_U256
g18364 nand P2_U3079 P2_U3492 ; P2_R1131_U257
g18365 not P2_R1131_U164 ; P2_R1131_U258
g18366 or P2_U3495 P2_U3074 ; P2_R1131_U259
g18367 nand P2_R1131_U259 P2_R1131_U164 ; P2_R1131_U260
g18368 nand P2_U3074 P2_U3495 ; P2_R1131_U261
g18369 not P2_R1131_U92 ; P2_R1131_U262
g18370 or P2_U3069 P2_U3501 ; P2_R1131_U263
g18371 or P2_U3073 P2_U3498 ; P2_R1131_U264
g18372 not P2_R1131_U59 ; P2_R1131_U265
g18373 nand P2_R1131_U60 P2_R1131_U59 ; P2_R1131_U266
g18374 nand P2_U3069 P2_R1131_U266 ; P2_R1131_U267
g18375 nand P2_U3501 P2_R1131_U265 ; P2_R1131_U268
g18376 nand P2_R1131_U8 P2_R1131_U92 ; P2_R1131_U269
g18377 not P2_R1131_U162 ; P2_R1131_U270
g18378 or P2_U3076 P2_U3976 ; P2_R1131_U271
g18379 or P2_U3081 P2_U3506 ; P2_R1131_U272
g18380 or P2_U3075 P2_U3975 ; P2_R1131_U273
g18381 not P2_R1131_U80 ; P2_R1131_U274
g18382 nand P2_U3976 P2_R1131_U274 ; P2_R1131_U275
g18383 nand P2_R1131_U275 P2_R1131_U90 ; P2_R1131_U276
g18384 nand P2_R1131_U80 P2_R1131_U81 ; P2_R1131_U277
g18385 nand P2_R1131_U277 P2_R1131_U276 ; P2_R1131_U278
g18386 nand P2_R1131_U175 P2_R1131_U9 ; P2_R1131_U279
g18387 nand P2_U3075 P2_U3975 ; P2_R1131_U280
g18388 nand P2_R1131_U278 P2_R1131_U279 ; P2_R1131_U281
g18389 or P2_U3504 P2_U3082 ; P2_R1131_U282
g18390 or P2_U3975 P2_U3075 ; P2_R1131_U283
g18391 nand P2_R1131_U162 P2_R1131_U131 ; P2_R1131_U284
g18392 nand P2_R1131_U283 P2_R1131_U281 ; P2_R1131_U285
g18393 not P2_R1131_U159 ; P2_R1131_U286
g18394 or P2_U3974 P2_U3061 ; P2_R1131_U287
g18395 nand P2_R1131_U287 P2_R1131_U159 ; P2_R1131_U288
g18396 nand P2_U3061 P2_U3974 ; P2_R1131_U289
g18397 not P2_R1131_U157 ; P2_R1131_U290
g18398 or P2_U3973 P2_U3066 ; P2_R1131_U291
g18399 nand P2_R1131_U291 P2_R1131_U157 ; P2_R1131_U292
g18400 nand P2_U3066 P2_U3973 ; P2_R1131_U293
g18401 not P2_R1131_U155 ; P2_R1131_U294
g18402 or P2_U3058 P2_U3971 ; P2_R1131_U295
g18403 nand P2_R1131_U176 P2_R1131_U173 ; P2_R1131_U296
g18404 not P2_R1131_U86 ; P2_R1131_U297
g18405 or P2_U3972 P2_U3065 ; P2_R1131_U298
g18406 nand P2_R1131_U155 P2_R1131_U298 P2_R1131_U168 ; P2_R1131_U299
g18407 not P2_R1131_U154 ; P2_R1131_U300
g18408 or P2_U3969 P2_U3053 ; P2_R1131_U301
g18409 nand P2_U3053 P2_U3969 ; P2_R1131_U302
g18410 not P2_R1131_U152 ; P2_R1131_U303
g18411 nand P2_U3968 P2_R1131_U152 ; P2_R1131_U304
g18412 not P2_R1131_U150 ; P2_R1131_U305
g18413 nand P2_R1131_U298 P2_R1131_U155 ; P2_R1131_U306
g18414 not P2_R1131_U89 ; P2_R1131_U307
g18415 or P2_U3971 P2_U3058 ; P2_R1131_U308
g18416 nand P2_R1131_U308 P2_R1131_U89 ; P2_R1131_U309
g18417 nand P2_R1131_U135 P2_R1131_U309 ; P2_R1131_U310
g18418 nand P2_R1131_U307 P2_R1131_U173 ; P2_R1131_U311
g18419 nand P2_U3970 P2_U3057 ; P2_R1131_U312
g18420 nand P2_R1131_U311 P2_R1131_U312 P2_R1131_U168 ; P2_R1131_U313
g18421 or P2_U3058 P2_U3971 ; P2_R1131_U314
g18422 nand P2_R1131_U282 P2_R1131_U162 ; P2_R1131_U315
g18423 not P2_R1131_U91 ; P2_R1131_U316
g18424 nand P2_R1131_U9 P2_R1131_U91 ; P2_R1131_U317
g18425 nand P2_R1131_U136 P2_R1131_U317 ; P2_R1131_U318
g18426 nand P2_R1131_U317 P2_R1131_U278 ; P2_R1131_U319
g18427 nand P2_R1131_U453 P2_R1131_U319 ; P2_R1131_U320
g18428 or P2_U3506 P2_U3081 ; P2_R1131_U321
g18429 nand P2_R1131_U321 P2_R1131_U91 ; P2_R1131_U322
g18430 nand P2_R1131_U137 P2_R1131_U322 ; P2_R1131_U323
g18431 nand P2_R1131_U316 P2_R1131_U80 ; P2_R1131_U324
g18432 nand P2_U3076 P2_U3976 ; P2_R1131_U325
g18433 nand P2_R1131_U138 P2_R1131_U324 ; P2_R1131_U326
g18434 or P2_U3453 P2_U3078 ; P2_R1131_U327
g18435 not P2_R1131_U161 ; P2_R1131_U328
g18436 or P2_U3081 P2_U3506 ; P2_R1131_U329
g18437 or P2_U3498 P2_U3073 ; P2_R1131_U330
g18438 nand P2_R1131_U330 P2_R1131_U92 ; P2_R1131_U331
g18439 nand P2_R1131_U139 P2_R1131_U331 ; P2_R1131_U332
g18440 nand P2_R1131_U262 P2_R1131_U59 ; P2_R1131_U333
g18441 nand P2_U3501 P2_U3069 ; P2_R1131_U334
g18442 nand P2_R1131_U140 P2_R1131_U333 ; P2_R1131_U335
g18443 or P2_U3073 P2_U3498 ; P2_R1131_U336
g18444 nand P2_R1131_U250 P2_R1131_U167 ; P2_R1131_U337
g18445 not P2_R1131_U93 ; P2_R1131_U338
g18446 or P2_U3486 P2_U3072 ; P2_R1131_U339
g18447 nand P2_R1131_U339 P2_R1131_U93 ; P2_R1131_U340
g18448 nand P2_R1131_U141 P2_R1131_U340 ; P2_R1131_U341
g18449 nand P2_R1131_U338 P2_R1131_U172 ; P2_R1131_U342
g18450 nand P2_U3080 P2_U3489 ; P2_R1131_U343
g18451 nand P2_R1131_U142 P2_R1131_U342 ; P2_R1131_U344
g18452 or P2_U3072 P2_U3486 ; P2_R1131_U345
g18453 or P2_U3477 P2_U3083 ; P2_R1131_U346
g18454 nand P2_R1131_U346 P2_R1131_U40 ; P2_R1131_U347
g18455 nand P2_R1131_U143 P2_R1131_U347 ; P2_R1131_U348
g18456 nand P2_R1131_U206 P2_R1131_U171 ; P2_R1131_U349
g18457 nand P2_U3062 P2_U3480 ; P2_R1131_U350
g18458 nand P2_R1131_U144 P2_R1131_U349 ; P2_R1131_U351
g18459 nand P2_R1131_U207 P2_R1131_U171 ; P2_R1131_U352
g18460 nand P2_R1131_U204 P2_R1131_U61 ; P2_R1131_U353
g18461 nand P2_R1131_U214 P2_R1131_U22 ; P2_R1131_U354
g18462 nand P2_R1131_U228 P2_R1131_U34 ; P2_R1131_U355
g18463 nand P2_R1131_U231 P2_R1131_U180 ; P2_R1131_U356
g18464 nand P2_R1131_U314 P2_R1131_U173 ; P2_R1131_U357
g18465 nand P2_R1131_U298 P2_R1131_U176 ; P2_R1131_U358
g18466 nand P2_R1131_U329 P2_R1131_U80 ; P2_R1131_U359
g18467 nand P2_R1131_U282 P2_R1131_U77 ; P2_R1131_U360
g18468 nand P2_R1131_U336 P2_R1131_U59 ; P2_R1131_U361
g18469 nand P2_R1131_U345 P2_R1131_U172 ; P2_R1131_U362
g18470 nand P2_R1131_U250 P2_R1131_U68 ; P2_R1131_U363
g18471 nand P2_U3968 P2_U3054 ; P2_R1131_U364
g18472 nand P2_R1131_U296 P2_R1131_U168 ; P2_R1131_U365
g18473 nand P2_U3057 P2_R1131_U295 ; P2_R1131_U366
g18474 nand P2_U3970 P2_R1131_U295 ; P2_R1131_U367
g18475 nand P2_R1131_U296 P2_R1131_U168 P2_R1131_U301 ; P2_R1131_U368
g18476 nand P2_R1131_U155 P2_R1131_U168 P2_R1131_U133 ; P2_R1131_U369
g18477 nand P2_R1131_U297 P2_R1131_U301 ; P2_R1131_U370
g18478 nand P2_U3083 P2_R1131_U39 ; P2_R1131_U371
g18479 nand P2_U3477 P2_R1131_U38 ; P2_R1131_U372
g18480 nand P2_R1131_U372 P2_R1131_U371 ; P2_R1131_U373
g18481 nand P2_R1131_U352 P2_R1131_U40 ; P2_R1131_U374
g18482 nand P2_R1131_U373 P2_R1131_U206 ; P2_R1131_U375
g18483 nand P2_U3084 P2_R1131_U36 ; P2_R1131_U376
g18484 nand P2_U3474 P2_R1131_U37 ; P2_R1131_U377
g18485 nand P2_R1131_U377 P2_R1131_U376 ; P2_R1131_U378
g18486 nand P2_R1131_U353 P2_R1131_U145 ; P2_R1131_U379
g18487 nand P2_R1131_U203 P2_R1131_U378 ; P2_R1131_U380
g18488 nand P2_U3070 P2_R1131_U23 ; P2_R1131_U381
g18489 nand P2_U3471 P2_R1131_U21 ; P2_R1131_U382
g18490 nand P2_U3071 P2_R1131_U19 ; P2_R1131_U383
g18491 nand P2_U3468 P2_R1131_U20 ; P2_R1131_U384
g18492 nand P2_R1131_U384 P2_R1131_U383 ; P2_R1131_U385
g18493 nand P2_R1131_U354 P2_R1131_U41 ; P2_R1131_U386
g18494 nand P2_R1131_U385 P2_R1131_U195 ; P2_R1131_U387
g18495 nand P2_U3067 P2_R1131_U35 ; P2_R1131_U388
g18496 nand P2_U3465 P2_R1131_U26 ; P2_R1131_U389
g18497 nand P2_U3060 P2_R1131_U24 ; P2_R1131_U390
g18498 nand P2_U3462 P2_R1131_U25 ; P2_R1131_U391
g18499 nand P2_R1131_U391 P2_R1131_U390 ; P2_R1131_U392
g18500 nand P2_R1131_U355 P2_R1131_U44 ; P2_R1131_U393
g18501 nand P2_R1131_U392 P2_R1131_U221 ; P2_R1131_U394
g18502 nand P2_U3064 P2_R1131_U32 ; P2_R1131_U395
g18503 nand P2_U3459 P2_R1131_U33 ; P2_R1131_U396
g18504 nand P2_R1131_U396 P2_R1131_U395 ; P2_R1131_U397
g18505 nand P2_R1131_U356 P2_R1131_U146 ; P2_R1131_U398
g18506 nand P2_R1131_U230 P2_R1131_U397 ; P2_R1131_U399
g18507 nand P2_U3068 P2_R1131_U27 ; P2_R1131_U400
g18508 nand P2_U3456 P2_R1131_U28 ; P2_R1131_U401
g18509 nand P2_U3055 P2_R1131_U148 ; P2_R1131_U402
g18510 nand P2_U3979 P2_R1131_U147 ; P2_R1131_U403
g18511 nand P2_U3055 P2_R1131_U148 ; P2_R1131_U404
g18512 nand P2_U3979 P2_R1131_U147 ; P2_R1131_U405
g18513 nand P2_R1131_U405 P2_R1131_U404 ; P2_R1131_U406
g18514 nand P2_R1131_U149 P2_R1131_U150 ; P2_R1131_U407
g18515 nand P2_R1131_U305 P2_R1131_U406 ; P2_R1131_U408
g18516 nand P2_U3054 P2_R1131_U88 ; P2_R1131_U409
g18517 nand P2_U3968 P2_R1131_U87 ; P2_R1131_U410
g18518 nand P2_U3054 P2_R1131_U88 ; P2_R1131_U411
g18519 nand P2_U3968 P2_R1131_U87 ; P2_R1131_U412
g18520 nand P2_R1131_U412 P2_R1131_U411 ; P2_R1131_U413
g18521 nand P2_R1131_U151 P2_R1131_U152 ; P2_R1131_U414
g18522 nand P2_R1131_U303 P2_R1131_U413 ; P2_R1131_U415
g18523 nand P2_U3053 P2_R1131_U46 ; P2_R1131_U416
g18524 nand P2_U3969 P2_R1131_U47 ; P2_R1131_U417
g18525 nand P2_U3053 P2_R1131_U46 ; P2_R1131_U418
g18526 nand P2_U3969 P2_R1131_U47 ; P2_R1131_U419
g18527 nand P2_R1131_U419 P2_R1131_U418 ; P2_R1131_U420
g18528 nand P2_R1131_U153 P2_R1131_U154 ; P2_R1131_U421
g18529 nand P2_R1131_U300 P2_R1131_U420 ; P2_R1131_U422
g18530 nand P2_U3057 P2_R1131_U49 ; P2_R1131_U423
g18531 nand P2_U3970 P2_R1131_U48 ; P2_R1131_U424
g18532 nand P2_U3058 P2_R1131_U50 ; P2_R1131_U425
g18533 nand P2_U3971 P2_R1131_U51 ; P2_R1131_U426
g18534 nand P2_R1131_U426 P2_R1131_U425 ; P2_R1131_U427
g18535 nand P2_R1131_U357 P2_R1131_U89 ; P2_R1131_U428
g18536 nand P2_R1131_U427 P2_R1131_U307 ; P2_R1131_U429
g18537 nand P2_U3065 P2_R1131_U52 ; P2_R1131_U430
g18538 nand P2_U3972 P2_R1131_U53 ; P2_R1131_U431
g18539 nand P2_R1131_U431 P2_R1131_U430 ; P2_R1131_U432
g18540 nand P2_R1131_U358 P2_R1131_U155 ; P2_R1131_U433
g18541 nand P2_R1131_U294 P2_R1131_U432 ; P2_R1131_U434
g18542 nand P2_U3066 P2_R1131_U84 ; P2_R1131_U435
g18543 nand P2_U3973 P2_R1131_U85 ; P2_R1131_U436
g18544 nand P2_U3066 P2_R1131_U84 ; P2_R1131_U437
g18545 nand P2_U3973 P2_R1131_U85 ; P2_R1131_U438
g18546 nand P2_R1131_U438 P2_R1131_U437 ; P2_R1131_U439
g18547 nand P2_R1131_U156 P2_R1131_U157 ; P2_R1131_U440
g18548 nand P2_R1131_U290 P2_R1131_U439 ; P2_R1131_U441
g18549 nand P2_U3061 P2_R1131_U82 ; P2_R1131_U442
g18550 nand P2_U3974 P2_R1131_U83 ; P2_R1131_U443
g18551 nand P2_U3061 P2_R1131_U82 ; P2_R1131_U444
g18552 nand P2_U3974 P2_R1131_U83 ; P2_R1131_U445
g18553 nand P2_R1131_U445 P2_R1131_U444 ; P2_R1131_U446
g18554 nand P2_R1131_U158 P2_R1131_U159 ; P2_R1131_U447
g18555 nand P2_R1131_U286 P2_R1131_U446 ; P2_R1131_U448
g18556 nand P2_U3075 P2_R1131_U54 ; P2_R1131_U449
g18557 nand P2_U3975 P2_R1131_U55 ; P2_R1131_U450
g18558 nand P2_U3075 P2_R1131_U54 ; P2_R1131_U451
g18559 nand P2_U3975 P2_R1131_U55 ; P2_R1131_U452
g18560 nand P2_R1131_U452 P2_R1131_U451 ; P2_R1131_U453
g18561 nand P2_U3076 P2_R1131_U81 ; P2_R1131_U454
g18562 nand P2_U3976 P2_R1131_U90 ; P2_R1131_U455
g18563 nand P2_R1131_U182 P2_R1131_U161 ; P2_R1131_U456
g18564 nand P2_R1131_U328 P2_R1131_U31 ; P2_R1131_U457
g18565 nand P2_U3081 P2_R1131_U78 ; P2_R1131_U458
g18566 nand P2_U3506 P2_R1131_U79 ; P2_R1131_U459
g18567 nand P2_R1131_U459 P2_R1131_U458 ; P2_R1131_U460
g18568 nand P2_R1131_U359 P2_R1131_U91 ; P2_R1131_U461
g18569 nand P2_R1131_U460 P2_R1131_U316 ; P2_R1131_U462
g18570 nand P2_U3082 P2_R1131_U75 ; P2_R1131_U463
g18571 nand P2_U3504 P2_R1131_U76 ; P2_R1131_U464
g18572 nand P2_R1131_U464 P2_R1131_U463 ; P2_R1131_U465
g18573 nand P2_R1131_U360 P2_R1131_U162 ; P2_R1131_U466
g18574 nand P2_R1131_U270 P2_R1131_U465 ; P2_R1131_U467
g18575 nand P2_U3069 P2_R1131_U60 ; P2_R1131_U468
g18576 nand P2_U3501 P2_R1131_U58 ; P2_R1131_U469
g18577 nand P2_U3073 P2_R1131_U56 ; P2_R1131_U470
g18578 nand P2_U3498 P2_R1131_U57 ; P2_R1131_U471
g18579 nand P2_R1131_U471 P2_R1131_U470 ; P2_R1131_U472
g18580 nand P2_R1131_U361 P2_R1131_U92 ; P2_R1131_U473
g18581 nand P2_R1131_U472 P2_R1131_U262 ; P2_R1131_U474
g18582 nand P2_U3074 P2_R1131_U73 ; P2_R1131_U475
g18583 nand P2_U3495 P2_R1131_U74 ; P2_R1131_U476
g18584 nand P2_U3074 P2_R1131_U73 ; P2_R1131_U477
g18585 nand P2_U3495 P2_R1131_U74 ; P2_R1131_U478
g18586 nand P2_R1131_U478 P2_R1131_U477 ; P2_R1131_U479
g18587 nand P2_R1131_U163 P2_R1131_U164 ; P2_R1131_U480
g18588 nand P2_R1131_U258 P2_R1131_U479 ; P2_R1131_U481
g18589 nand P2_U3079 P2_R1131_U71 ; P2_R1131_U482
g18590 nand P2_U3492 P2_R1131_U72 ; P2_R1131_U483
g18591 nand P2_U3079 P2_R1131_U71 ; P2_R1131_U484
g18592 nand P2_U3492 P2_R1131_U72 ; P2_R1131_U485
g18593 nand P2_R1131_U485 P2_R1131_U484 ; P2_R1131_U486
g18594 nand P2_R1131_U165 P2_R1131_U166 ; P2_R1131_U487
g18595 nand P2_R1131_U254 P2_R1131_U486 ; P2_R1131_U488
g18596 nand P2_U3080 P2_R1131_U69 ; P2_R1131_U489
g18597 nand P2_U3489 P2_R1131_U70 ; P2_R1131_U490
g18598 nand P2_U3072 P2_R1131_U64 ; P2_R1131_U491
g18599 nand P2_U3486 P2_R1131_U65 ; P2_R1131_U492
g18600 nand P2_R1131_U492 P2_R1131_U491 ; P2_R1131_U493
g18601 nand P2_R1131_U362 P2_R1131_U93 ; P2_R1131_U494
g18602 nand P2_R1131_U493 P2_R1131_U338 ; P2_R1131_U495
g18603 nand P2_U3063 P2_R1131_U66 ; P2_R1131_U496
g18604 nand P2_U3483 P2_R1131_U67 ; P2_R1131_U497
g18605 nand P2_R1131_U497 P2_R1131_U496 ; P2_R1131_U498
g18606 nand P2_R1131_U363 P2_R1131_U167 ; P2_R1131_U499
g18607 nand P2_R1131_U244 P2_R1131_U498 ; P2_R1131_U500
g18608 nand P2_U3062 P2_R1131_U62 ; P2_R1131_U501
g18609 nand P2_U3480 P2_R1131_U63 ; P2_R1131_U502
g18610 nand P2_U3077 P2_R1131_U29 ; P2_R1131_U503
g18611 nand P2_U3448 P2_R1131_U30 ; P2_R1131_U504
g18612 and P2_R1146_U205 P2_R1146_U204 ; P2_R1146_U6
g18613 and P2_R1146_U244 P2_R1146_U243 ; P2_R1146_U7
g18614 and P2_R1146_U261 P2_R1146_U260 ; P2_R1146_U8
g18615 and P2_R1146_U285 P2_R1146_U284 ; P2_R1146_U9
g18616 and P2_R1146_U384 P2_R1146_U383 ; P2_R1146_U10
g18617 nand P2_R1146_U340 P2_R1146_U343 ; P2_R1146_U11
g18618 nand P2_R1146_U329 P2_R1146_U332 ; P2_R1146_U12
g18619 nand P2_R1146_U318 P2_R1146_U321 ; P2_R1146_U13
g18620 nand P2_R1146_U310 P2_R1146_U312 ; P2_R1146_U14
g18621 nand P2_R1146_U349 P2_R1146_U177 P2_R1146_U156 ; P2_R1146_U15
g18622 nand P2_R1146_U238 P2_R1146_U240 ; P2_R1146_U16
g18623 nand P2_R1146_U230 P2_R1146_U233 ; P2_R1146_U17
g18624 nand P2_R1146_U222 P2_R1146_U224 ; P2_R1146_U18
g18625 nand P2_R1146_U166 P2_R1146_U346 ; P2_R1146_U19
g18626 not P2_U3471 ; P2_R1146_U20
g18627 not P2_U3465 ; P2_R1146_U21
g18628 not P2_U3456 ; P2_R1146_U22
g18629 not P2_U3448 ; P2_R1146_U23
g18630 not P2_U3078 ; P2_R1146_U24
g18631 not P2_U3459 ; P2_R1146_U25
g18632 not P2_U3068 ; P2_R1146_U26
g18633 nand P2_U3068 P2_R1146_U22 ; P2_R1146_U27
g18634 not P2_U3064 ; P2_R1146_U28
g18635 not P2_U3468 ; P2_R1146_U29
g18636 not P2_U3462 ; P2_R1146_U30
g18637 not P2_U3071 ; P2_R1146_U31
g18638 not P2_U3067 ; P2_R1146_U32
g18639 not P2_U3060 ; P2_R1146_U33
g18640 nand P2_U3060 P2_R1146_U30 ; P2_R1146_U34
g18641 not P2_U3474 ; P2_R1146_U35
g18642 not P2_U3070 ; P2_R1146_U36
g18643 nand P2_U3070 P2_R1146_U20 ; P2_R1146_U37
g18644 not P2_U3084 ; P2_R1146_U38
g18645 not P2_U3477 ; P2_R1146_U39
g18646 not P2_U3083 ; P2_R1146_U40
g18647 nand P2_R1146_U211 P2_R1146_U210 ; P2_R1146_U41
g18648 nand P2_R1146_U34 P2_R1146_U226 ; P2_R1146_U42
g18649 nand P2_R1146_U195 P2_R1146_U179 P2_R1146_U347 ; P2_R1146_U43
g18650 not P2_U3970 ; P2_R1146_U44
g18651 not P2_U3974 ; P2_R1146_U45
g18652 not P2_U3495 ; P2_R1146_U46
g18653 not P2_U3480 ; P2_R1146_U47
g18654 not P2_U3483 ; P2_R1146_U48
g18655 not P2_U3063 ; P2_R1146_U49
g18656 not P2_U3062 ; P2_R1146_U50
g18657 nand P2_U3083 P2_R1146_U39 ; P2_R1146_U51
g18658 not P2_U3486 ; P2_R1146_U52
g18659 not P2_U3072 ; P2_R1146_U53
g18660 not P2_U3489 ; P2_R1146_U54
g18661 not P2_U3080 ; P2_R1146_U55
g18662 not P2_U3498 ; P2_R1146_U56
g18663 not P2_U3492 ; P2_R1146_U57
g18664 not P2_U3073 ; P2_R1146_U58
g18665 not P2_U3074 ; P2_R1146_U59
g18666 not P2_U3079 ; P2_R1146_U60
g18667 nand P2_U3079 P2_R1146_U57 ; P2_R1146_U61
g18668 not P2_U3501 ; P2_R1146_U62
g18669 not P2_U3069 ; P2_R1146_U63
g18670 not P2_U3082 ; P2_R1146_U64
g18671 not P2_U3506 ; P2_R1146_U65
g18672 not P2_U3081 ; P2_R1146_U66
g18673 not P2_U3976 ; P2_R1146_U67
g18674 not P2_U3076 ; P2_R1146_U68
g18675 not P2_U3973 ; P2_R1146_U69
g18676 not P2_U3975 ; P2_R1146_U70
g18677 not P2_U3066 ; P2_R1146_U71
g18678 not P2_U3061 ; P2_R1146_U72
g18679 not P2_U3075 ; P2_R1146_U73
g18680 nand P2_U3075 P2_R1146_U70 ; P2_R1146_U74
g18681 not P2_U3972 ; P2_R1146_U75
g18682 not P2_U3065 ; P2_R1146_U76
g18683 not P2_U3971 ; P2_R1146_U77
g18684 not P2_U3058 ; P2_R1146_U78
g18685 not P2_U3969 ; P2_R1146_U79
g18686 not P2_U3057 ; P2_R1146_U80
g18687 nand P2_U3057 P2_R1146_U44 ; P2_R1146_U81
g18688 not P2_U3053 ; P2_R1146_U82
g18689 not P2_U3968 ; P2_R1146_U83
g18690 not P2_U3054 ; P2_R1146_U84
g18691 nand P2_R1146_U299 P2_R1146_U298 ; P2_R1146_U85
g18692 nand P2_R1146_U74 P2_R1146_U314 ; P2_R1146_U86
g18693 nand P2_R1146_U61 P2_R1146_U325 ; P2_R1146_U87
g18694 nand P2_R1146_U51 P2_R1146_U336 ; P2_R1146_U88
g18695 not P2_U3077 ; P2_R1146_U89
g18696 nand P2_R1146_U394 P2_R1146_U393 ; P2_R1146_U90
g18697 nand P2_R1146_U408 P2_R1146_U407 ; P2_R1146_U91
g18698 nand P2_R1146_U413 P2_R1146_U412 ; P2_R1146_U92
g18699 nand P2_R1146_U429 P2_R1146_U428 ; P2_R1146_U93
g18700 nand P2_R1146_U434 P2_R1146_U433 ; P2_R1146_U94
g18701 nand P2_R1146_U439 P2_R1146_U438 ; P2_R1146_U95
g18702 nand P2_R1146_U444 P2_R1146_U443 ; P2_R1146_U96
g18703 nand P2_R1146_U449 P2_R1146_U448 ; P2_R1146_U97
g18704 nand P2_R1146_U465 P2_R1146_U464 ; P2_R1146_U98
g18705 nand P2_R1146_U470 P2_R1146_U469 ; P2_R1146_U99
g18706 nand P2_R1146_U353 P2_R1146_U352 ; P2_R1146_U100
g18707 nand P2_R1146_U362 P2_R1146_U361 ; P2_R1146_U101
g18708 nand P2_R1146_U369 P2_R1146_U368 ; P2_R1146_U102
g18709 nand P2_R1146_U373 P2_R1146_U372 ; P2_R1146_U103
g18710 nand P2_R1146_U382 P2_R1146_U381 ; P2_R1146_U104
g18711 nand P2_R1146_U403 P2_R1146_U402 ; P2_R1146_U105
g18712 nand P2_R1146_U420 P2_R1146_U419 ; P2_R1146_U106
g18713 nand P2_R1146_U424 P2_R1146_U423 ; P2_R1146_U107
g18714 nand P2_R1146_U456 P2_R1146_U455 ; P2_R1146_U108
g18715 nand P2_R1146_U460 P2_R1146_U459 ; P2_R1146_U109
g18716 nand P2_R1146_U477 P2_R1146_U476 ; P2_R1146_U110
g18717 and P2_R1146_U197 P2_R1146_U187 ; P2_R1146_U111
g18718 and P2_R1146_U200 P2_R1146_U201 ; P2_R1146_U112
g18719 and P2_R1146_U208 P2_R1146_U203 P2_R1146_U188 ; P2_R1146_U113
g18720 and P2_R1146_U213 P2_R1146_U189 ; P2_R1146_U114
g18721 and P2_R1146_U216 P2_R1146_U217 ; P2_R1146_U115
g18722 and P2_R1146_U355 P2_R1146_U354 P2_R1146_U37 ; P2_R1146_U116
g18723 and P2_R1146_U358 P2_R1146_U189 ; P2_R1146_U117
g18724 and P2_R1146_U232 P2_R1146_U6 ; P2_R1146_U118
g18725 and P2_R1146_U365 P2_R1146_U188 ; P2_R1146_U119
g18726 and P2_R1146_U375 P2_R1146_U374 P2_R1146_U27 ; P2_R1146_U120
g18727 and P2_R1146_U378 P2_R1146_U187 ; P2_R1146_U121
g18728 and P2_R1146_U242 P2_R1146_U219 P2_R1146_U183 ; P2_R1146_U122
g18729 and P2_R1146_U264 P2_R1146_U184 P2_R1146_U259 ; P2_R1146_U123
g18730 and P2_R1146_U288 P2_R1146_U185 P2_R1146_U283 ; P2_R1146_U124
g18731 and P2_R1146_U301 P2_R1146_U186 ; P2_R1146_U125
g18732 and P2_R1146_U304 P2_R1146_U305 ; P2_R1146_U126
g18733 and P2_R1146_U304 P2_R1146_U305 ; P2_R1146_U127
g18734 and P2_R1146_U10 P2_R1146_U308 ; P2_R1146_U128
g18735 nand P2_R1146_U391 P2_R1146_U390 ; P2_R1146_U129
g18736 and P2_R1146_U396 P2_R1146_U395 P2_R1146_U81 ; P2_R1146_U130
g18737 and P2_R1146_U399 P2_R1146_U186 ; P2_R1146_U131
g18738 nand P2_R1146_U405 P2_R1146_U404 ; P2_R1146_U132
g18739 nand P2_R1146_U410 P2_R1146_U409 ; P2_R1146_U133
g18740 and P2_R1146_U320 P2_R1146_U9 ; P2_R1146_U134
g18741 and P2_R1146_U416 P2_R1146_U185 ; P2_R1146_U135
g18742 nand P2_R1146_U426 P2_R1146_U425 ; P2_R1146_U136
g18743 nand P2_R1146_U431 P2_R1146_U430 ; P2_R1146_U137
g18744 nand P2_R1146_U436 P2_R1146_U435 ; P2_R1146_U138
g18745 nand P2_R1146_U441 P2_R1146_U440 ; P2_R1146_U139
g18746 nand P2_R1146_U446 P2_R1146_U445 ; P2_R1146_U140
g18747 and P2_R1146_U331 P2_R1146_U8 ; P2_R1146_U141
g18748 and P2_R1146_U452 P2_R1146_U184 ; P2_R1146_U142
g18749 nand P2_R1146_U462 P2_R1146_U461 ; P2_R1146_U143
g18750 nand P2_R1146_U467 P2_R1146_U466 ; P2_R1146_U144
g18751 and P2_R1146_U342 P2_R1146_U7 ; P2_R1146_U145
g18752 and P2_R1146_U473 P2_R1146_U183 ; P2_R1146_U146
g18753 and P2_R1146_U351 P2_R1146_U350 ; P2_R1146_U147
g18754 nand P2_R1146_U115 P2_R1146_U214 ; P2_R1146_U148
g18755 and P2_R1146_U360 P2_R1146_U359 ; P2_R1146_U149
g18756 and P2_R1146_U367 P2_R1146_U366 ; P2_R1146_U150
g18757 and P2_R1146_U371 P2_R1146_U370 ; P2_R1146_U151
g18758 nand P2_R1146_U112 P2_R1146_U198 ; P2_R1146_U152
g18759 and P2_R1146_U380 P2_R1146_U379 ; P2_R1146_U153
g18760 not P2_U3979 ; P2_R1146_U154
g18761 not P2_U3055 ; P2_R1146_U155
g18762 and P2_R1146_U389 P2_R1146_U388 ; P2_R1146_U156
g18763 nand P2_R1146_U126 P2_R1146_U302 ; P2_R1146_U157
g18764 and P2_R1146_U401 P2_R1146_U400 ; P2_R1146_U158
g18765 nand P2_R1146_U295 P2_R1146_U294 ; P2_R1146_U159
g18766 nand P2_R1146_U291 P2_R1146_U290 ; P2_R1146_U160
g18767 and P2_R1146_U418 P2_R1146_U417 ; P2_R1146_U161
g18768 and P2_R1146_U422 P2_R1146_U421 ; P2_R1146_U162
g18769 nand P2_R1146_U281 P2_R1146_U280 ; P2_R1146_U163
g18770 nand P2_R1146_U277 P2_R1146_U276 ; P2_R1146_U164
g18771 not P2_U3453 ; P2_R1146_U165
g18772 nand P2_U3448 P2_R1146_U89 ; P2_R1146_U166
g18773 nand P2_R1146_U273 P2_R1146_U178 P2_R1146_U348 ; P2_R1146_U167
g18774 not P2_U3504 ; P2_R1146_U168
g18775 nand P2_R1146_U271 P2_R1146_U270 ; P2_R1146_U169
g18776 nand P2_R1146_U267 P2_R1146_U266 ; P2_R1146_U170
g18777 and P2_R1146_U454 P2_R1146_U453 ; P2_R1146_U171
g18778 and P2_R1146_U458 P2_R1146_U457 ; P2_R1146_U172
g18779 nand P2_R1146_U257 P2_R1146_U256 ; P2_R1146_U173
g18780 nand P2_R1146_U253 P2_R1146_U252 ; P2_R1146_U174
g18781 nand P2_R1146_U249 P2_R1146_U248 ; P2_R1146_U175
g18782 and P2_R1146_U475 P2_R1146_U474 ; P2_R1146_U176
g18783 nand P2_R1146_U307 P2_R1146_U157 P2_R1146_U387 ; P2_R1146_U177
g18784 nand P2_R1146_U169 P2_R1146_U168 ; P2_R1146_U178
g18785 nand P2_R1146_U166 P2_R1146_U165 ; P2_R1146_U179
g18786 not P2_R1146_U81 ; P2_R1146_U180
g18787 not P2_R1146_U27 ; P2_R1146_U181
g18788 not P2_R1146_U37 ; P2_R1146_U182
g18789 nand P2_U3480 P2_R1146_U50 ; P2_R1146_U183
g18790 nand P2_U3495 P2_R1146_U59 ; P2_R1146_U184
g18791 nand P2_U3974 P2_R1146_U72 ; P2_R1146_U185
g18792 nand P2_U3970 P2_R1146_U80 ; P2_R1146_U186
g18793 nand P2_U3456 P2_R1146_U26 ; P2_R1146_U187
g18794 nand P2_U3465 P2_R1146_U32 ; P2_R1146_U188
g18795 nand P2_U3471 P2_R1146_U36 ; P2_R1146_U189
g18796 not P2_R1146_U61 ; P2_R1146_U190
g18797 not P2_R1146_U74 ; P2_R1146_U191
g18798 not P2_R1146_U34 ; P2_R1146_U192
g18799 not P2_R1146_U51 ; P2_R1146_U193
g18800 not P2_R1146_U166 ; P2_R1146_U194
g18801 nand P2_U3078 P2_R1146_U166 ; P2_R1146_U195
g18802 not P2_R1146_U43 ; P2_R1146_U196
g18803 nand P2_U3459 P2_R1146_U28 ; P2_R1146_U197
g18804 nand P2_R1146_U111 P2_R1146_U43 ; P2_R1146_U198
g18805 nand P2_R1146_U28 P2_R1146_U27 ; P2_R1146_U199
g18806 nand P2_R1146_U199 P2_R1146_U25 ; P2_R1146_U200
g18807 nand P2_U3064 P2_R1146_U181 ; P2_R1146_U201
g18808 not P2_R1146_U152 ; P2_R1146_U202
g18809 nand P2_U3468 P2_R1146_U31 ; P2_R1146_U203
g18810 nand P2_U3071 P2_R1146_U29 ; P2_R1146_U204
g18811 nand P2_U3067 P2_R1146_U21 ; P2_R1146_U205
g18812 nand P2_R1146_U192 P2_R1146_U188 ; P2_R1146_U206
g18813 nand P2_R1146_U6 P2_R1146_U206 ; P2_R1146_U207
g18814 nand P2_U3462 P2_R1146_U33 ; P2_R1146_U208
g18815 nand P2_U3468 P2_R1146_U31 ; P2_R1146_U209
g18816 nand P2_R1146_U152 P2_R1146_U113 ; P2_R1146_U210
g18817 nand P2_R1146_U209 P2_R1146_U207 ; P2_R1146_U211
g18818 not P2_R1146_U41 ; P2_R1146_U212
g18819 nand P2_U3474 P2_R1146_U38 ; P2_R1146_U213
g18820 nand P2_R1146_U114 P2_R1146_U41 ; P2_R1146_U214
g18821 nand P2_R1146_U38 P2_R1146_U37 ; P2_R1146_U215
g18822 nand P2_R1146_U215 P2_R1146_U35 ; P2_R1146_U216
g18823 nand P2_U3084 P2_R1146_U182 ; P2_R1146_U217
g18824 not P2_R1146_U148 ; P2_R1146_U218
g18825 nand P2_U3477 P2_R1146_U40 ; P2_R1146_U219
g18826 nand P2_R1146_U219 P2_R1146_U51 ; P2_R1146_U220
g18827 nand P2_R1146_U212 P2_R1146_U37 ; P2_R1146_U221
g18828 nand P2_R1146_U117 P2_R1146_U221 ; P2_R1146_U222
g18829 nand P2_R1146_U41 P2_R1146_U189 ; P2_R1146_U223
g18830 nand P2_R1146_U116 P2_R1146_U223 ; P2_R1146_U224
g18831 nand P2_R1146_U37 P2_R1146_U189 ; P2_R1146_U225
g18832 nand P2_R1146_U208 P2_R1146_U152 ; P2_R1146_U226
g18833 not P2_R1146_U42 ; P2_R1146_U227
g18834 nand P2_U3067 P2_R1146_U21 ; P2_R1146_U228
g18835 nand P2_R1146_U227 P2_R1146_U228 ; P2_R1146_U229
g18836 nand P2_R1146_U119 P2_R1146_U229 ; P2_R1146_U230
g18837 nand P2_R1146_U42 P2_R1146_U188 ; P2_R1146_U231
g18838 nand P2_U3468 P2_R1146_U31 ; P2_R1146_U232
g18839 nand P2_R1146_U118 P2_R1146_U231 ; P2_R1146_U233
g18840 nand P2_U3067 P2_R1146_U21 ; P2_R1146_U234
g18841 nand P2_R1146_U188 P2_R1146_U234 ; P2_R1146_U235
g18842 nand P2_R1146_U208 P2_R1146_U34 ; P2_R1146_U236
g18843 nand P2_R1146_U196 P2_R1146_U27 ; P2_R1146_U237
g18844 nand P2_R1146_U121 P2_R1146_U237 ; P2_R1146_U238
g18845 nand P2_R1146_U43 P2_R1146_U187 ; P2_R1146_U239
g18846 nand P2_R1146_U120 P2_R1146_U239 ; P2_R1146_U240
g18847 nand P2_R1146_U27 P2_R1146_U187 ; P2_R1146_U241
g18848 nand P2_U3483 P2_R1146_U49 ; P2_R1146_U242
g18849 nand P2_U3063 P2_R1146_U48 ; P2_R1146_U243
g18850 nand P2_U3062 P2_R1146_U47 ; P2_R1146_U244
g18851 nand P2_R1146_U193 P2_R1146_U183 ; P2_R1146_U245
g18852 nand P2_R1146_U7 P2_R1146_U245 ; P2_R1146_U246
g18853 nand P2_U3483 P2_R1146_U49 ; P2_R1146_U247
g18854 nand P2_R1146_U148 P2_R1146_U122 ; P2_R1146_U248
g18855 nand P2_R1146_U247 P2_R1146_U246 ; P2_R1146_U249
g18856 not P2_R1146_U175 ; P2_R1146_U250
g18857 nand P2_U3486 P2_R1146_U53 ; P2_R1146_U251
g18858 nand P2_R1146_U251 P2_R1146_U175 ; P2_R1146_U252
g18859 nand P2_U3072 P2_R1146_U52 ; P2_R1146_U253
g18860 not P2_R1146_U174 ; P2_R1146_U254
g18861 nand P2_U3489 P2_R1146_U55 ; P2_R1146_U255
g18862 nand P2_R1146_U255 P2_R1146_U174 ; P2_R1146_U256
g18863 nand P2_U3080 P2_R1146_U54 ; P2_R1146_U257
g18864 not P2_R1146_U173 ; P2_R1146_U258
g18865 nand P2_U3498 P2_R1146_U58 ; P2_R1146_U259
g18866 nand P2_U3073 P2_R1146_U56 ; P2_R1146_U260
g18867 nand P2_U3074 P2_R1146_U46 ; P2_R1146_U261
g18868 nand P2_R1146_U190 P2_R1146_U184 ; P2_R1146_U262
g18869 nand P2_R1146_U8 P2_R1146_U262 ; P2_R1146_U263
g18870 nand P2_U3492 P2_R1146_U60 ; P2_R1146_U264
g18871 nand P2_U3498 P2_R1146_U58 ; P2_R1146_U265
g18872 nand P2_R1146_U173 P2_R1146_U123 ; P2_R1146_U266
g18873 nand P2_R1146_U265 P2_R1146_U263 ; P2_R1146_U267
g18874 not P2_R1146_U170 ; P2_R1146_U268
g18875 nand P2_U3501 P2_R1146_U63 ; P2_R1146_U269
g18876 nand P2_R1146_U269 P2_R1146_U170 ; P2_R1146_U270
g18877 nand P2_U3069 P2_R1146_U62 ; P2_R1146_U271
g18878 not P2_R1146_U169 ; P2_R1146_U272
g18879 nand P2_U3082 P2_R1146_U169 ; P2_R1146_U273
g18880 not P2_R1146_U167 ; P2_R1146_U274
g18881 nand P2_U3506 P2_R1146_U66 ; P2_R1146_U275
g18882 nand P2_R1146_U275 P2_R1146_U167 ; P2_R1146_U276
g18883 nand P2_U3081 P2_R1146_U65 ; P2_R1146_U277
g18884 not P2_R1146_U164 ; P2_R1146_U278
g18885 nand P2_U3976 P2_R1146_U68 ; P2_R1146_U279
g18886 nand P2_R1146_U279 P2_R1146_U164 ; P2_R1146_U280
g18887 nand P2_U3076 P2_R1146_U67 ; P2_R1146_U281
g18888 not P2_R1146_U163 ; P2_R1146_U282
g18889 nand P2_U3973 P2_R1146_U71 ; P2_R1146_U283
g18890 nand P2_U3066 P2_R1146_U69 ; P2_R1146_U284
g18891 nand P2_U3061 P2_R1146_U45 ; P2_R1146_U285
g18892 nand P2_R1146_U191 P2_R1146_U185 ; P2_R1146_U286
g18893 nand P2_R1146_U9 P2_R1146_U286 ; P2_R1146_U287
g18894 nand P2_U3975 P2_R1146_U73 ; P2_R1146_U288
g18895 nand P2_U3973 P2_R1146_U71 ; P2_R1146_U289
g18896 nand P2_R1146_U163 P2_R1146_U124 ; P2_R1146_U290
g18897 nand P2_R1146_U289 P2_R1146_U287 ; P2_R1146_U291
g18898 not P2_R1146_U160 ; P2_R1146_U292
g18899 nand P2_U3972 P2_R1146_U76 ; P2_R1146_U293
g18900 nand P2_R1146_U293 P2_R1146_U160 ; P2_R1146_U294
g18901 nand P2_U3065 P2_R1146_U75 ; P2_R1146_U295
g18902 not P2_R1146_U159 ; P2_R1146_U296
g18903 nand P2_U3971 P2_R1146_U78 ; P2_R1146_U297
g18904 nand P2_R1146_U297 P2_R1146_U159 ; P2_R1146_U298
g18905 nand P2_U3058 P2_R1146_U77 ; P2_R1146_U299
g18906 not P2_R1146_U85 ; P2_R1146_U300
g18907 nand P2_U3969 P2_R1146_U82 ; P2_R1146_U301
g18908 nand P2_R1146_U125 P2_R1146_U85 ; P2_R1146_U302
g18909 nand P2_R1146_U82 P2_R1146_U81 ; P2_R1146_U303
g18910 nand P2_R1146_U303 P2_R1146_U79 ; P2_R1146_U304
g18911 nand P2_U3053 P2_R1146_U180 ; P2_R1146_U305
g18912 not P2_R1146_U157 ; P2_R1146_U306
g18913 nand P2_U3968 P2_R1146_U84 ; P2_R1146_U307
g18914 nand P2_U3054 P2_R1146_U83 ; P2_R1146_U308
g18915 nand P2_R1146_U300 P2_R1146_U81 ; P2_R1146_U309
g18916 nand P2_R1146_U131 P2_R1146_U309 ; P2_R1146_U310
g18917 nand P2_R1146_U85 P2_R1146_U186 ; P2_R1146_U311
g18918 nand P2_R1146_U130 P2_R1146_U311 ; P2_R1146_U312
g18919 nand P2_R1146_U81 P2_R1146_U186 ; P2_R1146_U313
g18920 nand P2_R1146_U288 P2_R1146_U163 ; P2_R1146_U314
g18921 not P2_R1146_U86 ; P2_R1146_U315
g18922 nand P2_U3061 P2_R1146_U45 ; P2_R1146_U316
g18923 nand P2_R1146_U315 P2_R1146_U316 ; P2_R1146_U317
g18924 nand P2_R1146_U135 P2_R1146_U317 ; P2_R1146_U318
g18925 nand P2_R1146_U86 P2_R1146_U185 ; P2_R1146_U319
g18926 nand P2_U3973 P2_R1146_U71 ; P2_R1146_U320
g18927 nand P2_R1146_U134 P2_R1146_U319 ; P2_R1146_U321
g18928 nand P2_U3061 P2_R1146_U45 ; P2_R1146_U322
g18929 nand P2_R1146_U185 P2_R1146_U322 ; P2_R1146_U323
g18930 nand P2_R1146_U288 P2_R1146_U74 ; P2_R1146_U324
g18931 nand P2_R1146_U264 P2_R1146_U173 ; P2_R1146_U325
g18932 not P2_R1146_U87 ; P2_R1146_U326
g18933 nand P2_U3074 P2_R1146_U46 ; P2_R1146_U327
g18934 nand P2_R1146_U326 P2_R1146_U327 ; P2_R1146_U328
g18935 nand P2_R1146_U142 P2_R1146_U328 ; P2_R1146_U329
g18936 nand P2_R1146_U87 P2_R1146_U184 ; P2_R1146_U330
g18937 nand P2_U3498 P2_R1146_U58 ; P2_R1146_U331
g18938 nand P2_R1146_U141 P2_R1146_U330 ; P2_R1146_U332
g18939 nand P2_U3074 P2_R1146_U46 ; P2_R1146_U333
g18940 nand P2_R1146_U184 P2_R1146_U333 ; P2_R1146_U334
g18941 nand P2_R1146_U264 P2_R1146_U61 ; P2_R1146_U335
g18942 nand P2_R1146_U219 P2_R1146_U148 ; P2_R1146_U336
g18943 not P2_R1146_U88 ; P2_R1146_U337
g18944 nand P2_U3062 P2_R1146_U47 ; P2_R1146_U338
g18945 nand P2_R1146_U337 P2_R1146_U338 ; P2_R1146_U339
g18946 nand P2_R1146_U146 P2_R1146_U339 ; P2_R1146_U340
g18947 nand P2_R1146_U88 P2_R1146_U183 ; P2_R1146_U341
g18948 nand P2_U3483 P2_R1146_U49 ; P2_R1146_U342
g18949 nand P2_R1146_U145 P2_R1146_U341 ; P2_R1146_U343
g18950 nand P2_U3062 P2_R1146_U47 ; P2_R1146_U344
g18951 nand P2_R1146_U183 P2_R1146_U344 ; P2_R1146_U345
g18952 nand P2_U3077 P2_R1146_U23 ; P2_R1146_U346
g18953 nand P2_U3078 P2_R1146_U165 ; P2_R1146_U347
g18954 nand P2_U3082 P2_R1146_U168 ; P2_R1146_U348
g18955 nand P2_R1146_U127 P2_R1146_U302 P2_R1146_U128 ; P2_R1146_U349
g18956 nand P2_U3477 P2_R1146_U40 ; P2_R1146_U350
g18957 nand P2_U3083 P2_R1146_U39 ; P2_R1146_U351
g18958 nand P2_R1146_U220 P2_R1146_U148 ; P2_R1146_U352
g18959 nand P2_R1146_U218 P2_R1146_U147 ; P2_R1146_U353
g18960 nand P2_U3474 P2_R1146_U38 ; P2_R1146_U354
g18961 nand P2_U3084 P2_R1146_U35 ; P2_R1146_U355
g18962 nand P2_U3474 P2_R1146_U38 ; P2_R1146_U356
g18963 nand P2_U3084 P2_R1146_U35 ; P2_R1146_U357
g18964 nand P2_R1146_U357 P2_R1146_U356 ; P2_R1146_U358
g18965 nand P2_U3471 P2_R1146_U36 ; P2_R1146_U359
g18966 nand P2_U3070 P2_R1146_U20 ; P2_R1146_U360
g18967 nand P2_R1146_U225 P2_R1146_U41 ; P2_R1146_U361
g18968 nand P2_R1146_U149 P2_R1146_U212 ; P2_R1146_U362
g18969 nand P2_U3468 P2_R1146_U31 ; P2_R1146_U363
g18970 nand P2_U3071 P2_R1146_U29 ; P2_R1146_U364
g18971 nand P2_R1146_U364 P2_R1146_U363 ; P2_R1146_U365
g18972 nand P2_U3465 P2_R1146_U32 ; P2_R1146_U366
g18973 nand P2_U3067 P2_R1146_U21 ; P2_R1146_U367
g18974 nand P2_R1146_U235 P2_R1146_U42 ; P2_R1146_U368
g18975 nand P2_R1146_U150 P2_R1146_U227 ; P2_R1146_U369
g18976 nand P2_U3462 P2_R1146_U33 ; P2_R1146_U370
g18977 nand P2_U3060 P2_R1146_U30 ; P2_R1146_U371
g18978 nand P2_R1146_U236 P2_R1146_U152 ; P2_R1146_U372
g18979 nand P2_R1146_U202 P2_R1146_U151 ; P2_R1146_U373
g18980 nand P2_U3459 P2_R1146_U28 ; P2_R1146_U374
g18981 nand P2_U3064 P2_R1146_U25 ; P2_R1146_U375
g18982 nand P2_U3459 P2_R1146_U28 ; P2_R1146_U376
g18983 nand P2_U3064 P2_R1146_U25 ; P2_R1146_U377
g18984 nand P2_R1146_U377 P2_R1146_U376 ; P2_R1146_U378
g18985 nand P2_U3456 P2_R1146_U26 ; P2_R1146_U379
g18986 nand P2_U3068 P2_R1146_U22 ; P2_R1146_U380
g18987 nand P2_R1146_U241 P2_R1146_U43 ; P2_R1146_U381
g18988 nand P2_R1146_U153 P2_R1146_U196 ; P2_R1146_U382
g18989 nand P2_U3979 P2_R1146_U155 ; P2_R1146_U383
g18990 nand P2_U3055 P2_R1146_U154 ; P2_R1146_U384
g18991 nand P2_U3979 P2_R1146_U155 ; P2_R1146_U385
g18992 nand P2_U3055 P2_R1146_U154 ; P2_R1146_U386
g18993 nand P2_R1146_U386 P2_R1146_U385 ; P2_R1146_U387
g18994 nand P2_U3968 P2_R1146_U10 P2_R1146_U84 ; P2_R1146_U388
g18995 nand P2_R1146_U387 P2_R1146_U83 P2_U3054 ; P2_R1146_U389
g18996 nand P2_U3968 P2_R1146_U84 ; P2_R1146_U390
g18997 nand P2_U3054 P2_R1146_U83 ; P2_R1146_U391
g18998 not P2_R1146_U129 ; P2_R1146_U392
g18999 nand P2_R1146_U306 P2_R1146_U392 ; P2_R1146_U393
g19000 nand P2_R1146_U129 P2_R1146_U157 ; P2_R1146_U394
g19001 nand P2_U3969 P2_R1146_U82 ; P2_R1146_U395
g19002 nand P2_U3053 P2_R1146_U79 ; P2_R1146_U396
g19003 nand P2_U3969 P2_R1146_U82 ; P2_R1146_U397
g19004 nand P2_U3053 P2_R1146_U79 ; P2_R1146_U398
g19005 nand P2_R1146_U398 P2_R1146_U397 ; P2_R1146_U399
g19006 nand P2_U3970 P2_R1146_U80 ; P2_R1146_U400
g19007 nand P2_U3057 P2_R1146_U44 ; P2_R1146_U401
g19008 nand P2_R1146_U313 P2_R1146_U85 ; P2_R1146_U402
g19009 nand P2_R1146_U158 P2_R1146_U300 ; P2_R1146_U403
g19010 nand P2_U3971 P2_R1146_U78 ; P2_R1146_U404
g19011 nand P2_U3058 P2_R1146_U77 ; P2_R1146_U405
g19012 not P2_R1146_U132 ; P2_R1146_U406
g19013 nand P2_R1146_U296 P2_R1146_U406 ; P2_R1146_U407
g19014 nand P2_R1146_U132 P2_R1146_U159 ; P2_R1146_U408
g19015 nand P2_U3972 P2_R1146_U76 ; P2_R1146_U409
g19016 nand P2_U3065 P2_R1146_U75 ; P2_R1146_U410
g19017 not P2_R1146_U133 ; P2_R1146_U411
g19018 nand P2_R1146_U292 P2_R1146_U411 ; P2_R1146_U412
g19019 nand P2_R1146_U133 P2_R1146_U160 ; P2_R1146_U413
g19020 nand P2_U3973 P2_R1146_U71 ; P2_R1146_U414
g19021 nand P2_U3066 P2_R1146_U69 ; P2_R1146_U415
g19022 nand P2_R1146_U415 P2_R1146_U414 ; P2_R1146_U416
g19023 nand P2_U3974 P2_R1146_U72 ; P2_R1146_U417
g19024 nand P2_U3061 P2_R1146_U45 ; P2_R1146_U418
g19025 nand P2_R1146_U323 P2_R1146_U86 ; P2_R1146_U419
g19026 nand P2_R1146_U161 P2_R1146_U315 ; P2_R1146_U420
g19027 nand P2_U3975 P2_R1146_U73 ; P2_R1146_U421
g19028 nand P2_U3075 P2_R1146_U70 ; P2_R1146_U422
g19029 nand P2_R1146_U324 P2_R1146_U163 ; P2_R1146_U423
g19030 nand P2_R1146_U282 P2_R1146_U162 ; P2_R1146_U424
g19031 nand P2_U3976 P2_R1146_U68 ; P2_R1146_U425
g19032 nand P2_U3076 P2_R1146_U67 ; P2_R1146_U426
g19033 not P2_R1146_U136 ; P2_R1146_U427
g19034 nand P2_R1146_U278 P2_R1146_U427 ; P2_R1146_U428
g19035 nand P2_R1146_U136 P2_R1146_U164 ; P2_R1146_U429
g19036 nand P2_U3453 P2_R1146_U24 ; P2_R1146_U430
g19037 nand P2_U3078 P2_R1146_U165 ; P2_R1146_U431
g19038 not P2_R1146_U137 ; P2_R1146_U432
g19039 nand P2_R1146_U194 P2_R1146_U432 ; P2_R1146_U433
g19040 nand P2_R1146_U137 P2_R1146_U166 ; P2_R1146_U434
g19041 nand P2_U3506 P2_R1146_U66 ; P2_R1146_U435
g19042 nand P2_U3081 P2_R1146_U65 ; P2_R1146_U436
g19043 not P2_R1146_U138 ; P2_R1146_U437
g19044 nand P2_R1146_U274 P2_R1146_U437 ; P2_R1146_U438
g19045 nand P2_R1146_U138 P2_R1146_U167 ; P2_R1146_U439
g19046 nand P2_U3504 P2_R1146_U64 ; P2_R1146_U440
g19047 nand P2_U3082 P2_R1146_U168 ; P2_R1146_U441
g19048 not P2_R1146_U139 ; P2_R1146_U442
g19049 nand P2_R1146_U272 P2_R1146_U442 ; P2_R1146_U443
g19050 nand P2_R1146_U139 P2_R1146_U169 ; P2_R1146_U444
g19051 nand P2_U3501 P2_R1146_U63 ; P2_R1146_U445
g19052 nand P2_U3069 P2_R1146_U62 ; P2_R1146_U446
g19053 not P2_R1146_U140 ; P2_R1146_U447
g19054 nand P2_R1146_U268 P2_R1146_U447 ; P2_R1146_U448
g19055 nand P2_R1146_U140 P2_R1146_U170 ; P2_R1146_U449
g19056 nand P2_U3498 P2_R1146_U58 ; P2_R1146_U450
g19057 nand P2_U3073 P2_R1146_U56 ; P2_R1146_U451
g19058 nand P2_R1146_U451 P2_R1146_U450 ; P2_R1146_U452
g19059 nand P2_U3495 P2_R1146_U59 ; P2_R1146_U453
g19060 nand P2_U3074 P2_R1146_U46 ; P2_R1146_U454
g19061 nand P2_R1146_U334 P2_R1146_U87 ; P2_R1146_U455
g19062 nand P2_R1146_U171 P2_R1146_U326 ; P2_R1146_U456
g19063 nand P2_U3492 P2_R1146_U60 ; P2_R1146_U457
g19064 nand P2_U3079 P2_R1146_U57 ; P2_R1146_U458
g19065 nand P2_R1146_U335 P2_R1146_U173 ; P2_R1146_U459
g19066 nand P2_R1146_U258 P2_R1146_U172 ; P2_R1146_U460
g19067 nand P2_U3489 P2_R1146_U55 ; P2_R1146_U461
g19068 nand P2_U3080 P2_R1146_U54 ; P2_R1146_U462
g19069 not P2_R1146_U143 ; P2_R1146_U463
g19070 nand P2_R1146_U254 P2_R1146_U463 ; P2_R1146_U464
g19071 nand P2_R1146_U143 P2_R1146_U174 ; P2_R1146_U465
g19072 nand P2_U3486 P2_R1146_U53 ; P2_R1146_U466
g19073 nand P2_U3072 P2_R1146_U52 ; P2_R1146_U467
g19074 not P2_R1146_U144 ; P2_R1146_U468
g19075 nand P2_R1146_U250 P2_R1146_U468 ; P2_R1146_U469
g19076 nand P2_R1146_U144 P2_R1146_U175 ; P2_R1146_U470
g19077 nand P2_U3483 P2_R1146_U49 ; P2_R1146_U471
g19078 nand P2_U3063 P2_R1146_U48 ; P2_R1146_U472
g19079 nand P2_R1146_U472 P2_R1146_U471 ; P2_R1146_U473
g19080 nand P2_U3480 P2_R1146_U50 ; P2_R1146_U474
g19081 nand P2_U3062 P2_R1146_U47 ; P2_R1146_U475
g19082 nand P2_R1146_U345 P2_R1146_U88 ; P2_R1146_U476
g19083 nand P2_R1146_U176 P2_R1146_U337 ; P2_R1146_U477
g19084 and P2_R1203_U205 P2_R1203_U204 ; P2_R1203_U6
g19085 and P2_R1203_U244 P2_R1203_U243 ; P2_R1203_U7
g19086 and P2_R1203_U261 P2_R1203_U260 ; P2_R1203_U8
g19087 and P2_R1203_U285 P2_R1203_U284 ; P2_R1203_U9
g19088 and P2_R1203_U384 P2_R1203_U383 ; P2_R1203_U10
g19089 nand P2_R1203_U340 P2_R1203_U343 ; P2_R1203_U11
g19090 nand P2_R1203_U329 P2_R1203_U332 ; P2_R1203_U12
g19091 nand P2_R1203_U318 P2_R1203_U321 ; P2_R1203_U13
g19092 nand P2_R1203_U310 P2_R1203_U312 ; P2_R1203_U14
g19093 nand P2_R1203_U349 P2_R1203_U177 P2_R1203_U156 ; P2_R1203_U15
g19094 nand P2_R1203_U238 P2_R1203_U240 ; P2_R1203_U16
g19095 nand P2_R1203_U230 P2_R1203_U233 ; P2_R1203_U17
g19096 nand P2_R1203_U222 P2_R1203_U224 ; P2_R1203_U18
g19097 nand P2_R1203_U166 P2_R1203_U346 ; P2_R1203_U19
g19098 not P2_U3471 ; P2_R1203_U20
g19099 not P2_U3465 ; P2_R1203_U21
g19100 not P2_U3456 ; P2_R1203_U22
g19101 not P2_U3448 ; P2_R1203_U23
g19102 not P2_U3078 ; P2_R1203_U24
g19103 not P2_U3459 ; P2_R1203_U25
g19104 not P2_U3068 ; P2_R1203_U26
g19105 nand P2_U3068 P2_R1203_U22 ; P2_R1203_U27
g19106 not P2_U3064 ; P2_R1203_U28
g19107 not P2_U3468 ; P2_R1203_U29
g19108 not P2_U3462 ; P2_R1203_U30
g19109 not P2_U3071 ; P2_R1203_U31
g19110 not P2_U3067 ; P2_R1203_U32
g19111 not P2_U3060 ; P2_R1203_U33
g19112 nand P2_U3060 P2_R1203_U30 ; P2_R1203_U34
g19113 not P2_U3474 ; P2_R1203_U35
g19114 not P2_U3070 ; P2_R1203_U36
g19115 nand P2_U3070 P2_R1203_U20 ; P2_R1203_U37
g19116 not P2_U3084 ; P2_R1203_U38
g19117 not P2_U3477 ; P2_R1203_U39
g19118 not P2_U3083 ; P2_R1203_U40
g19119 nand P2_R1203_U211 P2_R1203_U210 ; P2_R1203_U41
g19120 nand P2_R1203_U34 P2_R1203_U226 ; P2_R1203_U42
g19121 nand P2_R1203_U195 P2_R1203_U179 P2_R1203_U347 ; P2_R1203_U43
g19122 not P2_U3970 ; P2_R1203_U44
g19123 not P2_U3974 ; P2_R1203_U45
g19124 not P2_U3495 ; P2_R1203_U46
g19125 not P2_U3480 ; P2_R1203_U47
g19126 not P2_U3483 ; P2_R1203_U48
g19127 not P2_U3063 ; P2_R1203_U49
g19128 not P2_U3062 ; P2_R1203_U50
g19129 nand P2_U3083 P2_R1203_U39 ; P2_R1203_U51
g19130 not P2_U3486 ; P2_R1203_U52
g19131 not P2_U3072 ; P2_R1203_U53
g19132 not P2_U3489 ; P2_R1203_U54
g19133 not P2_U3080 ; P2_R1203_U55
g19134 not P2_U3498 ; P2_R1203_U56
g19135 not P2_U3492 ; P2_R1203_U57
g19136 not P2_U3073 ; P2_R1203_U58
g19137 not P2_U3074 ; P2_R1203_U59
g19138 not P2_U3079 ; P2_R1203_U60
g19139 nand P2_U3079 P2_R1203_U57 ; P2_R1203_U61
g19140 not P2_U3501 ; P2_R1203_U62
g19141 not P2_U3069 ; P2_R1203_U63
g19142 not P2_U3082 ; P2_R1203_U64
g19143 not P2_U3506 ; P2_R1203_U65
g19144 not P2_U3081 ; P2_R1203_U66
g19145 not P2_U3976 ; P2_R1203_U67
g19146 not P2_U3076 ; P2_R1203_U68
g19147 not P2_U3973 ; P2_R1203_U69
g19148 not P2_U3975 ; P2_R1203_U70
g19149 not P2_U3066 ; P2_R1203_U71
g19150 not P2_U3061 ; P2_R1203_U72
g19151 not P2_U3075 ; P2_R1203_U73
g19152 nand P2_U3075 P2_R1203_U70 ; P2_R1203_U74
g19153 not P2_U3972 ; P2_R1203_U75
g19154 not P2_U3065 ; P2_R1203_U76
g19155 not P2_U3971 ; P2_R1203_U77
g19156 not P2_U3058 ; P2_R1203_U78
g19157 not P2_U3969 ; P2_R1203_U79
g19158 not P2_U3057 ; P2_R1203_U80
g19159 nand P2_U3057 P2_R1203_U44 ; P2_R1203_U81
g19160 not P2_U3053 ; P2_R1203_U82
g19161 not P2_U3968 ; P2_R1203_U83
g19162 not P2_U3054 ; P2_R1203_U84
g19163 nand P2_R1203_U299 P2_R1203_U298 ; P2_R1203_U85
g19164 nand P2_R1203_U74 P2_R1203_U314 ; P2_R1203_U86
g19165 nand P2_R1203_U61 P2_R1203_U325 ; P2_R1203_U87
g19166 nand P2_R1203_U51 P2_R1203_U336 ; P2_R1203_U88
g19167 not P2_U3077 ; P2_R1203_U89
g19168 nand P2_R1203_U394 P2_R1203_U393 ; P2_R1203_U90
g19169 nand P2_R1203_U408 P2_R1203_U407 ; P2_R1203_U91
g19170 nand P2_R1203_U413 P2_R1203_U412 ; P2_R1203_U92
g19171 nand P2_R1203_U429 P2_R1203_U428 ; P2_R1203_U93
g19172 nand P2_R1203_U434 P2_R1203_U433 ; P2_R1203_U94
g19173 nand P2_R1203_U439 P2_R1203_U438 ; P2_R1203_U95
g19174 nand P2_R1203_U444 P2_R1203_U443 ; P2_R1203_U96
g19175 nand P2_R1203_U449 P2_R1203_U448 ; P2_R1203_U97
g19176 nand P2_R1203_U465 P2_R1203_U464 ; P2_R1203_U98
g19177 nand P2_R1203_U470 P2_R1203_U469 ; P2_R1203_U99
g19178 nand P2_R1203_U353 P2_R1203_U352 ; P2_R1203_U100
g19179 nand P2_R1203_U362 P2_R1203_U361 ; P2_R1203_U101
g19180 nand P2_R1203_U369 P2_R1203_U368 ; P2_R1203_U102
g19181 nand P2_R1203_U373 P2_R1203_U372 ; P2_R1203_U103
g19182 nand P2_R1203_U382 P2_R1203_U381 ; P2_R1203_U104
g19183 nand P2_R1203_U403 P2_R1203_U402 ; P2_R1203_U105
g19184 nand P2_R1203_U420 P2_R1203_U419 ; P2_R1203_U106
g19185 nand P2_R1203_U424 P2_R1203_U423 ; P2_R1203_U107
g19186 nand P2_R1203_U456 P2_R1203_U455 ; P2_R1203_U108
g19187 nand P2_R1203_U460 P2_R1203_U459 ; P2_R1203_U109
g19188 nand P2_R1203_U477 P2_R1203_U476 ; P2_R1203_U110
g19189 and P2_R1203_U197 P2_R1203_U187 ; P2_R1203_U111
g19190 and P2_R1203_U200 P2_R1203_U201 ; P2_R1203_U112
g19191 and P2_R1203_U208 P2_R1203_U203 P2_R1203_U188 ; P2_R1203_U113
g19192 and P2_R1203_U213 P2_R1203_U189 ; P2_R1203_U114
g19193 and P2_R1203_U216 P2_R1203_U217 ; P2_R1203_U115
g19194 and P2_R1203_U355 P2_R1203_U354 P2_R1203_U37 ; P2_R1203_U116
g19195 and P2_R1203_U358 P2_R1203_U189 ; P2_R1203_U117
g19196 and P2_R1203_U232 P2_R1203_U6 ; P2_R1203_U118
g19197 and P2_R1203_U365 P2_R1203_U188 ; P2_R1203_U119
g19198 and P2_R1203_U375 P2_R1203_U374 P2_R1203_U27 ; P2_R1203_U120
g19199 and P2_R1203_U378 P2_R1203_U187 ; P2_R1203_U121
g19200 and P2_R1203_U242 P2_R1203_U219 P2_R1203_U183 ; P2_R1203_U122
g19201 and P2_R1203_U264 P2_R1203_U184 P2_R1203_U259 ; P2_R1203_U123
g19202 and P2_R1203_U288 P2_R1203_U185 P2_R1203_U283 ; P2_R1203_U124
g19203 and P2_R1203_U301 P2_R1203_U186 ; P2_R1203_U125
g19204 and P2_R1203_U304 P2_R1203_U305 ; P2_R1203_U126
g19205 and P2_R1203_U304 P2_R1203_U305 ; P2_R1203_U127
g19206 and P2_R1203_U10 P2_R1203_U308 ; P2_R1203_U128
g19207 nand P2_R1203_U391 P2_R1203_U390 ; P2_R1203_U129
g19208 and P2_R1203_U396 P2_R1203_U395 P2_R1203_U81 ; P2_R1203_U130
g19209 and P2_R1203_U399 P2_R1203_U186 ; P2_R1203_U131
g19210 nand P2_R1203_U405 P2_R1203_U404 ; P2_R1203_U132
g19211 nand P2_R1203_U410 P2_R1203_U409 ; P2_R1203_U133
g19212 and P2_R1203_U320 P2_R1203_U9 ; P2_R1203_U134
g19213 and P2_R1203_U416 P2_R1203_U185 ; P2_R1203_U135
g19214 nand P2_R1203_U426 P2_R1203_U425 ; P2_R1203_U136
g19215 nand P2_R1203_U431 P2_R1203_U430 ; P2_R1203_U137
g19216 nand P2_R1203_U436 P2_R1203_U435 ; P2_R1203_U138
g19217 nand P2_R1203_U441 P2_R1203_U440 ; P2_R1203_U139
g19218 nand P2_R1203_U446 P2_R1203_U445 ; P2_R1203_U140
g19219 and P2_R1203_U331 P2_R1203_U8 ; P2_R1203_U141
g19220 and P2_R1203_U452 P2_R1203_U184 ; P2_R1203_U142
g19221 nand P2_R1203_U462 P2_R1203_U461 ; P2_R1203_U143
g19222 nand P2_R1203_U467 P2_R1203_U466 ; P2_R1203_U144
g19223 and P2_R1203_U342 P2_R1203_U7 ; P2_R1203_U145
g19224 and P2_R1203_U473 P2_R1203_U183 ; P2_R1203_U146
g19225 and P2_R1203_U351 P2_R1203_U350 ; P2_R1203_U147
g19226 nand P2_R1203_U115 P2_R1203_U214 ; P2_R1203_U148
g19227 and P2_R1203_U360 P2_R1203_U359 ; P2_R1203_U149
g19228 and P2_R1203_U367 P2_R1203_U366 ; P2_R1203_U150
g19229 and P2_R1203_U371 P2_R1203_U370 ; P2_R1203_U151
g19230 nand P2_R1203_U112 P2_R1203_U198 ; P2_R1203_U152
g19231 and P2_R1203_U380 P2_R1203_U379 ; P2_R1203_U153
g19232 not P2_U3979 ; P2_R1203_U154
g19233 not P2_U3055 ; P2_R1203_U155
g19234 and P2_R1203_U389 P2_R1203_U388 ; P2_R1203_U156
g19235 nand P2_R1203_U126 P2_R1203_U302 ; P2_R1203_U157
g19236 and P2_R1203_U401 P2_R1203_U400 ; P2_R1203_U158
g19237 nand P2_R1203_U295 P2_R1203_U294 ; P2_R1203_U159
g19238 nand P2_R1203_U291 P2_R1203_U290 ; P2_R1203_U160
g19239 and P2_R1203_U418 P2_R1203_U417 ; P2_R1203_U161
g19240 and P2_R1203_U422 P2_R1203_U421 ; P2_R1203_U162
g19241 nand P2_R1203_U281 P2_R1203_U280 ; P2_R1203_U163
g19242 nand P2_R1203_U277 P2_R1203_U276 ; P2_R1203_U164
g19243 not P2_U3453 ; P2_R1203_U165
g19244 nand P2_U3448 P2_R1203_U89 ; P2_R1203_U166
g19245 nand P2_R1203_U273 P2_R1203_U178 P2_R1203_U348 ; P2_R1203_U167
g19246 not P2_U3504 ; P2_R1203_U168
g19247 nand P2_R1203_U271 P2_R1203_U270 ; P2_R1203_U169
g19248 nand P2_R1203_U267 P2_R1203_U266 ; P2_R1203_U170
g19249 and P2_R1203_U454 P2_R1203_U453 ; P2_R1203_U171
g19250 and P2_R1203_U458 P2_R1203_U457 ; P2_R1203_U172
g19251 nand P2_R1203_U257 P2_R1203_U256 ; P2_R1203_U173
g19252 nand P2_R1203_U253 P2_R1203_U252 ; P2_R1203_U174
g19253 nand P2_R1203_U249 P2_R1203_U248 ; P2_R1203_U175
g19254 and P2_R1203_U475 P2_R1203_U474 ; P2_R1203_U176
g19255 nand P2_R1203_U307 P2_R1203_U157 P2_R1203_U387 ; P2_R1203_U177
g19256 nand P2_R1203_U169 P2_R1203_U168 ; P2_R1203_U178
g19257 nand P2_R1203_U166 P2_R1203_U165 ; P2_R1203_U179
g19258 not P2_R1203_U81 ; P2_R1203_U180
g19259 not P2_R1203_U27 ; P2_R1203_U181
g19260 not P2_R1203_U37 ; P2_R1203_U182
g19261 nand P2_U3480 P2_R1203_U50 ; P2_R1203_U183
g19262 nand P2_U3495 P2_R1203_U59 ; P2_R1203_U184
g19263 nand P2_U3974 P2_R1203_U72 ; P2_R1203_U185
g19264 nand P2_U3970 P2_R1203_U80 ; P2_R1203_U186
g19265 nand P2_U3456 P2_R1203_U26 ; P2_R1203_U187
g19266 nand P2_U3465 P2_R1203_U32 ; P2_R1203_U188
g19267 nand P2_U3471 P2_R1203_U36 ; P2_R1203_U189
g19268 not P2_R1203_U61 ; P2_R1203_U190
g19269 not P2_R1203_U74 ; P2_R1203_U191
g19270 not P2_R1203_U34 ; P2_R1203_U192
g19271 not P2_R1203_U51 ; P2_R1203_U193
g19272 not P2_R1203_U166 ; P2_R1203_U194
g19273 nand P2_U3078 P2_R1203_U166 ; P2_R1203_U195
g19274 not P2_R1203_U43 ; P2_R1203_U196
g19275 nand P2_U3459 P2_R1203_U28 ; P2_R1203_U197
g19276 nand P2_R1203_U111 P2_R1203_U43 ; P2_R1203_U198
g19277 nand P2_R1203_U28 P2_R1203_U27 ; P2_R1203_U199
g19278 nand P2_R1203_U199 P2_R1203_U25 ; P2_R1203_U200
g19279 nand P2_U3064 P2_R1203_U181 ; P2_R1203_U201
g19280 not P2_R1203_U152 ; P2_R1203_U202
g19281 nand P2_U3468 P2_R1203_U31 ; P2_R1203_U203
g19282 nand P2_U3071 P2_R1203_U29 ; P2_R1203_U204
g19283 nand P2_U3067 P2_R1203_U21 ; P2_R1203_U205
g19284 nand P2_R1203_U192 P2_R1203_U188 ; P2_R1203_U206
g19285 nand P2_R1203_U6 P2_R1203_U206 ; P2_R1203_U207
g19286 nand P2_U3462 P2_R1203_U33 ; P2_R1203_U208
g19287 nand P2_U3468 P2_R1203_U31 ; P2_R1203_U209
g19288 nand P2_R1203_U152 P2_R1203_U113 ; P2_R1203_U210
g19289 nand P2_R1203_U209 P2_R1203_U207 ; P2_R1203_U211
g19290 not P2_R1203_U41 ; P2_R1203_U212
g19291 nand P2_U3474 P2_R1203_U38 ; P2_R1203_U213
g19292 nand P2_R1203_U114 P2_R1203_U41 ; P2_R1203_U214
g19293 nand P2_R1203_U38 P2_R1203_U37 ; P2_R1203_U215
g19294 nand P2_R1203_U215 P2_R1203_U35 ; P2_R1203_U216
g19295 nand P2_U3084 P2_R1203_U182 ; P2_R1203_U217
g19296 not P2_R1203_U148 ; P2_R1203_U218
g19297 nand P2_U3477 P2_R1203_U40 ; P2_R1203_U219
g19298 nand P2_R1203_U219 P2_R1203_U51 ; P2_R1203_U220
g19299 nand P2_R1203_U212 P2_R1203_U37 ; P2_R1203_U221
g19300 nand P2_R1203_U117 P2_R1203_U221 ; P2_R1203_U222
g19301 nand P2_R1203_U41 P2_R1203_U189 ; P2_R1203_U223
g19302 nand P2_R1203_U116 P2_R1203_U223 ; P2_R1203_U224
g19303 nand P2_R1203_U37 P2_R1203_U189 ; P2_R1203_U225
g19304 nand P2_R1203_U208 P2_R1203_U152 ; P2_R1203_U226
g19305 not P2_R1203_U42 ; P2_R1203_U227
g19306 nand P2_U3067 P2_R1203_U21 ; P2_R1203_U228
g19307 nand P2_R1203_U227 P2_R1203_U228 ; P2_R1203_U229
g19308 nand P2_R1203_U119 P2_R1203_U229 ; P2_R1203_U230
g19309 nand P2_R1203_U42 P2_R1203_U188 ; P2_R1203_U231
g19310 nand P2_U3468 P2_R1203_U31 ; P2_R1203_U232
g19311 nand P2_R1203_U118 P2_R1203_U231 ; P2_R1203_U233
g19312 nand P2_U3067 P2_R1203_U21 ; P2_R1203_U234
g19313 nand P2_R1203_U188 P2_R1203_U234 ; P2_R1203_U235
g19314 nand P2_R1203_U208 P2_R1203_U34 ; P2_R1203_U236
g19315 nand P2_R1203_U196 P2_R1203_U27 ; P2_R1203_U237
g19316 nand P2_R1203_U121 P2_R1203_U237 ; P2_R1203_U238
g19317 nand P2_R1203_U43 P2_R1203_U187 ; P2_R1203_U239
g19318 nand P2_R1203_U120 P2_R1203_U239 ; P2_R1203_U240
g19319 nand P2_R1203_U27 P2_R1203_U187 ; P2_R1203_U241
g19320 nand P2_U3483 P2_R1203_U49 ; P2_R1203_U242
g19321 nand P2_U3063 P2_R1203_U48 ; P2_R1203_U243
g19322 nand P2_U3062 P2_R1203_U47 ; P2_R1203_U244
g19323 nand P2_R1203_U193 P2_R1203_U183 ; P2_R1203_U245
g19324 nand P2_R1203_U7 P2_R1203_U245 ; P2_R1203_U246
g19325 nand P2_U3483 P2_R1203_U49 ; P2_R1203_U247
g19326 nand P2_R1203_U148 P2_R1203_U122 ; P2_R1203_U248
g19327 nand P2_R1203_U247 P2_R1203_U246 ; P2_R1203_U249
g19328 not P2_R1203_U175 ; P2_R1203_U250
g19329 nand P2_U3486 P2_R1203_U53 ; P2_R1203_U251
g19330 nand P2_R1203_U251 P2_R1203_U175 ; P2_R1203_U252
g19331 nand P2_U3072 P2_R1203_U52 ; P2_R1203_U253
g19332 not P2_R1203_U174 ; P2_R1203_U254
g19333 nand P2_U3489 P2_R1203_U55 ; P2_R1203_U255
g19334 nand P2_R1203_U255 P2_R1203_U174 ; P2_R1203_U256
g19335 nand P2_U3080 P2_R1203_U54 ; P2_R1203_U257
g19336 not P2_R1203_U173 ; P2_R1203_U258
g19337 nand P2_U3498 P2_R1203_U58 ; P2_R1203_U259
g19338 nand P2_U3073 P2_R1203_U56 ; P2_R1203_U260
g19339 nand P2_U3074 P2_R1203_U46 ; P2_R1203_U261
g19340 nand P2_R1203_U190 P2_R1203_U184 ; P2_R1203_U262
g19341 nand P2_R1203_U8 P2_R1203_U262 ; P2_R1203_U263
g19342 nand P2_U3492 P2_R1203_U60 ; P2_R1203_U264
g19343 nand P2_U3498 P2_R1203_U58 ; P2_R1203_U265
g19344 nand P2_R1203_U173 P2_R1203_U123 ; P2_R1203_U266
g19345 nand P2_R1203_U265 P2_R1203_U263 ; P2_R1203_U267
g19346 not P2_R1203_U170 ; P2_R1203_U268
g19347 nand P2_U3501 P2_R1203_U63 ; P2_R1203_U269
g19348 nand P2_R1203_U269 P2_R1203_U170 ; P2_R1203_U270
g19349 nand P2_U3069 P2_R1203_U62 ; P2_R1203_U271
g19350 not P2_R1203_U169 ; P2_R1203_U272
g19351 nand P2_U3082 P2_R1203_U169 ; P2_R1203_U273
g19352 not P2_R1203_U167 ; P2_R1203_U274
g19353 nand P2_U3506 P2_R1203_U66 ; P2_R1203_U275
g19354 nand P2_R1203_U275 P2_R1203_U167 ; P2_R1203_U276
g19355 nand P2_U3081 P2_R1203_U65 ; P2_R1203_U277
g19356 not P2_R1203_U164 ; P2_R1203_U278
g19357 nand P2_U3976 P2_R1203_U68 ; P2_R1203_U279
g19358 nand P2_R1203_U279 P2_R1203_U164 ; P2_R1203_U280
g19359 nand P2_U3076 P2_R1203_U67 ; P2_R1203_U281
g19360 not P2_R1203_U163 ; P2_R1203_U282
g19361 nand P2_U3973 P2_R1203_U71 ; P2_R1203_U283
g19362 nand P2_U3066 P2_R1203_U69 ; P2_R1203_U284
g19363 nand P2_U3061 P2_R1203_U45 ; P2_R1203_U285
g19364 nand P2_R1203_U191 P2_R1203_U185 ; P2_R1203_U286
g19365 nand P2_R1203_U9 P2_R1203_U286 ; P2_R1203_U287
g19366 nand P2_U3975 P2_R1203_U73 ; P2_R1203_U288
g19367 nand P2_U3973 P2_R1203_U71 ; P2_R1203_U289
g19368 nand P2_R1203_U163 P2_R1203_U124 ; P2_R1203_U290
g19369 nand P2_R1203_U289 P2_R1203_U287 ; P2_R1203_U291
g19370 not P2_R1203_U160 ; P2_R1203_U292
g19371 nand P2_U3972 P2_R1203_U76 ; P2_R1203_U293
g19372 nand P2_R1203_U293 P2_R1203_U160 ; P2_R1203_U294
g19373 nand P2_U3065 P2_R1203_U75 ; P2_R1203_U295
g19374 not P2_R1203_U159 ; P2_R1203_U296
g19375 nand P2_U3971 P2_R1203_U78 ; P2_R1203_U297
g19376 nand P2_R1203_U297 P2_R1203_U159 ; P2_R1203_U298
g19377 nand P2_U3058 P2_R1203_U77 ; P2_R1203_U299
g19378 not P2_R1203_U85 ; P2_R1203_U300
g19379 nand P2_U3969 P2_R1203_U82 ; P2_R1203_U301
g19380 nand P2_R1203_U125 P2_R1203_U85 ; P2_R1203_U302
g19381 nand P2_R1203_U82 P2_R1203_U81 ; P2_R1203_U303
g19382 nand P2_R1203_U303 P2_R1203_U79 ; P2_R1203_U304
g19383 nand P2_U3053 P2_R1203_U180 ; P2_R1203_U305
g19384 not P2_R1203_U157 ; P2_R1203_U306
g19385 nand P2_U3968 P2_R1203_U84 ; P2_R1203_U307
g19386 nand P2_U3054 P2_R1203_U83 ; P2_R1203_U308
g19387 nand P2_R1203_U300 P2_R1203_U81 ; P2_R1203_U309
g19388 nand P2_R1203_U131 P2_R1203_U309 ; P2_R1203_U310
g19389 nand P2_R1203_U85 P2_R1203_U186 ; P2_R1203_U311
g19390 nand P2_R1203_U130 P2_R1203_U311 ; P2_R1203_U312
g19391 nand P2_R1203_U81 P2_R1203_U186 ; P2_R1203_U313
g19392 nand P2_R1203_U288 P2_R1203_U163 ; P2_R1203_U314
g19393 not P2_R1203_U86 ; P2_R1203_U315
g19394 nand P2_U3061 P2_R1203_U45 ; P2_R1203_U316
g19395 nand P2_R1203_U315 P2_R1203_U316 ; P2_R1203_U317
g19396 nand P2_R1203_U135 P2_R1203_U317 ; P2_R1203_U318
g19397 nand P2_R1203_U86 P2_R1203_U185 ; P2_R1203_U319
g19398 nand P2_U3973 P2_R1203_U71 ; P2_R1203_U320
g19399 nand P2_R1203_U134 P2_R1203_U319 ; P2_R1203_U321
g19400 nand P2_U3061 P2_R1203_U45 ; P2_R1203_U322
g19401 nand P2_R1203_U185 P2_R1203_U322 ; P2_R1203_U323
g19402 nand P2_R1203_U288 P2_R1203_U74 ; P2_R1203_U324
g19403 nand P2_R1203_U264 P2_R1203_U173 ; P2_R1203_U325
g19404 not P2_R1203_U87 ; P2_R1203_U326
g19405 nand P2_U3074 P2_R1203_U46 ; P2_R1203_U327
g19406 nand P2_R1203_U326 P2_R1203_U327 ; P2_R1203_U328
g19407 nand P2_R1203_U142 P2_R1203_U328 ; P2_R1203_U329
g19408 nand P2_R1203_U87 P2_R1203_U184 ; P2_R1203_U330
g19409 nand P2_U3498 P2_R1203_U58 ; P2_R1203_U331
g19410 nand P2_R1203_U141 P2_R1203_U330 ; P2_R1203_U332
g19411 nand P2_U3074 P2_R1203_U46 ; P2_R1203_U333
g19412 nand P2_R1203_U184 P2_R1203_U333 ; P2_R1203_U334
g19413 nand P2_R1203_U264 P2_R1203_U61 ; P2_R1203_U335
g19414 nand P2_R1203_U219 P2_R1203_U148 ; P2_R1203_U336
g19415 not P2_R1203_U88 ; P2_R1203_U337
g19416 nand P2_U3062 P2_R1203_U47 ; P2_R1203_U338
g19417 nand P2_R1203_U337 P2_R1203_U338 ; P2_R1203_U339
g19418 nand P2_R1203_U146 P2_R1203_U339 ; P2_R1203_U340
g19419 nand P2_R1203_U88 P2_R1203_U183 ; P2_R1203_U341
g19420 nand P2_U3483 P2_R1203_U49 ; P2_R1203_U342
g19421 nand P2_R1203_U145 P2_R1203_U341 ; P2_R1203_U343
g19422 nand P2_U3062 P2_R1203_U47 ; P2_R1203_U344
g19423 nand P2_R1203_U183 P2_R1203_U344 ; P2_R1203_U345
g19424 nand P2_U3077 P2_R1203_U23 ; P2_R1203_U346
g19425 nand P2_U3078 P2_R1203_U165 ; P2_R1203_U347
g19426 nand P2_U3082 P2_R1203_U168 ; P2_R1203_U348
g19427 nand P2_R1203_U127 P2_R1203_U302 P2_R1203_U128 ; P2_R1203_U349
g19428 nand P2_U3477 P2_R1203_U40 ; P2_R1203_U350
g19429 nand P2_U3083 P2_R1203_U39 ; P2_R1203_U351
g19430 nand P2_R1203_U220 P2_R1203_U148 ; P2_R1203_U352
g19431 nand P2_R1203_U218 P2_R1203_U147 ; P2_R1203_U353
g19432 nand P2_U3474 P2_R1203_U38 ; P2_R1203_U354
g19433 nand P2_U3084 P2_R1203_U35 ; P2_R1203_U355
g19434 nand P2_U3474 P2_R1203_U38 ; P2_R1203_U356
g19435 nand P2_U3084 P2_R1203_U35 ; P2_R1203_U357
g19436 nand P2_R1203_U357 P2_R1203_U356 ; P2_R1203_U358
g19437 nand P2_U3471 P2_R1203_U36 ; P2_R1203_U359
g19438 nand P2_U3070 P2_R1203_U20 ; P2_R1203_U360
g19439 nand P2_R1203_U225 P2_R1203_U41 ; P2_R1203_U361
g19440 nand P2_R1203_U149 P2_R1203_U212 ; P2_R1203_U362
g19441 nand P2_U3468 P2_R1203_U31 ; P2_R1203_U363
g19442 nand P2_U3071 P2_R1203_U29 ; P2_R1203_U364
g19443 nand P2_R1203_U364 P2_R1203_U363 ; P2_R1203_U365
g19444 nand P2_U3465 P2_R1203_U32 ; P2_R1203_U366
g19445 nand P2_U3067 P2_R1203_U21 ; P2_R1203_U367
g19446 nand P2_R1203_U235 P2_R1203_U42 ; P2_R1203_U368
g19447 nand P2_R1203_U150 P2_R1203_U227 ; P2_R1203_U369
g19448 nand P2_U3462 P2_R1203_U33 ; P2_R1203_U370
g19449 nand P2_U3060 P2_R1203_U30 ; P2_R1203_U371
g19450 nand P2_R1203_U236 P2_R1203_U152 ; P2_R1203_U372
g19451 nand P2_R1203_U202 P2_R1203_U151 ; P2_R1203_U373
g19452 nand P2_U3459 P2_R1203_U28 ; P2_R1203_U374
g19453 nand P2_U3064 P2_R1203_U25 ; P2_R1203_U375
g19454 nand P2_U3459 P2_R1203_U28 ; P2_R1203_U376
g19455 nand P2_U3064 P2_R1203_U25 ; P2_R1203_U377
g19456 nand P2_R1203_U377 P2_R1203_U376 ; P2_R1203_U378
g19457 nand P2_U3456 P2_R1203_U26 ; P2_R1203_U379
g19458 nand P2_U3068 P2_R1203_U22 ; P2_R1203_U380
g19459 nand P2_R1203_U241 P2_R1203_U43 ; P2_R1203_U381
g19460 nand P2_R1203_U153 P2_R1203_U196 ; P2_R1203_U382
g19461 nand P2_U3979 P2_R1203_U155 ; P2_R1203_U383
g19462 nand P2_U3055 P2_R1203_U154 ; P2_R1203_U384
g19463 nand P2_U3979 P2_R1203_U155 ; P2_R1203_U385
g19464 nand P2_U3055 P2_R1203_U154 ; P2_R1203_U386
g19465 nand P2_R1203_U386 P2_R1203_U385 ; P2_R1203_U387
g19466 nand P2_U3968 P2_R1203_U10 P2_R1203_U84 ; P2_R1203_U388
g19467 nand P2_R1203_U387 P2_R1203_U83 P2_U3054 ; P2_R1203_U389
g19468 nand P2_U3968 P2_R1203_U84 ; P2_R1203_U390
g19469 nand P2_U3054 P2_R1203_U83 ; P2_R1203_U391
g19470 not P2_R1203_U129 ; P2_R1203_U392
g19471 nand P2_R1203_U306 P2_R1203_U392 ; P2_R1203_U393
g19472 nand P2_R1203_U129 P2_R1203_U157 ; P2_R1203_U394
g19473 nand P2_U3969 P2_R1203_U82 ; P2_R1203_U395
g19474 nand P2_U3053 P2_R1203_U79 ; P2_R1203_U396
g19475 nand P2_U3969 P2_R1203_U82 ; P2_R1203_U397
g19476 nand P2_U3053 P2_R1203_U79 ; P2_R1203_U398
g19477 nand P2_R1203_U398 P2_R1203_U397 ; P2_R1203_U399
g19478 nand P2_U3970 P2_R1203_U80 ; P2_R1203_U400
g19479 nand P2_U3057 P2_R1203_U44 ; P2_R1203_U401
g19480 nand P2_R1203_U313 P2_R1203_U85 ; P2_R1203_U402
g19481 nand P2_R1203_U158 P2_R1203_U300 ; P2_R1203_U403
g19482 nand P2_U3971 P2_R1203_U78 ; P2_R1203_U404
g19483 nand P2_U3058 P2_R1203_U77 ; P2_R1203_U405
g19484 not P2_R1203_U132 ; P2_R1203_U406
g19485 nand P2_R1203_U296 P2_R1203_U406 ; P2_R1203_U407
g19486 nand P2_R1203_U132 P2_R1203_U159 ; P2_R1203_U408
g19487 nand P2_U3972 P2_R1203_U76 ; P2_R1203_U409
g19488 nand P2_U3065 P2_R1203_U75 ; P2_R1203_U410
g19489 not P2_R1203_U133 ; P2_R1203_U411
g19490 nand P2_R1203_U292 P2_R1203_U411 ; P2_R1203_U412
g19491 nand P2_R1203_U133 P2_R1203_U160 ; P2_R1203_U413
g19492 nand P2_U3973 P2_R1203_U71 ; P2_R1203_U414
g19493 nand P2_U3066 P2_R1203_U69 ; P2_R1203_U415
g19494 nand P2_R1203_U415 P2_R1203_U414 ; P2_R1203_U416
g19495 nand P2_U3974 P2_R1203_U72 ; P2_R1203_U417
g19496 nand P2_U3061 P2_R1203_U45 ; P2_R1203_U418
g19497 nand P2_R1203_U323 P2_R1203_U86 ; P2_R1203_U419
g19498 nand P2_R1203_U161 P2_R1203_U315 ; P2_R1203_U420
g19499 nand P2_U3975 P2_R1203_U73 ; P2_R1203_U421
g19500 nand P2_U3075 P2_R1203_U70 ; P2_R1203_U422
g19501 nand P2_R1203_U324 P2_R1203_U163 ; P2_R1203_U423
g19502 nand P2_R1203_U282 P2_R1203_U162 ; P2_R1203_U424
g19503 nand P2_U3976 P2_R1203_U68 ; P2_R1203_U425
g19504 nand P2_U3076 P2_R1203_U67 ; P2_R1203_U426
g19505 not P2_R1203_U136 ; P2_R1203_U427
g19506 nand P2_R1203_U278 P2_R1203_U427 ; P2_R1203_U428
g19507 nand P2_R1203_U136 P2_R1203_U164 ; P2_R1203_U429
g19508 nand P2_U3453 P2_R1203_U24 ; P2_R1203_U430
g19509 nand P2_U3078 P2_R1203_U165 ; P2_R1203_U431
g19510 not P2_R1203_U137 ; P2_R1203_U432
g19511 nand P2_R1203_U194 P2_R1203_U432 ; P2_R1203_U433
g19512 nand P2_R1203_U137 P2_R1203_U166 ; P2_R1203_U434
g19513 nand P2_U3506 P2_R1203_U66 ; P2_R1203_U435
g19514 nand P2_U3081 P2_R1203_U65 ; P2_R1203_U436
g19515 not P2_R1203_U138 ; P2_R1203_U437
g19516 nand P2_R1203_U274 P2_R1203_U437 ; P2_R1203_U438
g19517 nand P2_R1203_U138 P2_R1203_U167 ; P2_R1203_U439
g19518 nand P2_U3504 P2_R1203_U64 ; P2_R1203_U440
g19519 nand P2_U3082 P2_R1203_U168 ; P2_R1203_U441
g19520 not P2_R1203_U139 ; P2_R1203_U442
g19521 nand P2_R1203_U272 P2_R1203_U442 ; P2_R1203_U443
g19522 nand P2_R1203_U139 P2_R1203_U169 ; P2_R1203_U444
g19523 nand P2_U3501 P2_R1203_U63 ; P2_R1203_U445
g19524 nand P2_U3069 P2_R1203_U62 ; P2_R1203_U446
g19525 not P2_R1203_U140 ; P2_R1203_U447
g19526 nand P2_R1203_U268 P2_R1203_U447 ; P2_R1203_U448
g19527 nand P2_R1203_U140 P2_R1203_U170 ; P2_R1203_U449
g19528 nand P2_U3498 P2_R1203_U58 ; P2_R1203_U450
g19529 nand P2_U3073 P2_R1203_U56 ; P2_R1203_U451
g19530 nand P2_R1203_U451 P2_R1203_U450 ; P2_R1203_U452
g19531 nand P2_U3495 P2_R1203_U59 ; P2_R1203_U453
g19532 nand P2_U3074 P2_R1203_U46 ; P2_R1203_U454
g19533 nand P2_R1203_U334 P2_R1203_U87 ; P2_R1203_U455
g19534 nand P2_R1203_U171 P2_R1203_U326 ; P2_R1203_U456
g19535 nand P2_U3492 P2_R1203_U60 ; P2_R1203_U457
g19536 nand P2_U3079 P2_R1203_U57 ; P2_R1203_U458
g19537 nand P2_R1203_U335 P2_R1203_U173 ; P2_R1203_U459
g19538 nand P2_R1203_U258 P2_R1203_U172 ; P2_R1203_U460
g19539 nand P2_U3489 P2_R1203_U55 ; P2_R1203_U461
g19540 nand P2_U3080 P2_R1203_U54 ; P2_R1203_U462
g19541 not P2_R1203_U143 ; P2_R1203_U463
g19542 nand P2_R1203_U254 P2_R1203_U463 ; P2_R1203_U464
g19543 nand P2_R1203_U143 P2_R1203_U174 ; P2_R1203_U465
g19544 nand P2_U3486 P2_R1203_U53 ; P2_R1203_U466
g19545 nand P2_U3072 P2_R1203_U52 ; P2_R1203_U467
g19546 not P2_R1203_U144 ; P2_R1203_U468
g19547 nand P2_R1203_U250 P2_R1203_U468 ; P2_R1203_U469
g19548 nand P2_R1203_U144 P2_R1203_U175 ; P2_R1203_U470
g19549 nand P2_U3483 P2_R1203_U49 ; P2_R1203_U471
g19550 nand P2_U3063 P2_R1203_U48 ; P2_R1203_U472
g19551 nand P2_R1203_U472 P2_R1203_U471 ; P2_R1203_U473
g19552 nand P2_U3480 P2_R1203_U50 ; P2_R1203_U474
g19553 nand P2_U3062 P2_R1203_U47 ; P2_R1203_U475
g19554 nand P2_R1203_U345 P2_R1203_U88 ; P2_R1203_U476
g19555 nand P2_R1203_U176 P2_R1203_U337 ; P2_R1203_U477
g19556 and P2_R1113_U205 P2_R1113_U204 ; P2_R1113_U6
g19557 and P2_R1113_U244 P2_R1113_U243 ; P2_R1113_U7
g19558 and P2_R1113_U261 P2_R1113_U260 ; P2_R1113_U8
g19559 and P2_R1113_U285 P2_R1113_U284 ; P2_R1113_U9
g19560 and P2_R1113_U384 P2_R1113_U383 ; P2_R1113_U10
g19561 nand P2_R1113_U340 P2_R1113_U343 ; P2_R1113_U11
g19562 nand P2_R1113_U329 P2_R1113_U332 ; P2_R1113_U12
g19563 nand P2_R1113_U318 P2_R1113_U321 ; P2_R1113_U13
g19564 nand P2_R1113_U310 P2_R1113_U312 ; P2_R1113_U14
g19565 nand P2_R1113_U349 P2_R1113_U177 P2_R1113_U156 ; P2_R1113_U15
g19566 nand P2_R1113_U238 P2_R1113_U240 ; P2_R1113_U16
g19567 nand P2_R1113_U230 P2_R1113_U233 ; P2_R1113_U17
g19568 nand P2_R1113_U222 P2_R1113_U224 ; P2_R1113_U18
g19569 nand P2_R1113_U166 P2_R1113_U346 ; P2_R1113_U19
g19570 not P2_U3471 ; P2_R1113_U20
g19571 not P2_U3465 ; P2_R1113_U21
g19572 not P2_U3456 ; P2_R1113_U22
g19573 not P2_U3448 ; P2_R1113_U23
g19574 not P2_U3078 ; P2_R1113_U24
g19575 not P2_U3459 ; P2_R1113_U25
g19576 not P2_U3068 ; P2_R1113_U26
g19577 nand P2_U3068 P2_R1113_U22 ; P2_R1113_U27
g19578 not P2_U3064 ; P2_R1113_U28
g19579 not P2_U3468 ; P2_R1113_U29
g19580 not P2_U3462 ; P2_R1113_U30
g19581 not P2_U3071 ; P2_R1113_U31
g19582 not P2_U3067 ; P2_R1113_U32
g19583 not P2_U3060 ; P2_R1113_U33
g19584 nand P2_U3060 P2_R1113_U30 ; P2_R1113_U34
g19585 not P2_U3474 ; P2_R1113_U35
g19586 not P2_U3070 ; P2_R1113_U36
g19587 nand P2_U3070 P2_R1113_U20 ; P2_R1113_U37
g19588 not P2_U3084 ; P2_R1113_U38
g19589 not P2_U3477 ; P2_R1113_U39
g19590 not P2_U3083 ; P2_R1113_U40
g19591 nand P2_R1113_U211 P2_R1113_U210 ; P2_R1113_U41
g19592 nand P2_R1113_U34 P2_R1113_U226 ; P2_R1113_U42
g19593 nand P2_R1113_U195 P2_R1113_U179 P2_R1113_U347 ; P2_R1113_U43
g19594 not P2_U3970 ; P2_R1113_U44
g19595 not P2_U3974 ; P2_R1113_U45
g19596 not P2_U3495 ; P2_R1113_U46
g19597 not P2_U3480 ; P2_R1113_U47
g19598 not P2_U3483 ; P2_R1113_U48
g19599 not P2_U3063 ; P2_R1113_U49
g19600 not P2_U3062 ; P2_R1113_U50
g19601 nand P2_U3083 P2_R1113_U39 ; P2_R1113_U51
g19602 not P2_U3486 ; P2_R1113_U52
g19603 not P2_U3072 ; P2_R1113_U53
g19604 not P2_U3489 ; P2_R1113_U54
g19605 not P2_U3080 ; P2_R1113_U55
g19606 not P2_U3498 ; P2_R1113_U56
g19607 not P2_U3492 ; P2_R1113_U57
g19608 not P2_U3073 ; P2_R1113_U58
g19609 not P2_U3074 ; P2_R1113_U59
g19610 not P2_U3079 ; P2_R1113_U60
g19611 nand P2_U3079 P2_R1113_U57 ; P2_R1113_U61
g19612 not P2_U3501 ; P2_R1113_U62
g19613 not P2_U3069 ; P2_R1113_U63
g19614 not P2_U3082 ; P2_R1113_U64
g19615 not P2_U3506 ; P2_R1113_U65
g19616 not P2_U3081 ; P2_R1113_U66
g19617 not P2_U3976 ; P2_R1113_U67
g19618 not P2_U3076 ; P2_R1113_U68
g19619 not P2_U3973 ; P2_R1113_U69
g19620 not P2_U3975 ; P2_R1113_U70
g19621 not P2_U3066 ; P2_R1113_U71
g19622 not P2_U3061 ; P2_R1113_U72
g19623 not P2_U3075 ; P2_R1113_U73
g19624 nand P2_U3075 P2_R1113_U70 ; P2_R1113_U74
g19625 not P2_U3972 ; P2_R1113_U75
g19626 not P2_U3065 ; P2_R1113_U76
g19627 not P2_U3971 ; P2_R1113_U77
g19628 not P2_U3058 ; P2_R1113_U78
g19629 not P2_U3969 ; P2_R1113_U79
g19630 not P2_U3057 ; P2_R1113_U80
g19631 nand P2_U3057 P2_R1113_U44 ; P2_R1113_U81
g19632 not P2_U3053 ; P2_R1113_U82
g19633 not P2_U3968 ; P2_R1113_U83
g19634 not P2_U3054 ; P2_R1113_U84
g19635 nand P2_R1113_U299 P2_R1113_U298 ; P2_R1113_U85
g19636 nand P2_R1113_U74 P2_R1113_U314 ; P2_R1113_U86
g19637 nand P2_R1113_U61 P2_R1113_U325 ; P2_R1113_U87
g19638 nand P2_R1113_U51 P2_R1113_U336 ; P2_R1113_U88
g19639 not P2_U3077 ; P2_R1113_U89
g19640 nand P2_R1113_U394 P2_R1113_U393 ; P2_R1113_U90
g19641 nand P2_R1113_U408 P2_R1113_U407 ; P2_R1113_U91
g19642 nand P2_R1113_U413 P2_R1113_U412 ; P2_R1113_U92
g19643 nand P2_R1113_U429 P2_R1113_U428 ; P2_R1113_U93
g19644 nand P2_R1113_U434 P2_R1113_U433 ; P2_R1113_U94
g19645 nand P2_R1113_U439 P2_R1113_U438 ; P2_R1113_U95
g19646 nand P2_R1113_U444 P2_R1113_U443 ; P2_R1113_U96
g19647 nand P2_R1113_U449 P2_R1113_U448 ; P2_R1113_U97
g19648 nand P2_R1113_U465 P2_R1113_U464 ; P2_R1113_U98
g19649 nand P2_R1113_U470 P2_R1113_U469 ; P2_R1113_U99
g19650 nand P2_R1113_U353 P2_R1113_U352 ; P2_R1113_U100
g19651 nand P2_R1113_U362 P2_R1113_U361 ; P2_R1113_U101
g19652 nand P2_R1113_U369 P2_R1113_U368 ; P2_R1113_U102
g19653 nand P2_R1113_U373 P2_R1113_U372 ; P2_R1113_U103
g19654 nand P2_R1113_U382 P2_R1113_U381 ; P2_R1113_U104
g19655 nand P2_R1113_U403 P2_R1113_U402 ; P2_R1113_U105
g19656 nand P2_R1113_U420 P2_R1113_U419 ; P2_R1113_U106
g19657 nand P2_R1113_U424 P2_R1113_U423 ; P2_R1113_U107
g19658 nand P2_R1113_U456 P2_R1113_U455 ; P2_R1113_U108
g19659 nand P2_R1113_U460 P2_R1113_U459 ; P2_R1113_U109
g19660 nand P2_R1113_U477 P2_R1113_U476 ; P2_R1113_U110
g19661 and P2_R1113_U197 P2_R1113_U187 ; P2_R1113_U111
g19662 and P2_R1113_U200 P2_R1113_U201 ; P2_R1113_U112
g19663 and P2_R1113_U208 P2_R1113_U203 P2_R1113_U188 ; P2_R1113_U113
g19664 and P2_R1113_U213 P2_R1113_U189 ; P2_R1113_U114
g19665 and P2_R1113_U216 P2_R1113_U217 ; P2_R1113_U115
g19666 and P2_R1113_U355 P2_R1113_U354 P2_R1113_U37 ; P2_R1113_U116
g19667 and P2_R1113_U358 P2_R1113_U189 ; P2_R1113_U117
g19668 and P2_R1113_U232 P2_R1113_U6 ; P2_R1113_U118
g19669 and P2_R1113_U365 P2_R1113_U188 ; P2_R1113_U119
g19670 and P2_R1113_U375 P2_R1113_U374 P2_R1113_U27 ; P2_R1113_U120
g19671 and P2_R1113_U378 P2_R1113_U187 ; P2_R1113_U121
g19672 and P2_R1113_U242 P2_R1113_U219 P2_R1113_U183 ; P2_R1113_U122
g19673 and P2_R1113_U264 P2_R1113_U184 P2_R1113_U259 ; P2_R1113_U123
g19674 and P2_R1113_U288 P2_R1113_U185 P2_R1113_U283 ; P2_R1113_U124
g19675 and P2_R1113_U301 P2_R1113_U186 ; P2_R1113_U125
g19676 and P2_R1113_U304 P2_R1113_U305 ; P2_R1113_U126
g19677 and P2_R1113_U304 P2_R1113_U305 ; P2_R1113_U127
g19678 and P2_R1113_U10 P2_R1113_U308 ; P2_R1113_U128
g19679 nand P2_R1113_U391 P2_R1113_U390 ; P2_R1113_U129
g19680 and P2_R1113_U396 P2_R1113_U395 P2_R1113_U81 ; P2_R1113_U130
g19681 and P2_R1113_U399 P2_R1113_U186 ; P2_R1113_U131
g19682 nand P2_R1113_U405 P2_R1113_U404 ; P2_R1113_U132
g19683 nand P2_R1113_U410 P2_R1113_U409 ; P2_R1113_U133
g19684 and P2_R1113_U320 P2_R1113_U9 ; P2_R1113_U134
g19685 and P2_R1113_U416 P2_R1113_U185 ; P2_R1113_U135
g19686 nand P2_R1113_U426 P2_R1113_U425 ; P2_R1113_U136
g19687 nand P2_R1113_U431 P2_R1113_U430 ; P2_R1113_U137
g19688 nand P2_R1113_U436 P2_R1113_U435 ; P2_R1113_U138
g19689 nand P2_R1113_U441 P2_R1113_U440 ; P2_R1113_U139
g19690 nand P2_R1113_U446 P2_R1113_U445 ; P2_R1113_U140
g19691 and P2_R1113_U331 P2_R1113_U8 ; P2_R1113_U141
g19692 and P2_R1113_U452 P2_R1113_U184 ; P2_R1113_U142
g19693 nand P2_R1113_U462 P2_R1113_U461 ; P2_R1113_U143
g19694 nand P2_R1113_U467 P2_R1113_U466 ; P2_R1113_U144
g19695 and P2_R1113_U342 P2_R1113_U7 ; P2_R1113_U145
g19696 and P2_R1113_U473 P2_R1113_U183 ; P2_R1113_U146
g19697 and P2_R1113_U351 P2_R1113_U350 ; P2_R1113_U147
g19698 nand P2_R1113_U115 P2_R1113_U214 ; P2_R1113_U148
g19699 and P2_R1113_U360 P2_R1113_U359 ; P2_R1113_U149
g19700 and P2_R1113_U367 P2_R1113_U366 ; P2_R1113_U150
g19701 and P2_R1113_U371 P2_R1113_U370 ; P2_R1113_U151
g19702 nand P2_R1113_U112 P2_R1113_U198 ; P2_R1113_U152
g19703 and P2_R1113_U380 P2_R1113_U379 ; P2_R1113_U153
g19704 not P2_U3979 ; P2_R1113_U154
g19705 not P2_U3055 ; P2_R1113_U155
g19706 and P2_R1113_U389 P2_R1113_U388 ; P2_R1113_U156
g19707 nand P2_R1113_U126 P2_R1113_U302 ; P2_R1113_U157
g19708 and P2_R1113_U401 P2_R1113_U400 ; P2_R1113_U158
g19709 nand P2_R1113_U295 P2_R1113_U294 ; P2_R1113_U159
g19710 nand P2_R1113_U291 P2_R1113_U290 ; P2_R1113_U160
g19711 and P2_R1113_U418 P2_R1113_U417 ; P2_R1113_U161
g19712 and P2_R1113_U422 P2_R1113_U421 ; P2_R1113_U162
g19713 nand P2_R1113_U281 P2_R1113_U280 ; P2_R1113_U163
g19714 nand P2_R1113_U277 P2_R1113_U276 ; P2_R1113_U164
g19715 not P2_U3453 ; P2_R1113_U165
g19716 nand P2_U3448 P2_R1113_U89 ; P2_R1113_U166
g19717 nand P2_R1113_U273 P2_R1113_U178 P2_R1113_U348 ; P2_R1113_U167
g19718 not P2_U3504 ; P2_R1113_U168
g19719 nand P2_R1113_U271 P2_R1113_U270 ; P2_R1113_U169
g19720 nand P2_R1113_U267 P2_R1113_U266 ; P2_R1113_U170
g19721 and P2_R1113_U454 P2_R1113_U453 ; P2_R1113_U171
g19722 and P2_R1113_U458 P2_R1113_U457 ; P2_R1113_U172
g19723 nand P2_R1113_U257 P2_R1113_U256 ; P2_R1113_U173
g19724 nand P2_R1113_U253 P2_R1113_U252 ; P2_R1113_U174
g19725 nand P2_R1113_U249 P2_R1113_U248 ; P2_R1113_U175
g19726 and P2_R1113_U475 P2_R1113_U474 ; P2_R1113_U176
g19727 nand P2_R1113_U307 P2_R1113_U157 P2_R1113_U387 ; P2_R1113_U177
g19728 nand P2_R1113_U169 P2_R1113_U168 ; P2_R1113_U178
g19729 nand P2_R1113_U166 P2_R1113_U165 ; P2_R1113_U179
g19730 not P2_R1113_U81 ; P2_R1113_U180
g19731 not P2_R1113_U27 ; P2_R1113_U181
g19732 not P2_R1113_U37 ; P2_R1113_U182
g19733 nand P2_U3480 P2_R1113_U50 ; P2_R1113_U183
g19734 nand P2_U3495 P2_R1113_U59 ; P2_R1113_U184
g19735 nand P2_U3974 P2_R1113_U72 ; P2_R1113_U185
g19736 nand P2_U3970 P2_R1113_U80 ; P2_R1113_U186
g19737 nand P2_U3456 P2_R1113_U26 ; P2_R1113_U187
g19738 nand P2_U3465 P2_R1113_U32 ; P2_R1113_U188
g19739 nand P2_U3471 P2_R1113_U36 ; P2_R1113_U189
g19740 not P2_R1113_U61 ; P2_R1113_U190
g19741 not P2_R1113_U74 ; P2_R1113_U191
g19742 not P2_R1113_U34 ; P2_R1113_U192
g19743 not P2_R1113_U51 ; P2_R1113_U193
g19744 not P2_R1113_U166 ; P2_R1113_U194
g19745 nand P2_U3078 P2_R1113_U166 ; P2_R1113_U195
g19746 not P2_R1113_U43 ; P2_R1113_U196
g19747 nand P2_U3459 P2_R1113_U28 ; P2_R1113_U197
g19748 nand P2_R1113_U111 P2_R1113_U43 ; P2_R1113_U198
g19749 nand P2_R1113_U28 P2_R1113_U27 ; P2_R1113_U199
g19750 nand P2_R1113_U199 P2_R1113_U25 ; P2_R1113_U200
g19751 nand P2_U3064 P2_R1113_U181 ; P2_R1113_U201
g19752 not P2_R1113_U152 ; P2_R1113_U202
g19753 nand P2_U3468 P2_R1113_U31 ; P2_R1113_U203
g19754 nand P2_U3071 P2_R1113_U29 ; P2_R1113_U204
g19755 nand P2_U3067 P2_R1113_U21 ; P2_R1113_U205
g19756 nand P2_R1113_U192 P2_R1113_U188 ; P2_R1113_U206
g19757 nand P2_R1113_U6 P2_R1113_U206 ; P2_R1113_U207
g19758 nand P2_U3462 P2_R1113_U33 ; P2_R1113_U208
g19759 nand P2_U3468 P2_R1113_U31 ; P2_R1113_U209
g19760 nand P2_R1113_U152 P2_R1113_U113 ; P2_R1113_U210
g19761 nand P2_R1113_U209 P2_R1113_U207 ; P2_R1113_U211
g19762 not P2_R1113_U41 ; P2_R1113_U212
g19763 nand P2_U3474 P2_R1113_U38 ; P2_R1113_U213
g19764 nand P2_R1113_U114 P2_R1113_U41 ; P2_R1113_U214
g19765 nand P2_R1113_U38 P2_R1113_U37 ; P2_R1113_U215
g19766 nand P2_R1113_U215 P2_R1113_U35 ; P2_R1113_U216
g19767 nand P2_U3084 P2_R1113_U182 ; P2_R1113_U217
g19768 not P2_R1113_U148 ; P2_R1113_U218
g19769 nand P2_U3477 P2_R1113_U40 ; P2_R1113_U219
g19770 nand P2_R1113_U219 P2_R1113_U51 ; P2_R1113_U220
g19771 nand P2_R1113_U212 P2_R1113_U37 ; P2_R1113_U221
g19772 nand P2_R1113_U117 P2_R1113_U221 ; P2_R1113_U222
g19773 nand P2_R1113_U41 P2_R1113_U189 ; P2_R1113_U223
g19774 nand P2_R1113_U116 P2_R1113_U223 ; P2_R1113_U224
g19775 nand P2_R1113_U37 P2_R1113_U189 ; P2_R1113_U225
g19776 nand P2_R1113_U208 P2_R1113_U152 ; P2_R1113_U226
g19777 not P2_R1113_U42 ; P2_R1113_U227
g19778 nand P2_U3067 P2_R1113_U21 ; P2_R1113_U228
g19779 nand P2_R1113_U227 P2_R1113_U228 ; P2_R1113_U229
g19780 nand P2_R1113_U119 P2_R1113_U229 ; P2_R1113_U230
g19781 nand P2_R1113_U42 P2_R1113_U188 ; P2_R1113_U231
g19782 nand P2_U3468 P2_R1113_U31 ; P2_R1113_U232
g19783 nand P2_R1113_U118 P2_R1113_U231 ; P2_R1113_U233
g19784 nand P2_U3067 P2_R1113_U21 ; P2_R1113_U234
g19785 nand P2_R1113_U188 P2_R1113_U234 ; P2_R1113_U235
g19786 nand P2_R1113_U208 P2_R1113_U34 ; P2_R1113_U236
g19787 nand P2_R1113_U196 P2_R1113_U27 ; P2_R1113_U237
g19788 nand P2_R1113_U121 P2_R1113_U237 ; P2_R1113_U238
g19789 nand P2_R1113_U43 P2_R1113_U187 ; P2_R1113_U239
g19790 nand P2_R1113_U120 P2_R1113_U239 ; P2_R1113_U240
g19791 nand P2_R1113_U27 P2_R1113_U187 ; P2_R1113_U241
g19792 nand P2_U3483 P2_R1113_U49 ; P2_R1113_U242
g19793 nand P2_U3063 P2_R1113_U48 ; P2_R1113_U243
g19794 nand P2_U3062 P2_R1113_U47 ; P2_R1113_U244
g19795 nand P2_R1113_U193 P2_R1113_U183 ; P2_R1113_U245
g19796 nand P2_R1113_U7 P2_R1113_U245 ; P2_R1113_U246
g19797 nand P2_U3483 P2_R1113_U49 ; P2_R1113_U247
g19798 nand P2_R1113_U148 P2_R1113_U122 ; P2_R1113_U248
g19799 nand P2_R1113_U247 P2_R1113_U246 ; P2_R1113_U249
g19800 not P2_R1113_U175 ; P2_R1113_U250
g19801 nand P2_U3486 P2_R1113_U53 ; P2_R1113_U251
g19802 nand P2_R1113_U251 P2_R1113_U175 ; P2_R1113_U252
g19803 nand P2_U3072 P2_R1113_U52 ; P2_R1113_U253
g19804 not P2_R1113_U174 ; P2_R1113_U254
g19805 nand P2_U3489 P2_R1113_U55 ; P2_R1113_U255
g19806 nand P2_R1113_U255 P2_R1113_U174 ; P2_R1113_U256
g19807 nand P2_U3080 P2_R1113_U54 ; P2_R1113_U257
g19808 not P2_R1113_U173 ; P2_R1113_U258
g19809 nand P2_U3498 P2_R1113_U58 ; P2_R1113_U259
g19810 nand P2_U3073 P2_R1113_U56 ; P2_R1113_U260
g19811 nand P2_U3074 P2_R1113_U46 ; P2_R1113_U261
g19812 nand P2_R1113_U190 P2_R1113_U184 ; P2_R1113_U262
g19813 nand P2_R1113_U8 P2_R1113_U262 ; P2_R1113_U263
g19814 nand P2_U3492 P2_R1113_U60 ; P2_R1113_U264
g19815 nand P2_U3498 P2_R1113_U58 ; P2_R1113_U265
g19816 nand P2_R1113_U173 P2_R1113_U123 ; P2_R1113_U266
g19817 nand P2_R1113_U265 P2_R1113_U263 ; P2_R1113_U267
g19818 not P2_R1113_U170 ; P2_R1113_U268
g19819 nand P2_U3501 P2_R1113_U63 ; P2_R1113_U269
g19820 nand P2_R1113_U269 P2_R1113_U170 ; P2_R1113_U270
g19821 nand P2_U3069 P2_R1113_U62 ; P2_R1113_U271
g19822 not P2_R1113_U169 ; P2_R1113_U272
g19823 nand P2_U3082 P2_R1113_U169 ; P2_R1113_U273
g19824 not P2_R1113_U167 ; P2_R1113_U274
g19825 nand P2_U3506 P2_R1113_U66 ; P2_R1113_U275
g19826 nand P2_R1113_U275 P2_R1113_U167 ; P2_R1113_U276
g19827 nand P2_U3081 P2_R1113_U65 ; P2_R1113_U277
g19828 not P2_R1113_U164 ; P2_R1113_U278
g19829 nand P2_U3976 P2_R1113_U68 ; P2_R1113_U279
g19830 nand P2_R1113_U279 P2_R1113_U164 ; P2_R1113_U280
g19831 nand P2_U3076 P2_R1113_U67 ; P2_R1113_U281
g19832 not P2_R1113_U163 ; P2_R1113_U282
g19833 nand P2_U3973 P2_R1113_U71 ; P2_R1113_U283
g19834 nand P2_U3066 P2_R1113_U69 ; P2_R1113_U284
g19835 nand P2_U3061 P2_R1113_U45 ; P2_R1113_U285
g19836 nand P2_R1113_U191 P2_R1113_U185 ; P2_R1113_U286
g19837 nand P2_R1113_U9 P2_R1113_U286 ; P2_R1113_U287
g19838 nand P2_U3975 P2_R1113_U73 ; P2_R1113_U288
g19839 nand P2_U3973 P2_R1113_U71 ; P2_R1113_U289
g19840 nand P2_R1113_U163 P2_R1113_U124 ; P2_R1113_U290
g19841 nand P2_R1113_U289 P2_R1113_U287 ; P2_R1113_U291
g19842 not P2_R1113_U160 ; P2_R1113_U292
g19843 nand P2_U3972 P2_R1113_U76 ; P2_R1113_U293
g19844 nand P2_R1113_U293 P2_R1113_U160 ; P2_R1113_U294
g19845 nand P2_U3065 P2_R1113_U75 ; P2_R1113_U295
g19846 not P2_R1113_U159 ; P2_R1113_U296
g19847 nand P2_U3971 P2_R1113_U78 ; P2_R1113_U297
g19848 nand P2_R1113_U297 P2_R1113_U159 ; P2_R1113_U298
g19849 nand P2_U3058 P2_R1113_U77 ; P2_R1113_U299
g19850 not P2_R1113_U85 ; P2_R1113_U300
g19851 nand P2_U3969 P2_R1113_U82 ; P2_R1113_U301
g19852 nand P2_R1113_U125 P2_R1113_U85 ; P2_R1113_U302
g19853 nand P2_R1113_U82 P2_R1113_U81 ; P2_R1113_U303
g19854 nand P2_R1113_U303 P2_R1113_U79 ; P2_R1113_U304
g19855 nand P2_U3053 P2_R1113_U180 ; P2_R1113_U305
g19856 not P2_R1113_U157 ; P2_R1113_U306
g19857 nand P2_U3968 P2_R1113_U84 ; P2_R1113_U307
g19858 nand P2_U3054 P2_R1113_U83 ; P2_R1113_U308
g19859 nand P2_R1113_U300 P2_R1113_U81 ; P2_R1113_U309
g19860 nand P2_R1113_U131 P2_R1113_U309 ; P2_R1113_U310
g19861 nand P2_R1113_U85 P2_R1113_U186 ; P2_R1113_U311
g19862 nand P2_R1113_U130 P2_R1113_U311 ; P2_R1113_U312
g19863 nand P2_R1113_U81 P2_R1113_U186 ; P2_R1113_U313
g19864 nand P2_R1113_U288 P2_R1113_U163 ; P2_R1113_U314
g19865 not P2_R1113_U86 ; P2_R1113_U315
g19866 nand P2_U3061 P2_R1113_U45 ; P2_R1113_U316
g19867 nand P2_R1113_U315 P2_R1113_U316 ; P2_R1113_U317
g19868 nand P2_R1113_U135 P2_R1113_U317 ; P2_R1113_U318
g19869 nand P2_R1113_U86 P2_R1113_U185 ; P2_R1113_U319
g19870 nand P2_U3973 P2_R1113_U71 ; P2_R1113_U320
g19871 nand P2_R1113_U134 P2_R1113_U319 ; P2_R1113_U321
g19872 nand P2_U3061 P2_R1113_U45 ; P2_R1113_U322
g19873 nand P2_R1113_U185 P2_R1113_U322 ; P2_R1113_U323
g19874 nand P2_R1113_U288 P2_R1113_U74 ; P2_R1113_U324
g19875 nand P2_R1113_U264 P2_R1113_U173 ; P2_R1113_U325
g19876 not P2_R1113_U87 ; P2_R1113_U326
g19877 nand P2_U3074 P2_R1113_U46 ; P2_R1113_U327
g19878 nand P2_R1113_U326 P2_R1113_U327 ; P2_R1113_U328
g19879 nand P2_R1113_U142 P2_R1113_U328 ; P2_R1113_U329
g19880 nand P2_R1113_U87 P2_R1113_U184 ; P2_R1113_U330
g19881 nand P2_U3498 P2_R1113_U58 ; P2_R1113_U331
g19882 nand P2_R1113_U141 P2_R1113_U330 ; P2_R1113_U332
g19883 nand P2_U3074 P2_R1113_U46 ; P2_R1113_U333
g19884 nand P2_R1113_U184 P2_R1113_U333 ; P2_R1113_U334
g19885 nand P2_R1113_U264 P2_R1113_U61 ; P2_R1113_U335
g19886 nand P2_R1113_U219 P2_R1113_U148 ; P2_R1113_U336
g19887 not P2_R1113_U88 ; P2_R1113_U337
g19888 nand P2_U3062 P2_R1113_U47 ; P2_R1113_U338
g19889 nand P2_R1113_U337 P2_R1113_U338 ; P2_R1113_U339
g19890 nand P2_R1113_U146 P2_R1113_U339 ; P2_R1113_U340
g19891 nand P2_R1113_U88 P2_R1113_U183 ; P2_R1113_U341
g19892 nand P2_U3483 P2_R1113_U49 ; P2_R1113_U342
g19893 nand P2_R1113_U145 P2_R1113_U341 ; P2_R1113_U343
g19894 nand P2_U3062 P2_R1113_U47 ; P2_R1113_U344
g19895 nand P2_R1113_U183 P2_R1113_U344 ; P2_R1113_U345
g19896 nand P2_U3077 P2_R1113_U23 ; P2_R1113_U346
g19897 nand P2_U3078 P2_R1113_U165 ; P2_R1113_U347
g19898 nand P2_U3082 P2_R1113_U168 ; P2_R1113_U348
g19899 nand P2_R1113_U127 P2_R1113_U302 P2_R1113_U128 ; P2_R1113_U349
g19900 nand P2_U3477 P2_R1113_U40 ; P2_R1113_U350
g19901 nand P2_U3083 P2_R1113_U39 ; P2_R1113_U351
g19902 nand P2_R1113_U220 P2_R1113_U148 ; P2_R1113_U352
g19903 nand P2_R1113_U218 P2_R1113_U147 ; P2_R1113_U353
g19904 nand P2_U3474 P2_R1113_U38 ; P2_R1113_U354
g19905 nand P2_U3084 P2_R1113_U35 ; P2_R1113_U355
g19906 nand P2_U3474 P2_R1113_U38 ; P2_R1113_U356
g19907 nand P2_U3084 P2_R1113_U35 ; P2_R1113_U357
g19908 nand P2_R1113_U357 P2_R1113_U356 ; P2_R1113_U358
g19909 nand P2_U3471 P2_R1113_U36 ; P2_R1113_U359
g19910 nand P2_U3070 P2_R1113_U20 ; P2_R1113_U360
g19911 nand P2_R1113_U225 P2_R1113_U41 ; P2_R1113_U361
g19912 nand P2_R1113_U149 P2_R1113_U212 ; P2_R1113_U362
g19913 nand P2_U3468 P2_R1113_U31 ; P2_R1113_U363
g19914 nand P2_U3071 P2_R1113_U29 ; P2_R1113_U364
g19915 nand P2_R1113_U364 P2_R1113_U363 ; P2_R1113_U365
g19916 nand P2_U3465 P2_R1113_U32 ; P2_R1113_U366
g19917 nand P2_U3067 P2_R1113_U21 ; P2_R1113_U367
g19918 nand P2_R1113_U235 P2_R1113_U42 ; P2_R1113_U368
g19919 nand P2_R1113_U150 P2_R1113_U227 ; P2_R1113_U369
g19920 nand P2_U3462 P2_R1113_U33 ; P2_R1113_U370
g19921 nand P2_U3060 P2_R1113_U30 ; P2_R1113_U371
g19922 nand P2_R1113_U236 P2_R1113_U152 ; P2_R1113_U372
g19923 nand P2_R1113_U202 P2_R1113_U151 ; P2_R1113_U373
g19924 nand P2_U3459 P2_R1113_U28 ; P2_R1113_U374
g19925 nand P2_U3064 P2_R1113_U25 ; P2_R1113_U375
g19926 nand P2_U3459 P2_R1113_U28 ; P2_R1113_U376
g19927 nand P2_U3064 P2_R1113_U25 ; P2_R1113_U377
g19928 nand P2_R1113_U377 P2_R1113_U376 ; P2_R1113_U378
g19929 nand P2_U3456 P2_R1113_U26 ; P2_R1113_U379
g19930 nand P2_U3068 P2_R1113_U22 ; P2_R1113_U380
g19931 nand P2_R1113_U241 P2_R1113_U43 ; P2_R1113_U381
g19932 nand P2_R1113_U153 P2_R1113_U196 ; P2_R1113_U382
g19933 nand P2_U3979 P2_R1113_U155 ; P2_R1113_U383
g19934 nand P2_U3055 P2_R1113_U154 ; P2_R1113_U384
g19935 nand P2_U3979 P2_R1113_U155 ; P2_R1113_U385
g19936 nand P2_U3055 P2_R1113_U154 ; P2_R1113_U386
g19937 nand P2_R1113_U386 P2_R1113_U385 ; P2_R1113_U387
g19938 nand P2_U3968 P2_R1113_U10 P2_R1113_U84 ; P2_R1113_U388
g19939 nand P2_R1113_U387 P2_R1113_U83 P2_U3054 ; P2_R1113_U389
g19940 nand P2_U3968 P2_R1113_U84 ; P2_R1113_U390
g19941 nand P2_U3054 P2_R1113_U83 ; P2_R1113_U391
g19942 not P2_R1113_U129 ; P2_R1113_U392
g19943 nand P2_R1113_U306 P2_R1113_U392 ; P2_R1113_U393
g19944 nand P2_R1113_U129 P2_R1113_U157 ; P2_R1113_U394
g19945 nand P2_U3969 P2_R1113_U82 ; P2_R1113_U395
g19946 nand P2_U3053 P2_R1113_U79 ; P2_R1113_U396
g19947 nand P2_U3969 P2_R1113_U82 ; P2_R1113_U397
g19948 nand P2_U3053 P2_R1113_U79 ; P2_R1113_U398
g19949 nand P2_R1113_U398 P2_R1113_U397 ; P2_R1113_U399
g19950 nand P2_U3970 P2_R1113_U80 ; P2_R1113_U400
g19951 nand P2_U3057 P2_R1113_U44 ; P2_R1113_U401
g19952 nand P2_R1113_U313 P2_R1113_U85 ; P2_R1113_U402
g19953 nand P2_R1113_U158 P2_R1113_U300 ; P2_R1113_U403
g19954 nand P2_U3971 P2_R1113_U78 ; P2_R1113_U404
g19955 nand P2_U3058 P2_R1113_U77 ; P2_R1113_U405
g19956 not P2_R1113_U132 ; P2_R1113_U406
g19957 nand P2_R1113_U296 P2_R1113_U406 ; P2_R1113_U407
g19958 nand P2_R1113_U132 P2_R1113_U159 ; P2_R1113_U408
g19959 nand P2_U3972 P2_R1113_U76 ; P2_R1113_U409
g19960 nand P2_U3065 P2_R1113_U75 ; P2_R1113_U410
g19961 not P2_R1113_U133 ; P2_R1113_U411
g19962 nand P2_R1113_U292 P2_R1113_U411 ; P2_R1113_U412
g19963 nand P2_R1113_U133 P2_R1113_U160 ; P2_R1113_U413
g19964 nand P2_U3973 P2_R1113_U71 ; P2_R1113_U414
g19965 nand P2_U3066 P2_R1113_U69 ; P2_R1113_U415
g19966 nand P2_R1113_U415 P2_R1113_U414 ; P2_R1113_U416
g19967 nand P2_U3974 P2_R1113_U72 ; P2_R1113_U417
g19968 nand P2_U3061 P2_R1113_U45 ; P2_R1113_U418
g19969 nand P2_R1113_U323 P2_R1113_U86 ; P2_R1113_U419
g19970 nand P2_R1113_U161 P2_R1113_U315 ; P2_R1113_U420
g19971 nand P2_U3975 P2_R1113_U73 ; P2_R1113_U421
g19972 nand P2_U3075 P2_R1113_U70 ; P2_R1113_U422
g19973 nand P2_R1113_U324 P2_R1113_U163 ; P2_R1113_U423
g19974 nand P2_R1113_U282 P2_R1113_U162 ; P2_R1113_U424
g19975 nand P2_U3976 P2_R1113_U68 ; P2_R1113_U425
g19976 nand P2_U3076 P2_R1113_U67 ; P2_R1113_U426
g19977 not P2_R1113_U136 ; P2_R1113_U427
g19978 nand P2_R1113_U278 P2_R1113_U427 ; P2_R1113_U428
g19979 nand P2_R1113_U136 P2_R1113_U164 ; P2_R1113_U429
g19980 nand P2_U3453 P2_R1113_U24 ; P2_R1113_U430
g19981 nand P2_U3078 P2_R1113_U165 ; P2_R1113_U431
g19982 not P2_R1113_U137 ; P2_R1113_U432
g19983 nand P2_R1113_U194 P2_R1113_U432 ; P2_R1113_U433
g19984 nand P2_R1113_U137 P2_R1113_U166 ; P2_R1113_U434
g19985 nand P2_U3506 P2_R1113_U66 ; P2_R1113_U435
g19986 nand P2_U3081 P2_R1113_U65 ; P2_R1113_U436
g19987 not P2_R1113_U138 ; P2_R1113_U437
g19988 nand P2_R1113_U274 P2_R1113_U437 ; P2_R1113_U438
g19989 nand P2_R1113_U138 P2_R1113_U167 ; P2_R1113_U439
g19990 nand P2_U3504 P2_R1113_U64 ; P2_R1113_U440
g19991 nand P2_U3082 P2_R1113_U168 ; P2_R1113_U441
g19992 not P2_R1113_U139 ; P2_R1113_U442
g19993 nand P2_R1113_U272 P2_R1113_U442 ; P2_R1113_U443
g19994 nand P2_R1113_U139 P2_R1113_U169 ; P2_R1113_U444
g19995 nand P2_U3501 P2_R1113_U63 ; P2_R1113_U445
g19996 nand P2_U3069 P2_R1113_U62 ; P2_R1113_U446
g19997 not P2_R1113_U140 ; P2_R1113_U447
g19998 nand P2_R1113_U268 P2_R1113_U447 ; P2_R1113_U448
g19999 nand P2_R1113_U140 P2_R1113_U170 ; P2_R1113_U449
g20000 nand P2_U3498 P2_R1113_U58 ; P2_R1113_U450
g20001 nand P2_U3073 P2_R1113_U56 ; P2_R1113_U451
g20002 nand P2_R1113_U451 P2_R1113_U450 ; P2_R1113_U452
g20003 nand P2_U3495 P2_R1113_U59 ; P2_R1113_U453
g20004 nand P2_U3074 P2_R1113_U46 ; P2_R1113_U454
g20005 nand P2_R1113_U334 P2_R1113_U87 ; P2_R1113_U455
g20006 nand P2_R1113_U171 P2_R1113_U326 ; P2_R1113_U456
g20007 nand P2_U3492 P2_R1113_U60 ; P2_R1113_U457
g20008 nand P2_U3079 P2_R1113_U57 ; P2_R1113_U458
g20009 nand P2_R1113_U335 P2_R1113_U173 ; P2_R1113_U459
g20010 nand P2_R1113_U258 P2_R1113_U172 ; P2_R1113_U460
g20011 nand P2_U3489 P2_R1113_U55 ; P2_R1113_U461
g20012 nand P2_U3080 P2_R1113_U54 ; P2_R1113_U462
g20013 not P2_R1113_U143 ; P2_R1113_U463
g20014 nand P2_R1113_U254 P2_R1113_U463 ; P2_R1113_U464
g20015 nand P2_R1113_U143 P2_R1113_U174 ; P2_R1113_U465
g20016 nand P2_U3486 P2_R1113_U53 ; P2_R1113_U466
g20017 nand P2_U3072 P2_R1113_U52 ; P2_R1113_U467
g20018 not P2_R1113_U144 ; P2_R1113_U468
g20019 nand P2_R1113_U250 P2_R1113_U468 ; P2_R1113_U469
g20020 nand P2_R1113_U144 P2_R1113_U175 ; P2_R1113_U470
g20021 nand P2_U3483 P2_R1113_U49 ; P2_R1113_U471
g20022 nand P2_U3063 P2_R1113_U48 ; P2_R1113_U472
g20023 nand P2_R1113_U472 P2_R1113_U471 ; P2_R1113_U473
g20024 nand P2_U3480 P2_R1113_U50 ; P2_R1113_U474
g20025 nand P2_U3062 P2_R1113_U47 ; P2_R1113_U475
g20026 nand P2_R1113_U345 P2_R1113_U88 ; P2_R1113_U476
g20027 nand P2_R1113_U176 P2_R1113_U337 ; P2_R1113_U477
