i P3_WR_REG_SCAN_IN
i SI_31_
i SI_30_
i SI_29_
i SI_28_
i SI_27_
i SI_26_
i SI_25_
i SI_24_
i SI_23_
i SI_22_
i SI_21_
i SI_20_
i SI_19_
i SI_18_
i SI_17_
i SI_16_
i SI_15_
i SI_14_
i SI_13_
i SI_12_
i SI_11_
i SI_10_
i SI_9_
i SI_8_
i SI_7_
i SI_6_
i SI_5_
i SI_4_
i SI_3_
i SI_2_
i SI_1_
i SI_0_
i P3_RD_REG_SCAN_IN
i P3_STATE_REG_SCAN_IN
i P3_REG3_REG_7__SCAN_IN
i P3_REG3_REG_27__SCAN_IN
i P3_REG3_REG_14__SCAN_IN
i P3_REG3_REG_23__SCAN_IN
i P3_REG3_REG_10__SCAN_IN
i P3_REG3_REG_3__SCAN_IN
i P3_REG3_REG_19__SCAN_IN
i P3_REG3_REG_28__SCAN_IN
i P3_REG3_REG_8__SCAN_IN
i P3_REG3_REG_1__SCAN_IN
i P3_REG3_REG_21__SCAN_IN
i P3_REG3_REG_12__SCAN_IN
i P3_REG3_REG_25__SCAN_IN
i P3_REG3_REG_16__SCAN_IN
i P3_REG3_REG_5__SCAN_IN
i P3_REG3_REG_17__SCAN_IN
i P3_REG3_REG_24__SCAN_IN
i P3_REG3_REG_4__SCAN_IN
i P3_REG3_REG_9__SCAN_IN
i P3_REG3_REG_0__SCAN_IN
i P3_REG3_REG_20__SCAN_IN
i P3_REG3_REG_13__SCAN_IN
i P3_REG3_REG_22__SCAN_IN
i P3_REG3_REG_11__SCAN_IN
i P3_REG3_REG_2__SCAN_IN
i P3_REG3_REG_18__SCAN_IN
i P3_REG3_REG_6__SCAN_IN
i P3_REG3_REG_26__SCAN_IN
i P3_REG3_REG_15__SCAN_IN
i P3_B_REG_SCAN_IN
i P3_DATAO_REG_31__SCAN_IN
i P3_DATAO_REG_30__SCAN_IN
i P3_DATAO_REG_29__SCAN_IN
i P3_DATAO_REG_28__SCAN_IN
i P3_DATAO_REG_27__SCAN_IN
i P3_DATAO_REG_26__SCAN_IN
i P3_DATAO_REG_25__SCAN_IN
i P3_DATAO_REG_24__SCAN_IN
i P3_DATAO_REG_23__SCAN_IN
i P3_DATAO_REG_22__SCAN_IN
i P3_DATAO_REG_21__SCAN_IN
i P3_DATAO_REG_20__SCAN_IN
i P3_DATAO_REG_19__SCAN_IN
i P3_DATAO_REG_18__SCAN_IN
i P3_DATAO_REG_17__SCAN_IN
i P3_DATAO_REG_16__SCAN_IN
i P3_DATAO_REG_15__SCAN_IN
i P3_DATAO_REG_14__SCAN_IN
i P3_DATAO_REG_13__SCAN_IN
i P3_DATAO_REG_12__SCAN_IN
i P3_DATAO_REG_11__SCAN_IN
i P3_DATAO_REG_10__SCAN_IN
i P3_DATAO_REG_9__SCAN_IN
i P3_DATAO_REG_8__SCAN_IN
i P3_DATAO_REG_7__SCAN_IN
i P3_DATAO_REG_6__SCAN_IN
i P3_DATAO_REG_5__SCAN_IN
i P3_DATAO_REG_4__SCAN_IN
i P3_DATAO_REG_3__SCAN_IN
i P3_DATAO_REG_2__SCAN_IN
i P3_DATAO_REG_1__SCAN_IN
i P3_DATAO_REG_0__SCAN_IN
i P3_ADDR_REG_0__SCAN_IN
i P3_ADDR_REG_1__SCAN_IN
i P3_ADDR_REG_2__SCAN_IN
i P3_ADDR_REG_3__SCAN_IN
i P3_ADDR_REG_4__SCAN_IN
i P3_ADDR_REG_5__SCAN_IN
i P3_ADDR_REG_6__SCAN_IN
i P3_ADDR_REG_7__SCAN_IN
i P3_ADDR_REG_8__SCAN_IN
i P3_ADDR_REG_9__SCAN_IN
i P1_IR_REG_0__SCAN_IN
i P1_IR_REG_1__SCAN_IN
i P1_IR_REG_2__SCAN_IN
i P1_IR_REG_3__SCAN_IN
i P1_IR_REG_4__SCAN_IN
i P1_IR_REG_5__SCAN_IN
i P1_IR_REG_6__SCAN_IN
i P1_IR_REG_7__SCAN_IN
i P1_IR_REG_8__SCAN_IN
i P1_IR_REG_9__SCAN_IN
i P1_IR_REG_10__SCAN_IN
i P1_IR_REG_11__SCAN_IN
i P1_IR_REG_12__SCAN_IN
i P1_IR_REG_13__SCAN_IN
i P1_IR_REG_14__SCAN_IN
i P1_IR_REG_15__SCAN_IN
i P1_IR_REG_16__SCAN_IN
i P1_IR_REG_17__SCAN_IN
i P1_IR_REG_18__SCAN_IN
i P1_IR_REG_19__SCAN_IN
i P1_IR_REG_20__SCAN_IN
i P1_IR_REG_21__SCAN_IN
i P1_IR_REG_22__SCAN_IN
i P1_IR_REG_23__SCAN_IN
i P1_IR_REG_24__SCAN_IN
i P1_IR_REG_25__SCAN_IN
i P1_IR_REG_26__SCAN_IN
i P1_IR_REG_27__SCAN_IN
i P1_IR_REG_28__SCAN_IN
i P1_IR_REG_29__SCAN_IN
i P1_IR_REG_30__SCAN_IN
i P1_IR_REG_31__SCAN_IN
i P1_D_REG_0__SCAN_IN
i P1_D_REG_1__SCAN_IN
i P1_D_REG_2__SCAN_IN
i P1_D_REG_3__SCAN_IN
i P1_D_REG_4__SCAN_IN
i P1_D_REG_5__SCAN_IN
i P1_D_REG_6__SCAN_IN
i P1_D_REG_7__SCAN_IN
i P1_D_REG_8__SCAN_IN
i P1_D_REG_9__SCAN_IN
i P1_D_REG_10__SCAN_IN
i P1_D_REG_11__SCAN_IN
i P1_D_REG_12__SCAN_IN
i P1_D_REG_13__SCAN_IN
i P1_D_REG_14__SCAN_IN
i P1_D_REG_15__SCAN_IN
i P1_D_REG_16__SCAN_IN
i P1_D_REG_17__SCAN_IN
i P1_D_REG_18__SCAN_IN
i P1_D_REG_19__SCAN_IN
i P1_D_REG_20__SCAN_IN
i P1_D_REG_21__SCAN_IN
i P1_D_REG_22__SCAN_IN
i P1_D_REG_23__SCAN_IN
i P1_D_REG_24__SCAN_IN
i P1_D_REG_25__SCAN_IN
i P1_D_REG_26__SCAN_IN
i P1_D_REG_27__SCAN_IN
i P1_D_REG_28__SCAN_IN
i P1_D_REG_29__SCAN_IN
i P1_D_REG_30__SCAN_IN
i P1_D_REG_31__SCAN_IN
i P1_REG0_REG_0__SCAN_IN
i P1_REG0_REG_1__SCAN_IN
i P1_REG0_REG_2__SCAN_IN
i P1_REG0_REG_3__SCAN_IN
i P1_REG0_REG_4__SCAN_IN
i P1_REG0_REG_5__SCAN_IN
i P1_REG0_REG_6__SCAN_IN
i P1_REG0_REG_7__SCAN_IN
i P1_REG0_REG_8__SCAN_IN
i P1_REG0_REG_9__SCAN_IN
i P1_REG0_REG_10__SCAN_IN
i P1_REG0_REG_11__SCAN_IN
i P1_REG0_REG_12__SCAN_IN
i P1_REG0_REG_13__SCAN_IN
i P1_REG0_REG_14__SCAN_IN
i P1_REG0_REG_15__SCAN_IN
i P1_REG0_REG_16__SCAN_IN
i P1_REG0_REG_17__SCAN_IN
i P1_REG0_REG_18__SCAN_IN
i P1_REG0_REG_19__SCAN_IN
i P1_REG0_REG_20__SCAN_IN
i P1_REG0_REG_21__SCAN_IN
i P1_REG0_REG_22__SCAN_IN
i P1_REG0_REG_23__SCAN_IN
i P1_REG0_REG_24__SCAN_IN
i P1_REG0_REG_25__SCAN_IN
i P1_REG0_REG_26__SCAN_IN
i P1_REG0_REG_27__SCAN_IN
i P1_REG0_REG_28__SCAN_IN
i P1_REG0_REG_29__SCAN_IN
i P1_REG0_REG_30__SCAN_IN
i P1_REG0_REG_31__SCAN_IN
i P1_REG1_REG_0__SCAN_IN
i P1_REG1_REG_1__SCAN_IN
i P1_REG1_REG_2__SCAN_IN
i P1_REG1_REG_3__SCAN_IN
i P1_REG1_REG_4__SCAN_IN
i P1_REG1_REG_5__SCAN_IN
i P1_REG1_REG_6__SCAN_IN
i P1_REG1_REG_7__SCAN_IN
i P1_REG1_REG_8__SCAN_IN
i P1_REG1_REG_9__SCAN_IN
i P1_REG1_REG_10__SCAN_IN
i P1_REG1_REG_11__SCAN_IN
i P1_REG1_REG_12__SCAN_IN
i P1_REG1_REG_13__SCAN_IN
i P1_REG1_REG_14__SCAN_IN
i P1_REG1_REG_15__SCAN_IN
i P1_REG1_REG_16__SCAN_IN
i P1_REG1_REG_17__SCAN_IN
i P1_REG1_REG_18__SCAN_IN
i P1_REG1_REG_19__SCAN_IN
i P1_REG1_REG_20__SCAN_IN
i P1_REG1_REG_21__SCAN_IN
i P1_REG1_REG_22__SCAN_IN
i P1_REG1_REG_23__SCAN_IN
i P1_REG1_REG_24__SCAN_IN
i P1_REG1_REG_25__SCAN_IN
i P1_REG1_REG_26__SCAN_IN
i P1_REG1_REG_27__SCAN_IN
i P1_REG1_REG_28__SCAN_IN
i P1_REG1_REG_29__SCAN_IN
i P1_REG1_REG_30__SCAN_IN
i P1_REG1_REG_31__SCAN_IN
i P1_REG2_REG_0__SCAN_IN
i P1_REG2_REG_1__SCAN_IN
i P1_REG2_REG_2__SCAN_IN
i P1_REG2_REG_3__SCAN_IN
i P1_REG2_REG_4__SCAN_IN
i P1_REG2_REG_5__SCAN_IN
i P1_REG2_REG_6__SCAN_IN
i P1_REG2_REG_7__SCAN_IN
i P1_REG2_REG_8__SCAN_IN
i P1_REG2_REG_9__SCAN_IN
i P1_REG2_REG_10__SCAN_IN
i P1_REG2_REG_11__SCAN_IN
i P1_REG2_REG_12__SCAN_IN
i P1_REG2_REG_13__SCAN_IN
i P1_REG2_REG_14__SCAN_IN
i P1_REG2_REG_15__SCAN_IN
i P1_REG2_REG_16__SCAN_IN
i P1_REG2_REG_17__SCAN_IN
i P1_REG2_REG_18__SCAN_IN
i P1_REG2_REG_19__SCAN_IN
i P1_REG2_REG_20__SCAN_IN
i P1_REG2_REG_21__SCAN_IN
i P1_REG2_REG_22__SCAN_IN
i P1_REG2_REG_23__SCAN_IN
i P1_REG2_REG_24__SCAN_IN
i P1_REG2_REG_25__SCAN_IN
i P1_REG2_REG_26__SCAN_IN
i P1_REG2_REG_27__SCAN_IN
i P1_REG2_REG_28__SCAN_IN
i P1_REG2_REG_29__SCAN_IN
i P1_REG2_REG_30__SCAN_IN
i P1_REG2_REG_31__SCAN_IN
i P1_ADDR_REG_19__SCAN_IN
i P1_ADDR_REG_18__SCAN_IN
i P1_ADDR_REG_17__SCAN_IN
i P1_ADDR_REG_16__SCAN_IN
i P1_ADDR_REG_15__SCAN_IN
i P1_ADDR_REG_14__SCAN_IN
i P1_ADDR_REG_13__SCAN_IN
i P1_ADDR_REG_12__SCAN_IN
i P1_ADDR_REG_11__SCAN_IN
i P1_ADDR_REG_10__SCAN_IN
i P1_ADDR_REG_9__SCAN_IN
i P1_ADDR_REG_8__SCAN_IN
i P1_ADDR_REG_7__SCAN_IN
i P1_ADDR_REG_6__SCAN_IN
i P1_ADDR_REG_5__SCAN_IN
i P1_ADDR_REG_4__SCAN_IN
i P1_ADDR_REG_3__SCAN_IN
i P1_ADDR_REG_2__SCAN_IN
i P1_ADDR_REG_1__SCAN_IN
i P1_ADDR_REG_0__SCAN_IN
i P1_DATAO_REG_0__SCAN_IN
i P1_DATAO_REG_1__SCAN_IN
i P1_DATAO_REG_2__SCAN_IN
i P1_DATAO_REG_3__SCAN_IN
i P1_DATAO_REG_4__SCAN_IN
i P1_DATAO_REG_5__SCAN_IN
i P1_DATAO_REG_6__SCAN_IN
i P1_DATAO_REG_7__SCAN_IN
i P1_DATAO_REG_8__SCAN_IN
i P1_DATAO_REG_9__SCAN_IN
i P1_DATAO_REG_10__SCAN_IN
i P1_DATAO_REG_11__SCAN_IN
i P1_DATAO_REG_12__SCAN_IN
i P1_DATAO_REG_13__SCAN_IN
i P1_DATAO_REG_14__SCAN_IN
i P1_DATAO_REG_15__SCAN_IN
i P1_DATAO_REG_16__SCAN_IN
i P1_DATAO_REG_17__SCAN_IN
i P1_DATAO_REG_18__SCAN_IN
i P1_DATAO_REG_19__SCAN_IN
i P1_DATAO_REG_20__SCAN_IN
i P1_DATAO_REG_21__SCAN_IN
i P1_DATAO_REG_22__SCAN_IN
i P1_DATAO_REG_23__SCAN_IN
i P1_DATAO_REG_24__SCAN_IN
i P1_DATAO_REG_25__SCAN_IN
i P1_DATAO_REG_26__SCAN_IN
i P1_DATAO_REG_27__SCAN_IN
i P1_DATAO_REG_28__SCAN_IN
i P1_DATAO_REG_29__SCAN_IN
i P1_DATAO_REG_30__SCAN_IN
i P1_DATAO_REG_31__SCAN_IN
i P1_B_REG_SCAN_IN
i P1_REG3_REG_15__SCAN_IN
i P1_REG3_REG_26__SCAN_IN
i P1_REG3_REG_6__SCAN_IN
i P1_REG3_REG_18__SCAN_IN
i P1_REG3_REG_2__SCAN_IN
i P1_REG3_REG_11__SCAN_IN
i P1_REG3_REG_22__SCAN_IN
i P1_REG3_REG_13__SCAN_IN
i P1_REG3_REG_20__SCAN_IN
i P1_REG3_REG_0__SCAN_IN
i P1_REG3_REG_9__SCAN_IN
i P1_REG3_REG_4__SCAN_IN
i P1_REG3_REG_24__SCAN_IN
i P1_REG3_REG_17__SCAN_IN
i P1_REG3_REG_5__SCAN_IN
i P1_REG3_REG_16__SCAN_IN
i P1_REG3_REG_25__SCAN_IN
i P1_REG3_REG_12__SCAN_IN
i P1_REG3_REG_21__SCAN_IN
i P1_REG3_REG_1__SCAN_IN
i P1_REG3_REG_8__SCAN_IN
i P1_REG3_REG_28__SCAN_IN
i P1_REG3_REG_19__SCAN_IN
i P1_REG3_REG_3__SCAN_IN
i P1_REG3_REG_10__SCAN_IN
i P1_REG3_REG_23__SCAN_IN
i P1_REG3_REG_14__SCAN_IN
i P1_REG3_REG_27__SCAN_IN
i P1_REG3_REG_7__SCAN_IN
i P1_STATE_REG_SCAN_IN
i P1_RD_REG_SCAN_IN
i P1_WR_REG_SCAN_IN
i P2_IR_REG_0__SCAN_IN
i P2_IR_REG_1__SCAN_IN
i P2_IR_REG_2__SCAN_IN
i P2_IR_REG_3__SCAN_IN
i P2_IR_REG_4__SCAN_IN
i P2_IR_REG_5__SCAN_IN
i P2_IR_REG_6__SCAN_IN
i P2_IR_REG_7__SCAN_IN
i P2_IR_REG_8__SCAN_IN
i P2_IR_REG_9__SCAN_IN
i P2_IR_REG_10__SCAN_IN
i P2_IR_REG_11__SCAN_IN
i P2_IR_REG_12__SCAN_IN
i P2_IR_REG_13__SCAN_IN
i P2_IR_REG_14__SCAN_IN
i P2_IR_REG_15__SCAN_IN
i P2_IR_REG_16__SCAN_IN
i P2_IR_REG_17__SCAN_IN
i P2_IR_REG_18__SCAN_IN
i P2_IR_REG_19__SCAN_IN
i P2_IR_REG_20__SCAN_IN
i P2_IR_REG_21__SCAN_IN
i P2_IR_REG_22__SCAN_IN
i P2_IR_REG_23__SCAN_IN
i P2_IR_REG_24__SCAN_IN
i P2_IR_REG_25__SCAN_IN
i P2_IR_REG_26__SCAN_IN
i P2_IR_REG_27__SCAN_IN
i P2_IR_REG_28__SCAN_IN
i P2_IR_REG_29__SCAN_IN
i P2_IR_REG_30__SCAN_IN
i P2_IR_REG_31__SCAN_IN
i P2_D_REG_0__SCAN_IN
i P2_D_REG_1__SCAN_IN
i P2_D_REG_2__SCAN_IN
i P2_D_REG_3__SCAN_IN
i P2_D_REG_4__SCAN_IN
i P2_D_REG_5__SCAN_IN
i P2_D_REG_6__SCAN_IN
i P2_D_REG_7__SCAN_IN
i P2_D_REG_8__SCAN_IN
i P2_D_REG_9__SCAN_IN
i P2_D_REG_10__SCAN_IN
i P2_D_REG_11__SCAN_IN
i P2_D_REG_12__SCAN_IN
i P2_D_REG_13__SCAN_IN
i P2_D_REG_14__SCAN_IN
i P2_D_REG_15__SCAN_IN
i P2_D_REG_16__SCAN_IN
i P2_D_REG_17__SCAN_IN
i P2_D_REG_18__SCAN_IN
i P2_D_REG_19__SCAN_IN
i P2_D_REG_20__SCAN_IN
i P2_D_REG_21__SCAN_IN
i P2_D_REG_22__SCAN_IN
i P2_D_REG_23__SCAN_IN
i P2_D_REG_24__SCAN_IN
i P2_D_REG_25__SCAN_IN
i P2_D_REG_26__SCAN_IN
i P2_D_REG_27__SCAN_IN
i P2_D_REG_28__SCAN_IN
i P2_D_REG_29__SCAN_IN
i P2_D_REG_30__SCAN_IN
i P2_D_REG_31__SCAN_IN
i P2_REG0_REG_0__SCAN_IN
i P2_REG0_REG_1__SCAN_IN
i P2_REG0_REG_2__SCAN_IN
i P2_REG0_REG_3__SCAN_IN
i P2_REG0_REG_4__SCAN_IN
i P2_REG0_REG_5__SCAN_IN
i P2_REG0_REG_6__SCAN_IN
i P2_REG0_REG_7__SCAN_IN
i P2_REG0_REG_8__SCAN_IN
i P2_REG0_REG_9__SCAN_IN
i P2_REG0_REG_10__SCAN_IN
i P2_REG0_REG_11__SCAN_IN
i P2_REG0_REG_12__SCAN_IN
i P2_REG0_REG_13__SCAN_IN
i P2_REG0_REG_14__SCAN_IN
i P2_REG0_REG_15__SCAN_IN
i P2_REG0_REG_16__SCAN_IN
i P2_REG0_REG_17__SCAN_IN
i P2_REG0_REG_18__SCAN_IN
i P2_REG0_REG_19__SCAN_IN
i P2_REG0_REG_20__SCAN_IN
i P2_REG0_REG_21__SCAN_IN
i P2_REG0_REG_22__SCAN_IN
i P2_REG0_REG_23__SCAN_IN
i P2_REG0_REG_24__SCAN_IN
i P2_REG0_REG_25__SCAN_IN
i P2_REG0_REG_26__SCAN_IN
i P2_REG0_REG_27__SCAN_IN
i P2_REG0_REG_28__SCAN_IN
i P2_REG0_REG_29__SCAN_IN
i P2_REG0_REG_30__SCAN_IN
i P2_REG0_REG_31__SCAN_IN
i P2_REG1_REG_0__SCAN_IN
i P2_REG1_REG_1__SCAN_IN
i P2_REG1_REG_2__SCAN_IN
i P2_REG1_REG_3__SCAN_IN
i P2_REG1_REG_4__SCAN_IN
i P2_REG1_REG_5__SCAN_IN
i P2_REG1_REG_6__SCAN_IN
i P2_REG1_REG_7__SCAN_IN
i P2_REG1_REG_8__SCAN_IN
i P2_REG1_REG_9__SCAN_IN
i P2_REG1_REG_10__SCAN_IN
i P2_REG1_REG_11__SCAN_IN
i P2_REG1_REG_12__SCAN_IN
i P2_REG1_REG_13__SCAN_IN
i P2_REG1_REG_14__SCAN_IN
i P2_REG1_REG_15__SCAN_IN
i P2_REG1_REG_16__SCAN_IN
i P2_REG1_REG_17__SCAN_IN
i P2_REG1_REG_18__SCAN_IN
i P2_REG1_REG_19__SCAN_IN
i P2_REG1_REG_20__SCAN_IN
i P2_REG1_REG_21__SCAN_IN
i P2_REG1_REG_22__SCAN_IN
i P2_REG1_REG_23__SCAN_IN
i P2_REG1_REG_24__SCAN_IN
i P2_REG1_REG_25__SCAN_IN
i P2_REG1_REG_26__SCAN_IN
i P2_REG1_REG_27__SCAN_IN
i P2_REG1_REG_28__SCAN_IN
i P2_REG1_REG_29__SCAN_IN
i P2_REG1_REG_30__SCAN_IN
i P2_REG1_REG_31__SCAN_IN
i P2_REG2_REG_0__SCAN_IN
i P2_REG2_REG_1__SCAN_IN
i P2_REG2_REG_2__SCAN_IN
i P2_REG2_REG_3__SCAN_IN
i P2_REG2_REG_4__SCAN_IN
i P2_REG2_REG_5__SCAN_IN
i P2_REG2_REG_6__SCAN_IN
i P2_REG2_REG_7__SCAN_IN
i P2_REG2_REG_8__SCAN_IN
i P2_REG2_REG_9__SCAN_IN
i P2_REG2_REG_10__SCAN_IN
i P2_REG2_REG_11__SCAN_IN
i P2_REG2_REG_12__SCAN_IN
i P2_REG2_REG_13__SCAN_IN
i P2_REG2_REG_14__SCAN_IN
i P2_REG2_REG_15__SCAN_IN
i P2_REG2_REG_16__SCAN_IN
i P2_REG2_REG_17__SCAN_IN
i P2_REG2_REG_18__SCAN_IN
i P2_REG2_REG_19__SCAN_IN
i P2_REG2_REG_20__SCAN_IN
i P2_REG2_REG_21__SCAN_IN
i P2_REG2_REG_22__SCAN_IN
i P2_REG2_REG_23__SCAN_IN
i P2_REG2_REG_24__SCAN_IN
i P2_REG2_REG_25__SCAN_IN
i P2_REG2_REG_26__SCAN_IN
i P2_REG2_REG_27__SCAN_IN
i P2_REG2_REG_28__SCAN_IN
i P2_REG2_REG_29__SCAN_IN
i P2_REG2_REG_30__SCAN_IN
i P2_REG2_REG_31__SCAN_IN
i P2_ADDR_REG_19__SCAN_IN
i P2_ADDR_REG_18__SCAN_IN
i P2_ADDR_REG_17__SCAN_IN
i P2_ADDR_REG_16__SCAN_IN
i P2_ADDR_REG_15__SCAN_IN
i P2_ADDR_REG_14__SCAN_IN
i P2_ADDR_REG_13__SCAN_IN
i P2_ADDR_REG_12__SCAN_IN
i P2_ADDR_REG_11__SCAN_IN
i P2_ADDR_REG_10__SCAN_IN
i P2_ADDR_REG_9__SCAN_IN
i P2_ADDR_REG_8__SCAN_IN
i P2_ADDR_REG_7__SCAN_IN
i P2_ADDR_REG_6__SCAN_IN
i P2_ADDR_REG_5__SCAN_IN
i P2_ADDR_REG_4__SCAN_IN
i P2_ADDR_REG_3__SCAN_IN
i P2_ADDR_REG_2__SCAN_IN
i P2_ADDR_REG_1__SCAN_IN
i P2_ADDR_REG_0__SCAN_IN
i P2_DATAO_REG_0__SCAN_IN
i P2_DATAO_REG_1__SCAN_IN
i P2_DATAO_REG_2__SCAN_IN
i P2_DATAO_REG_3__SCAN_IN
i P2_DATAO_REG_4__SCAN_IN
i P2_DATAO_REG_5__SCAN_IN
i P2_DATAO_REG_6__SCAN_IN
i P2_DATAO_REG_7__SCAN_IN
i P2_DATAO_REG_8__SCAN_IN
i P2_DATAO_REG_9__SCAN_IN
i P2_DATAO_REG_10__SCAN_IN
i P2_DATAO_REG_11__SCAN_IN
i P2_DATAO_REG_12__SCAN_IN
i P2_DATAO_REG_13__SCAN_IN
i P2_DATAO_REG_14__SCAN_IN
i P2_DATAO_REG_15__SCAN_IN
i P2_DATAO_REG_16__SCAN_IN
i P2_DATAO_REG_17__SCAN_IN
i P2_DATAO_REG_18__SCAN_IN
i P2_DATAO_REG_19__SCAN_IN
i P2_DATAO_REG_20__SCAN_IN
i P2_DATAO_REG_21__SCAN_IN
i P2_DATAO_REG_22__SCAN_IN
i P2_DATAO_REG_23__SCAN_IN
i P2_DATAO_REG_24__SCAN_IN
i P2_DATAO_REG_25__SCAN_IN
i P2_DATAO_REG_26__SCAN_IN
i P2_DATAO_REG_27__SCAN_IN
i P2_DATAO_REG_28__SCAN_IN
i P2_DATAO_REG_29__SCAN_IN
i P2_DATAO_REG_30__SCAN_IN
i P2_DATAO_REG_31__SCAN_IN
i P2_B_REG_SCAN_IN
i P2_REG3_REG_15__SCAN_IN
i P2_REG3_REG_26__SCAN_IN
i P2_REG3_REG_6__SCAN_IN
i P2_REG3_REG_18__SCAN_IN
i P2_REG3_REG_2__SCAN_IN
i P2_REG3_REG_11__SCAN_IN
i P2_REG3_REG_22__SCAN_IN
i P2_REG3_REG_13__SCAN_IN
i P2_REG3_REG_20__SCAN_IN
i P2_REG3_REG_0__SCAN_IN
i P2_REG3_REG_9__SCAN_IN
i P2_REG3_REG_4__SCAN_IN
i P2_REG3_REG_24__SCAN_IN
i P2_REG3_REG_17__SCAN_IN
i P2_REG3_REG_5__SCAN_IN
i P2_REG3_REG_16__SCAN_IN
i P2_REG3_REG_25__SCAN_IN
i P2_REG3_REG_12__SCAN_IN
i P2_REG3_REG_21__SCAN_IN
i P2_REG3_REG_1__SCAN_IN
i P2_REG3_REG_8__SCAN_IN
i P2_REG3_REG_28__SCAN_IN
i P2_REG3_REG_19__SCAN_IN
i P2_REG3_REG_3__SCAN_IN
i P2_REG3_REG_10__SCAN_IN
i P2_REG3_REG_23__SCAN_IN
i P2_REG3_REG_14__SCAN_IN
i P2_REG3_REG_27__SCAN_IN
i P2_REG3_REG_7__SCAN_IN
i P2_STATE_REG_SCAN_IN
i P2_RD_REG_SCAN_IN
i P2_WR_REG_SCAN_IN
i P3_IR_REG_0__SCAN_IN
i P3_IR_REG_1__SCAN_IN
i P3_IR_REG_2__SCAN_IN
i P3_IR_REG_3__SCAN_IN
i P3_IR_REG_4__SCAN_IN
i P3_IR_REG_5__SCAN_IN
i P3_IR_REG_6__SCAN_IN
i P3_IR_REG_7__SCAN_IN
i P3_IR_REG_8__SCAN_IN
i P3_IR_REG_9__SCAN_IN
i P3_IR_REG_10__SCAN_IN
i P3_IR_REG_11__SCAN_IN
i P3_IR_REG_12__SCAN_IN
i P3_IR_REG_13__SCAN_IN
i P3_IR_REG_14__SCAN_IN
i P3_IR_REG_15__SCAN_IN
i P3_IR_REG_16__SCAN_IN
i P3_IR_REG_17__SCAN_IN
i P3_IR_REG_18__SCAN_IN
i P3_IR_REG_19__SCAN_IN
i P3_IR_REG_20__SCAN_IN
i P3_IR_REG_21__SCAN_IN
i P3_IR_REG_22__SCAN_IN
i P3_IR_REG_23__SCAN_IN
i P3_IR_REG_24__SCAN_IN
i P3_IR_REG_25__SCAN_IN
i P3_IR_REG_26__SCAN_IN
i P3_IR_REG_27__SCAN_IN
i P3_IR_REG_28__SCAN_IN
i P3_IR_REG_29__SCAN_IN
i P3_IR_REG_30__SCAN_IN
i P3_IR_REG_31__SCAN_IN
i P3_D_REG_0__SCAN_IN
i P3_D_REG_1__SCAN_IN
i P3_D_REG_2__SCAN_IN
i P3_D_REG_3__SCAN_IN
i P3_D_REG_4__SCAN_IN
i P3_D_REG_5__SCAN_IN
i P3_D_REG_6__SCAN_IN
i P3_D_REG_7__SCAN_IN
i P3_D_REG_8__SCAN_IN
i P3_D_REG_9__SCAN_IN
i P3_D_REG_10__SCAN_IN
i P3_D_REG_11__SCAN_IN
i P3_D_REG_12__SCAN_IN
i P3_D_REG_13__SCAN_IN
i P3_D_REG_14__SCAN_IN
i P3_D_REG_15__SCAN_IN
i P3_D_REG_16__SCAN_IN
i P3_D_REG_17__SCAN_IN
i P3_D_REG_18__SCAN_IN
i P3_D_REG_19__SCAN_IN
i P3_D_REG_20__SCAN_IN
i P3_D_REG_21__SCAN_IN
i P3_D_REG_22__SCAN_IN
i P3_D_REG_23__SCAN_IN
i P3_D_REG_24__SCAN_IN
i P3_D_REG_25__SCAN_IN
i P3_D_REG_26__SCAN_IN
i P3_D_REG_27__SCAN_IN
i P3_D_REG_28__SCAN_IN
i P3_D_REG_29__SCAN_IN
i P3_D_REG_30__SCAN_IN
i P3_D_REG_31__SCAN_IN
i P3_REG0_REG_0__SCAN_IN
i P3_REG0_REG_1__SCAN_IN
i P3_REG0_REG_2__SCAN_IN
i P3_REG0_REG_3__SCAN_IN
i P3_REG0_REG_4__SCAN_IN
i P3_REG0_REG_5__SCAN_IN
i P3_REG0_REG_6__SCAN_IN
i P3_REG0_REG_7__SCAN_IN
i P3_REG0_REG_8__SCAN_IN
i P3_REG0_REG_9__SCAN_IN
i P3_REG0_REG_10__SCAN_IN
i P3_REG0_REG_11__SCAN_IN
i P3_REG0_REG_12__SCAN_IN
i P3_REG0_REG_13__SCAN_IN
i P3_REG0_REG_14__SCAN_IN
i P3_REG0_REG_15__SCAN_IN
i P3_REG0_REG_16__SCAN_IN
i P3_REG0_REG_17__SCAN_IN
i P3_REG0_REG_18__SCAN_IN
i P3_REG0_REG_19__SCAN_IN
i P3_REG0_REG_20__SCAN_IN
i P3_REG0_REG_21__SCAN_IN
i P3_REG0_REG_22__SCAN_IN
i P3_REG0_REG_23__SCAN_IN
i P3_REG0_REG_24__SCAN_IN
i P3_REG0_REG_25__SCAN_IN
i P3_REG0_REG_26__SCAN_IN
i P3_REG0_REG_27__SCAN_IN
i P3_REG0_REG_28__SCAN_IN
i P3_REG0_REG_29__SCAN_IN
i P3_REG0_REG_30__SCAN_IN
i P3_REG0_REG_31__SCAN_IN
i P3_REG1_REG_0__SCAN_IN
i P3_REG1_REG_1__SCAN_IN
i P3_REG1_REG_2__SCAN_IN
i P3_REG1_REG_3__SCAN_IN
i P3_REG1_REG_4__SCAN_IN
i P3_REG1_REG_5__SCAN_IN
i P3_REG1_REG_6__SCAN_IN
i P3_REG1_REG_7__SCAN_IN
i P3_REG1_REG_8__SCAN_IN
i P3_REG1_REG_9__SCAN_IN
i P3_REG1_REG_10__SCAN_IN
i P3_REG1_REG_11__SCAN_IN
i P3_REG1_REG_12__SCAN_IN
i P3_REG1_REG_13__SCAN_IN
i P3_REG1_REG_14__SCAN_IN
i P3_REG1_REG_15__SCAN_IN
i P3_REG1_REG_16__SCAN_IN
i P3_REG1_REG_17__SCAN_IN
i P3_REG1_REG_18__SCAN_IN
i P3_REG1_REG_19__SCAN_IN
i P3_REG1_REG_20__SCAN_IN
i P3_REG1_REG_21__SCAN_IN
i P3_REG1_REG_22__SCAN_IN
i P3_REG1_REG_23__SCAN_IN
i P3_REG1_REG_24__SCAN_IN
i P3_REG1_REG_25__SCAN_IN
i P3_REG1_REG_26__SCAN_IN
i P3_REG1_REG_27__SCAN_IN
i P3_REG1_REG_28__SCAN_IN
i P3_REG1_REG_29__SCAN_IN
i P3_REG1_REG_30__SCAN_IN
i P3_REG1_REG_31__SCAN_IN
i P3_REG2_REG_0__SCAN_IN
i P3_REG2_REG_1__SCAN_IN
i P3_REG2_REG_2__SCAN_IN
i P3_REG2_REG_3__SCAN_IN
i P3_REG2_REG_4__SCAN_IN
i P3_REG2_REG_5__SCAN_IN
i P3_REG2_REG_6__SCAN_IN
i P3_REG2_REG_7__SCAN_IN
i P3_REG2_REG_8__SCAN_IN
i P3_REG2_REG_9__SCAN_IN
i P3_REG2_REG_10__SCAN_IN
i P3_REG2_REG_11__SCAN_IN
i P3_REG2_REG_12__SCAN_IN
i P3_REG2_REG_13__SCAN_IN
i P3_REG2_REG_14__SCAN_IN
i P3_REG2_REG_15__SCAN_IN
i P3_REG2_REG_16__SCAN_IN
i P3_REG2_REG_17__SCAN_IN
i P3_REG2_REG_18__SCAN_IN
i P3_REG2_REG_19__SCAN_IN
i P3_REG2_REG_20__SCAN_IN
i P3_REG2_REG_21__SCAN_IN
i P3_REG2_REG_22__SCAN_IN
i P3_REG2_REG_23__SCAN_IN
i P3_REG2_REG_24__SCAN_IN
i P3_REG2_REG_25__SCAN_IN
i P3_REG2_REG_26__SCAN_IN
i P3_REG2_REG_27__SCAN_IN
i P3_REG2_REG_28__SCAN_IN
i P3_REG2_REG_29__SCAN_IN
i P3_REG2_REG_30__SCAN_IN
i P3_REG2_REG_31__SCAN_IN
i P3_ADDR_REG_19__SCAN_IN
i P3_ADDR_REG_18__SCAN_IN
i P3_ADDR_REG_17__SCAN_IN
i P3_ADDR_REG_16__SCAN_IN
i P3_ADDR_REG_15__SCAN_IN
i P3_ADDR_REG_14__SCAN_IN
i P3_ADDR_REG_13__SCAN_IN
i P3_ADDR_REG_12__SCAN_IN
i P3_ADDR_REG_11__SCAN_IN
i P3_ADDR_REG_10__SCAN_IN
o SUB_1596_U4
o SUB_1596_U62
o SUB_1596_U63
o SUB_1596_U64
o SUB_1596_U65
o SUB_1596_U66
o SUB_1596_U67
o SUB_1596_U68
o SUB_1596_U69
o SUB_1596_U70
o SUB_1596_U54
o SUB_1596_U55
o SUB_1596_U56
o SUB_1596_U57
o SUB_1596_U58
o SUB_1596_U59
o SUB_1596_U60
o SUB_1596_U61
o SUB_1596_U5
o SUB_1596_U53
o U29
o U28
o P1_U3355
o P1_U3354
o P1_U3353
o P1_U3352
o P1_U3351
o P1_U3350
o P1_U3349
o P1_U3348
o P1_U3347
o P1_U3346
o P1_U3345
o P1_U3344
o P1_U3343
o P1_U3342
o P1_U3341
o P1_U3340
o P1_U3339
o P1_U3338
o P1_U3337
o P1_U3336
o P1_U3335
o P1_U3334
o P1_U3333
o P1_U3332
o P1_U3331
o P1_U3330
o P1_U3329
o P1_U3328
o P1_U3327
o P1_U3326
o P1_U3325
o P1_U3324
o P1_U3445
o P1_U3446
o P1_U3323
o P1_U3322
o P1_U3321
o P1_U3320
o P1_U3319
o P1_U3318
o P1_U3317
o P1_U3316
o P1_U3315
o P1_U3314
o P1_U3313
o P1_U3312
o P1_U3311
o P1_U3310
o P1_U3309
o P1_U3308
o P1_U3307
o P1_U3306
o P1_U3305
o P1_U3304
o P1_U3303
o P1_U3302
o P1_U3301
o P1_U3300
o P1_U3299
o P1_U3298
o P1_U3297
o P1_U3296
o P1_U3295
o P1_U3294
o P1_U3459
o P1_U3462
o P1_U3465
o P1_U3468
o P1_U3471
o P1_U3474
o P1_U3477
o P1_U3480
o P1_U3483
o P1_U3486
o P1_U3489
o P1_U3492
o P1_U3495
o P1_U3498
o P1_U3501
o P1_U3504
o P1_U3507
o P1_U3510
o P1_U3513
o P1_U3515
o P1_U3516
o P1_U3517
o P1_U3518
o P1_U3519
o P1_U3520
o P1_U3521
o P1_U3522
o P1_U3523
o P1_U3524
o P1_U3525
o P1_U3526
o P1_U3527
o P1_U3528
o P1_U3529
o P1_U3530
o P1_U3531
o P1_U3532
o P1_U3533
o P1_U3534
o P1_U3535
o P1_U3536
o P1_U3537
o P1_U3538
o P1_U3539
o P1_U3540
o P1_U3541
o P1_U3542
o P1_U3543
o P1_U3544
o P1_U3545
o P1_U3546
o P1_U3547
o P1_U3548
o P1_U3549
o P1_U3550
o P1_U3551
o P1_U3552
o P1_U3553
o P1_U3554
o P1_U3555
o P1_U3556
o P1_U3557
o P1_U3558
o P1_U3559
o P1_U3293
o P1_U3292
o P1_U3291
o P1_U3290
o P1_U3289
o P1_U3288
o P1_U3287
o P1_U3286
o P1_U3285
o P1_U3284
o P1_U3283
o P1_U3282
o P1_U3281
o P1_U3280
o P1_U3279
o P1_U3278
o P1_U3277
o P1_U3276
o P1_U3275
o P1_U3274
o P1_U3273
o P1_U3272
o P1_U3271
o P1_U3270
o P1_U3269
o P1_U3268
o P1_U3267
o P1_U3266
o P1_U3265
o P1_U3356
o P1_U3264
o P1_U3263
o P1_U3262
o P1_U3261
o P1_U3260
o P1_U3259
o P1_U3258
o P1_U3257
o P1_U3256
o P1_U3255
o P1_U3254
o P1_U3253
o P1_U3252
o P1_U3251
o P1_U3250
o P1_U3249
o P1_U3248
o P1_U3247
o P1_U3246
o P1_U3245
o P1_U3244
o P1_U3243
o P1_U3560
o P1_U3561
o P1_U3562
o P1_U3563
o P1_U3564
o P1_U3565
o P1_U3566
o P1_U3567
o P1_U3568
o P1_U3569
o P1_U3570
o P1_U3571
o P1_U3572
o P1_U3573
o P1_U3574
o P1_U3575
o P1_U3576
o P1_U3577
o P1_U3578
o P1_U3579
o P1_U3580
o P1_U3581
o P1_U3582
o P1_U3583
o P1_U3584
o P1_U3585
o P1_U3586
o P1_U3587
o P1_U3588
o P1_U3589
o P1_U3590
o P1_U3591
o P1_U3242
o P1_U3241
o P1_U3240
o P1_U3239
o P1_U3238
o P1_U3237
o P1_U3236
o P1_U3235
o P1_U3234
o P1_U3233
o P1_U3232
o P1_U3231
o P1_U3230
o P1_U3229
o P1_U3228
o P1_U3227
o P1_U3226
o P1_U3225
o P1_U3224
o P1_U3223
o P1_U3222
o P1_U3221
o P1_U3220
o P1_U3219
o P1_U3218
o P1_U3217
o P1_U3216
o P1_U3215
o P1_U3214
o P1_U3213
o P1_U3086
o P1_U3085
o P1_U4016
o P2_U3327
o P2_U3326
o P2_U3325
o P2_U3324
o P2_U3323
o P2_U3322
o P2_U3321
o P2_U3320
o P2_U3319
o P2_U3318
o P2_U3317
o P2_U3316
o P2_U3315
o P2_U3314
o P2_U3313
o P2_U3312
o P2_U3311
o P2_U3310
o P2_U3309
o P2_U3308
o P2_U3307
o P2_U3306
o P2_U3305
o P2_U3304
o P2_U3303
o P2_U3302
o P2_U3301
o P2_U3300
o P2_U3299
o P2_U3298
o P2_U3297
o P2_U3296
o P2_U3416
o P2_U3417
o P2_U3295
o P2_U3294
o P2_U3293
o P2_U3292
o P2_U3291
o P2_U3290
o P2_U3289
o P2_U3288
o P2_U3287
o P2_U3286
o P2_U3285
o P2_U3284
o P2_U3283
o P2_U3282
o P2_U3281
o P2_U3280
o P2_U3279
o P2_U3278
o P2_U3277
o P2_U3276
o P2_U3275
o P2_U3274
o P2_U3273
o P2_U3272
o P2_U3271
o P2_U3270
o P2_U3269
o P2_U3268
o P2_U3267
o P2_U3266
o P2_U3430
o P2_U3433
o P2_U3436
o P2_U3439
o P2_U3442
o P2_U3445
o P2_U3448
o P2_U3451
o P2_U3454
o P2_U3457
o P2_U3460
o P2_U3463
o P2_U3466
o P2_U3469
o P2_U3472
o P2_U3475
o P2_U3478
o P2_U3481
o P2_U3484
o P2_U3486
o P2_U3487
o P2_U3488
o P2_U3489
o P2_U3490
o P2_U3491
o P2_U3492
o P2_U3493
o P2_U3494
o P2_U3495
o P2_U3496
o P2_U3497
o P2_U3498
o P2_U3499
o P2_U3500
o P2_U3501
o P2_U3502
o P2_U3503
o P2_U3504
o P2_U3505
o P2_U3506
o P2_U3507
o P2_U3508
o P2_U3509
o P2_U3510
o P2_U3511
o P2_U3512
o P2_U3513
o P2_U3514
o P2_U3515
o P2_U3516
o P2_U3517
o P2_U3518
o P2_U3519
o P2_U3520
o P2_U3521
o P2_U3522
o P2_U3523
o P2_U3524
o P2_U3525
o P2_U3526
o P2_U3527
o P2_U3528
o P2_U3529
o P2_U3530
o P2_U3265
o P2_U3264
o P2_U3263
o P2_U3262
o P2_U3261
o P2_U3260
o P2_U3259
o P2_U3258
o P2_U3257
o P2_U3256
o P2_U3255
o P2_U3254
o P2_U3253
o P2_U3252
o P2_U3251
o P2_U3250
o P2_U3249
o P2_U3248
o P2_U3247
o P2_U3246
o P2_U3245
o P2_U3244
o P2_U3243
o P2_U3242
o P2_U3241
o P2_U3240
o P2_U3239
o P2_U3238
o P2_U3237
o P2_U3236
o P2_U3235
o P2_U3234
o P2_U3233
o P2_U3232
o P2_U3231
o P2_U3230
o P2_U3229
o P2_U3228
o P2_U3227
o P2_U3226
o P2_U3225
o P2_U3224
o P2_U3223
o P2_U3222
o P2_U3221
o P2_U3220
o P2_U3219
o P2_U3218
o P2_U3217
o P2_U3216
o P2_U3215
o P2_U3214
o P2_U3531
o P2_U3532
o P2_U3533
o P2_U3534
o P2_U3535
o P2_U3536
o P2_U3537
o P2_U3538
o P2_U3539
o P2_U3540
o P2_U3541
o P2_U3542
o P2_U3543
o P2_U3544
o P2_U3545
o P2_U3546
o P2_U3547
o P2_U3548
o P2_U3549
o P2_U3550
o P2_U3551
o P2_U3552
o P2_U3553
o P2_U3554
o P2_U3555
o P2_U3556
o P2_U3557
o P2_U3558
o P2_U3559
o P2_U3560
o P2_U3561
o P2_U3562
o P2_U3328
o P2_U3213
o P2_U3212
o P2_U3211
o P2_U3210
o P2_U3209
o P2_U3208
o P2_U3207
o P2_U3206
o P2_U3205
o P2_U3204
o P2_U3203
o P2_U3202
o P2_U3201
o P2_U3200
o P2_U3199
o P2_U3198
o P2_U3197
o P2_U3196
o P2_U3195
o P2_U3194
o P2_U3193
o P2_U3192
o P2_U3191
o P2_U3190
o P2_U3189
o P2_U3188
o P2_U3187
o P2_U3186
o P2_U3185
o P2_U3088
o P2_U3087
o P2_U3947
o P3_U3295
o P3_U3294
o P3_U3293
o P3_U3292
o P3_U3291
o P3_U3290
o P3_U3289
o P3_U3288
o P3_U3287
o P3_U3286
o P3_U3285
o P3_U3284
o P3_U3283
o P3_U3282
o P3_U3281
o P3_U3280
o P3_U3279
o P3_U3278
o P3_U3277
o P3_U3276
o P3_U3275
o P3_U3274
o P3_U3273
o P3_U3272
o P3_U3271
o P3_U3270
o P3_U3269
o P3_U3268
o P3_U3267
o P3_U3266
o P3_U3265
o P3_U3264
o P3_U3376
o P3_U3377
o P3_U3263
o P3_U3262
o P3_U3261
o P3_U3260
o P3_U3259
o P3_U3258
o P3_U3257
o P3_U3256
o P3_U3255
o P3_U3254
o P3_U3253
o P3_U3252
o P3_U3251
o P3_U3250
o P3_U3249
o P3_U3248
o P3_U3247
o P3_U3246
o P3_U3245
o P3_U3244
o P3_U3243
o P3_U3242
o P3_U3241
o P3_U3240
o P3_U3239
o P3_U3238
o P3_U3237
o P3_U3236
o P3_U3235
o P3_U3234
o P3_U3390
o P3_U3393
o P3_U3396
o P3_U3399
o P3_U3402
o P3_U3405
o P3_U3408
o P3_U3411
o P3_U3414
o P3_U3417
o P3_U3420
o P3_U3423
o P3_U3426
o P3_U3429
o P3_U3432
o P3_U3435
o P3_U3438
o P3_U3441
o P3_U3444
o P3_U3446
o P3_U3447
o P3_U3448
o P3_U3449
o P3_U3450
o P3_U3451
o P3_U3452
o P3_U3453
o P3_U3454
o P3_U3455
o P3_U3456
o P3_U3457
o P3_U3458
o P3_U3459
o P3_U3460
o P3_U3461
o P3_U3462
o P3_U3463
o P3_U3464
o P3_U3465
o P3_U3466
o P3_U3467
o P3_U3468
o P3_U3469
o P3_U3470
o P3_U3471
o P3_U3472
o P3_U3473
o P3_U3474
o P3_U3475
o P3_U3476
o P3_U3477
o P3_U3478
o P3_U3479
o P3_U3480
o P3_U3481
o P3_U3482
o P3_U3483
o P3_U3484
o P3_U3485
o P3_U3486
o P3_U3487
o P3_U3488
o P3_U3489
o P3_U3490
o P3_U3233
o P3_U3232
o P3_U3231
o P3_U3230
o P3_U3229
o P3_U3228
o P3_U3227
o P3_U3226
o P3_U3225
o P3_U3224
o P3_U3223
o P3_U3222
o P3_U3221
o P3_U3220
o P3_U3219
o P3_U3218
o P3_U3217
o P3_U3216
o P3_U3215
o P3_U3214
o P3_U3213
o P3_U3212
o P3_U3211
o P3_U3210
o P3_U3209
o P3_U3208
o P3_U3207
o P3_U3206
o P3_U3205
o P3_U3204
o P3_U3203
o P3_U3202
o P3_U3201
o P3_U3200
o P3_U3199
o P3_U3198
o P3_U3197
o P3_U3196
o P3_U3195
o P3_U3194
o P3_U3193
o P3_U3192
o P3_U3191
o P3_U3190
o P3_U3189
o P3_U3188
o P3_U3187
o P3_U3186
o P3_U3185
o P3_U3184
o P3_U3183
o P3_U3182
o P3_U3491
o P3_U3492
o P3_U3493
o P3_U3494
o P3_U3495
o P3_U3496
o P3_U3497
o P3_U3498
o P3_U3499
o P3_U3500
o P3_U3501
o P3_U3502
o P3_U3503
o P3_U3504
o P3_U3505
o P3_U3506
o P3_U3507
o P3_U3508
o P3_U3509
o P3_U3510
o P3_U3511
o P3_U3512
o P3_U3513
o P3_U3514
o P3_U3515
o P3_U3516
o P3_U3517
o P3_U3518
o P3_U3519
o P3_U3520
o P3_U3521
o P3_U3522
o P3_U3296
o P3_U3181
o P3_U3180
o P3_U3179
o P3_U3178
o P3_U3177
o P3_U3176
o P3_U3175
o P3_U3174
o P3_U3173
o P3_U3172
o P3_U3171
o P3_U3170
o P3_U3169
o P3_U3168
o P3_U3167
o P3_U3166
o P3_U3165
o P3_U3164
o P3_U3163
o P3_U3162
o P3_U3161
o P3_U3160
o P3_U3159
o P3_U3158
o P3_U3157
o P3_U3156
o P3_U3155
o P3_U3154
o P3_U3153
o P3_U3151
o P3_U3150
o P3_U3897
g1 or U160 P3_WR_REG_SCAN_IN ; U28
g2 or U163 P3_RD_REG_SCAN_IN ; U29
g3 nand U173 U172 ; U30
g4 nand U175 U174 ; U31
g5 nand U177 U176 ; U32
g6 nand U179 U178 ; U33
g7 nand U181 U180 ; U34
g8 nand U183 U182 ; U35
g9 nand U185 U184 ; U36
g10 nand U187 U186 ; U37
g11 nand U189 U188 ; U38
g12 nand U191 U190 ; U39
g13 nand U193 U192 ; U40
g14 nand U195 U194 ; U41
g15 nand U197 U196 ; U42
g16 nand U199 U198 ; U43
g17 nand U201 U200 ; U44
g18 nand U203 U202 ; U45
g19 nand U205 U204 ; U46
g20 nand U207 U206 ; U47
g21 nand U209 U208 ; U48
g22 nand U211 U210 ; U49
g23 nand U213 U212 ; U50
g24 nand U215 U214 ; U51
g25 nand U217 U216 ; U52
g26 nand U219 U218 ; U53
g27 nand U221 U220 ; U54
g28 nand U223 U222 ; U55
g29 nand U225 U224 ; U56
g30 nand U227 U226 ; U57
g31 nand U229 U228 ; U58
g32 nand U231 U230 ; U59
g33 nand U233 U232 ; U60
g34 nand U235 U234 ; U61
g35 nand U237 U236 ; U62
g36 nand U239 U238 ; U63
g37 nand U241 U240 ; U64
g38 nand U243 U242 ; U65
g39 nand U245 U244 ; U66
g40 nand U247 U246 ; U67
g41 nand U249 U248 ; U68
g42 nand U251 U250 ; U69
g43 nand U253 U252 ; U70
g44 nand U255 U254 ; U71
g45 nand U257 U256 ; U72
g46 nand U259 U258 ; U73
g47 nand U261 U260 ; U74
g48 nand U263 U262 ; U75
g49 nand U265 U264 ; U76
g50 nand U267 U266 ; U77
g51 nand U269 U268 ; U78
g52 nand U271 U270 ; U79
g53 nand U273 U272 ; U80
g54 nand U275 U274 ; U81
g55 nand U277 U276 ; U82
g56 nand U279 U278 ; U83
g57 nand U281 U280 ; U84
g58 nand U283 U282 ; U85
g59 nand U285 U284 ; U86
g60 nand U287 U286 ; U87
g61 nand U289 U288 ; U88
g62 nand U291 U290 ; U89
g63 nand U293 U292 ; U90
g64 nand U295 U294 ; U91
g65 nand U297 U296 ; U92
g66 nand U299 U298 ; U93
g67 nand U301 U300 ; U94
g68 nand U303 U302 ; U95
g69 nand U305 U304 ; U96
g70 nand U307 U306 ; U97
g71 nand U309 U308 ; U98
g72 nand U311 U310 ; U99
g73 nand U313 U312 ; U100
g74 nand U315 U314 ; U101
g75 nand U317 U316 ; U102
g76 nand U319 U318 ; U103
g77 nand U321 U320 ; U104
g78 nand U323 U322 ; U105
g79 nand U325 U324 ; U106
g80 nand U327 U326 ; U107
g81 nand U329 U328 ; U108
g82 nand U331 U330 ; U109
g83 nand U333 U332 ; U110
g84 nand U335 U334 ; U111
g85 nand U337 U336 ; U112
g86 nand U339 U338 ; U113
g87 nand U341 U340 ; U114
g88 nand U343 U342 ; U115
g89 nand U345 U344 ; U116
g90 nand U347 U346 ; U117
g91 nand U349 U348 ; U118
g92 nand U351 U350 ; U119
g93 nand U353 U352 ; U120
g94 nand U355 U354 ; U121
g95 nand U357 U356 ; U122
g96 nand U359 U358 ; U123
g97 nand U361 U360 ; U124
g98 nand U363 U362 ; U125
g99 nand U365 U364 ; U126
g100 nand U367 U366 ; U127
g101 nand U369 U368 ; U128
g102 nand U371 U370 ; U129
g103 nand U373 U372 ; U130
g104 nand U375 U374 ; U131
g105 nand U377 U376 ; U132
g106 nand U379 U378 ; U133
g107 nand U381 U380 ; U134
g108 nand U383 U382 ; U135
g109 nand U385 U384 ; U136
g110 nand U387 U386 ; U137
g111 nand U389 U388 ; U138
g112 nand U391 U390 ; U139
g113 nand U393 U392 ; U140
g114 nand U395 U394 ; U141
g115 nand U397 U396 ; U142
g116 nand U399 U398 ; U143
g117 nand U401 U400 ; U144
g118 nand U403 U402 ; U145
g119 nand U405 U404 ; U146
g120 nand U407 U406 ; U147
g121 nand U409 U408 ; U148
g122 nand U411 U410 ; U149
g123 nand U413 U412 ; U150
g124 nand U415 U414 ; U151
g125 nand U417 U416 ; U152
g126 nand U419 U418 ; U153
g127 nand U421 U420 ; U154
g128 nand U423 U422 ; U155
g129 nand U425 U424 ; U156
g130 nand U427 U426 ; U157
g131 not P2_WR_REG_SCAN_IN ; U158
g132 not P1_WR_REG_SCAN_IN ; U159
g133 and U169 U168 ; U160
g134 not P2_RD_REG_SCAN_IN ; U161
g135 not P1_RD_REG_SCAN_IN ; U162
g136 and U171 U170 ; U163
g137 nand U166 U165 ; U164
g138 nand LT_1602_U6 U161 P1_ADDR_REG_19__SCAN_IN P2_ADDR_REG_19__SCAN_IN ; U165
g139 nand LT_1601_U6 LT_1601_21_U6 U162 P3_ADDR_REG_19__SCAN_IN ; U166
g140 not U164 ; U167
g141 nand U159 P2_WR_REG_SCAN_IN ; U168
g142 nand U158 P1_WR_REG_SCAN_IN ; U169
g143 nand U162 P2_RD_REG_SCAN_IN ; U170
g144 nand U161 P1_RD_REG_SCAN_IN ; U171
g145 nand SUB_1605_U79 U164 ; U172
g146 nand SI_9_ U167 ; U173
g147 nand SUB_1605_U80 U164 ; U174
g148 nand SI_8_ U167 ; U175
g149 nand SUB_1605_U81 U164 ; U176
g150 nand SI_7_ U167 ; U177
g151 nand SUB_1605_U82 U164 ; U178
g152 nand SI_6_ U167 ; U179
g153 nand SUB_1605_U83 U164 ; U180
g154 nand SI_5_ U167 ; U181
g155 nand SUB_1605_U84 U164 ; U182
g156 nand SI_4_ U167 ; U183
g157 nand SUB_1605_U85 U164 ; U184
g158 nand SI_3_ U167 ; U185
g159 nand SUB_1605_U12 U164 ; U186
g160 nand SI_31_ U167 ; U187
g161 nand SUB_1605_U86 U164 ; U188
g162 nand SI_30_ U167 ; U189
g163 nand SUB_1605_U87 U164 ; U190
g164 nand SI_2_ U167 ; U191
g165 nand SUB_1605_U88 U164 ; U192
g166 nand SI_29_ U167 ; U193
g167 nand SUB_1605_U89 U164 ; U194
g168 nand SI_28_ U167 ; U195
g169 nand SUB_1605_U90 U164 ; U196
g170 nand SI_27_ U167 ; U197
g171 nand SUB_1605_U91 U164 ; U198
g172 nand SI_26_ U167 ; U199
g173 nand SUB_1605_U92 U164 ; U200
g174 nand SI_25_ U167 ; U201
g175 nand SUB_1605_U93 U164 ; U202
g176 nand SI_24_ U167 ; U203
g177 nand SUB_1605_U94 U164 ; U204
g178 nand SI_23_ U167 ; U205
g179 nand SUB_1605_U95 U164 ; U206
g180 nand SI_22_ U167 ; U207
g181 nand SUB_1605_U96 U164 ; U208
g182 nand SI_21_ U167 ; U209
g183 nand SUB_1605_U97 U164 ; U210
g184 nand SI_20_ U167 ; U211
g185 nand SUB_1605_U98 U164 ; U212
g186 nand SI_1_ U167 ; U213
g187 nand SUB_1605_U99 U164 ; U214
g188 nand SI_19_ U167 ; U215
g189 nand SUB_1605_U100 U164 ; U216
g190 nand SI_18_ U167 ; U217
g191 nand SUB_1605_U101 U164 ; U218
g192 nand SI_17_ U167 ; U219
g193 nand SUB_1605_U102 U164 ; U220
g194 nand SI_16_ U167 ; U221
g195 nand SUB_1605_U103 U164 ; U222
g196 nand SI_15_ U167 ; U223
g197 nand SUB_1605_U104 U164 ; U224
g198 nand SI_14_ U167 ; U225
g199 nand SUB_1605_U105 U164 ; U226
g200 nand SI_13_ U167 ; U227
g201 nand SUB_1605_U106 U164 ; U228
g202 nand SI_12_ U167 ; U229
g203 nand SUB_1605_U107 U164 ; U230
g204 nand SI_11_ U167 ; U231
g205 nand SUB_1605_U108 U164 ; U232
g206 nand SI_10_ U167 ; U233
g207 nand SUB_1605_U13 U164 ; U234
g208 nand SI_0_ U167 ; U235
g209 nand U164 P1_DATAO_REG_9__SCAN_IN ; U236
g210 nand R152_U85 U167 ; U237
g211 nand U164 P1_DATAO_REG_8__SCAN_IN ; U238
g212 nand R152_U86 U167 ; U239
g213 nand U164 P1_DATAO_REG_7__SCAN_IN ; U240
g214 nand R152_U87 U167 ; U241
g215 nand U164 P1_DATAO_REG_6__SCAN_IN ; U242
g216 nand R152_U88 U167 ; U243
g217 nand U164 P1_DATAO_REG_5__SCAN_IN ; U244
g218 nand R152_U89 U167 ; U245
g219 nand U164 P1_DATAO_REG_4__SCAN_IN ; U246
g220 nand R152_U90 U167 ; U247
g221 nand U164 P1_DATAO_REG_3__SCAN_IN ; U248
g222 nand R152_U91 U167 ; U249
g223 nand U164 P1_DATAO_REG_31__SCAN_IN ; U250
g224 nand R152_U12 U167 ; U251
g225 nand U164 P1_DATAO_REG_30__SCAN_IN ; U252
g226 nand R152_U92 U167 ; U253
g227 nand U164 P1_DATAO_REG_2__SCAN_IN ; U254
g228 nand R152_U93 U167 ; U255
g229 nand U164 P1_DATAO_REG_29__SCAN_IN ; U256
g230 nand R152_U94 U167 ; U257
g231 nand U164 P1_DATAO_REG_28__SCAN_IN ; U258
g232 nand R152_U95 U167 ; U259
g233 nand U164 P1_DATAO_REG_27__SCAN_IN ; U260
g234 nand R152_U96 U167 ; U261
g235 nand U164 P1_DATAO_REG_26__SCAN_IN ; U262
g236 nand R152_U97 U167 ; U263
g237 nand U164 P1_DATAO_REG_25__SCAN_IN ; U264
g238 nand R152_U98 U167 ; U265
g239 nand U164 P1_DATAO_REG_24__SCAN_IN ; U266
g240 nand R152_U99 U167 ; U267
g241 nand U164 P1_DATAO_REG_23__SCAN_IN ; U268
g242 nand R152_U100 U167 ; U269
g243 nand U164 P1_DATAO_REG_22__SCAN_IN ; U270
g244 nand R152_U101 U167 ; U271
g245 nand U164 P1_DATAO_REG_21__SCAN_IN ; U272
g246 nand R152_U102 U167 ; U273
g247 nand U164 P1_DATAO_REG_20__SCAN_IN ; U274
g248 nand R152_U103 U167 ; U275
g249 nand U164 P1_DATAO_REG_1__SCAN_IN ; U276
g250 nand R152_U13 U167 ; U277
g251 nand U164 P1_DATAO_REG_19__SCAN_IN ; U278
g252 nand R152_U104 U167 ; U279
g253 nand U164 P1_DATAO_REG_18__SCAN_IN ; U280
g254 nand R152_U105 U167 ; U281
g255 nand U164 P1_DATAO_REG_17__SCAN_IN ; U282
g256 nand R152_U106 U167 ; U283
g257 nand U164 P1_DATAO_REG_16__SCAN_IN ; U284
g258 nand R152_U107 U167 ; U285
g259 nand U164 P1_DATAO_REG_15__SCAN_IN ; U286
g260 nand R152_U108 U167 ; U287
g261 nand U164 P1_DATAO_REG_14__SCAN_IN ; U288
g262 nand R152_U109 U167 ; U289
g263 nand U164 P1_DATAO_REG_13__SCAN_IN ; U290
g264 nand R152_U110 U167 ; U291
g265 nand U164 P1_DATAO_REG_12__SCAN_IN ; U292
g266 nand R152_U111 U167 ; U293
g267 nand U164 P1_DATAO_REG_11__SCAN_IN ; U294
g268 nand R152_U112 U167 ; U295
g269 nand U164 P1_DATAO_REG_10__SCAN_IN ; U296
g270 nand R152_U113 U167 ; U297
g271 nand U164 P1_DATAO_REG_0__SCAN_IN ; U298
g272 nand R152_U84 U167 ; U299
g273 nand R152_U85 U164 ; U300
g274 nand U167 P2_DATAO_REG_9__SCAN_IN ; U301
g275 nand R152_U86 U164 ; U302
g276 nand U167 P2_DATAO_REG_8__SCAN_IN ; U303
g277 nand R152_U87 U164 ; U304
g278 nand U167 P2_DATAO_REG_7__SCAN_IN ; U305
g279 nand R152_U88 U164 ; U306
g280 nand U167 P2_DATAO_REG_6__SCAN_IN ; U307
g281 nand R152_U89 U164 ; U308
g282 nand U167 P2_DATAO_REG_5__SCAN_IN ; U309
g283 nand R152_U90 U164 ; U310
g284 nand U167 P2_DATAO_REG_4__SCAN_IN ; U311
g285 nand R152_U91 U164 ; U312
g286 nand U167 P2_DATAO_REG_3__SCAN_IN ; U313
g287 nand R152_U12 U164 ; U314
g288 nand U167 P2_DATAO_REG_31__SCAN_IN ; U315
g289 nand R152_U92 U164 ; U316
g290 nand U167 P2_DATAO_REG_30__SCAN_IN ; U317
g291 nand R152_U93 U164 ; U318
g292 nand U167 P2_DATAO_REG_2__SCAN_IN ; U319
g293 nand R152_U94 U164 ; U320
g294 nand U167 P2_DATAO_REG_29__SCAN_IN ; U321
g295 nand R152_U95 U164 ; U322
g296 nand U167 P2_DATAO_REG_28__SCAN_IN ; U323
g297 nand R152_U96 U164 ; U324
g298 nand U167 P2_DATAO_REG_27__SCAN_IN ; U325
g299 nand R152_U97 U164 ; U326
g300 nand U167 P2_DATAO_REG_26__SCAN_IN ; U327
g301 nand R152_U98 U164 ; U328
g302 nand U167 P2_DATAO_REG_25__SCAN_IN ; U329
g303 nand R152_U99 U164 ; U330
g304 nand U167 P2_DATAO_REG_24__SCAN_IN ; U331
g305 nand R152_U100 U164 ; U332
g306 nand U167 P2_DATAO_REG_23__SCAN_IN ; U333
g307 nand R152_U101 U164 ; U334
g308 nand U167 P2_DATAO_REG_22__SCAN_IN ; U335
g309 nand R152_U102 U164 ; U336
g310 nand U167 P2_DATAO_REG_21__SCAN_IN ; U337
g311 nand R152_U103 U164 ; U338
g312 nand U167 P2_DATAO_REG_20__SCAN_IN ; U339
g313 nand R152_U13 U164 ; U340
g314 nand U167 P2_DATAO_REG_1__SCAN_IN ; U341
g315 nand R152_U104 U164 ; U342
g316 nand U167 P2_DATAO_REG_19__SCAN_IN ; U343
g317 nand R152_U105 U164 ; U344
g318 nand U167 P2_DATAO_REG_18__SCAN_IN ; U345
g319 nand R152_U106 U164 ; U346
g320 nand U167 P2_DATAO_REG_17__SCAN_IN ; U347
g321 nand R152_U107 U164 ; U348
g322 nand U167 P2_DATAO_REG_16__SCAN_IN ; U349
g323 nand R152_U108 U164 ; U350
g324 nand U167 P2_DATAO_REG_15__SCAN_IN ; U351
g325 nand R152_U109 U164 ; U352
g326 nand U167 P2_DATAO_REG_14__SCAN_IN ; U353
g327 nand R152_U110 U164 ; U354
g328 nand U167 P2_DATAO_REG_13__SCAN_IN ; U355
g329 nand R152_U111 U164 ; U356
g330 nand U167 P2_DATAO_REG_12__SCAN_IN ; U357
g331 nand R152_U112 U164 ; U358
g332 nand U167 P2_DATAO_REG_11__SCAN_IN ; U359
g333 nand R152_U113 U164 ; U360
g334 nand U167 P2_DATAO_REG_10__SCAN_IN ; U361
g335 nand R152_U84 U164 ; U362
g336 nand U167 P2_DATAO_REG_0__SCAN_IN ; U363
g337 nand U164 P2_DATAO_REG_9__SCAN_IN ; U364
g338 nand U167 P1_DATAO_REG_9__SCAN_IN ; U365
g339 nand U164 P2_DATAO_REG_8__SCAN_IN ; U366
g340 nand U167 P1_DATAO_REG_8__SCAN_IN ; U367
g341 nand U164 P2_DATAO_REG_7__SCAN_IN ; U368
g342 nand U167 P1_DATAO_REG_7__SCAN_IN ; U369
g343 nand U164 P2_DATAO_REG_6__SCAN_IN ; U370
g344 nand U167 P1_DATAO_REG_6__SCAN_IN ; U371
g345 nand U164 P2_DATAO_REG_5__SCAN_IN ; U372
g346 nand U167 P1_DATAO_REG_5__SCAN_IN ; U373
g347 nand U164 P2_DATAO_REG_4__SCAN_IN ; U374
g348 nand U167 P1_DATAO_REG_4__SCAN_IN ; U375
g349 nand U164 P2_DATAO_REG_31__SCAN_IN ; U376
g350 nand U167 P1_DATAO_REG_31__SCAN_IN ; U377
g351 nand U164 P2_DATAO_REG_30__SCAN_IN ; U378
g352 nand U167 P1_DATAO_REG_30__SCAN_IN ; U379
g353 nand U164 P2_DATAO_REG_3__SCAN_IN ; U380
g354 nand U167 P1_DATAO_REG_3__SCAN_IN ; U381
g355 nand U164 P2_DATAO_REG_29__SCAN_IN ; U382
g356 nand U167 P1_DATAO_REG_29__SCAN_IN ; U383
g357 nand U164 P2_DATAO_REG_28__SCAN_IN ; U384
g358 nand U167 P1_DATAO_REG_28__SCAN_IN ; U385
g359 nand U164 P2_DATAO_REG_27__SCAN_IN ; U386
g360 nand U167 P1_DATAO_REG_27__SCAN_IN ; U387
g361 nand U164 P2_DATAO_REG_26__SCAN_IN ; U388
g362 nand U167 P1_DATAO_REG_26__SCAN_IN ; U389
g363 nand U164 P2_DATAO_REG_25__SCAN_IN ; U390
g364 nand U167 P1_DATAO_REG_25__SCAN_IN ; U391
g365 nand U164 P2_DATAO_REG_24__SCAN_IN ; U392
g366 nand U167 P1_DATAO_REG_24__SCAN_IN ; U393
g367 nand U164 P2_DATAO_REG_23__SCAN_IN ; U394
g368 nand U167 P1_DATAO_REG_23__SCAN_IN ; U395
g369 nand U164 P2_DATAO_REG_22__SCAN_IN ; U396
g370 nand U167 P1_DATAO_REG_22__SCAN_IN ; U397
g371 nand U164 P2_DATAO_REG_21__SCAN_IN ; U398
g372 nand U167 P1_DATAO_REG_21__SCAN_IN ; U399
g373 nand U164 P2_DATAO_REG_20__SCAN_IN ; U400
g374 nand U167 P1_DATAO_REG_20__SCAN_IN ; U401
g375 nand U164 P2_DATAO_REG_2__SCAN_IN ; U402
g376 nand U167 P1_DATAO_REG_2__SCAN_IN ; U403
g377 nand U164 P2_DATAO_REG_19__SCAN_IN ; U404
g378 nand U167 P1_DATAO_REG_19__SCAN_IN ; U405
g379 nand U164 P2_DATAO_REG_18__SCAN_IN ; U406
g380 nand U167 P1_DATAO_REG_18__SCAN_IN ; U407
g381 nand U164 P2_DATAO_REG_17__SCAN_IN ; U408
g382 nand U167 P1_DATAO_REG_17__SCAN_IN ; U409
g383 nand U164 P2_DATAO_REG_16__SCAN_IN ; U410
g384 nand U167 P1_DATAO_REG_16__SCAN_IN ; U411
g385 nand U164 P2_DATAO_REG_15__SCAN_IN ; U412
g386 nand U167 P1_DATAO_REG_15__SCAN_IN ; U413
g387 nand U164 P2_DATAO_REG_14__SCAN_IN ; U414
g388 nand U167 P1_DATAO_REG_14__SCAN_IN ; U415
g389 nand U164 P2_DATAO_REG_13__SCAN_IN ; U416
g390 nand U167 P1_DATAO_REG_13__SCAN_IN ; U417
g391 nand U164 P2_DATAO_REG_12__SCAN_IN ; U418
g392 nand U167 P1_DATAO_REG_12__SCAN_IN ; U419
g393 nand U164 P2_DATAO_REG_11__SCAN_IN ; U420
g394 nand U167 P1_DATAO_REG_11__SCAN_IN ; U421
g395 nand U164 P2_DATAO_REG_10__SCAN_IN ; U422
g396 nand U167 P1_DATAO_REG_10__SCAN_IN ; U423
g397 nand U164 P2_DATAO_REG_1__SCAN_IN ; U424
g398 nand U167 P1_DATAO_REG_1__SCAN_IN ; U425
g399 nand U164 P2_DATAO_REG_0__SCAN_IN ; U426
g400 nand U167 P1_DATAO_REG_0__SCAN_IN ; U427
g401 and P1_U4002 P1_U3451 ; P1_U3014
g402 and P1_U3455 P1_U3449 ; P1_U3015
g403 and P1_U3605 P1_U3600 ; P1_U3016
g404 and P1_U3447 P1_U3448 ; P1_U3017
g405 and P1_U5808 P1_U3447 ; P1_U3018
g406 and P1_U5805 P1_U3448 ; P1_U3019
g407 and P1_U5805 P1_U5808 ; P1_U3020
g408 and P1_U5412 P1_U3425 ; P1_U3021
g409 and P1_U3592 P1_U3425 ; P1_U3022
g410 and P1_U4043 P1_U3428 ; P1_U3023
g411 and P1_U3048 P1_U5793 ; P1_U3024
g412 and P1_U4030 P1_U5811 ; P1_U3025
g413 and P1_U3851 P1_U4015 ; P1_U3026
g414 and P1_R1352_U6 P1_U3437 ; P1_U3027
g415 and P1_R1352_U6 P1_U3440 ; P1_U3028
g416 and P1_U3357 P1_STATE_REG_SCAN_IN ; P1_U3029
g417 and P1_U4008 P1_U4031 ; P1_U3030
g418 and P1_U4031 P1_U3426 ; P1_U3031
g419 and P1_U4003 P1_U4031 ; P1_U3032
g420 and P1_U4009 P1_U4031 ; P1_U3033
g421 and P1_U4030 P1_U3449 ; P1_U3034
g422 and P1_U4015 P1_U5811 ; P1_U3035
g423 and P1_U4031 P1_U3025 ; P1_U3036
g424 and P1_U4015 P1_U3449 ; P1_U3037
g425 and P1_U5817 P1_U4923 ; P1_U3038
g426 and P1_U3023 P1_U5817 ; P1_U3039
g427 and P1_U5811 P1_U4923 ; P1_U3040
g428 and P1_U3023 P1_U5811 ; P1_U3041
g429 and P1_U3015 P1_U4923 ; P1_U3042
g430 and P1_U3023 P1_U3015 ; P1_U3043
g431 and P1_U3022 P1_U3428 ; P1_U3044
g432 and P1_U3022 P1_U5159 ; P1_U3045
g433 and P1_U3606 P1_U3016 ; P1_U3046
g434 and P1_U3452 P1_U3453 ; P1_U3047
g435 and P1_U5799 P1_U3452 ; P1_U3048
g436 and P1_U5802 P1_U5796 ; P1_U3049
g437 and P1_U3850 P1_U5148 ; P1_U3050
g438 and P1_U3419 P1_U3367 ; P1_U3051
g439 and P1_U5541 P1_U3422 P1_U3879 ; P1_U3052
g440 nand P1_U4680 P1_U4681 P1_U4679 P1_U4682 ; P1_U3053
g441 nand P1_U4699 P1_U4700 P1_U4698 P1_U4701 ; P1_U3054
g442 nand P1_U4720 P1_U4719 P1_U4718 P1_U4717 ; P1_U3055
g443 nand P1_U4757 P1_U4758 P1_U4756 ; P1_U3056
g444 nand P1_U4661 P1_U4662 P1_U4660 P1_U4663 ; P1_U3057
g445 nand P1_U4642 P1_U4643 P1_U4641 P1_U4644 ; P1_U3058
g446 nand P1_U4737 P1_U4738 P1_U4736 ; P1_U3059
g447 nand P1_U4245 P1_U4244 P1_U4243 P1_U4242 ; P1_U3060
g448 nand P1_U4585 P1_U4586 P1_U4584 P1_U4587 ; P1_U3061
g449 nand P1_U4357 P1_U4358 P1_U4356 P1_U4359 ; P1_U3062
g450 nand P1_U4376 P1_U4377 P1_U4375 P1_U4378 ; P1_U3063
g451 nand P1_U4226 P1_U4225 P1_U4224 P1_U4223 ; P1_U3064
g452 nand P1_U4623 P1_U4624 P1_U4622 P1_U4625 ; P1_U3065
g453 nand P1_U4604 P1_U4605 P1_U4603 P1_U4606 ; P1_U3066
g454 nand P1_U4264 P1_U4263 P1_U4262 P1_U4261 ; P1_U3067
g455 nand P1_U4202 P1_U4201 P1_U4200 P1_U4199 ; P1_U3068
g456 nand P1_U4490 P1_U4491 P1_U4489 P1_U4492 ; P1_U3069
g457 nand P1_U4302 P1_U4301 P1_U4300 P1_U4299 ; P1_U3070
g458 nand P1_U4283 P1_U4282 P1_U4281 P1_U4280 ; P1_U3071
g459 nand P1_U4395 P1_U4396 P1_U4394 P1_U4397 ; P1_U3072
g460 nand P1_U4471 P1_U4472 P1_U4470 P1_U4473 ; P1_U3073
g461 nand P1_U4452 P1_U4453 P1_U4451 P1_U4454 ; P1_U3074
g462 nand P1_U4566 P1_U4567 P1_U4565 P1_U4568 ; P1_U3075
g463 nand P1_U4547 P1_U4548 P1_U4546 P1_U4549 ; P1_U3076
g464 nand P1_U4207 P1_U4206 P1_U4205 P1_U4204 ; P1_U3077
g465 nand P1_U4183 P1_U4182 P1_U4181 P1_U4180 ; P1_U3078
g466 nand P1_U4433 P1_U4434 P1_U4432 P1_U4435 ; P1_U3079
g467 nand P1_U4414 P1_U4415 P1_U4413 P1_U4416 ; P1_U3080
g468 nand P1_U4528 P1_U4529 P1_U4527 P1_U4530 ; P1_U3081
g469 nand P1_U4509 P1_U4510 P1_U4508 P1_U4511 ; P1_U3082
g470 nand P1_U4338 P1_U4339 P1_U4337 P1_U4340 ; P1_U3083
g471 nand P1_U4321 P1_U4320 P1_U4319 P1_U4318 ; P1_U3084
g472 nand P1_U4930 P1_STATE_REG_SCAN_IN ; P1_U3085
g473 not P1_STATE_REG_SCAN_IN ; P1_U3086
g474 nand P1_U5668 P1_U5666 P1_U5667 ; P1_U3087
g475 nand P1_U5671 P1_U5669 P1_U5670 ; P1_U3088
g476 nand P1_U3929 P1_U5678 P1_U5679 ; P1_U3089
g477 nand P1_U5683 P1_U5682 P1_U3930 ; P1_U3090
g478 nand P1_U5687 P1_U5686 P1_U3931 ; P1_U3091
g479 nand P1_U5691 P1_U5690 P1_U3932 ; P1_U3092
g480 nand P1_U5695 P1_U5694 P1_U3933 ; P1_U3093
g481 nand P1_U5699 P1_U5698 P1_U3934 ; P1_U3094
g482 nand P1_U5703 P1_U5702 P1_U3935 ; P1_U3095
g483 nand P1_U5707 P1_U5706 P1_U3936 ; P1_U3096
g484 nand P1_U5711 P1_U5710 P1_U3937 ; P1_U3097
g485 nand P1_U5715 P1_U5714 P1_U3938 ; P1_U3098
g486 nand P1_U5723 P1_U5722 P1_U3940 ; P1_U3099
g487 nand P1_U5727 P1_U5726 P1_U3941 ; P1_U3100
g488 nand P1_U5731 P1_U5730 P1_U3942 ; P1_U3101
g489 nand P1_U5735 P1_U5734 P1_U3943 ; P1_U3102
g490 nand P1_U5739 P1_U5738 P1_U3944 ; P1_U3103
g491 nand P1_U5743 P1_U5742 P1_U3945 ; P1_U3104
g492 nand P1_U5747 P1_U5746 P1_U3946 ; P1_U3105
g493 nand P1_U5751 P1_U5750 P1_U3947 ; P1_U3106
g494 nand P1_U5755 P1_U5754 P1_U3948 ; P1_U3107
g495 nand P1_U5759 P1_U5758 P1_U3949 ; P1_U3108
g496 nand P1_U3922 P1_U5644 P1_U5643 ; P1_U3109
g497 nand P1_U3923 P1_U5648 P1_U5647 ; P1_U3110
g498 nand P1_U5653 P1_U5652 P1_U3924 ; P1_U3111
g499 nand P1_U5657 P1_U5656 P1_U3925 ; P1_U3112
g500 nand P1_U5661 P1_U5660 P1_U3926 ; P1_U3113
g501 nand P1_U5665 P1_U5664 P1_U3927 ; P1_U3114
g502 nand P1_U3928 P1_U5674 ; P1_U3115
g503 nand P1_U3939 P1_U5718 ; P1_U3116
g504 nand P1_U3950 P1_U5762 ; P1_U3117
g505 nand P1_U3951 P1_U5766 ; P1_U3118
g506 nand P1_U3892 P1_U5563 ; P1_U3119
g507 nand P1_U3893 P1_U5566 ; P1_U3120
g508 nand P1_U5572 P1_U5571 P1_U3896 ; P1_U3121
g509 nand P1_U5575 P1_U5574 P1_U3897 ; P1_U3122
g510 nand P1_U5578 P1_U5577 P1_U3898 ; P1_U3123
g511 nand P1_U5581 P1_U5580 P1_U3899 ; P1_U3124
g512 nand P1_U5584 P1_U5583 P1_U3900 ; P1_U3125
g513 nand P1_U5587 P1_U5586 P1_U3901 ; P1_U3126
g514 nand P1_U5590 P1_U5589 P1_U3902 ; P1_U3127
g515 nand P1_U5593 P1_U5592 P1_U3903 ; P1_U3128
g516 nand P1_U5596 P1_U5595 P1_U3904 ; P1_U3129
g517 nand P1_U5599 P1_U5598 P1_U3905 ; P1_U3130
g518 nand P1_U5605 P1_U5604 P1_U3908 ; P1_U3131
g519 nand P1_U5608 P1_U5607 P1_U3909 ; P1_U3132
g520 nand P1_U5611 P1_U5610 P1_U3910 ; P1_U3133
g521 nand P1_U5614 P1_U5613 P1_U3911 ; P1_U3134
g522 nand P1_U5617 P1_U5616 P1_U3912 ; P1_U3135
g523 nand P1_U5620 P1_U5619 P1_U3913 ; P1_U3136
g524 nand P1_U5623 P1_U5622 P1_U3914 ; P1_U3137
g525 nand P1_U5626 P1_U5625 P1_U3915 ; P1_U3138
g526 nand P1_U5629 P1_U5628 P1_U3916 ; P1_U3139
g527 nand P1_U5632 P1_U5631 P1_U3917 ; P1_U3140
g528 nand P1_U5545 P1_U3880 ; P1_U3141
g529 nand P1_U5548 P1_U3882 ; P1_U3142
g530 nand P1_U5551 P1_U3884 ; P1_U3143
g531 nand P1_U5554 P1_U3886 ; P1_U3144
g532 nand P1_U5557 P1_U3888 ; P1_U3145
g533 nand P1_U5560 P1_U3890 ; P1_U3146
g534 nand P1_U5569 P1_U3894 ; P1_U3147
g535 nand P1_U5602 P1_U3906 ; P1_U3148
g536 nand P1_U5635 P1_U3918 ; P1_U3149
g537 nand P1_U5638 P1_U3920 ; P1_U3150
g538 nand P1_U3877 P1_U5537 ; P1_U3151
g539 nand P1_U3014 P1_U5786 ; P1_U3152
g540 nand P1_U5492 P1_U5491 ; P1_U3153
g541 nand P1_U5494 P1_U5493 ; P1_U3154
g542 nand P1_U5496 P1_U5495 ; P1_U3155
g543 nand P1_U5498 P1_U5497 ; P1_U3156
g544 nand P1_U5500 P1_U5499 ; P1_U3157
g545 nand P1_U5502 P1_U5501 ; P1_U3158
g546 nand P1_U5504 P1_U5503 ; P1_U3159
g547 nand P1_U5506 P1_U5505 ; P1_U3160
g548 nand P1_U5508 P1_U5507 ; P1_U3161
g549 nand P1_U5512 P1_U5511 ; P1_U3162
g550 nand P1_U5514 P1_U5513 ; P1_U3163
g551 nand P1_U5516 P1_U5515 ; P1_U3164
g552 nand P1_U5518 P1_U5517 ; P1_U3165
g553 nand P1_U5520 P1_U5519 ; P1_U3166
g554 nand P1_U5522 P1_U5521 ; P1_U3167
g555 nand P1_U5524 P1_U5523 ; P1_U3168
g556 nand P1_U5526 P1_U5525 ; P1_U3169
g557 nand P1_U5528 P1_U5527 ; P1_U3170
g558 nand P1_U5530 P1_U5529 ; P1_U3171
g559 nand P1_U5478 P1_U5477 ; P1_U3172
g560 nand P1_U5480 P1_U5479 ; P1_U3173
g561 nand P1_U5482 P1_U5481 ; P1_U3174
g562 nand P1_U5484 P1_U5483 ; P1_U3175
g563 nand P1_U5486 P1_U5485 ; P1_U3176
g564 nand P1_U5488 P1_U5487 ; P1_U3177
g565 nand P1_U5490 P1_U5489 ; P1_U3178
g566 nand P1_U5510 P1_U5509 ; P1_U3179
g567 nand P1_U5532 P1_U5531 ; P1_U3180
g568 nand P1_U3876 P1_U5534 ; P1_U3181
g569 nand P1_U5433 P1_U5432 ; P1_U3182
g570 nand P1_U5435 P1_U5434 ; P1_U3183
g571 nand P1_U5437 P1_U5436 ; P1_U3184
g572 nand P1_U5439 P1_U5438 ; P1_U3185
g573 nand P1_U5441 P1_U5440 ; P1_U3186
g574 nand P1_U5443 P1_U5442 ; P1_U3187
g575 nand P1_U5445 P1_U5444 ; P1_U3188
g576 nand P1_U5447 P1_U5446 ; P1_U3189
g577 nand P1_U5449 P1_U5448 ; P1_U3190
g578 nand P1_U5453 P1_U5452 ; P1_U3191
g579 nand P1_U5455 P1_U5454 ; P1_U3192
g580 nand P1_U5457 P1_U5456 ; P1_U3193
g581 nand P1_U5459 P1_U5458 ; P1_U3194
g582 nand P1_U5461 P1_U5460 ; P1_U3195
g583 nand P1_U5463 P1_U5462 ; P1_U3196
g584 nand P1_U5465 P1_U5464 ; P1_U3197
g585 nand P1_U5467 P1_U5466 ; P1_U3198
g586 nand P1_U5469 P1_U5468 ; P1_U3199
g587 nand P1_U5471 P1_U5470 ; P1_U3200
g588 nand P1_U5419 P1_U5418 ; P1_U3201
g589 nand P1_U5421 P1_U5420 ; P1_U3202
g590 nand P1_U5423 P1_U5422 ; P1_U3203
g591 nand P1_U5425 P1_U5424 ; P1_U3204
g592 nand P1_U5427 P1_U5426 ; P1_U3205
g593 nand P1_U5429 P1_U5428 ; P1_U3206
g594 nand P1_U5431 P1_U5430 ; P1_U3207
g595 nand P1_U5451 P1_U5450 ; P1_U3208
g596 nand P1_U5473 P1_U5472 ; P1_U3209
g597 nand P1_U3875 P1_U5474 ; P1_U3210
g598 and P1_U5411 P1_U3425 ; P1_U3211
g599 nand P1_U6285 P1_U6284 P1_U5409 ; P1_U3212
g600 nand P1_U5403 P1_U5402 P1_U3872 P1_U5404 ; P1_U3213
g601 nand P1_U5394 P1_U5393 P1_U5397 P1_U5396 P1_U5395 ; P1_U3214
g602 nand P1_U5385 P1_U5384 P1_U5388 P1_U5387 P1_U5386 ; P1_U3215
g603 nand P1_U5376 P1_U5375 P1_U5379 P1_U5378 P1_U5377 ; P1_U3216
g604 nand P1_U5367 P1_U5366 P1_U3871 P1_U5368 ; P1_U3217
g605 nand P1_U3869 P1_U5358 P1_U3870 ; P1_U3218
g606 nand P1_U5349 P1_U5348 P1_U5352 P1_U5351 P1_U5350 ; P1_U3219
g607 nand P1_U5340 P1_U5339 P1_U5343 P1_U5342 P1_U5341 ; P1_U3220
g608 nand P1_U5331 P1_U5330 P1_U3868 P1_U5332 ; P1_U3221
g609 nand P1_U3866 P1_U5322 P1_U3867 ; P1_U3222
g610 nand P1_U5313 P1_U5312 P1_U5316 P1_U5315 P1_U5314 ; P1_U3223
g611 nand P1_U5304 P1_U5303 P1_U3865 P1_U5305 ; P1_U3224
g612 nand P1_U5295 P1_U5294 P1_U5298 P1_U5297 P1_U5296 ; P1_U3225
g613 nand P1_U5286 P1_U5285 P1_U5289 P1_U5288 P1_U5287 ; P1_U3226
g614 nand P1_U5277 P1_U5276 P1_U5278 P1_U3864 ; P1_U3227
g615 nand P1_U5268 P1_U5267 P1_U5271 P1_U5270 P1_U5269 ; P1_U3228
g616 nand P1_U5259 P1_U5258 P1_U5262 P1_U5261 P1_U5260 ; P1_U3229
g617 nand P1_U3862 P1_U5250 P1_U3863 ; P1_U3230
g618 nand P1_U5241 P1_U5240 P1_U3861 P1_U5242 ; P1_U3231
g619 nand P1_U5233 P1_U3859 ; P1_U3232
g620 nand P1_U5224 P1_U5223 P1_U5227 P1_U5226 P1_U5225 ; P1_U3233
g621 nand P1_U5215 P1_U5214 P1_U3857 P1_U5216 ; P1_U3234
g622 nand P1_U5206 P1_U5205 P1_U5209 P1_U5208 P1_U5207 ; P1_U3235
g623 nand P1_U5197 P1_U5196 P1_U3856 P1_U5198 ; P1_U3236
g624 nand P1_U3854 P1_U5188 P1_U3855 ; P1_U3237
g625 nand P1_U5179 P1_U5178 P1_U5182 P1_U5181 P1_U5180 ; P1_U3238
g626 nand P1_U5170 P1_U5169 P1_U3853 P1_U5171 ; P1_U3239
g627 nand P1_U5161 P1_U5160 P1_U5164 P1_U5163 P1_U5162 ; P1_U3240
g628 nand P1_U5150 P1_U5149 P1_U5153 P1_U5152 P1_U5151 ; P1_U3241
g629 nand P1_U3846 P1_U5137 ; P1_U3242
g630 nand P1_U3830 P1_U5123 P1_U3831 ; P1_U3243
g631 nand P1_U3828 P1_U5113 P1_U3829 ; P1_U3244
g632 nand P1_U5103 P1_U3825 P1_U3827 ; P1_U3245
g633 nand P1_U3823 P1_U5093 P1_U3824 ; P1_U3246
g634 nand P1_U5083 P1_U3820 P1_U3822 ; P1_U3247
g635 nand P1_U3818 P1_U5073 P1_U3819 ; P1_U3248
g636 nand P1_U3816 P1_U3817 P1_U5063 ; P1_U3249
g637 nand P1_U3814 P1_U3815 P1_U5053 ; P1_U3250
g638 nand P1_U3812 P1_U3813 P1_U5043 ; P1_U3251
g639 nand P1_U3810 P1_U3811 P1_U5033 ; P1_U3252
g640 nand P1_U3808 P1_U3809 P1_U5023 ; P1_U3253
g641 nand P1_U3806 P1_U3807 P1_U5013 ; P1_U3254
g642 nand P1_U3804 P1_U3805 P1_U5003 ; P1_U3255
g643 nand P1_U3802 P1_U3803 P1_U4993 ; P1_U3256
g644 nand P1_U3800 P1_U3801 P1_U4983 ; P1_U3257
g645 nand P1_U3798 P1_U3799 P1_U4973 ; P1_U3258
g646 nand P1_U3796 P1_U3797 P1_U4963 ; P1_U3259
g647 nand P1_U3794 P1_U3795 P1_U4953 ; P1_U3260
g648 nand P1_U3792 P1_U3793 P1_U4943 ; P1_U3261
g649 nand P1_U3790 P1_U3791 P1_U4933 ; P1_U3262
g650 nand P1_U3989 P1_U4921 P1_U4922 ; P1_U3263
g651 nand P1_U3988 P1_U4919 P1_U4920 ; P1_U3264
g652 nand P1_U3784 P1_U3785 P1_U4912 P1_U3985 ; P1_U3265
g653 nand P1_U3782 P1_U3783 P1_U4907 P1_U3984 ; P1_U3266
g654 nand P1_U3780 P1_U3781 P1_U4902 P1_U3983 ; P1_U3267
g655 nand P1_U3778 P1_U3779 P1_U4897 P1_U3982 ; P1_U3268
g656 nand P1_U3776 P1_U3777 P1_U4892 P1_U3981 ; P1_U3269
g657 nand P1_U3774 P1_U3775 P1_U4887 P1_U3980 ; P1_U3270
g658 nand P1_U3772 P1_U3773 P1_U4882 P1_U3979 ; P1_U3271
g659 nand P1_U3770 P1_U3771 P1_U4877 P1_U3978 ; P1_U3272
g660 nand P1_U3768 P1_U3769 P1_U4872 P1_U3977 ; P1_U3273
g661 nand P1_U3766 P1_U3767 P1_U4867 P1_U3976 ; P1_U3274
g662 nand P1_U3765 P1_U3764 P1_U3975 ; P1_U3275
g663 nand P1_U3763 P1_U3762 P1_U3974 ; P1_U3276
g664 nand P1_U3760 P1_U3761 P1_U4852 P1_U3973 ; P1_U3277
g665 nand P1_U3758 P1_U3759 P1_U4847 P1_U3972 ; P1_U3278
g666 nand P1_U3757 P1_U3756 P1_U3971 ; P1_U3279
g667 nand P1_U3755 P1_U3754 P1_U3970 ; P1_U3280
g668 nand P1_U3753 P1_U3752 P1_U3969 ; P1_U3281
g669 nand P1_U3751 P1_U3750 P1_U3968 ; P1_U3282
g670 nand P1_U3748 P1_U3749 P1_U4822 P1_U3967 ; P1_U3283
g671 nand P1_U3746 P1_U3747 P1_U4817 P1_U3966 ; P1_U3284
g672 nand P1_U3745 P1_U3744 P1_U3965 ; P1_U3285
g673 nand P1_U3743 P1_U3742 P1_U3964 ; P1_U3286
g674 nand P1_U3741 P1_U3740 P1_U3963 ; P1_U3287
g675 nand P1_U3739 P1_U3738 P1_U3962 ; P1_U3288
g676 nand P1_U3737 P1_U3736 ; P1_U3289
g677 nand P1_U3735 P1_U3734 ; P1_U3290
g678 nand P1_U3733 P1_U3732 ; P1_U3291
g679 nand P1_U3731 P1_U3730 ; P1_U3292
g680 nand P1_U3729 P1_U3728 ; P1_U3293
g681 and P1_U3953 P1_D_REG_31__SCAN_IN ; P1_U3294
g682 and P1_U3953 P1_D_REG_30__SCAN_IN ; P1_U3295
g683 and P1_U3953 P1_D_REG_29__SCAN_IN ; P1_U3296
g684 and P1_U3953 P1_D_REG_28__SCAN_IN ; P1_U3297
g685 and P1_U3953 P1_D_REG_27__SCAN_IN ; P1_U3298
g686 and P1_U3953 P1_D_REG_26__SCAN_IN ; P1_U3299
g687 and P1_U3953 P1_D_REG_25__SCAN_IN ; P1_U3300
g688 and P1_U3953 P1_D_REG_24__SCAN_IN ; P1_U3301
g689 and P1_U3953 P1_D_REG_23__SCAN_IN ; P1_U3302
g690 and P1_U3953 P1_D_REG_22__SCAN_IN ; P1_U3303
g691 and P1_U3953 P1_D_REG_21__SCAN_IN ; P1_U3304
g692 and P1_U3953 P1_D_REG_20__SCAN_IN ; P1_U3305
g693 and P1_U3953 P1_D_REG_19__SCAN_IN ; P1_U3306
g694 and P1_U3953 P1_D_REG_18__SCAN_IN ; P1_U3307
g695 and P1_U3953 P1_D_REG_17__SCAN_IN ; P1_U3308
g696 and P1_U3953 P1_D_REG_16__SCAN_IN ; P1_U3309
g697 and P1_U3953 P1_D_REG_15__SCAN_IN ; P1_U3310
g698 and P1_U3953 P1_D_REG_14__SCAN_IN ; P1_U3311
g699 and P1_U3953 P1_D_REG_13__SCAN_IN ; P1_U3312
g700 and P1_U3953 P1_D_REG_12__SCAN_IN ; P1_U3313
g701 and P1_U3953 P1_D_REG_11__SCAN_IN ; P1_U3314
g702 and P1_U3953 P1_D_REG_10__SCAN_IN ; P1_U3315
g703 and P1_U3953 P1_D_REG_9__SCAN_IN ; P1_U3316
g704 and P1_U3953 P1_D_REG_8__SCAN_IN ; P1_U3317
g705 and P1_U3953 P1_D_REG_7__SCAN_IN ; P1_U3318
g706 and P1_U3953 P1_D_REG_6__SCAN_IN ; P1_U3319
g707 and P1_U3953 P1_D_REG_5__SCAN_IN ; P1_U3320
g708 and P1_U3953 P1_D_REG_4__SCAN_IN ; P1_U3321
g709 and P1_U3953 P1_D_REG_3__SCAN_IN ; P1_U3322
g710 and P1_U3953 P1_D_REG_2__SCAN_IN ; P1_U3323
g711 nand P1_U4142 P1_U4143 P1_U4141 ; P1_U3324
g712 nand P1_U4139 P1_U4140 P1_U4138 ; P1_U3325
g713 nand P1_U4136 P1_U4137 P1_U4135 ; P1_U3326
g714 nand P1_U4133 P1_U4134 P1_U4132 ; P1_U3327
g715 nand P1_U4130 P1_U4131 P1_U4129 ; P1_U3328
g716 nand P1_U4127 P1_U4128 P1_U4126 ; P1_U3329
g717 nand P1_U4124 P1_U4125 P1_U4123 ; P1_U3330
g718 nand P1_U4121 P1_U4122 P1_U4120 ; P1_U3331
g719 nand P1_U4118 P1_U4119 P1_U4117 ; P1_U3332
g720 nand P1_U4115 P1_U4116 P1_U4114 ; P1_U3333
g721 nand P1_U4112 P1_U4113 P1_U4111 ; P1_U3334
g722 nand P1_U4109 P1_U4110 P1_U4108 ; P1_U3335
g723 nand P1_U4106 P1_U4107 P1_U4105 ; P1_U3336
g724 nand P1_U4103 P1_U4104 P1_U4102 ; P1_U3337
g725 nand P1_U4100 P1_U4101 P1_U4099 ; P1_U3338
g726 nand P1_U4097 P1_U4098 P1_U4096 ; P1_U3339
g727 nand P1_U4094 P1_U4095 P1_U4093 ; P1_U3340
g728 nand P1_U4091 P1_U4092 P1_U4090 ; P1_U3341
g729 nand P1_U4088 P1_U4089 P1_U4087 ; P1_U3342
g730 nand P1_U4085 P1_U4086 P1_U4084 ; P1_U3343
g731 nand P1_U4082 P1_U4083 P1_U4081 ; P1_U3344
g732 nand P1_U4079 P1_U4080 P1_U4078 ; P1_U3345
g733 nand P1_U4076 P1_U4077 P1_U4075 ; P1_U3346
g734 nand P1_U4073 P1_U4074 P1_U4072 ; P1_U3347
g735 nand P1_U4070 P1_U4071 P1_U4069 ; P1_U3348
g736 nand P1_U4067 P1_U4068 P1_U4066 ; P1_U3349
g737 nand P1_U4064 P1_U4065 P1_U4063 ; P1_U3350
g738 nand P1_U4061 P1_U4062 P1_U4060 ; P1_U3351
g739 nand P1_U4058 P1_U4059 P1_U4057 ; P1_U3352
g740 nand P1_U4055 P1_U4056 P1_U4054 ; P1_U3353
g741 nand P1_U4052 P1_U4053 P1_U4051 ; P1_U3354
g742 nand P1_U4049 P1_U4050 P1_U4048 ; P1_U3355
g743 nand P1_U4917 P1_U4915 P1_U4918 P1_U4916 P1_U3986 ; P1_U3356
g744 nand P1_U3952 P1_STATE_REG_SCAN_IN ; P1_U3357
g745 nand P1_U3443 P1_U5778 ; P1_U3358
g746 not P1_B_REG_SCAN_IN ; P1_U3359
g747 nand P1_U5783 P1_U5782 P1_U3443 ; P1_U3360
g748 nand P1_U3048 P1_U3451 ; P1_U3361
g749 nand P1_U3047 P1_U3451 ; P1_U3362
g750 nand P1_U3453 P1_U5796 ; P1_U3363
g751 nand P1_U4042 P1_U3451 ; P1_U3364
g752 nand P1_U3047 P1_U3450 ; P1_U3365
g753 nand P1_U4042 P1_U3450 ; P1_U3366
g754 nand P1_U3049 P1_U3451 ; P1_U3367
g755 nand P1_U4001 P1_U5799 ; P1_U3368
g756 nand P1_U5799 P1_U5796 ; P1_U3369
g757 nand P1_U4044 P1_U3450 ; P1_U3370
g758 nand P1_U4002 P1_U5793 ; P1_U3371
g759 nand P1_U3451 P1_U3450 ; P1_U3372
g760 nand P1_U5799 P1_U5793 P1_U5802 ; P1_U3373
g761 nand P1_U3049 P1_U5793 ; P1_U3374
g762 nand P1_U5802 P1_U3452 ; P1_U3375
g763 nand P1_U4191 P1_U4190 P1_U4192 P1_U3594 P1_U3593 ; P1_U3376
g764 not P1_REG2_REG_0__SCAN_IN ; P1_U3377
g765 nand P1_U4210 P1_U4209 P1_U3608 P1_U3610 ; P1_U3378
g766 nand P1_U4229 P1_U4228 P1_U3612 P1_U3614 ; P1_U3379
g767 nand P1_U4248 P1_U4247 P1_U3616 P1_U3618 ; P1_U3380
g768 nand P1_U4267 P1_U4266 P1_U3620 P1_U3622 ; P1_U3381
g769 nand P1_U4286 P1_U4285 P1_U3624 P1_U3626 ; P1_U3382
g770 nand P1_U4305 P1_U4304 P1_U3628 P1_U3630 ; P1_U3383
g771 nand P1_U4324 P1_U4323 P1_U3632 P1_U3634 ; P1_U3384
g772 nand P1_U4343 P1_U4342 P1_U3636 P1_U3638 ; P1_U3385
g773 nand P1_U4362 P1_U4361 P1_U3640 P1_U3642 ; P1_U3386
g774 nand P1_U4381 P1_U4380 P1_U3644 P1_U3646 ; P1_U3387
g775 nand P1_U4400 P1_U4399 P1_U3648 P1_U3650 ; P1_U3388
g776 nand P1_U4419 P1_U4418 P1_U3652 P1_U3654 ; P1_U3389
g777 nand P1_U4438 P1_U4437 P1_U3656 P1_U3658 ; P1_U3390
g778 nand P1_U4457 P1_U4456 P1_U3660 P1_U3662 ; P1_U3391
g779 nand P1_U4476 P1_U4475 P1_U3664 P1_U3666 ; P1_U3392
g780 nand P1_U4495 P1_U4494 P1_U3668 P1_U3670 ; P1_U3393
g781 nand P1_U4514 P1_U4513 P1_U3672 P1_U3674 ; P1_U3394
g782 nand P1_U4533 P1_U4532 P1_U3676 P1_U3678 ; P1_U3395
g783 nand P1_U4552 P1_U4551 P1_U3680 P1_U3682 ; P1_U3396
g784 nand U113 P1_U3954 ; P1_U3397
g785 nand P1_U4571 P1_U4570 P1_U3684 P1_U3686 ; P1_U3398
g786 nand U112 P1_U3954 ; P1_U3399
g787 nand P1_U4590 P1_U4589 P1_U3688 P1_U3690 ; P1_U3400
g788 nand U111 P1_U3954 ; P1_U3401
g789 nand P1_U4609 P1_U4608 P1_U3692 P1_U3694 ; P1_U3402
g790 nand U110 P1_U3954 ; P1_U3403
g791 nand P1_U4628 P1_U4627 P1_U3696 P1_U3698 ; P1_U3404
g792 nand U109 P1_U3954 ; P1_U3405
g793 nand P1_U4647 P1_U4646 P1_U3700 P1_U3702 ; P1_U3406
g794 nand U108 P1_U3954 ; P1_U3407
g795 nand P1_U4666 P1_U4665 P1_U3704 P1_U3706 ; P1_U3408
g796 nand U107 P1_U3954 ; P1_U3409
g797 nand P1_U4685 P1_U4684 P1_U3708 P1_U3710 ; P1_U3410
g798 nand U106 P1_U3954 ; P1_U3411
g799 nand P1_U4704 P1_U4703 P1_U3712 P1_U3714 ; P1_U3412
g800 nand U105 P1_U3954 ; P1_U3413
g801 nand P1_U4723 P1_U4722 P1_U3716 P1_U3718 ; P1_U3414
g802 nand U104 P1_U3954 ; P1_U3415
g803 nand P1_U3723 P1_U3721 ; P1_U3416
g804 nand U102 P1_U3954 ; P1_U3417
g805 nand U101 P1_U3954 ; P1_U3418
g806 nand P1_U4041 P1_U5793 ; P1_U3419
g807 nand P1_U3022 P1_U4767 ; P1_U3420
g808 nand P1_U3998 P1_U5799 ; P1_U3421
g809 nand P1_U3048 P1_U3450 ; P1_U3422
g810 nand P1_U3047 P1_U5793 ; P1_U3423
g811 nand P1_U3993 P1_U5799 ; P1_U3424
g812 nand P1_U3441 P1_U3443 P1_U3442 ; P1_U3425
g813 nand P1_U4010 P1_U4768 ; P1_U3426
g814 nand P1_U3444 P1_STATE_REG_SCAN_IN ; P1_U3427
g815 nand P1_U3429 P1_U4931 ; P1_U3428
g816 nand P1_U4145 P1_U5786 ; P1_U3429
g817 nand P1_U4045 P1_STATE_REG_SCAN_IN ; P1_U3430
g818 nand P1_U3014 P1_U3015 ; P1_U3431
g819 not P1_R1375_U9 ; P1_U3432
g820 nand P1_U3022 P1_U3426 ; P1_U3433
g821 nand P1_U3847 P1_U3016 ; P1_U3434
g822 nand P1_U3852 P1_U5143 ; P1_U3435
g823 nand P1_U5415 P1_U5414 ; P1_U3436
g824 nand P1_U3999 P1_U3362 ; P1_U3437
g825 nand P1_U5536 P1_U3051 ; P1_U3438
g826 not P1_R1352_U6 ; P1_U3439
g827 nand P1_U3364 P1_U3423 ; P1_U3440
g828 nand P1_U5774 P1_U5773 ; P1_U3441
g829 nand P1_U5777 P1_U5776 ; P1_U3442
g830 nand P1_U5780 P1_U5779 ; P1_U3443
g831 nand P1_U5785 P1_U5784 ; P1_U3444
g832 nand P1_U5788 P1_U5787 ; P1_U3445
g833 nand P1_U5790 P1_U5789 ; P1_U3446
g834 nand P1_U5804 P1_U5803 ; P1_U3447
g835 nand P1_U5807 P1_U5806 ; P1_U3448
g836 nand P1_U5810 P1_U5809 ; P1_U3449
g837 nand P1_U5801 P1_U5800 ; P1_U3450
g838 nand P1_U5792 P1_U5791 ; P1_U3451
g839 nand P1_U5795 P1_U5794 ; P1_U3452
g840 nand P1_U5798 P1_U5797 ; P1_U3453
g841 nand P1_U5813 P1_U5812 ; P1_U3454
g842 nand P1_U5816 P1_U5815 ; P1_U3455
g843 nand P1_U5819 P1_U5818 ; P1_U3456
g844 nand P1_U5827 P1_U5826 ; P1_U3457
g845 nand P1_U5824 P1_U5823 ; P1_U3458
g846 nand P1_U5830 P1_U5829 ; P1_U3459
g847 nand P1_U5832 P1_U5831 ; P1_U3460
g848 nand P1_U5834 P1_U5833 ; P1_U3461
g849 nand P1_U5837 P1_U5836 ; P1_U3462
g850 nand P1_U5839 P1_U5838 ; P1_U3463
g851 nand P1_U5841 P1_U5840 ; P1_U3464
g852 nand P1_U5844 P1_U5843 ; P1_U3465
g853 nand P1_U5846 P1_U5845 ; P1_U3466
g854 nand P1_U5848 P1_U5847 ; P1_U3467
g855 nand P1_U5851 P1_U5850 ; P1_U3468
g856 nand P1_U5853 P1_U5852 ; P1_U3469
g857 nand P1_U5855 P1_U5854 ; P1_U3470
g858 nand P1_U5858 P1_U5857 ; P1_U3471
g859 nand P1_U5860 P1_U5859 ; P1_U3472
g860 nand P1_U5862 P1_U5861 ; P1_U3473
g861 nand P1_U5865 P1_U5864 ; P1_U3474
g862 nand P1_U5867 P1_U5866 ; P1_U3475
g863 nand P1_U5869 P1_U5868 ; P1_U3476
g864 nand P1_U5872 P1_U5871 ; P1_U3477
g865 nand P1_U5874 P1_U5873 ; P1_U3478
g866 nand P1_U5876 P1_U5875 ; P1_U3479
g867 nand P1_U5879 P1_U5878 ; P1_U3480
g868 nand P1_U5881 P1_U5880 ; P1_U3481
g869 nand P1_U5883 P1_U5882 ; P1_U3482
g870 nand P1_U5886 P1_U5885 ; P1_U3483
g871 nand P1_U5888 P1_U5887 ; P1_U3484
g872 nand P1_U5890 P1_U5889 ; P1_U3485
g873 nand P1_U5893 P1_U5892 ; P1_U3486
g874 nand P1_U5895 P1_U5894 ; P1_U3487
g875 nand P1_U5897 P1_U5896 ; P1_U3488
g876 nand P1_U5900 P1_U5899 ; P1_U3489
g877 nand P1_U5902 P1_U5901 ; P1_U3490
g878 nand P1_U5904 P1_U5903 ; P1_U3491
g879 nand P1_U5907 P1_U5906 ; P1_U3492
g880 nand P1_U5909 P1_U5908 ; P1_U3493
g881 nand P1_U5911 P1_U5910 ; P1_U3494
g882 nand P1_U5914 P1_U5913 ; P1_U3495
g883 nand P1_U5916 P1_U5915 ; P1_U3496
g884 nand P1_U5918 P1_U5917 ; P1_U3497
g885 nand P1_U5921 P1_U5920 ; P1_U3498
g886 nand P1_U5923 P1_U5922 ; P1_U3499
g887 nand P1_U5925 P1_U5924 ; P1_U3500
g888 nand P1_U5928 P1_U5927 ; P1_U3501
g889 nand P1_U5930 P1_U5929 ; P1_U3502
g890 nand P1_U5932 P1_U5931 ; P1_U3503
g891 nand P1_U5935 P1_U5934 ; P1_U3504
g892 nand P1_U5937 P1_U5936 ; P1_U3505
g893 nand P1_U5939 P1_U5938 ; P1_U3506
g894 nand P1_U5942 P1_U5941 ; P1_U3507
g895 nand P1_U5944 P1_U5943 ; P1_U3508
g896 nand P1_U5946 P1_U5945 ; P1_U3509
g897 nand P1_U5949 P1_U5948 ; P1_U3510
g898 nand P1_U5951 P1_U5950 ; P1_U3511
g899 nand P1_U5953 P1_U5952 ; P1_U3512
g900 nand P1_U5956 P1_U5955 ; P1_U3513
g901 nand P1_U5958 P1_U5957 ; P1_U3514
g902 nand P1_U5961 P1_U5960 ; P1_U3515
g903 nand P1_U5963 P1_U5962 ; P1_U3516
g904 nand P1_U5965 P1_U5964 ; P1_U3517
g905 nand P1_U5967 P1_U5966 ; P1_U3518
g906 nand P1_U5969 P1_U5968 ; P1_U3519
g907 nand P1_U5971 P1_U5970 ; P1_U3520
g908 nand P1_U5973 P1_U5972 ; P1_U3521
g909 nand P1_U5975 P1_U5974 ; P1_U3522
g910 nand P1_U5977 P1_U5976 ; P1_U3523
g911 nand P1_U5979 P1_U5978 ; P1_U3524
g912 nand P1_U5981 P1_U5980 ; P1_U3525
g913 nand P1_U5983 P1_U5982 ; P1_U3526
g914 nand P1_U5985 P1_U5984 ; P1_U3527
g915 nand P1_U5987 P1_U5986 ; P1_U3528
g916 nand P1_U5989 P1_U5988 ; P1_U3529
g917 nand P1_U5991 P1_U5990 ; P1_U3530
g918 nand P1_U5993 P1_U5992 ; P1_U3531
g919 nand P1_U5995 P1_U5994 ; P1_U3532
g920 nand P1_U5997 P1_U5996 ; P1_U3533
g921 nand P1_U5999 P1_U5998 ; P1_U3534
g922 nand P1_U6001 P1_U6000 ; P1_U3535
g923 nand P1_U6003 P1_U6002 ; P1_U3536
g924 nand P1_U6005 P1_U6004 ; P1_U3537
g925 nand P1_U6007 P1_U6006 ; P1_U3538
g926 nand P1_U6009 P1_U6008 ; P1_U3539
g927 nand P1_U6011 P1_U6010 ; P1_U3540
g928 nand P1_U6013 P1_U6012 ; P1_U3541
g929 nand P1_U6015 P1_U6014 ; P1_U3542
g930 nand P1_U6017 P1_U6016 ; P1_U3543
g931 nand P1_U6019 P1_U6018 ; P1_U3544
g932 nand P1_U6021 P1_U6020 ; P1_U3545
g933 nand P1_U6023 P1_U6022 ; P1_U3546
g934 nand P1_U6025 P1_U6024 ; P1_U3547
g935 nand P1_U6027 P1_U6026 ; P1_U3548
g936 nand P1_U6029 P1_U6028 ; P1_U3549
g937 nand P1_U6031 P1_U6030 ; P1_U3550
g938 nand P1_U6033 P1_U6032 ; P1_U3551
g939 nand P1_U6035 P1_U6034 ; P1_U3552
g940 nand P1_U6037 P1_U6036 ; P1_U3553
g941 nand P1_U6039 P1_U6038 ; P1_U3554
g942 nand P1_U6041 P1_U6040 ; P1_U3555
g943 nand P1_U6043 P1_U6042 ; P1_U3556
g944 nand P1_U6045 P1_U6044 ; P1_U3557
g945 nand P1_U6047 P1_U6046 ; P1_U3558
g946 nand P1_U6049 P1_U6048 ; P1_U3559
g947 nand P1_U6115 P1_U6114 ; P1_U3560
g948 nand P1_U6117 P1_U6116 ; P1_U3561
g949 nand P1_U6119 P1_U6118 ; P1_U3562
g950 nand P1_U6121 P1_U6120 ; P1_U3563
g951 nand P1_U6123 P1_U6122 ; P1_U3564
g952 nand P1_U6125 P1_U6124 ; P1_U3565
g953 nand P1_U6127 P1_U6126 ; P1_U3566
g954 nand P1_U6129 P1_U6128 ; P1_U3567
g955 nand P1_U6131 P1_U6130 ; P1_U3568
g956 nand P1_U6133 P1_U6132 ; P1_U3569
g957 nand P1_U6135 P1_U6134 ; P1_U3570
g958 nand P1_U6137 P1_U6136 ; P1_U3571
g959 nand P1_U6139 P1_U6138 ; P1_U3572
g960 nand P1_U6141 P1_U6140 ; P1_U3573
g961 nand P1_U6143 P1_U6142 ; P1_U3574
g962 nand P1_U6145 P1_U6144 ; P1_U3575
g963 nand P1_U6147 P1_U6146 ; P1_U3576
g964 nand P1_U6149 P1_U6148 ; P1_U3577
g965 nand P1_U6151 P1_U6150 ; P1_U3578
g966 nand P1_U6153 P1_U6152 ; P1_U3579
g967 nand P1_U6155 P1_U6154 ; P1_U3580
g968 nand P1_U6157 P1_U6156 ; P1_U3581
g969 nand P1_U6159 P1_U6158 ; P1_U3582
g970 nand P1_U6161 P1_U6160 ; P1_U3583
g971 nand P1_U6163 P1_U6162 ; P1_U3584
g972 nand P1_U6165 P1_U6164 ; P1_U3585
g973 nand P1_U6167 P1_U6166 ; P1_U3586
g974 nand P1_U6169 P1_U6168 ; P1_U3587
g975 nand P1_U6171 P1_U6170 ; P1_U3588
g976 nand P1_U6173 P1_U6172 ; P1_U3589
g977 nand P1_U6175 P1_U6174 ; P1_U3590
g978 nand P1_U6177 P1_U6176 ; P1_U3591
g979 and P1_U5786 P1_STATE_REG_SCAN_IN ; P1_U3592
g980 and P1_U4187 P1_U4186 ; P1_U3593
g981 and P1_U4189 P1_U4188 ; P1_U3594
g982 and P1_U4195 P1_U4196 ; P1_U3595
g983 and P1_U4151 P1_U4150 P1_U4149 P1_U4148 ; P1_U3596
g984 and P1_U4155 P1_U4154 P1_U4153 P1_U4152 ; P1_U3597
g985 and P1_U4159 P1_U4158 P1_U4157 P1_U4156 ; P1_U3598
g986 and P1_U4161 P1_U4160 P1_U4162 ; P1_U3599
g987 and P1_U3599 P1_U3598 P1_U3597 P1_U3596 ; P1_U3600
g988 and P1_U4166 P1_U4165 P1_U4164 P1_U4163 ; P1_U3601
g989 and P1_U4170 P1_U4169 P1_U4168 P1_U4167 ; P1_U3602
g990 and P1_U4174 P1_U4173 P1_U4172 P1_U4171 ; P1_U3603
g991 and P1_U4176 P1_U4175 P1_U4177 ; P1_U3604
g992 and P1_U3604 P1_U3603 P1_U3602 P1_U3601 ; P1_U3605
g993 and P1_U5825 P1_U4179 ; P1_U3606
g994 and P1_U5828 P1_U3022 ; P1_U3607
g995 and P1_U4212 P1_U4211 ; P1_U3608
g996 and P1_U4214 P1_U4213 ; P1_U3609
g997 and P1_U4216 P1_U4215 P1_U3609 ; P1_U3610
g998 and P1_U4220 P1_U4218 P1_U4221 P1_U4219 ; P1_U3611
g999 and P1_U4231 P1_U4230 ; P1_U3612
g1000 and P1_U4233 P1_U4232 ; P1_U3613
g1001 and P1_U4235 P1_U4234 P1_U3613 ; P1_U3614
g1002 and P1_U4239 P1_U4237 P1_U4240 P1_U4238 ; P1_U3615
g1003 and P1_U4250 P1_U4249 ; P1_U3616
g1004 and P1_U4252 P1_U4251 ; P1_U3617
g1005 and P1_U4254 P1_U4253 P1_U3617 ; P1_U3618
g1006 and P1_U4258 P1_U4256 P1_U4259 P1_U4257 ; P1_U3619
g1007 and P1_U4269 P1_U4268 ; P1_U3620
g1008 and P1_U4271 P1_U4270 ; P1_U3621
g1009 and P1_U4273 P1_U4272 P1_U3621 ; P1_U3622
g1010 and P1_U4277 P1_U4275 P1_U4278 P1_U4276 ; P1_U3623
g1011 and P1_U4288 P1_U4287 ; P1_U3624
g1012 and P1_U4290 P1_U4289 ; P1_U3625
g1013 and P1_U4292 P1_U4291 P1_U3625 ; P1_U3626
g1014 and P1_U4296 P1_U4294 P1_U4297 P1_U4295 ; P1_U3627
g1015 and P1_U4307 P1_U4306 ; P1_U3628
g1016 and P1_U4309 P1_U4308 ; P1_U3629
g1017 and P1_U4311 P1_U4310 P1_U3629 ; P1_U3630
g1018 and P1_U4315 P1_U4313 P1_U4316 P1_U4314 ; P1_U3631
g1019 and P1_U4326 P1_U4325 ; P1_U3632
g1020 and P1_U4328 P1_U4327 ; P1_U3633
g1021 and P1_U4330 P1_U4329 P1_U3633 ; P1_U3634
g1022 and P1_U4334 P1_U4332 P1_U4335 P1_U4333 ; P1_U3635
g1023 and P1_U4345 P1_U4344 ; P1_U3636
g1024 and P1_U4347 P1_U4346 ; P1_U3637
g1025 and P1_U4349 P1_U4348 P1_U3637 ; P1_U3638
g1026 and P1_U4353 P1_U4351 P1_U4354 P1_U4352 ; P1_U3639
g1027 and P1_U4364 P1_U4363 ; P1_U3640
g1028 and P1_U4366 P1_U4365 ; P1_U3641
g1029 and P1_U4368 P1_U4367 P1_U3641 ; P1_U3642
g1030 and P1_U4372 P1_U4370 P1_U4373 P1_U4371 ; P1_U3643
g1031 and P1_U4383 P1_U4382 ; P1_U3644
g1032 and P1_U4385 P1_U4384 ; P1_U3645
g1033 and P1_U4387 P1_U4386 P1_U3645 ; P1_U3646
g1034 and P1_U4391 P1_U4389 P1_U4392 P1_U4390 ; P1_U3647
g1035 and P1_U4402 P1_U4401 ; P1_U3648
g1036 and P1_U4404 P1_U4403 ; P1_U3649
g1037 and P1_U4406 P1_U4405 P1_U3649 ; P1_U3650
g1038 and P1_U4411 P1_U4410 P1_U4409 P1_U4408 ; P1_U3651
g1039 and P1_U4421 P1_U4420 ; P1_U3652
g1040 and P1_U4423 P1_U4422 ; P1_U3653
g1041 and P1_U4425 P1_U4424 P1_U3653 ; P1_U3654
g1042 and P1_U4430 P1_U4428 P1_U4429 P1_U4427 ; P1_U3655
g1043 and P1_U4440 P1_U4439 ; P1_U3656
g1044 and P1_U4442 P1_U4441 ; P1_U3657
g1045 and P1_U4444 P1_U4443 P1_U3657 ; P1_U3658
g1046 and P1_U4449 P1_U4448 P1_U4447 P1_U4446 ; P1_U3659
g1047 and P1_U4459 P1_U4458 ; P1_U3660
g1048 and P1_U4461 P1_U4460 ; P1_U3661
g1049 and P1_U4463 P1_U4462 P1_U3661 ; P1_U3662
g1050 and P1_U4468 P1_U4466 P1_U4467 P1_U4465 ; P1_U3663
g1051 and P1_U4478 P1_U4477 ; P1_U3664
g1052 and P1_U4480 P1_U4479 ; P1_U3665
g1053 and P1_U4482 P1_U4481 P1_U3665 ; P1_U3666
g1054 and P1_U4486 P1_U4484 P1_U4487 P1_U4485 ; P1_U3667
g1055 and P1_U4497 P1_U4496 ; P1_U3668
g1056 and P1_U4499 P1_U4498 ; P1_U3669
g1057 and P1_U4501 P1_U4500 P1_U3669 ; P1_U3670
g1058 and P1_U4505 P1_U4503 P1_U4506 P1_U4504 ; P1_U3671
g1059 and P1_U4516 P1_U4515 ; P1_U3672
g1060 and P1_U4518 P1_U4517 ; P1_U3673
g1061 and P1_U4520 P1_U4519 P1_U3673 ; P1_U3674
g1062 and P1_U4525 P1_U4523 P1_U4524 P1_U4522 ; P1_U3675
g1063 and P1_U4535 P1_U4534 ; P1_U3676
g1064 and P1_U4537 P1_U4536 ; P1_U3677
g1065 and P1_U4539 P1_U4538 P1_U3677 ; P1_U3678
g1066 and P1_U4544 P1_U4542 P1_U4543 P1_U4541 ; P1_U3679
g1067 and P1_U4554 P1_U4553 ; P1_U3680
g1068 and P1_U4556 P1_U4555 ; P1_U3681
g1069 and P1_U4558 P1_U4557 P1_U3681 ; P1_U3682
g1070 and P1_U4562 P1_U4560 P1_U4563 P1_U4561 ; P1_U3683
g1071 and P1_U4573 P1_U4572 ; P1_U3684
g1072 and P1_U4575 P1_U4574 ; P1_U3685
g1073 and P1_U4577 P1_U4576 P1_U3685 ; P1_U3686
g1074 and P1_U4581 P1_U4579 P1_U4582 P1_U4580 ; P1_U3687
g1075 and P1_U4592 P1_U4591 ; P1_U3688
g1076 and P1_U4594 P1_U4593 ; P1_U3689
g1077 and P1_U4596 P1_U4595 P1_U3689 ; P1_U3690
g1078 and P1_U4600 P1_U4598 P1_U4601 P1_U4599 ; P1_U3691
g1079 and P1_U4611 P1_U4610 ; P1_U3692
g1080 and P1_U4613 P1_U4612 ; P1_U3693
g1081 and P1_U4615 P1_U4614 P1_U3693 ; P1_U3694
g1082 and P1_U4619 P1_U4617 P1_U4620 P1_U4618 ; P1_U3695
g1083 and P1_U4630 P1_U4629 ; P1_U3696
g1084 and P1_U4632 P1_U4631 ; P1_U3697
g1085 and P1_U4634 P1_U4633 P1_U3697 ; P1_U3698
g1086 and P1_U4638 P1_U4636 P1_U4639 P1_U4637 ; P1_U3699
g1087 and P1_U4649 P1_U4648 ; P1_U3700
g1088 and P1_U4651 P1_U4650 ; P1_U3701
g1089 and P1_U4653 P1_U4652 P1_U3701 ; P1_U3702
g1090 and P1_U4657 P1_U4655 P1_U4658 P1_U4656 ; P1_U3703
g1091 and P1_U4668 P1_U4667 ; P1_U3704
g1092 and P1_U4670 P1_U4669 ; P1_U3705
g1093 and P1_U4672 P1_U4671 P1_U3705 ; P1_U3706
g1094 and P1_U4676 P1_U4674 P1_U4677 P1_U4675 ; P1_U3707
g1095 and P1_U4687 P1_U4686 ; P1_U3708
g1096 and P1_U4689 P1_U4688 ; P1_U3709
g1097 and P1_U4691 P1_U4690 P1_U3709 ; P1_U3710
g1098 and P1_U4695 P1_U4693 P1_U4696 P1_U4694 ; P1_U3711
g1099 and P1_U4706 P1_U4705 ; P1_U3712
g1100 and P1_U4708 P1_U4707 ; P1_U3713
g1101 and P1_U4710 P1_U4709 P1_U3713 ; P1_U3714
g1102 and P1_U4714 P1_U4712 P1_U4715 P1_U4713 ; P1_U3715
g1103 and P1_U4725 P1_U4724 ; P1_U3716
g1104 and P1_U4727 P1_U4726 ; P1_U3717
g1105 and P1_U4729 P1_U4728 P1_U3717 ; P1_U3718
g1106 and P1_U4733 P1_U4731 P1_U4734 P1_U4732 ; P1_U3719
g1107 and P1_U4741 P1_U4030 ; P1_U3720
g1108 and P1_U4743 P1_U4742 P1_U4744 P1_U4745 P1_U4746 ; P1_U3721
g1109 and P1_U4748 P1_U4747 ; P1_U3722
g1110 and P1_U4750 P1_U4749 P1_U3722 ; P1_U3723
g1111 and P1_U4753 P1_U4754 P1_U4752 ; P1_U3724
g1112 and P1_U4030 P1_U4741 ; P1_U3725
g1113 and P1_U3022 P1_U3457 ; P1_U3726
g1114 and P1_U5828 P1_U4012 P1_U3458 ; P1_U3727
g1115 and P1_U4771 P1_U4770 P1_U4772 ; P1_U3728
g1116 and P1_U4774 P1_U4773 P1_U3957 ; P1_U3729
g1117 and P1_U4776 P1_U4775 P1_U4777 ; P1_U3730
g1118 and P1_U4779 P1_U4778 P1_U3958 ; P1_U3731
g1119 and P1_U4781 P1_U4780 P1_U4782 ; P1_U3732
g1120 and P1_U4784 P1_U4783 P1_U3959 ; P1_U3733
g1121 and P1_U4786 P1_U4785 P1_U4787 ; P1_U3734
g1122 and P1_U4789 P1_U4788 P1_U3960 ; P1_U3735
g1123 and P1_U4791 P1_U4790 P1_U4792 ; P1_U3736
g1124 and P1_U4794 P1_U4793 P1_U3961 ; P1_U3737
g1125 and P1_U4796 P1_U4795 P1_U4797 ; P1_U3738
g1126 and P1_U4799 P1_U4798 ; P1_U3739
g1127 and P1_U4801 P1_U4800 P1_U4802 ; P1_U3740
g1128 and P1_U4804 P1_U4803 ; P1_U3741
g1129 and P1_U4806 P1_U4805 P1_U4807 ; P1_U3742
g1130 and P1_U4809 P1_U4808 ; P1_U3743
g1131 and P1_U4811 P1_U4810 P1_U4812 ; P1_U3744
g1132 and P1_U4814 P1_U4813 ; P1_U3745
g1133 and P1_U4816 P1_U4815 ; P1_U3746
g1134 and P1_U4819 P1_U4818 ; P1_U3747
g1135 and P1_U4821 P1_U4820 ; P1_U3748
g1136 and P1_U4824 P1_U4823 ; P1_U3749
g1137 and P1_U4826 P1_U4825 P1_U4827 ; P1_U3750
g1138 and P1_U4829 P1_U4828 ; P1_U3751
g1139 and P1_U4831 P1_U4830 P1_U4832 ; P1_U3752
g1140 and P1_U4834 P1_U4833 ; P1_U3753
g1141 and P1_U4836 P1_U4835 P1_U4837 ; P1_U3754
g1142 and P1_U4839 P1_U4838 ; P1_U3755
g1143 and P1_U4841 P1_U4840 P1_U4842 ; P1_U3756
g1144 and P1_U4844 P1_U4843 ; P1_U3757
g1145 and P1_U4846 P1_U4845 ; P1_U3758
g1146 and P1_U4849 P1_U4848 ; P1_U3759
g1147 and P1_U4851 P1_U4850 ; P1_U3760
g1148 and P1_U4854 P1_U4853 ; P1_U3761
g1149 and P1_U4856 P1_U4855 P1_U4857 ; P1_U3762
g1150 and P1_U4859 P1_U4858 ; P1_U3763
g1151 and P1_U4861 P1_U4860 P1_U4862 ; P1_U3764
g1152 and P1_U4864 P1_U4863 ; P1_U3765
g1153 and P1_U4866 P1_U4865 ; P1_U3766
g1154 and P1_U4869 P1_U4868 ; P1_U3767
g1155 and P1_U4871 P1_U4870 ; P1_U3768
g1156 and P1_U4874 P1_U4873 ; P1_U3769
g1157 and P1_U4876 P1_U4875 ; P1_U3770
g1158 and P1_U4879 P1_U4878 ; P1_U3771
g1159 and P1_U4881 P1_U4880 ; P1_U3772
g1160 and P1_U4884 P1_U4883 ; P1_U3773
g1161 and P1_U4886 P1_U4885 ; P1_U3774
g1162 and P1_U4889 P1_U4888 ; P1_U3775
g1163 and P1_U4891 P1_U4890 ; P1_U3776
g1164 and P1_U4894 P1_U4893 ; P1_U3777
g1165 and P1_U4896 P1_U4895 ; P1_U3778
g1166 and P1_U4899 P1_U4898 ; P1_U3779
g1167 and P1_U4901 P1_U4900 ; P1_U3780
g1168 and P1_U4904 P1_U4903 ; P1_U3781
g1169 and P1_U4906 P1_U4905 ; P1_U3782
g1170 and P1_U4909 P1_U4908 ; P1_U3783
g1171 and P1_U4911 P1_U4910 ; P1_U3784
g1172 and P1_U4914 P1_U4913 ; P1_U3785
g1173 and P1_U3362 P1_U3364 P1_U3370 ; P1_U3786
g1174 and P1_U3366 P1_U3422 P1_U3365 ; P1_U3787
g1175 and P1_U3361 P1_U4006 ; P1_U3788
g1176 and P1_U3788 P1_U3424 ; P1_U3789
g1177 and P1_U4934 P1_U4935 ; P1_U3790
g1178 and P1_U4938 P1_U4936 P1_U4937 ; P1_U3791
g1179 and P1_U4944 P1_U4945 ; P1_U3792
g1180 and P1_U4948 P1_U4946 P1_U4947 ; P1_U3793
g1181 and P1_U4954 P1_U4955 ; P1_U3794
g1182 and P1_U4958 P1_U4956 P1_U4957 ; P1_U3795
g1183 and P1_U4964 P1_U4965 ; P1_U3796
g1184 and P1_U4968 P1_U4966 P1_U4967 ; P1_U3797
g1185 and P1_U4974 P1_U4975 ; P1_U3798
g1186 and P1_U4978 P1_U4976 P1_U4977 ; P1_U3799
g1187 and P1_U4984 P1_U4985 ; P1_U3800
g1188 and P1_U4988 P1_U4986 P1_U4987 ; P1_U3801
g1189 and P1_U4994 P1_U4995 ; P1_U3802
g1190 and P1_U4998 P1_U4996 P1_U4997 ; P1_U3803
g1191 and P1_U5004 P1_U5005 ; P1_U3804
g1192 and P1_U5008 P1_U5006 P1_U5007 ; P1_U3805
g1193 and P1_U5014 P1_U5015 ; P1_U3806
g1194 and P1_U5018 P1_U5016 P1_U5017 ; P1_U3807
g1195 and P1_U5024 P1_U5025 ; P1_U3808
g1196 and P1_U5028 P1_U5026 P1_U5027 ; P1_U3809
g1197 and P1_U5034 P1_U5035 ; P1_U3810
g1198 and P1_U5038 P1_U5036 P1_U5037 ; P1_U3811
g1199 and P1_U5044 P1_U5045 ; P1_U3812
g1200 and P1_U5048 P1_U5046 P1_U5047 ; P1_U3813
g1201 and P1_U5054 P1_U5055 ; P1_U3814
g1202 and P1_U5058 P1_U5056 P1_U5057 ; P1_U3815
g1203 and P1_U5064 P1_U5065 ; P1_U3816
g1204 and P1_U5067 P1_U5066 P1_U5068 ; P1_U3817
g1205 and P1_U5074 P1_U5075 ; P1_U3818
g1206 and P1_U5077 P1_U5076 P1_U5078 ; P1_U3819
g1207 and P1_U3821 P1_U5084 ; P1_U3820
g1208 and P1_U5085 P1_U4040 ; P1_U3821
g1209 and P1_U5087 P1_U5086 P1_U5088 ; P1_U3822
g1210 and P1_U5094 P1_U5095 ; P1_U3823
g1211 and P1_U5097 P1_U5096 P1_U5098 ; P1_U3824
g1212 and P1_U3826 P1_U5104 ; P1_U3825
g1213 and P1_U5105 P1_U4040 ; P1_U3826
g1214 and P1_U5107 P1_U5106 P1_U5108 ; P1_U3827
g1215 and P1_U5114 P1_U5115 ; P1_U3828
g1216 and P1_U5117 P1_U5116 P1_U5118 ; P1_U3829
g1217 and P1_U5124 P1_U5125 ; P1_U3830
g1218 and P1_U5127 P1_U5126 P1_U5128 ; P1_U3831
g1219 and P1_U6218 P1_U6215 P1_U6221 ; P1_U3832
g1220 and P1_U3834 P1_U3832 P1_U6233 ; P1_U3833
g1221 and P1_U6230 P1_U6227 P1_U6224 ; P1_U3834
g1222 and P1_U6242 P1_U6239 P1_U6245 ; P1_U3835
g1223 and P1_U6251 P1_U6248 P1_U6254 ; P1_U3836
g1224 and P1_U3836 P1_U3835 P1_U6236 ; P1_U3837
g1225 and P1_U6188 P1_U6185 P1_U6191 ; P1_U3838
g1226 and P1_U6203 P1_U6200 P1_U6197 P1_U6194 P1_U6206 ; P1_U3839
g1227 and P1_U6269 P1_U6266 P1_U6263 P1_U6260 ; P1_U3840
g1228 and P1_U6275 P1_U6272 ; P1_U3841
g1229 and P1_U3841 P1_U3840 ; P1_U3842
g1230 and P1_U3837 P1_U3833 P1_U6212 P1_U6257 P1_U6209 ; P1_U3843
g1231 and P1_U3839 P1_U3838 P1_U6182 ; P1_U3844
g1232 and P1_U3429 P1_STATE_REG_SCAN_IN ; P1_U3845
g1233 and P1_U5138 P1_U5136 ; P1_U3846
g1234 and P1_U3457 P1_U3458 ; P1_U3847
g1235 and P1_U3997 P1_U3371 P1_U3996 ; P1_U3848
g1236 and P1_U3368 P1_U3424 ; P1_U3849
g1237 and P1_U3427 P1_U3430 ; P1_U3850
g1238 and P1_U3022 P1_U5145 ; P1_U3851
g1239 and P1_U3425 P1_STATE_REG_SCAN_IN ; P1_U3852
g1240 and P1_U5173 P1_U5172 ; P1_U3853
g1241 and P1_U5189 P1_U5187 ; P1_U3854
g1242 and P1_U5191 P1_U5190 ; P1_U3855
g1243 and P1_U5200 P1_U5199 ; P1_U3856
g1244 and P1_U5218 P1_U5217 ; P1_U3857
g1245 and P1_U4037 P1_U3078 ; P1_U3858
g1246 and P1_U5232 P1_U5231 P1_U3860 ; P1_U3859
g1247 and P1_U5235 P1_U5234 ; P1_U3860
g1248 and P1_U5244 P1_U5243 ; P1_U3861
g1249 and P1_U5251 P1_U5249 ; P1_U3862
g1250 and P1_U5253 P1_U5252 ; P1_U3863
g1251 and P1_U5280 P1_U5279 ; P1_U3864
g1252 and P1_U5307 P1_U5306 ; P1_U3865
g1253 and P1_U5323 P1_U5321 ; P1_U3866
g1254 and P1_U5325 P1_U5324 ; P1_U3867
g1255 and P1_U5334 P1_U5333 ; P1_U3868
g1256 and P1_U5359 P1_U5357 ; P1_U3869
g1257 and P1_U5361 P1_U5360 ; P1_U3870
g1258 and P1_U5370 P1_U5369 ; P1_U3871
g1259 and P1_U5406 P1_U5405 ; P1_U3872
g1260 and P1_U5802 P1_U5793 ; P1_U3873
g1261 and P1_U3375 P1_U5410 ; P1_U3874
g1262 and P1_U5475 P1_U5476 ; P1_U3875
g1263 and P1_U5535 P1_U5533 ; P1_U3876
g1264 and P1_U3444 P1_U5538 ; P1_U3877
g1265 and P1_U3374 P1_U3997 ; P1_U3878
g1266 and P1_U3878 P1_U3371 ; P1_U3879
g1267 and P1_U3881 P1_U5546 ; P1_U3880
g1268 and P1_U3444 P1_U5544 ; P1_U3881
g1269 and P1_U3883 P1_U5549 ; P1_U3882
g1270 and P1_U3444 P1_U5547 ; P1_U3883
g1271 and P1_U3885 P1_U5552 ; P1_U3884
g1272 and P1_U3444 P1_U5550 ; P1_U3885
g1273 and P1_U3887 P1_U5555 ; P1_U3886
g1274 and P1_U3444 P1_U5553 ; P1_U3887
g1275 and P1_U3889 P1_U5558 ; P1_U3888
g1276 and P1_U3444 P1_U5556 ; P1_U3889
g1277 and P1_U3891 P1_U5561 ; P1_U3890
g1278 and P1_U3444 P1_U5559 ; P1_U3891
g1279 and P1_U5564 P1_U5562 ; P1_U3892
g1280 and P1_U5567 P1_U5565 ; P1_U3893
g1281 and P1_U3895 P1_U5570 ; P1_U3894
g1282 and P1_U3444 P1_U5568 ; P1_U3895
g1283 and P1_U3444 P1_U5573 ; P1_U3896
g1284 and P1_U3444 P1_U5576 ; P1_U3897
g1285 and P1_U3444 P1_U5579 ; P1_U3898
g1286 and P1_U3444 P1_U5582 ; P1_U3899
g1287 and P1_U3444 P1_U5585 ; P1_U3900
g1288 and P1_U3444 P1_U5588 ; P1_U3901
g1289 and P1_U3444 P1_U5591 ; P1_U3902
g1290 and P1_U3444 P1_U5594 ; P1_U3903
g1291 and P1_U3444 P1_U5597 ; P1_U3904
g1292 and P1_U3444 P1_U5600 ; P1_U3905
g1293 and P1_U3907 P1_U5603 ; P1_U3906
g1294 and P1_U3444 P1_U5601 ; P1_U3907
g1295 and P1_U3444 P1_U5606 ; P1_U3908
g1296 and P1_U3444 P1_U5609 ; P1_U3909
g1297 and P1_U3444 P1_U5612 ; P1_U3910
g1298 and P1_U3444 P1_U5615 ; P1_U3911
g1299 and P1_U3444 P1_U5618 ; P1_U3912
g1300 and P1_U3444 P1_U5621 ; P1_U3913
g1301 and P1_U3444 P1_U5624 ; P1_U3914
g1302 and P1_U3444 P1_U5627 ; P1_U3915
g1303 and P1_U3444 P1_U5630 ; P1_U3916
g1304 and P1_U3444 P1_U5633 ; P1_U3917
g1305 and P1_U3919 P1_U5636 ; P1_U3918
g1306 and P1_U3444 P1_U5634 ; P1_U3919
g1307 and P1_U3921 P1_U5639 ; P1_U3920
g1308 and P1_U3444 P1_U5637 ; P1_U3921
g1309 and P1_U5645 P1_U5642 ; P1_U3922
g1310 and P1_U5649 P1_U5646 ; P1_U3923
g1311 and P1_U5651 P1_U5650 ; P1_U3924
g1312 and P1_U5655 P1_U5654 ; P1_U3925
g1313 and P1_U5659 P1_U5658 ; P1_U3926
g1314 and P1_U5663 P1_U5662 ; P1_U3927
g1315 and P1_U5673 P1_U5672 P1_U5675 ; P1_U3928
g1316 and P1_U5677 P1_U5676 ; P1_U3929
g1317 and P1_U5681 P1_U5680 ; P1_U3930
g1318 and P1_U5685 P1_U5684 ; P1_U3931
g1319 and P1_U5689 P1_U5688 ; P1_U3932
g1320 and P1_U5693 P1_U5692 ; P1_U3933
g1321 and P1_U5697 P1_U5696 ; P1_U3934
g1322 and P1_U5701 P1_U5700 ; P1_U3935
g1323 and P1_U5705 P1_U5704 ; P1_U3936
g1324 and P1_U5709 P1_U5708 ; P1_U3937
g1325 and P1_U5713 P1_U5712 ; P1_U3938
g1326 and P1_U5717 P1_U5716 P1_U5719 ; P1_U3939
g1327 and P1_U5721 P1_U5720 ; P1_U3940
g1328 and P1_U5725 P1_U5724 ; P1_U3941
g1329 and P1_U5729 P1_U5728 ; P1_U3942
g1330 and P1_U5733 P1_U5732 ; P1_U3943
g1331 and P1_U5737 P1_U5736 ; P1_U3944
g1332 and P1_U5741 P1_U5740 ; P1_U3945
g1333 and P1_U5745 P1_U5744 ; P1_U3946
g1334 and P1_U5749 P1_U5748 ; P1_U3947
g1335 and P1_U5753 P1_U5752 ; P1_U3948
g1336 and P1_U5757 P1_U5756 ; P1_U3949
g1337 and P1_U5761 P1_U5760 P1_U5763 ; P1_U3950
g1338 and P1_U5765 P1_U5764 ; P1_U3951
g1339 not P1_IR_REG_31__SCAN_IN ; P1_U3952
g1340 nand P1_U3022 P1_U3360 ; P1_U3953
g1341 nand P1_U5817 P1_U5811 ; P1_U3954
g1342 nand P1_U3607 P1_U3046 ; P1_U3955
g1343 nand P1_U3726 P1_U3046 ; P1_U3956
g1344 and P1_U6051 P1_U6050 ; P1_U3957
g1345 and P1_U6053 P1_U6052 ; P1_U3958
g1346 and P1_U6055 P1_U6054 ; P1_U3959
g1347 and P1_U6057 P1_U6056 ; P1_U3960
g1348 and P1_U6059 P1_U6058 ; P1_U3961
g1349 and P1_U6061 P1_U6060 ; P1_U3962
g1350 and P1_U6063 P1_U6062 ; P1_U3963
g1351 and P1_U6065 P1_U6064 ; P1_U3964
g1352 and P1_U6067 P1_U6066 ; P1_U3965
g1353 and P1_U6069 P1_U6068 ; P1_U3966
g1354 and P1_U6071 P1_U6070 ; P1_U3967
g1355 and P1_U6073 P1_U6072 ; P1_U3968
g1356 and P1_U6075 P1_U6074 ; P1_U3969
g1357 and P1_U6077 P1_U6076 ; P1_U3970
g1358 and P1_U6079 P1_U6078 ; P1_U3971
g1359 and P1_U6081 P1_U6080 ; P1_U3972
g1360 and P1_U6083 P1_U6082 ; P1_U3973
g1361 and P1_U6085 P1_U6084 ; P1_U3974
g1362 and P1_U6087 P1_U6086 ; P1_U3975
g1363 and P1_U6089 P1_U6088 ; P1_U3976
g1364 and P1_U6091 P1_U6090 ; P1_U3977
g1365 and P1_U6093 P1_U6092 ; P1_U3978
g1366 and P1_U6095 P1_U6094 ; P1_U3979
g1367 and P1_U6097 P1_U6096 ; P1_U3980
g1368 and P1_U6099 P1_U6098 ; P1_U3981
g1369 and P1_U6101 P1_U6100 ; P1_U3982
g1370 and P1_U6103 P1_U6102 ; P1_U3983
g1371 and P1_U6105 P1_U6104 ; P1_U3984
g1372 and P1_U6107 P1_U6106 ; P1_U3985
g1373 and P1_U6109 P1_U6108 ; P1_U3986
g1374 nand P1_U3725 P1_U3056 ; P1_U3987
g1375 and P1_U6111 P1_U6110 ; P1_U3988
g1376 and P1_U6113 P1_U6112 ; P1_U3989
g1377 and P1_U6179 P1_U6178 ; P1_U3990
g1378 nand P1_U3842 P1_U3843 P1_U3844 ; P1_U3991
g1379 not P1_U3371 ; P1_U3992
g1380 not P1_U3374 ; P1_U3993
g1381 not P1_U3364 ; P1_U3994
g1382 not P1_U3423 ; P1_U3995
g1383 nand P1_U4003 P1_U5793 ; P1_U3996
g1384 nand P1_U4041 P1_U3451 ; P1_U3997
g1385 not P1_U3419 ; P1_U3998
g1386 nand P1_U4042 P1_U5793 ; P1_U3999
g1387 not P1_U3362 ; P1_U4000
g1388 not P1_U3367 ; P1_U4001
g1389 not P1_U3370 ; P1_U4002
g1390 not P1_U3422 ; P1_U4003
g1391 not P1_U3366 ; P1_U4004
g1392 not P1_U3365 ; P1_U4005
g1393 nand P1_U4044 P1_U3451 ; P1_U4006
g1394 not P1_U3361 ; P1_U4007
g1395 not P1_U3424 ; P1_U4008
g1396 not P1_U3421 ; P1_U4009
g1397 nand P1_U3993 P1_U3453 ; P1_U4010
g1398 not P1_U3368 ; P1_U4011
g1399 nand P1_U4030 P1_U3369 ; P1_U4012
g1400 nand P1_U3873 P1_U3425 ; P1_U4013
g1401 not P1_U3954 ; P1_U4014
g1402 not P1_U3434 ; P1_U4015
g1403 not P1_U3430 ; P1_U4016
g1404 not P1_U3413 ; P1_U4017
g1405 not P1_U3411 ; P1_U4018
g1406 not P1_U3409 ; P1_U4019
g1407 not P1_U3407 ; P1_U4020
g1408 not P1_U3405 ; P1_U4021
g1409 not P1_U3403 ; P1_U4022
g1410 not P1_U3401 ; P1_U4023
g1411 not P1_U3399 ; P1_U4024
g1412 not P1_U3397 ; P1_U4025
g1413 not P1_U3418 ; P1_U4026
g1414 not P1_U3417 ; P1_U4027
g1415 not P1_U3415 ; P1_U4028
g1416 not P1_U3431 ; P1_U4029
g1417 not P1_U3372 ; P1_U4030
g1418 not P1_U3420 ; P1_U4031
g1419 not P1_U3956 ; P1_U4032
g1420 not P1_U3955 ; P1_U4033
g1421 not P1_U3953 ; P1_U4034
g1422 not P1_U3987 ; P1_U4035
g1423 not P1_U3373 ; P1_U4036
g1424 not P1_U3435 ; P1_U4037
g1425 not P1_U3433 ; P1_U4038
g1426 nand P1_U4009 P1_U3022 ; P1_U4039
g1427 nand P1_U4016 P1_U3212 ; P1_U4040
g1428 not P1_U3375 ; P1_U4041
g1429 not P1_U3363 ; P1_U4042
g1430 not P1_U3427 ; P1_U4043
g1431 not P1_U3369 ; P1_U4044
g1432 not P1_U3429 ; P1_U4045
g1433 not P1_U3358 ; P1_U4046
g1434 not P1_U3357 ; P1_U4047
g1435 nand U125 P1_U3086 ; P1_U4048
g1436 nand P1_U3029 P1_IR_REG_0__SCAN_IN ; P1_U4049
g1437 nand P1_U4047 P1_IR_REG_0__SCAN_IN ; P1_U4050
g1438 nand U114 P1_U3086 ; P1_U4051
g1439 nand P1_SUB_88_U40 P1_U3029 ; P1_U4052
g1440 nand P1_U4047 P1_IR_REG_1__SCAN_IN ; P1_U4053
g1441 nand U103 P1_U3086 ; P1_U4054
g1442 nand P1_SUB_88_U21 P1_U3029 ; P1_U4055
g1443 nand P1_U4047 P1_IR_REG_2__SCAN_IN ; P1_U4056
g1444 nand U100 P1_U3086 ; P1_U4057
g1445 nand P1_SUB_88_U22 P1_U3029 ; P1_U4058
g1446 nand P1_U4047 P1_IR_REG_3__SCAN_IN ; P1_U4059
g1447 nand U99 P1_U3086 ; P1_U4060
g1448 nand P1_SUB_88_U23 P1_U3029 ; P1_U4061
g1449 nand P1_U4047 P1_IR_REG_4__SCAN_IN ; P1_U4062
g1450 nand U98 P1_U3086 ; P1_U4063
g1451 nand P1_SUB_88_U162 P1_U3029 ; P1_U4064
g1452 nand P1_U4047 P1_IR_REG_5__SCAN_IN ; P1_U4065
g1453 nand U97 P1_U3086 ; P1_U4066
g1454 nand P1_SUB_88_U24 P1_U3029 ; P1_U4067
g1455 nand P1_U4047 P1_IR_REG_6__SCAN_IN ; P1_U4068
g1456 nand U96 P1_U3086 ; P1_U4069
g1457 nand P1_SUB_88_U25 P1_U3029 ; P1_U4070
g1458 nand P1_U4047 P1_IR_REG_7__SCAN_IN ; P1_U4071
g1459 nand U95 P1_U3086 ; P1_U4072
g1460 nand P1_SUB_88_U26 P1_U3029 ; P1_U4073
g1461 nand P1_U4047 P1_IR_REG_8__SCAN_IN ; P1_U4074
g1462 nand U94 P1_U3086 ; P1_U4075
g1463 nand P1_SUB_88_U160 P1_U3029 ; P1_U4076
g1464 nand P1_U4047 P1_IR_REG_9__SCAN_IN ; P1_U4077
g1465 nand U124 P1_U3086 ; P1_U4078
g1466 nand P1_SUB_88_U6 P1_U3029 ; P1_U4079
g1467 nand P1_U4047 P1_IR_REG_10__SCAN_IN ; P1_U4080
g1468 nand U123 P1_U3086 ; P1_U4081
g1469 nand P1_SUB_88_U7 P1_U3029 ; P1_U4082
g1470 nand P1_U4047 P1_IR_REG_11__SCAN_IN ; P1_U4083
g1471 nand U122 P1_U3086 ; P1_U4084
g1472 nand P1_SUB_88_U8 P1_U3029 ; P1_U4085
g1473 nand P1_U4047 P1_IR_REG_12__SCAN_IN ; P1_U4086
g1474 nand U121 P1_U3086 ; P1_U4087
g1475 nand P1_SUB_88_U179 P1_U3029 ; P1_U4088
g1476 nand P1_U4047 P1_IR_REG_13__SCAN_IN ; P1_U4089
g1477 nand U120 P1_U3086 ; P1_U4090
g1478 nand P1_SUB_88_U9 P1_U3029 ; P1_U4091
g1479 nand P1_U4047 P1_IR_REG_14__SCAN_IN ; P1_U4092
g1480 nand U119 P1_U3086 ; P1_U4093
g1481 nand P1_SUB_88_U10 P1_U3029 ; P1_U4094
g1482 nand P1_U4047 P1_IR_REG_15__SCAN_IN ; P1_U4095
g1483 nand U118 P1_U3086 ; P1_U4096
g1484 nand P1_SUB_88_U11 P1_U3029 ; P1_U4097
g1485 nand P1_U4047 P1_IR_REG_16__SCAN_IN ; P1_U4098
g1486 nand U117 P1_U3086 ; P1_U4099
g1487 nand P1_SUB_88_U177 P1_U3029 ; P1_U4100
g1488 nand P1_U4047 P1_IR_REG_17__SCAN_IN ; P1_U4101
g1489 nand U116 P1_U3086 ; P1_U4102
g1490 nand P1_SUB_88_U12 P1_U3029 ; P1_U4103
g1491 nand P1_U4047 P1_IR_REG_18__SCAN_IN ; P1_U4104
g1492 nand U115 P1_U3086 ; P1_U4105
g1493 nand P1_SUB_88_U13 P1_U3029 ; P1_U4106
g1494 nand P1_U4047 P1_IR_REG_19__SCAN_IN ; P1_U4107
g1495 nand U113 P1_U3086 ; P1_U4108
g1496 nand P1_SUB_88_U14 P1_U3029 ; P1_U4109
g1497 nand P1_U4047 P1_IR_REG_20__SCAN_IN ; P1_U4110
g1498 nand U112 P1_U3086 ; P1_U4111
g1499 nand P1_SUB_88_U173 P1_U3029 ; P1_U4112
g1500 nand P1_U4047 P1_IR_REG_21__SCAN_IN ; P1_U4113
g1501 nand U111 P1_U3086 ; P1_U4114
g1502 nand P1_SUB_88_U15 P1_U3029 ; P1_U4115
g1503 nand P1_U4047 P1_IR_REG_22__SCAN_IN ; P1_U4116
g1504 nand U110 P1_U3086 ; P1_U4117
g1505 nand P1_SUB_88_U16 P1_U3029 ; P1_U4118
g1506 nand P1_U4047 P1_IR_REG_23__SCAN_IN ; P1_U4119
g1507 nand U109 P1_U3086 ; P1_U4120
g1508 nand P1_SUB_88_U17 P1_U3029 ; P1_U4121
g1509 nand P1_U4047 P1_IR_REG_24__SCAN_IN ; P1_U4122
g1510 nand U108 P1_U3086 ; P1_U4123
g1511 nand P1_SUB_88_U170 P1_U3029 ; P1_U4124
g1512 nand P1_U4047 P1_IR_REG_25__SCAN_IN ; P1_U4125
g1513 nand U107 P1_U3086 ; P1_U4126
g1514 nand P1_SUB_88_U18 P1_U3029 ; P1_U4127
g1515 nand P1_U4047 P1_IR_REG_26__SCAN_IN ; P1_U4128
g1516 nand U106 P1_U3086 ; P1_U4129
g1517 nand P1_SUB_88_U42 P1_U3029 ; P1_U4130
g1518 nand P1_U4047 P1_IR_REG_27__SCAN_IN ; P1_U4131
g1519 nand U105 P1_U3086 ; P1_U4132
g1520 nand P1_SUB_88_U19 P1_U3029 ; P1_U4133
g1521 nand P1_U4047 P1_IR_REG_28__SCAN_IN ; P1_U4134
g1522 nand U104 P1_U3086 ; P1_U4135
g1523 nand P1_SUB_88_U20 P1_U3029 ; P1_U4136
g1524 nand P1_U4047 P1_IR_REG_29__SCAN_IN ; P1_U4137
g1525 nand U102 P1_U3086 ; P1_U4138
g1526 nand P1_SUB_88_U165 P1_U3029 ; P1_U4139
g1527 nand P1_U4047 P1_IR_REG_30__SCAN_IN ; P1_U4140
g1528 nand U101 P1_U3086 ; P1_U4141
g1529 nand P1_SUB_88_U41 P1_U3029 ; P1_U4142
g1530 nand P1_U4047 P1_IR_REG_31__SCAN_IN ; P1_U4143
g1531 not P1_U3360 ; P1_U4144
g1532 not P1_U3425 ; P1_U4145
g1533 nand P1_U3358 P1_U5775 ; P1_U4146
g1534 nand P1_U3358 P1_U5778 ; P1_U4147
g1535 nand P1_U4144 P1_D_REG_10__SCAN_IN ; P1_U4148
g1536 nand P1_U4144 P1_D_REG_11__SCAN_IN ; P1_U4149
g1537 nand P1_U4144 P1_D_REG_12__SCAN_IN ; P1_U4150
g1538 nand P1_U4144 P1_D_REG_13__SCAN_IN ; P1_U4151
g1539 nand P1_U4144 P1_D_REG_14__SCAN_IN ; P1_U4152
g1540 nand P1_U4144 P1_D_REG_15__SCAN_IN ; P1_U4153
g1541 nand P1_U4144 P1_D_REG_16__SCAN_IN ; P1_U4154
g1542 nand P1_U4144 P1_D_REG_17__SCAN_IN ; P1_U4155
g1543 nand P1_U4144 P1_D_REG_18__SCAN_IN ; P1_U4156
g1544 nand P1_U4144 P1_D_REG_19__SCAN_IN ; P1_U4157
g1545 nand P1_U4144 P1_D_REG_20__SCAN_IN ; P1_U4158
g1546 nand P1_U4144 P1_D_REG_21__SCAN_IN ; P1_U4159
g1547 nand P1_U4144 P1_D_REG_22__SCAN_IN ; P1_U4160
g1548 nand P1_U4144 P1_D_REG_23__SCAN_IN ; P1_U4161
g1549 nand P1_U4144 P1_D_REG_24__SCAN_IN ; P1_U4162
g1550 nand P1_U4144 P1_D_REG_25__SCAN_IN ; P1_U4163
g1551 nand P1_U4144 P1_D_REG_26__SCAN_IN ; P1_U4164
g1552 nand P1_U4144 P1_D_REG_27__SCAN_IN ; P1_U4165
g1553 nand P1_U4144 P1_D_REG_28__SCAN_IN ; P1_U4166
g1554 nand P1_U4144 P1_D_REG_29__SCAN_IN ; P1_U4167
g1555 nand P1_U4144 P1_D_REG_2__SCAN_IN ; P1_U4168
g1556 nand P1_U4144 P1_D_REG_30__SCAN_IN ; P1_U4169
g1557 nand P1_U4144 P1_D_REG_31__SCAN_IN ; P1_U4170
g1558 nand P1_U4144 P1_D_REG_3__SCAN_IN ; P1_U4171
g1559 nand P1_U4144 P1_D_REG_4__SCAN_IN ; P1_U4172
g1560 nand P1_U4144 P1_D_REG_5__SCAN_IN ; P1_U4173
g1561 nand P1_U4144 P1_D_REG_6__SCAN_IN ; P1_U4174
g1562 nand P1_U4144 P1_D_REG_7__SCAN_IN ; P1_U4175
g1563 nand P1_U4144 P1_D_REG_8__SCAN_IN ; P1_U4176
g1564 nand P1_U4144 P1_D_REG_9__SCAN_IN ; P1_U4177
g1565 nand P1_U5802 P1_U5799 ; P1_U4178
g1566 nand P1_U5822 P1_U5821 P1_U3369 ; P1_U4179
g1567 nand P1_U3018 P1_REG2_REG_1__SCAN_IN ; P1_U4180
g1568 nand P1_U3019 P1_REG1_REG_1__SCAN_IN ; P1_U4181
g1569 nand P1_U3020 P1_REG0_REG_1__SCAN_IN ; P1_U4182
g1570 nand P1_U3017 P1_REG3_REG_1__SCAN_IN ; P1_U4183
g1571 not P1_U3078 ; P1_U4184
g1572 nand P1_U3419 P1_U4010 ; P1_U4185
g1573 nand P1_U4007 P1_R1150_U21 ; P1_U4186
g1574 nand P1_U4000 P1_R1117_U21 ; P1_U4187
g1575 nand P1_U3994 P1_R1138_U96 ; P1_U4188
g1576 nand P1_U4005 P1_R1192_U21 ; P1_U4189
g1577 nand P1_U4004 P1_R1207_U21 ; P1_U4190
g1578 nand P1_U4011 P1_R1171_U96 ; P1_U4191
g1579 nand P1_U3992 P1_R1240_U96 ; P1_U4192
g1580 not P1_U3376 ; P1_U4193
g1581 nand P1_U3025 P1_U3078 ; P1_U4194
g1582 nand P1_R1222_U96 P1_U3024 ; P1_U4195
g1583 nand P1_U3456 P1_U4036 ; P1_U4196
g1584 nand P1_U3456 P1_U4185 ; P1_U4197
g1585 nand P1_U4197 P1_U4194 P1_U3595 P1_U4193 ; P1_U4198
g1586 nand P1_U3018 P1_REG2_REG_2__SCAN_IN ; P1_U4199
g1587 nand P1_U3019 P1_REG1_REG_2__SCAN_IN ; P1_U4200
g1588 nand P1_U3020 P1_REG0_REG_2__SCAN_IN ; P1_U4201
g1589 nand P1_U3017 P1_REG3_REG_2__SCAN_IN ; P1_U4202
g1590 not P1_U3068 ; P1_U4203
g1591 nand P1_U3020 P1_REG0_REG_0__SCAN_IN ; P1_U4204
g1592 nand P1_U3019 P1_REG1_REG_0__SCAN_IN ; P1_U4205
g1593 nand P1_U3018 P1_REG2_REG_0__SCAN_IN ; P1_U4206
g1594 nand P1_U3017 P1_REG3_REG_0__SCAN_IN ; P1_U4207
g1595 not P1_U3077 ; P1_U4208
g1596 nand P1_U3034 P1_U3077 ; P1_U4209
g1597 nand P1_R1150_U98 P1_U4007 ; P1_U4210
g1598 nand P1_R1117_U98 P1_U4000 ; P1_U4211
g1599 nand P1_R1138_U95 P1_U3994 ; P1_U4212
g1600 nand P1_R1192_U98 P1_U4005 ; P1_U4213
g1601 nand P1_R1207_U98 P1_U4004 ; P1_U4214
g1602 nand P1_R1171_U95 P1_U4011 ; P1_U4215
g1603 nand P1_R1240_U95 P1_U3992 ; P1_U4216
g1604 not P1_U3378 ; P1_U4217
g1605 nand P1_U3025 P1_U3068 ; P1_U4218
g1606 nand P1_R1222_U95 P1_U3024 ; P1_U4219
g1607 nand P1_R1282_U56 P1_U4036 ; P1_U4220
g1608 nand P1_U3461 P1_U4185 ; P1_U4221
g1609 nand P1_U3611 P1_U4217 ; P1_U4222
g1610 nand P1_U3018 P1_REG2_REG_3__SCAN_IN ; P1_U4223
g1611 nand P1_U3019 P1_REG1_REG_3__SCAN_IN ; P1_U4224
g1612 nand P1_U3020 P1_REG0_REG_3__SCAN_IN ; P1_U4225
g1613 nand P1_ADD_99_U4 P1_U3017 ; P1_U4226
g1614 not P1_U3064 ; P1_U4227
g1615 nand P1_U3034 P1_U3078 ; P1_U4228
g1616 nand P1_R1150_U108 P1_U4007 ; P1_U4229
g1617 nand P1_R1117_U108 P1_U4000 ; P1_U4230
g1618 nand P1_R1138_U17 P1_U3994 ; P1_U4231
g1619 nand P1_R1192_U108 P1_U4005 ; P1_U4232
g1620 nand P1_R1207_U108 P1_U4004 ; P1_U4233
g1621 nand P1_R1171_U17 P1_U4011 ; P1_U4234
g1622 nand P1_R1240_U17 P1_U3992 ; P1_U4235
g1623 not P1_U3379 ; P1_U4236
g1624 nand P1_U3025 P1_U3064 ; P1_U4237
g1625 nand P1_R1222_U17 P1_U3024 ; P1_U4238
g1626 nand P1_R1282_U18 P1_U4036 ; P1_U4239
g1627 nand P1_U3464 P1_U4185 ; P1_U4240
g1628 nand P1_U3615 P1_U4236 ; P1_U4241
g1629 nand P1_U3018 P1_REG2_REG_4__SCAN_IN ; P1_U4242
g1630 nand P1_U3019 P1_REG1_REG_4__SCAN_IN ; P1_U4243
g1631 nand P1_U3020 P1_REG0_REG_4__SCAN_IN ; P1_U4244
g1632 nand P1_ADD_99_U59 P1_U3017 ; P1_U4245
g1633 not P1_U3060 ; P1_U4246
g1634 nand P1_U3034 P1_U3068 ; P1_U4247
g1635 nand P1_R1150_U18 P1_U4007 ; P1_U4248
g1636 nand P1_R1117_U18 P1_U4000 ; P1_U4249
g1637 nand P1_R1138_U101 P1_U3994 ; P1_U4250
g1638 nand P1_R1192_U18 P1_U4005 ; P1_U4251
g1639 nand P1_R1207_U18 P1_U4004 ; P1_U4252
g1640 nand P1_R1171_U101 P1_U4011 ; P1_U4253
g1641 nand P1_R1240_U101 P1_U3992 ; P1_U4254
g1642 not P1_U3380 ; P1_U4255
g1643 nand P1_U3025 P1_U3060 ; P1_U4256
g1644 nand P1_R1222_U101 P1_U3024 ; P1_U4257
g1645 nand P1_R1282_U20 P1_U4036 ; P1_U4258
g1646 nand P1_U3467 P1_U4185 ; P1_U4259
g1647 nand P1_U3619 P1_U4255 ; P1_U4260
g1648 nand P1_U3018 P1_REG2_REG_5__SCAN_IN ; P1_U4261
g1649 nand P1_U3019 P1_REG1_REG_5__SCAN_IN ; P1_U4262
g1650 nand P1_U3020 P1_REG0_REG_5__SCAN_IN ; P1_U4263
g1651 nand P1_ADD_99_U58 P1_U3017 ; P1_U4264
g1652 not P1_U3067 ; P1_U4265
g1653 nand P1_U3034 P1_U3064 ; P1_U4266
g1654 nand P1_R1150_U107 P1_U4007 ; P1_U4267
g1655 nand P1_R1117_U107 P1_U4000 ; P1_U4268
g1656 nand P1_R1138_U100 P1_U3994 ; P1_U4269
g1657 nand P1_R1192_U107 P1_U4005 ; P1_U4270
g1658 nand P1_R1207_U107 P1_U4004 ; P1_U4271
g1659 nand P1_R1171_U100 P1_U4011 ; P1_U4272
g1660 nand P1_R1240_U100 P1_U3992 ; P1_U4273
g1661 not P1_U3381 ; P1_U4274
g1662 nand P1_U3025 P1_U3067 ; P1_U4275
g1663 nand P1_R1222_U100 P1_U3024 ; P1_U4276
g1664 nand P1_R1282_U21 P1_U4036 ; P1_U4277
g1665 nand P1_U3470 P1_U4185 ; P1_U4278
g1666 nand P1_U3623 P1_U4274 ; P1_U4279
g1667 nand P1_U3018 P1_REG2_REG_6__SCAN_IN ; P1_U4280
g1668 nand P1_U3019 P1_REG1_REG_6__SCAN_IN ; P1_U4281
g1669 nand P1_U3020 P1_REG0_REG_6__SCAN_IN ; P1_U4282
g1670 nand P1_ADD_99_U57 P1_U3017 ; P1_U4283
g1671 not P1_U3071 ; P1_U4284
g1672 nand P1_U3034 P1_U3060 ; P1_U4285
g1673 nand P1_R1150_U106 P1_U4007 ; P1_U4286
g1674 nand P1_R1117_U106 P1_U4000 ; P1_U4287
g1675 nand P1_R1138_U18 P1_U3994 ; P1_U4288
g1676 nand P1_R1192_U106 P1_U4005 ; P1_U4289
g1677 nand P1_R1207_U106 P1_U4004 ; P1_U4290
g1678 nand P1_R1171_U18 P1_U4011 ; P1_U4291
g1679 nand P1_R1240_U18 P1_U3992 ; P1_U4292
g1680 not P1_U3382 ; P1_U4293
g1681 nand P1_U3025 P1_U3071 ; P1_U4294
g1682 nand P1_R1222_U18 P1_U3024 ; P1_U4295
g1683 nand P1_R1282_U65 P1_U4036 ; P1_U4296
g1684 nand P1_U3473 P1_U4185 ; P1_U4297
g1685 nand P1_U3627 P1_U4293 ; P1_U4298
g1686 nand P1_U3018 P1_REG2_REG_7__SCAN_IN ; P1_U4299
g1687 nand P1_U3019 P1_REG1_REG_7__SCAN_IN ; P1_U4300
g1688 nand P1_U3020 P1_REG0_REG_7__SCAN_IN ; P1_U4301
g1689 nand P1_ADD_99_U56 P1_U3017 ; P1_U4302
g1690 not P1_U3070 ; P1_U4303
g1691 nand P1_U3034 P1_U3067 ; P1_U4304
g1692 nand P1_R1150_U19 P1_U4007 ; P1_U4305
g1693 nand P1_R1117_U19 P1_U4000 ; P1_U4306
g1694 nand P1_R1138_U99 P1_U3994 ; P1_U4307
g1695 nand P1_R1192_U19 P1_U4005 ; P1_U4308
g1696 nand P1_R1207_U19 P1_U4004 ; P1_U4309
g1697 nand P1_R1171_U99 P1_U4011 ; P1_U4310
g1698 nand P1_R1240_U99 P1_U3992 ; P1_U4311
g1699 not P1_U3383 ; P1_U4312
g1700 nand P1_U3025 P1_U3070 ; P1_U4313
g1701 nand P1_R1222_U99 P1_U3024 ; P1_U4314
g1702 nand P1_R1282_U22 P1_U4036 ; P1_U4315
g1703 nand P1_U3476 P1_U4185 ; P1_U4316
g1704 nand P1_U3631 P1_U4312 ; P1_U4317
g1705 nand P1_U3018 P1_REG2_REG_8__SCAN_IN ; P1_U4318
g1706 nand P1_U3019 P1_REG1_REG_8__SCAN_IN ; P1_U4319
g1707 nand P1_U3020 P1_REG0_REG_8__SCAN_IN ; P1_U4320
g1708 nand P1_ADD_99_U55 P1_U3017 ; P1_U4321
g1709 not P1_U3084 ; P1_U4322
g1710 nand P1_U3034 P1_U3071 ; P1_U4323
g1711 nand P1_R1150_U105 P1_U4007 ; P1_U4324
g1712 nand P1_R1117_U105 P1_U4000 ; P1_U4325
g1713 nand P1_R1138_U19 P1_U3994 ; P1_U4326
g1714 nand P1_R1192_U105 P1_U4005 ; P1_U4327
g1715 nand P1_R1207_U105 P1_U4004 ; P1_U4328
g1716 nand P1_R1171_U19 P1_U4011 ; P1_U4329
g1717 nand P1_R1240_U19 P1_U3992 ; P1_U4330
g1718 not P1_U3384 ; P1_U4331
g1719 nand P1_U3025 P1_U3084 ; P1_U4332
g1720 nand P1_R1222_U19 P1_U3024 ; P1_U4333
g1721 nand P1_R1282_U23 P1_U4036 ; P1_U4334
g1722 nand P1_U3479 P1_U4185 ; P1_U4335
g1723 nand P1_U3635 P1_U4331 ; P1_U4336
g1724 nand P1_U3018 P1_REG2_REG_9__SCAN_IN ; P1_U4337
g1725 nand P1_U3019 P1_REG1_REG_9__SCAN_IN ; P1_U4338
g1726 nand P1_U3020 P1_REG0_REG_9__SCAN_IN ; P1_U4339
g1727 nand P1_ADD_99_U54 P1_U3017 ; P1_U4340
g1728 not P1_U3083 ; P1_U4341
g1729 nand P1_U3034 P1_U3070 ; P1_U4342
g1730 nand P1_R1150_U20 P1_U4007 ; P1_U4343
g1731 nand P1_R1117_U20 P1_U4000 ; P1_U4344
g1732 nand P1_R1138_U98 P1_U3994 ; P1_U4345
g1733 nand P1_R1192_U20 P1_U4005 ; P1_U4346
g1734 nand P1_R1207_U20 P1_U4004 ; P1_U4347
g1735 nand P1_R1171_U98 P1_U4011 ; P1_U4348
g1736 nand P1_R1240_U98 P1_U3992 ; P1_U4349
g1737 not P1_U3385 ; P1_U4350
g1738 nand P1_U3025 P1_U3083 ; P1_U4351
g1739 nand P1_R1222_U98 P1_U3024 ; P1_U4352
g1740 nand P1_R1282_U24 P1_U4036 ; P1_U4353
g1741 nand P1_U3482 P1_U4185 ; P1_U4354
g1742 nand P1_U3639 P1_U4350 ; P1_U4355
g1743 nand P1_U3018 P1_REG2_REG_10__SCAN_IN ; P1_U4356
g1744 nand P1_U3019 P1_REG1_REG_10__SCAN_IN ; P1_U4357
g1745 nand P1_U3020 P1_REG0_REG_10__SCAN_IN ; P1_U4358
g1746 nand P1_ADD_99_U78 P1_U3017 ; P1_U4359
g1747 not P1_U3062 ; P1_U4360
g1748 nand P1_U3034 P1_U3084 ; P1_U4361
g1749 nand P1_R1150_U104 P1_U4007 ; P1_U4362
g1750 nand P1_R1117_U104 P1_U4000 ; P1_U4363
g1751 nand P1_R1138_U97 P1_U3994 ; P1_U4364
g1752 nand P1_R1192_U104 P1_U4005 ; P1_U4365
g1753 nand P1_R1207_U104 P1_U4004 ; P1_U4366
g1754 nand P1_R1171_U97 P1_U4011 ; P1_U4367
g1755 nand P1_R1240_U97 P1_U3992 ; P1_U4368
g1756 not P1_U3386 ; P1_U4369
g1757 nand P1_U3025 P1_U3062 ; P1_U4370
g1758 nand P1_R1222_U97 P1_U3024 ; P1_U4371
g1759 nand P1_R1282_U63 P1_U4036 ; P1_U4372
g1760 nand P1_U3485 P1_U4185 ; P1_U4373
g1761 nand P1_U3643 P1_U4369 ; P1_U4374
g1762 nand P1_U3018 P1_REG2_REG_11__SCAN_IN ; P1_U4375
g1763 nand P1_U3019 P1_REG1_REG_11__SCAN_IN ; P1_U4376
g1764 nand P1_U3020 P1_REG0_REG_11__SCAN_IN ; P1_U4377
g1765 nand P1_ADD_99_U77 P1_U3017 ; P1_U4378
g1766 not P1_U3063 ; P1_U4379
g1767 nand P1_U3034 P1_U3083 ; P1_U4380
g1768 nand P1_R1150_U114 P1_U4007 ; P1_U4381
g1769 nand P1_R1117_U114 P1_U4000 ; P1_U4382
g1770 nand P1_R1138_U11 P1_U3994 ; P1_U4383
g1771 nand P1_R1192_U114 P1_U4005 ; P1_U4384
g1772 nand P1_R1207_U114 P1_U4004 ; P1_U4385
g1773 nand P1_R1171_U11 P1_U4011 ; P1_U4386
g1774 nand P1_R1240_U11 P1_U3992 ; P1_U4387
g1775 not P1_U3387 ; P1_U4388
g1776 nand P1_U3025 P1_U3063 ; P1_U4389
g1777 nand P1_R1222_U11 P1_U3024 ; P1_U4390
g1778 nand P1_R1282_U6 P1_U4036 ; P1_U4391
g1779 nand P1_U3488 P1_U4185 ; P1_U4392
g1780 nand P1_U3647 P1_U4388 ; P1_U4393
g1781 nand P1_U3018 P1_REG2_REG_12__SCAN_IN ; P1_U4394
g1782 nand P1_U3019 P1_REG1_REG_12__SCAN_IN ; P1_U4395
g1783 nand P1_U3020 P1_REG0_REG_12__SCAN_IN ; P1_U4396
g1784 nand P1_ADD_99_U76 P1_U3017 ; P1_U4397
g1785 not P1_U3072 ; P1_U4398
g1786 nand P1_U3034 P1_U3062 ; P1_U4399
g1787 nand P1_R1150_U13 P1_U4007 ; P1_U4400
g1788 nand P1_R1117_U13 P1_U4000 ; P1_U4401
g1789 nand P1_R1138_U115 P1_U3994 ; P1_U4402
g1790 nand P1_R1192_U13 P1_U4005 ; P1_U4403
g1791 nand P1_R1207_U13 P1_U4004 ; P1_U4404
g1792 nand P1_R1171_U115 P1_U4011 ; P1_U4405
g1793 nand P1_R1240_U115 P1_U3992 ; P1_U4406
g1794 not P1_U3388 ; P1_U4407
g1795 nand P1_U3025 P1_U3072 ; P1_U4408
g1796 nand P1_R1222_U115 P1_U3024 ; P1_U4409
g1797 nand P1_R1282_U7 P1_U4036 ; P1_U4410
g1798 nand P1_U3491 P1_U4185 ; P1_U4411
g1799 nand P1_U3651 P1_U4407 ; P1_U4412
g1800 nand P1_U3018 P1_REG2_REG_13__SCAN_IN ; P1_U4413
g1801 nand P1_U3019 P1_REG1_REG_13__SCAN_IN ; P1_U4414
g1802 nand P1_U3020 P1_REG0_REG_13__SCAN_IN ; P1_U4415
g1803 nand P1_ADD_99_U75 P1_U3017 ; P1_U4416
g1804 not P1_U3080 ; P1_U4417
g1805 nand P1_U3034 P1_U3063 ; P1_U4418
g1806 nand P1_R1150_U103 P1_U4007 ; P1_U4419
g1807 nand P1_R1117_U103 P1_U4000 ; P1_U4420
g1808 nand P1_R1138_U114 P1_U3994 ; P1_U4421
g1809 nand P1_R1192_U103 P1_U4005 ; P1_U4422
g1810 nand P1_R1207_U103 P1_U4004 ; P1_U4423
g1811 nand P1_R1171_U114 P1_U4011 ; P1_U4424
g1812 nand P1_R1240_U114 P1_U3992 ; P1_U4425
g1813 not P1_U3389 ; P1_U4426
g1814 nand P1_U3025 P1_U3080 ; P1_U4427
g1815 nand P1_R1222_U114 P1_U3024 ; P1_U4428
g1816 nand P1_R1282_U8 P1_U4036 ; P1_U4429
g1817 nand P1_U3494 P1_U4185 ; P1_U4430
g1818 nand P1_U3655 P1_U4426 ; P1_U4431
g1819 nand P1_U3018 P1_REG2_REG_14__SCAN_IN ; P1_U4432
g1820 nand P1_U3019 P1_REG1_REG_14__SCAN_IN ; P1_U4433
g1821 nand P1_U3020 P1_REG0_REG_14__SCAN_IN ; P1_U4434
g1822 nand P1_ADD_99_U74 P1_U3017 ; P1_U4435
g1823 not P1_U3079 ; P1_U4436
g1824 nand P1_U3034 P1_U3072 ; P1_U4437
g1825 nand P1_R1150_U102 P1_U4007 ; P1_U4438
g1826 nand P1_R1117_U102 P1_U4000 ; P1_U4439
g1827 nand P1_R1138_U12 P1_U3994 ; P1_U4440
g1828 nand P1_R1192_U102 P1_U4005 ; P1_U4441
g1829 nand P1_R1207_U102 P1_U4004 ; P1_U4442
g1830 nand P1_R1171_U12 P1_U4011 ; P1_U4443
g1831 nand P1_R1240_U12 P1_U3992 ; P1_U4444
g1832 not P1_U3390 ; P1_U4445
g1833 nand P1_U3025 P1_U3079 ; P1_U4446
g1834 nand P1_R1222_U12 P1_U3024 ; P1_U4447
g1835 nand P1_R1282_U86 P1_U4036 ; P1_U4448
g1836 nand P1_U3497 P1_U4185 ; P1_U4449
g1837 nand P1_U3659 P1_U4445 ; P1_U4450
g1838 nand P1_U3018 P1_REG2_REG_15__SCAN_IN ; P1_U4451
g1839 nand P1_U3019 P1_REG1_REG_15__SCAN_IN ; P1_U4452
g1840 nand P1_U3020 P1_REG0_REG_15__SCAN_IN ; P1_U4453
g1841 nand P1_ADD_99_U73 P1_U3017 ; P1_U4454
g1842 not P1_U3074 ; P1_U4455
g1843 nand P1_U3034 P1_U3080 ; P1_U4456
g1844 nand P1_R1150_U113 P1_U4007 ; P1_U4457
g1845 nand P1_R1117_U113 P1_U4000 ; P1_U4458
g1846 nand P1_R1138_U113 P1_U3994 ; P1_U4459
g1847 nand P1_R1192_U113 P1_U4005 ; P1_U4460
g1848 nand P1_R1207_U113 P1_U4004 ; P1_U4461
g1849 nand P1_R1171_U113 P1_U4011 ; P1_U4462
g1850 nand P1_R1240_U113 P1_U3992 ; P1_U4463
g1851 not P1_U3391 ; P1_U4464
g1852 nand P1_U3025 P1_U3074 ; P1_U4465
g1853 nand P1_R1222_U113 P1_U3024 ; P1_U4466
g1854 nand P1_R1282_U9 P1_U4036 ; P1_U4467
g1855 nand P1_U3500 P1_U4185 ; P1_U4468
g1856 nand P1_U3663 P1_U4464 ; P1_U4469
g1857 nand P1_U3018 P1_REG2_REG_16__SCAN_IN ; P1_U4470
g1858 nand P1_U3019 P1_REG1_REG_16__SCAN_IN ; P1_U4471
g1859 nand P1_U3020 P1_REG0_REG_16__SCAN_IN ; P1_U4472
g1860 nand P1_ADD_99_U72 P1_U3017 ; P1_U4473
g1861 not P1_U3073 ; P1_U4474
g1862 nand P1_U3034 P1_U3079 ; P1_U4475
g1863 nand P1_R1150_U112 P1_U4007 ; P1_U4476
g1864 nand P1_R1117_U112 P1_U4000 ; P1_U4477
g1865 nand P1_R1138_U112 P1_U3994 ; P1_U4478
g1866 nand P1_R1192_U112 P1_U4005 ; P1_U4479
g1867 nand P1_R1207_U112 P1_U4004 ; P1_U4480
g1868 nand P1_R1171_U112 P1_U4011 ; P1_U4481
g1869 nand P1_R1240_U112 P1_U3992 ; P1_U4482
g1870 not P1_U3392 ; P1_U4483
g1871 nand P1_U3025 P1_U3073 ; P1_U4484
g1872 nand P1_R1222_U112 P1_U3024 ; P1_U4485
g1873 nand P1_R1282_U10 P1_U4036 ; P1_U4486
g1874 nand P1_U3503 P1_U4185 ; P1_U4487
g1875 nand P1_U3667 P1_U4483 ; P1_U4488
g1876 nand P1_U3018 P1_REG2_REG_17__SCAN_IN ; P1_U4489
g1877 nand P1_U3019 P1_REG1_REG_17__SCAN_IN ; P1_U4490
g1878 nand P1_U3020 P1_REG0_REG_17__SCAN_IN ; P1_U4491
g1879 nand P1_ADD_99_U71 P1_U3017 ; P1_U4492
g1880 not P1_U3069 ; P1_U4493
g1881 nand P1_U3034 P1_U3074 ; P1_U4494
g1882 nand P1_R1150_U14 P1_U4007 ; P1_U4495
g1883 nand P1_R1117_U14 P1_U4000 ; P1_U4496
g1884 nand P1_R1138_U111 P1_U3994 ; P1_U4497
g1885 nand P1_R1192_U14 P1_U4005 ; P1_U4498
g1886 nand P1_R1207_U14 P1_U4004 ; P1_U4499
g1887 nand P1_R1171_U111 P1_U4011 ; P1_U4500
g1888 nand P1_R1240_U111 P1_U3992 ; P1_U4501
g1889 not P1_U3393 ; P1_U4502
g1890 nand P1_U3025 P1_U3069 ; P1_U4503
g1891 nand P1_R1222_U111 P1_U3024 ; P1_U4504
g1892 nand P1_R1282_U11 P1_U4036 ; P1_U4505
g1893 nand P1_U3506 P1_U4185 ; P1_U4506
g1894 nand P1_U3671 P1_U4502 ; P1_U4507
g1895 nand P1_U3018 P1_REG2_REG_18__SCAN_IN ; P1_U4508
g1896 nand P1_U3019 P1_REG1_REG_18__SCAN_IN ; P1_U4509
g1897 nand P1_U3020 P1_REG0_REG_18__SCAN_IN ; P1_U4510
g1898 nand P1_ADD_99_U70 P1_U3017 ; P1_U4511
g1899 not P1_U3082 ; P1_U4512
g1900 nand P1_U3034 P1_U3073 ; P1_U4513
g1901 nand P1_R1150_U101 P1_U4007 ; P1_U4514
g1902 nand P1_R1117_U101 P1_U4000 ; P1_U4515
g1903 nand P1_R1138_U13 P1_U3994 ; P1_U4516
g1904 nand P1_R1192_U101 P1_U4005 ; P1_U4517
g1905 nand P1_R1207_U101 P1_U4004 ; P1_U4518
g1906 nand P1_R1171_U13 P1_U4011 ; P1_U4519
g1907 nand P1_R1240_U13 P1_U3992 ; P1_U4520
g1908 not P1_U3394 ; P1_U4521
g1909 nand P1_U3025 P1_U3082 ; P1_U4522
g1910 nand P1_R1222_U13 P1_U3024 ; P1_U4523
g1911 nand P1_R1282_U84 P1_U4036 ; P1_U4524
g1912 nand P1_U3509 P1_U4185 ; P1_U4525
g1913 nand P1_U3675 P1_U4521 ; P1_U4526
g1914 nand P1_U3018 P1_REG2_REG_19__SCAN_IN ; P1_U4527
g1915 nand P1_U3019 P1_REG1_REG_19__SCAN_IN ; P1_U4528
g1916 nand P1_U3020 P1_REG0_REG_19__SCAN_IN ; P1_U4529
g1917 nand P1_ADD_99_U69 P1_U3017 ; P1_U4530
g1918 not P1_U3081 ; P1_U4531
g1919 nand P1_U3034 P1_U3069 ; P1_U4532
g1920 nand P1_R1150_U100 P1_U4007 ; P1_U4533
g1921 nand P1_R1117_U100 P1_U4000 ; P1_U4534
g1922 nand P1_R1138_U110 P1_U3994 ; P1_U4535
g1923 nand P1_R1192_U100 P1_U4005 ; P1_U4536
g1924 nand P1_R1207_U100 P1_U4004 ; P1_U4537
g1925 nand P1_R1171_U110 P1_U4011 ; P1_U4538
g1926 nand P1_R1240_U110 P1_U3992 ; P1_U4539
g1927 not P1_U3395 ; P1_U4540
g1928 nand P1_U3025 P1_U3081 ; P1_U4541
g1929 nand P1_R1222_U110 P1_U3024 ; P1_U4542
g1930 nand P1_R1282_U12 P1_U4036 ; P1_U4543
g1931 nand P1_U3512 P1_U4185 ; P1_U4544
g1932 nand P1_U3679 P1_U4540 ; P1_U4545
g1933 nand P1_U3018 P1_REG2_REG_20__SCAN_IN ; P1_U4546
g1934 nand P1_U3019 P1_REG1_REG_20__SCAN_IN ; P1_U4547
g1935 nand P1_U3020 P1_REG0_REG_20__SCAN_IN ; P1_U4548
g1936 nand P1_ADD_99_U68 P1_U3017 ; P1_U4549
g1937 not P1_U3076 ; P1_U4550
g1938 nand P1_U3034 P1_U3082 ; P1_U4551
g1939 nand P1_R1150_U99 P1_U4007 ; P1_U4552
g1940 nand P1_R1117_U99 P1_U4000 ; P1_U4553
g1941 nand P1_R1138_U109 P1_U3994 ; P1_U4554
g1942 nand P1_R1192_U99 P1_U4005 ; P1_U4555
g1943 nand P1_R1207_U99 P1_U4004 ; P1_U4556
g1944 nand P1_R1171_U109 P1_U4011 ; P1_U4557
g1945 nand P1_R1240_U109 P1_U3992 ; P1_U4558
g1946 not P1_U3396 ; P1_U4559
g1947 nand P1_U3025 P1_U3076 ; P1_U4560
g1948 nand P1_R1222_U109 P1_U3024 ; P1_U4561
g1949 nand P1_R1282_U82 P1_U4036 ; P1_U4562
g1950 nand P1_U3514 P1_U4185 ; P1_U4563
g1951 nand P1_U3683 P1_U4559 ; P1_U4564
g1952 nand P1_U3018 P1_REG2_REG_21__SCAN_IN ; P1_U4565
g1953 nand P1_U3019 P1_REG1_REG_21__SCAN_IN ; P1_U4566
g1954 nand P1_U3020 P1_REG0_REG_21__SCAN_IN ; P1_U4567
g1955 nand P1_ADD_99_U67 P1_U3017 ; P1_U4568
g1956 not P1_U3075 ; P1_U4569
g1957 nand P1_U3034 P1_U3081 ; P1_U4570
g1958 nand P1_R1150_U97 P1_U4007 ; P1_U4571
g1959 nand P1_R1117_U97 P1_U4000 ; P1_U4572
g1960 nand P1_R1138_U14 P1_U3994 ; P1_U4573
g1961 nand P1_R1192_U97 P1_U4005 ; P1_U4574
g1962 nand P1_R1207_U97 P1_U4004 ; P1_U4575
g1963 nand P1_R1171_U14 P1_U4011 ; P1_U4576
g1964 nand P1_R1240_U14 P1_U3992 ; P1_U4577
g1965 not P1_U3398 ; P1_U4578
g1966 nand P1_U3025 P1_U3075 ; P1_U4579
g1967 nand P1_R1222_U14 P1_U3024 ; P1_U4580
g1968 nand P1_R1282_U13 P1_U4036 ; P1_U4581
g1969 nand P1_U4025 P1_U4185 ; P1_U4582
g1970 nand P1_U3687 P1_U4578 ; P1_U4583
g1971 nand P1_U3018 P1_REG2_REG_22__SCAN_IN ; P1_U4584
g1972 nand P1_U3019 P1_REG1_REG_22__SCAN_IN ; P1_U4585
g1973 nand P1_U3020 P1_REG0_REG_22__SCAN_IN ; P1_U4586
g1974 nand P1_ADD_99_U66 P1_U3017 ; P1_U4587
g1975 not P1_U3061 ; P1_U4588
g1976 nand P1_U3034 P1_U3076 ; P1_U4589
g1977 nand P1_R1150_U111 P1_U4007 ; P1_U4590
g1978 nand P1_R1117_U111 P1_U4000 ; P1_U4591
g1979 nand P1_R1138_U15 P1_U3994 ; P1_U4592
g1980 nand P1_R1192_U111 P1_U4005 ; P1_U4593
g1981 nand P1_R1207_U111 P1_U4004 ; P1_U4594
g1982 nand P1_R1171_U15 P1_U4011 ; P1_U4595
g1983 nand P1_R1240_U15 P1_U3992 ; P1_U4596
g1984 not P1_U3400 ; P1_U4597
g1985 nand P1_U3025 P1_U3061 ; P1_U4598
g1986 nand P1_R1222_U15 P1_U3024 ; P1_U4599
g1987 nand P1_R1282_U78 P1_U4036 ; P1_U4600
g1988 nand P1_U4024 P1_U4185 ; P1_U4601
g1989 nand P1_U3691 P1_U4597 ; P1_U4602
g1990 nand P1_U3018 P1_REG2_REG_23__SCAN_IN ; P1_U4603
g1991 nand P1_U3019 P1_REG1_REG_23__SCAN_IN ; P1_U4604
g1992 nand P1_U3020 P1_REG0_REG_23__SCAN_IN ; P1_U4605
g1993 nand P1_ADD_99_U65 P1_U3017 ; P1_U4606
g1994 not P1_U3066 ; P1_U4607
g1995 nand P1_U3034 P1_U3075 ; P1_U4608
g1996 nand P1_R1150_U110 P1_U4007 ; P1_U4609
g1997 nand P1_R1117_U110 P1_U4000 ; P1_U4610
g1998 nand P1_R1138_U108 P1_U3994 ; P1_U4611
g1999 nand P1_R1192_U110 P1_U4005 ; P1_U4612
g2000 nand P1_R1207_U110 P1_U4004 ; P1_U4613
g2001 nand P1_R1171_U108 P1_U4011 ; P1_U4614
g2002 nand P1_R1240_U108 P1_U3992 ; P1_U4615
g2003 not P1_U3402 ; P1_U4616
g2004 nand P1_U3025 P1_U3066 ; P1_U4617
g2005 nand P1_R1222_U108 P1_U3024 ; P1_U4618
g2006 nand P1_R1282_U14 P1_U4036 ; P1_U4619
g2007 nand P1_U4023 P1_U4185 ; P1_U4620
g2008 nand P1_U3695 P1_U4616 ; P1_U4621
g2009 nand P1_U3018 P1_REG2_REG_24__SCAN_IN ; P1_U4622
g2010 nand P1_U3019 P1_REG1_REG_24__SCAN_IN ; P1_U4623
g2011 nand P1_U3020 P1_REG0_REG_24__SCAN_IN ; P1_U4624
g2012 nand P1_ADD_99_U64 P1_U3017 ; P1_U4625
g2013 not P1_U3065 ; P1_U4626
g2014 nand P1_U3034 P1_U3061 ; P1_U4627
g2015 nand P1_R1150_U15 P1_U4007 ; P1_U4628
g2016 nand P1_R1117_U15 P1_U4000 ; P1_U4629
g2017 nand P1_R1138_U107 P1_U3994 ; P1_U4630
g2018 nand P1_R1192_U15 P1_U4005 ; P1_U4631
g2019 nand P1_R1207_U15 P1_U4004 ; P1_U4632
g2020 nand P1_R1171_U107 P1_U4011 ; P1_U4633
g2021 nand P1_R1240_U107 P1_U3992 ; P1_U4634
g2022 not P1_U3404 ; P1_U4635
g2023 nand P1_U3025 P1_U3065 ; P1_U4636
g2024 nand P1_R1222_U107 P1_U3024 ; P1_U4637
g2025 nand P1_R1282_U76 P1_U4036 ; P1_U4638
g2026 nand P1_U4022 P1_U4185 ; P1_U4639
g2027 nand P1_U3699 P1_U4635 ; P1_U4640
g2028 nand P1_U3018 P1_REG2_REG_25__SCAN_IN ; P1_U4641
g2029 nand P1_U3019 P1_REG1_REG_25__SCAN_IN ; P1_U4642
g2030 nand P1_U3020 P1_REG0_REG_25__SCAN_IN ; P1_U4643
g2031 nand P1_ADD_99_U63 P1_U3017 ; P1_U4644
g2032 not P1_U3058 ; P1_U4645
g2033 nand P1_U3034 P1_U3066 ; P1_U4646
g2034 nand P1_R1150_U96 P1_U4007 ; P1_U4647
g2035 nand P1_R1117_U96 P1_U4000 ; P1_U4648
g2036 nand P1_R1138_U106 P1_U3994 ; P1_U4649
g2037 nand P1_R1192_U96 P1_U4005 ; P1_U4650
g2038 nand P1_R1207_U96 P1_U4004 ; P1_U4651
g2039 nand P1_R1171_U106 P1_U4011 ; P1_U4652
g2040 nand P1_R1240_U106 P1_U3992 ; P1_U4653
g2041 not P1_U3406 ; P1_U4654
g2042 nand P1_U3025 P1_U3058 ; P1_U4655
g2043 nand P1_R1222_U106 P1_U3024 ; P1_U4656
g2044 nand P1_R1282_U15 P1_U4036 ; P1_U4657
g2045 nand P1_U4021 P1_U4185 ; P1_U4658
g2046 nand P1_U3703 P1_U4654 ; P1_U4659
g2047 nand P1_U3018 P1_REG2_REG_26__SCAN_IN ; P1_U4660
g2048 nand P1_U3019 P1_REG1_REG_26__SCAN_IN ; P1_U4661
g2049 nand P1_U3020 P1_REG0_REG_26__SCAN_IN ; P1_U4662
g2050 nand P1_ADD_99_U62 P1_U3017 ; P1_U4663
g2051 not P1_U3057 ; P1_U4664
g2052 nand P1_U3034 P1_U3065 ; P1_U4665
g2053 nand P1_R1150_U95 P1_U4007 ; P1_U4666
g2054 nand P1_R1117_U95 P1_U4000 ; P1_U4667
g2055 nand P1_R1138_U105 P1_U3994 ; P1_U4668
g2056 nand P1_R1192_U95 P1_U4005 ; P1_U4669
g2057 nand P1_R1207_U95 P1_U4004 ; P1_U4670
g2058 nand P1_R1171_U105 P1_U4011 ; P1_U4671
g2059 nand P1_R1240_U105 P1_U3992 ; P1_U4672
g2060 not P1_U3408 ; P1_U4673
g2061 nand P1_U3025 P1_U3057 ; P1_U4674
g2062 nand P1_R1222_U105 P1_U3024 ; P1_U4675
g2063 nand P1_R1282_U74 P1_U4036 ; P1_U4676
g2064 nand P1_U4020 P1_U4185 ; P1_U4677
g2065 nand P1_U3707 P1_U4673 ; P1_U4678
g2066 nand P1_U3018 P1_REG2_REG_27__SCAN_IN ; P1_U4679
g2067 nand P1_U3019 P1_REG1_REG_27__SCAN_IN ; P1_U4680
g2068 nand P1_U3020 P1_REG0_REG_27__SCAN_IN ; P1_U4681
g2069 nand P1_ADD_99_U61 P1_U3017 ; P1_U4682
g2070 not P1_U3053 ; P1_U4683
g2071 nand P1_U3034 P1_U3058 ; P1_U4684
g2072 nand P1_R1150_U109 P1_U4007 ; P1_U4685
g2073 nand P1_R1117_U109 P1_U4000 ; P1_U4686
g2074 nand P1_R1138_U16 P1_U3994 ; P1_U4687
g2075 nand P1_R1192_U109 P1_U4005 ; P1_U4688
g2076 nand P1_R1207_U109 P1_U4004 ; P1_U4689
g2077 nand P1_R1171_U16 P1_U4011 ; P1_U4690
g2078 nand P1_R1240_U16 P1_U3992 ; P1_U4691
g2079 not P1_U3410 ; P1_U4692
g2080 nand P1_U3025 P1_U3053 ; P1_U4693
g2081 nand P1_R1222_U16 P1_U3024 ; P1_U4694
g2082 nand P1_R1282_U16 P1_U4036 ; P1_U4695
g2083 nand P1_U4019 P1_U4185 ; P1_U4696
g2084 nand P1_U3711 P1_U4692 ; P1_U4697
g2085 nand P1_U3018 P1_REG2_REG_28__SCAN_IN ; P1_U4698
g2086 nand P1_U3019 P1_REG1_REG_28__SCAN_IN ; P1_U4699
g2087 nand P1_U3020 P1_REG0_REG_28__SCAN_IN ; P1_U4700
g2088 nand P1_ADD_99_U60 P1_U3017 ; P1_U4701
g2089 not P1_U3054 ; P1_U4702
g2090 nand P1_U3034 P1_U3057 ; P1_U4703
g2091 nand P1_R1150_U16 P1_U4007 ; P1_U4704
g2092 nand P1_R1117_U16 P1_U4000 ; P1_U4705
g2093 nand P1_R1138_U104 P1_U3994 ; P1_U4706
g2094 nand P1_R1192_U16 P1_U4005 ; P1_U4707
g2095 nand P1_R1207_U16 P1_U4004 ; P1_U4708
g2096 nand P1_R1171_U104 P1_U4011 ; P1_U4709
g2097 nand P1_R1240_U104 P1_U3992 ; P1_U4710
g2098 not P1_U3412 ; P1_U4711
g2099 nand P1_U3025 P1_U3054 ; P1_U4712
g2100 nand P1_R1222_U104 P1_U3024 ; P1_U4713
g2101 nand P1_R1282_U72 P1_U4036 ; P1_U4714
g2102 nand P1_U4018 P1_U4185 ; P1_U4715
g2103 nand P1_U3715 P1_U4711 ; P1_U4716
g2104 nand P1_ADD_99_U5 P1_U3017 ; P1_U4717
g2105 nand P1_U3018 P1_REG2_REG_29__SCAN_IN ; P1_U4718
g2106 nand P1_U3019 P1_REG1_REG_29__SCAN_IN ; P1_U4719
g2107 nand P1_U3020 P1_REG0_REG_29__SCAN_IN ; P1_U4720
g2108 not P1_U3055 ; P1_U4721
g2109 nand P1_U3034 P1_U3053 ; P1_U4722
g2110 nand P1_R1150_U94 P1_U4007 ; P1_U4723
g2111 nand P1_R1117_U94 P1_U4000 ; P1_U4724
g2112 nand P1_R1138_U103 P1_U3994 ; P1_U4725
g2113 nand P1_R1192_U94 P1_U4005 ; P1_U4726
g2114 nand P1_R1207_U94 P1_U4004 ; P1_U4727
g2115 nand P1_R1171_U103 P1_U4011 ; P1_U4728
g2116 nand P1_R1240_U103 P1_U3992 ; P1_U4729
g2117 not P1_U3414 ; P1_U4730
g2118 nand P1_U3025 P1_U3055 ; P1_U4731
g2119 nand P1_R1222_U103 P1_U3024 ; P1_U4732
g2120 nand P1_R1282_U17 P1_U4036 ; P1_U4733
g2121 nand P1_U4017 P1_U4185 ; P1_U4734
g2122 nand P1_U3719 P1_U4730 ; P1_U4735
g2123 nand P1_U3018 P1_REG2_REG_30__SCAN_IN ; P1_U4736
g2124 nand P1_U3019 P1_REG1_REG_30__SCAN_IN ; P1_U4737
g2125 nand P1_U3020 P1_REG0_REG_30__SCAN_IN ; P1_U4738
g2126 not P1_U3059 ; P1_U4739
g2127 nand P1_U5811 P1_U3359 ; P1_U4740
g2128 nand P1_U3954 P1_U4740 ; P1_U4741
g2129 nand P1_U3720 P1_U3059 ; P1_U4742
g2130 nand P1_U3034 P1_U3054 ; P1_U4743
g2131 nand P1_R1150_U17 P1_U4007 ; P1_U4744
g2132 nand P1_R1117_U17 P1_U4000 ; P1_U4745
g2133 nand P1_R1138_U102 P1_U3994 ; P1_U4746
g2134 nand P1_R1192_U17 P1_U4005 ; P1_U4747
g2135 nand P1_R1207_U17 P1_U4004 ; P1_U4748
g2136 nand P1_R1171_U102 P1_U4011 ; P1_U4749
g2137 nand P1_R1240_U102 P1_U3992 ; P1_U4750
g2138 not P1_U3416 ; P1_U4751
g2139 nand P1_R1222_U102 P1_U3024 ; P1_U4752
g2140 nand P1_R1282_U70 P1_U4036 ; P1_U4753
g2141 nand P1_U4028 P1_U4185 ; P1_U4754
g2142 nand P1_U3724 P1_U4751 ; P1_U4755
g2143 nand P1_U3018 P1_REG2_REG_31__SCAN_IN ; P1_U4756
g2144 nand P1_U3019 P1_REG1_REG_31__SCAN_IN ; P1_U4757
g2145 nand P1_U3020 P1_REG0_REG_31__SCAN_IN ; P1_U4758
g2146 not P1_U3056 ; P1_U4759
g2147 nand P1_R1282_U19 P1_U4036 ; P1_U4760
g2148 nand P1_U4027 P1_U4185 ; P1_U4761
g2149 nand P1_U4761 P1_U3987 P1_U4760 ; P1_U4762
g2150 nand P1_R1282_U68 P1_U4036 ; P1_U4763
g2151 nand P1_U4026 P1_U4185 ; P1_U4764
g2152 nand P1_U4764 P1_U3987 P1_U4763 ; P1_U4765
g2153 nand P1_U3727 P1_U3016 ; P1_U4766
g2154 nand P1_U3421 P1_U4766 ; P1_U4767
g2155 nand P1_U3995 P1_U5802 ; P1_U4768
g2156 not P1_U3426 ; P1_U4769
g2157 nand P1_U3036 P1_U3078 ; P1_U4770
g2158 nand P1_U3033 P1_REG3_REG_0__SCAN_IN ; P1_U4771
g2159 nand P1_U3032 P1_R1222_U96 ; P1_U4772
g2160 nand P1_U3031 P1_U3456 ; P1_U4773
g2161 nand P1_U3030 P1_U3456 ; P1_U4774
g2162 nand P1_U3036 P1_U3068 ; P1_U4775
g2163 nand P1_U3033 P1_REG3_REG_1__SCAN_IN ; P1_U4776
g2164 nand P1_U3032 P1_R1222_U95 ; P1_U4777
g2165 nand P1_U3031 P1_U3461 ; P1_U4778
g2166 nand P1_U3030 P1_R1282_U56 ; P1_U4779
g2167 nand P1_U3036 P1_U3064 ; P1_U4780
g2168 nand P1_U3033 P1_REG3_REG_2__SCAN_IN ; P1_U4781
g2169 nand P1_U3032 P1_R1222_U17 ; P1_U4782
g2170 nand P1_U3031 P1_U3464 ; P1_U4783
g2171 nand P1_U3030 P1_R1282_U18 ; P1_U4784
g2172 nand P1_U3036 P1_U3060 ; P1_U4785
g2173 nand P1_U3033 P1_ADD_99_U4 ; P1_U4786
g2174 nand P1_U3032 P1_R1222_U101 ; P1_U4787
g2175 nand P1_U3031 P1_U3467 ; P1_U4788
g2176 nand P1_U3030 P1_R1282_U20 ; P1_U4789
g2177 nand P1_U3036 P1_U3067 ; P1_U4790
g2178 nand P1_U3033 P1_ADD_99_U59 ; P1_U4791
g2179 nand P1_U3032 P1_R1222_U100 ; P1_U4792
g2180 nand P1_U3031 P1_U3470 ; P1_U4793
g2181 nand P1_U3030 P1_R1282_U21 ; P1_U4794
g2182 nand P1_U3036 P1_U3071 ; P1_U4795
g2183 nand P1_U3033 P1_ADD_99_U58 ; P1_U4796
g2184 nand P1_U3032 P1_R1222_U18 ; P1_U4797
g2185 nand P1_U3031 P1_U3473 ; P1_U4798
g2186 nand P1_U3030 P1_R1282_U65 ; P1_U4799
g2187 nand P1_U3036 P1_U3070 ; P1_U4800
g2188 nand P1_U3033 P1_ADD_99_U57 ; P1_U4801
g2189 nand P1_U3032 P1_R1222_U99 ; P1_U4802
g2190 nand P1_U3031 P1_U3476 ; P1_U4803
g2191 nand P1_U3030 P1_R1282_U22 ; P1_U4804
g2192 nand P1_U3036 P1_U3084 ; P1_U4805
g2193 nand P1_U3033 P1_ADD_99_U56 ; P1_U4806
g2194 nand P1_U3032 P1_R1222_U19 ; P1_U4807
g2195 nand P1_U3031 P1_U3479 ; P1_U4808
g2196 nand P1_U3030 P1_R1282_U23 ; P1_U4809
g2197 nand P1_U3036 P1_U3083 ; P1_U4810
g2198 nand P1_U3033 P1_ADD_99_U55 ; P1_U4811
g2199 nand P1_U3032 P1_R1222_U98 ; P1_U4812
g2200 nand P1_U3031 P1_U3482 ; P1_U4813
g2201 nand P1_U3030 P1_R1282_U24 ; P1_U4814
g2202 nand P1_U3036 P1_U3062 ; P1_U4815
g2203 nand P1_U3033 P1_ADD_99_U54 ; P1_U4816
g2204 nand P1_U3032 P1_R1222_U97 ; P1_U4817
g2205 nand P1_U3031 P1_U3485 ; P1_U4818
g2206 nand P1_U3030 P1_R1282_U63 ; P1_U4819
g2207 nand P1_U3036 P1_U3063 ; P1_U4820
g2208 nand P1_U3033 P1_ADD_99_U78 ; P1_U4821
g2209 nand P1_U3032 P1_R1222_U11 ; P1_U4822
g2210 nand P1_U3031 P1_U3488 ; P1_U4823
g2211 nand P1_U3030 P1_R1282_U6 ; P1_U4824
g2212 nand P1_U3036 P1_U3072 ; P1_U4825
g2213 nand P1_U3033 P1_ADD_99_U77 ; P1_U4826
g2214 nand P1_U3032 P1_R1222_U115 ; P1_U4827
g2215 nand P1_U3031 P1_U3491 ; P1_U4828
g2216 nand P1_U3030 P1_R1282_U7 ; P1_U4829
g2217 nand P1_U3036 P1_U3080 ; P1_U4830
g2218 nand P1_U3033 P1_ADD_99_U76 ; P1_U4831
g2219 nand P1_U3032 P1_R1222_U114 ; P1_U4832
g2220 nand P1_U3031 P1_U3494 ; P1_U4833
g2221 nand P1_U3030 P1_R1282_U8 ; P1_U4834
g2222 nand P1_U3036 P1_U3079 ; P1_U4835
g2223 nand P1_U3033 P1_ADD_99_U75 ; P1_U4836
g2224 nand P1_U3032 P1_R1222_U12 ; P1_U4837
g2225 nand P1_U3031 P1_U3497 ; P1_U4838
g2226 nand P1_U3030 P1_R1282_U86 ; P1_U4839
g2227 nand P1_U3036 P1_U3074 ; P1_U4840
g2228 nand P1_U3033 P1_ADD_99_U74 ; P1_U4841
g2229 nand P1_U3032 P1_R1222_U113 ; P1_U4842
g2230 nand P1_U3031 P1_U3500 ; P1_U4843
g2231 nand P1_U3030 P1_R1282_U9 ; P1_U4844
g2232 nand P1_U3036 P1_U3073 ; P1_U4845
g2233 nand P1_U3033 P1_ADD_99_U73 ; P1_U4846
g2234 nand P1_U3032 P1_R1222_U112 ; P1_U4847
g2235 nand P1_U3031 P1_U3503 ; P1_U4848
g2236 nand P1_U3030 P1_R1282_U10 ; P1_U4849
g2237 nand P1_U3036 P1_U3069 ; P1_U4850
g2238 nand P1_U3033 P1_ADD_99_U72 ; P1_U4851
g2239 nand P1_U3032 P1_R1222_U111 ; P1_U4852
g2240 nand P1_U3031 P1_U3506 ; P1_U4853
g2241 nand P1_U3030 P1_R1282_U11 ; P1_U4854
g2242 nand P1_U3036 P1_U3082 ; P1_U4855
g2243 nand P1_U3033 P1_ADD_99_U71 ; P1_U4856
g2244 nand P1_U3032 P1_R1222_U13 ; P1_U4857
g2245 nand P1_U3031 P1_U3509 ; P1_U4858
g2246 nand P1_U3030 P1_R1282_U84 ; P1_U4859
g2247 nand P1_U3036 P1_U3081 ; P1_U4860
g2248 nand P1_U3033 P1_ADD_99_U70 ; P1_U4861
g2249 nand P1_U3032 P1_R1222_U110 ; P1_U4862
g2250 nand P1_U3031 P1_U3512 ; P1_U4863
g2251 nand P1_U3030 P1_R1282_U12 ; P1_U4864
g2252 nand P1_U3036 P1_U3076 ; P1_U4865
g2253 nand P1_U3033 P1_ADD_99_U69 ; P1_U4866
g2254 nand P1_U3032 P1_R1222_U109 ; P1_U4867
g2255 nand P1_U3031 P1_U3514 ; P1_U4868
g2256 nand P1_U3030 P1_R1282_U82 ; P1_U4869
g2257 nand P1_U3036 P1_U3075 ; P1_U4870
g2258 nand P1_U3033 P1_ADD_99_U68 ; P1_U4871
g2259 nand P1_U3032 P1_R1222_U14 ; P1_U4872
g2260 nand P1_U3031 P1_U4025 ; P1_U4873
g2261 nand P1_U3030 P1_R1282_U13 ; P1_U4874
g2262 nand P1_U3036 P1_U3061 ; P1_U4875
g2263 nand P1_U3033 P1_ADD_99_U67 ; P1_U4876
g2264 nand P1_U3032 P1_R1222_U15 ; P1_U4877
g2265 nand P1_U3031 P1_U4024 ; P1_U4878
g2266 nand P1_U3030 P1_R1282_U78 ; P1_U4879
g2267 nand P1_U3036 P1_U3066 ; P1_U4880
g2268 nand P1_U3033 P1_ADD_99_U66 ; P1_U4881
g2269 nand P1_U3032 P1_R1222_U108 ; P1_U4882
g2270 nand P1_U3031 P1_U4023 ; P1_U4883
g2271 nand P1_U3030 P1_R1282_U14 ; P1_U4884
g2272 nand P1_U3036 P1_U3065 ; P1_U4885
g2273 nand P1_U3033 P1_ADD_99_U65 ; P1_U4886
g2274 nand P1_U3032 P1_R1222_U107 ; P1_U4887
g2275 nand P1_U3031 P1_U4022 ; P1_U4888
g2276 nand P1_U3030 P1_R1282_U76 ; P1_U4889
g2277 nand P1_U3036 P1_U3058 ; P1_U4890
g2278 nand P1_U3033 P1_ADD_99_U64 ; P1_U4891
g2279 nand P1_U3032 P1_R1222_U106 ; P1_U4892
g2280 nand P1_U3031 P1_U4021 ; P1_U4893
g2281 nand P1_U3030 P1_R1282_U15 ; P1_U4894
g2282 nand P1_U3036 P1_U3057 ; P1_U4895
g2283 nand P1_U3033 P1_ADD_99_U63 ; P1_U4896
g2284 nand P1_U3032 P1_R1222_U105 ; P1_U4897
g2285 nand P1_U3031 P1_U4020 ; P1_U4898
g2286 nand P1_U3030 P1_R1282_U74 ; P1_U4899
g2287 nand P1_U3036 P1_U3053 ; P1_U4900
g2288 nand P1_U3033 P1_ADD_99_U62 ; P1_U4901
g2289 nand P1_U3032 P1_R1222_U16 ; P1_U4902
g2290 nand P1_U3031 P1_U4019 ; P1_U4903
g2291 nand P1_U3030 P1_R1282_U16 ; P1_U4904
g2292 nand P1_U3036 P1_U3054 ; P1_U4905
g2293 nand P1_U3033 P1_ADD_99_U61 ; P1_U4906
g2294 nand P1_U3032 P1_R1222_U104 ; P1_U4907
g2295 nand P1_U3031 P1_U4018 ; P1_U4908
g2296 nand P1_U3030 P1_R1282_U72 ; P1_U4909
g2297 nand P1_U3036 P1_U3055 ; P1_U4910
g2298 nand P1_U3033 P1_ADD_99_U60 ; P1_U4911
g2299 nand P1_U3032 P1_R1222_U103 ; P1_U4912
g2300 nand P1_U3031 P1_U4017 ; P1_U4913
g2301 nand P1_U3030 P1_R1282_U17 ; P1_U4914
g2302 nand P1_U3033 P1_ADD_99_U5 ; P1_U4915
g2303 nand P1_U3032 P1_R1222_U102 ; P1_U4916
g2304 nand P1_U3031 P1_U4028 ; P1_U4917
g2305 nand P1_U3030 P1_R1282_U70 ; P1_U4918
g2306 nand P1_U3031 P1_U4027 ; P1_U4919
g2307 nand P1_U3030 P1_R1282_U19 ; P1_U4920
g2308 nand P1_U3031 P1_U4026 ; P1_U4921
g2309 nand P1_U3030 P1_R1282_U68 ; P1_U4922
g2310 nand P1_U3787 P1_U3786 P1_U3789 P1_U4769 P1_U3421 ; P1_U4923
g2311 nand P1_R1105_U13 P1_U3042 ; P1_U4924
g2312 nand P1_U3040 P1_U3452 ; P1_U4925
g2313 nand P1_R1162_U13 P1_U3038 ; P1_U4926
g2314 nand P1_U4925 P1_U4924 P1_U4926 ; P1_U4927
g2315 nand P1_U3425 P1_U3372 ; P1_U4928
g2316 nand P1_U5786 P1_U4928 ; P1_U4929
g2317 nand P1_U4929 P1_U3954 ; P1_U4930
g2318 not P1_U3085 ; P1_U4931
g2319 not P1_U3428 ; P1_U4932
g2320 nand P1_U3044 P1_U4927 ; P1_U4933
g2321 nand P1_U3043 P1_R1105_U13 ; P1_U4934
g2322 nand P1_U3086 P1_REG3_REG_19__SCAN_IN ; P1_U4935
g2323 nand P1_U3041 P1_U3452 ; P1_U4936
g2324 nand P1_U3039 P1_R1162_U13 ; P1_U4937
g2325 nand P1_U4932 P1_ADDR_REG_19__SCAN_IN ; P1_U4938
g2326 nand P1_R1105_U75 P1_U3042 ; P1_U4939
g2327 nand P1_U3040 P1_U3511 ; P1_U4940
g2328 nand P1_R1162_U75 P1_U3038 ; P1_U4941
g2329 nand P1_U4940 P1_U4939 P1_U4941 ; P1_U4942
g2330 nand P1_U3044 P1_U4942 ; P1_U4943
g2331 nand P1_R1105_U75 P1_U3043 ; P1_U4944
g2332 nand P1_U3086 P1_REG3_REG_18__SCAN_IN ; P1_U4945
g2333 nand P1_U3041 P1_U3511 ; P1_U4946
g2334 nand P1_R1162_U75 P1_U3039 ; P1_U4947
g2335 nand P1_U4932 P1_ADDR_REG_18__SCAN_IN ; P1_U4948
g2336 nand P1_R1105_U12 P1_U3042 ; P1_U4949
g2337 nand P1_U3040 P1_U3508 ; P1_U4950
g2338 nand P1_R1162_U12 P1_U3038 ; P1_U4951
g2339 nand P1_U4950 P1_U4949 P1_U4951 ; P1_U4952
g2340 nand P1_U3044 P1_U4952 ; P1_U4953
g2341 nand P1_R1105_U12 P1_U3043 ; P1_U4954
g2342 nand P1_U3086 P1_REG3_REG_17__SCAN_IN ; P1_U4955
g2343 nand P1_U3041 P1_U3508 ; P1_U4956
g2344 nand P1_R1162_U12 P1_U3039 ; P1_U4957
g2345 nand P1_U4932 P1_ADDR_REG_17__SCAN_IN ; P1_U4958
g2346 nand P1_R1105_U76 P1_U3042 ; P1_U4959
g2347 nand P1_U3040 P1_U3505 ; P1_U4960
g2348 nand P1_R1162_U76 P1_U3038 ; P1_U4961
g2349 nand P1_U4960 P1_U4959 P1_U4961 ; P1_U4962
g2350 nand P1_U3044 P1_U4962 ; P1_U4963
g2351 nand P1_R1105_U76 P1_U3043 ; P1_U4964
g2352 nand P1_U3086 P1_REG3_REG_16__SCAN_IN ; P1_U4965
g2353 nand P1_U3041 P1_U3505 ; P1_U4966
g2354 nand P1_R1162_U76 P1_U3039 ; P1_U4967
g2355 nand P1_U4932 P1_ADDR_REG_16__SCAN_IN ; P1_U4968
g2356 nand P1_R1105_U77 P1_U3042 ; P1_U4969
g2357 nand P1_U3040 P1_U3502 ; P1_U4970
g2358 nand P1_R1162_U77 P1_U3038 ; P1_U4971
g2359 nand P1_U4970 P1_U4969 P1_U4971 ; P1_U4972
g2360 nand P1_U3044 P1_U4972 ; P1_U4973
g2361 nand P1_R1105_U77 P1_U3043 ; P1_U4974
g2362 nand P1_U3086 P1_REG3_REG_15__SCAN_IN ; P1_U4975
g2363 nand P1_U3041 P1_U3502 ; P1_U4976
g2364 nand P1_R1162_U77 P1_U3039 ; P1_U4977
g2365 nand P1_U4932 P1_ADDR_REG_15__SCAN_IN ; P1_U4978
g2366 nand P1_R1105_U78 P1_U3042 ; P1_U4979
g2367 nand P1_U3040 P1_U3499 ; P1_U4980
g2368 nand P1_R1162_U78 P1_U3038 ; P1_U4981
g2369 nand P1_U4980 P1_U4979 P1_U4981 ; P1_U4982
g2370 nand P1_U3044 P1_U4982 ; P1_U4983
g2371 nand P1_R1105_U78 P1_U3043 ; P1_U4984
g2372 nand P1_U3086 P1_REG3_REG_14__SCAN_IN ; P1_U4985
g2373 nand P1_U3041 P1_U3499 ; P1_U4986
g2374 nand P1_R1162_U78 P1_U3039 ; P1_U4987
g2375 nand P1_U4932 P1_ADDR_REG_14__SCAN_IN ; P1_U4988
g2376 nand P1_R1105_U11 P1_U3042 ; P1_U4989
g2377 nand P1_U3040 P1_U3496 ; P1_U4990
g2378 nand P1_R1162_U11 P1_U3038 ; P1_U4991
g2379 nand P1_U4990 P1_U4989 P1_U4991 ; P1_U4992
g2380 nand P1_U3044 P1_U4992 ; P1_U4993
g2381 nand P1_R1105_U11 P1_U3043 ; P1_U4994
g2382 nand P1_U3086 P1_REG3_REG_13__SCAN_IN ; P1_U4995
g2383 nand P1_U3041 P1_U3496 ; P1_U4996
g2384 nand P1_R1162_U11 P1_U3039 ; P1_U4997
g2385 nand P1_U4932 P1_ADDR_REG_13__SCAN_IN ; P1_U4998
g2386 nand P1_R1105_U79 P1_U3042 ; P1_U4999
g2387 nand P1_U3040 P1_U3493 ; P1_U5000
g2388 nand P1_R1162_U79 P1_U3038 ; P1_U5001
g2389 nand P1_U5000 P1_U4999 P1_U5001 ; P1_U5002
g2390 nand P1_U3044 P1_U5002 ; P1_U5003
g2391 nand P1_R1105_U79 P1_U3043 ; P1_U5004
g2392 nand P1_U3086 P1_REG3_REG_12__SCAN_IN ; P1_U5005
g2393 nand P1_U3041 P1_U3493 ; P1_U5006
g2394 nand P1_R1162_U79 P1_U3039 ; P1_U5007
g2395 nand P1_U4932 P1_ADDR_REG_12__SCAN_IN ; P1_U5008
g2396 nand P1_R1105_U80 P1_U3042 ; P1_U5009
g2397 nand P1_U3040 P1_U3490 ; P1_U5010
g2398 nand P1_R1162_U80 P1_U3038 ; P1_U5011
g2399 nand P1_U5010 P1_U5009 P1_U5011 ; P1_U5012
g2400 nand P1_U3044 P1_U5012 ; P1_U5013
g2401 nand P1_R1105_U80 P1_U3043 ; P1_U5014
g2402 nand P1_U3086 P1_REG3_REG_11__SCAN_IN ; P1_U5015
g2403 nand P1_U3041 P1_U3490 ; P1_U5016
g2404 nand P1_R1162_U80 P1_U3039 ; P1_U5017
g2405 nand P1_U4932 P1_ADDR_REG_11__SCAN_IN ; P1_U5018
g2406 nand P1_R1105_U10 P1_U3042 ; P1_U5019
g2407 nand P1_U3040 P1_U3487 ; P1_U5020
g2408 nand P1_R1162_U10 P1_U3038 ; P1_U5021
g2409 nand P1_U5020 P1_U5019 P1_U5021 ; P1_U5022
g2410 nand P1_U3044 P1_U5022 ; P1_U5023
g2411 nand P1_R1105_U10 P1_U3043 ; P1_U5024
g2412 nand P1_U3086 P1_REG3_REG_10__SCAN_IN ; P1_U5025
g2413 nand P1_U3041 P1_U3487 ; P1_U5026
g2414 nand P1_R1162_U10 P1_U3039 ; P1_U5027
g2415 nand P1_U4932 P1_ADDR_REG_10__SCAN_IN ; P1_U5028
g2416 nand P1_R1105_U70 P1_U3042 ; P1_U5029
g2417 nand P1_U3040 P1_U3484 ; P1_U5030
g2418 nand P1_R1162_U70 P1_U3038 ; P1_U5031
g2419 nand P1_U5030 P1_U5029 P1_U5031 ; P1_U5032
g2420 nand P1_U3044 P1_U5032 ; P1_U5033
g2421 nand P1_R1105_U70 P1_U3043 ; P1_U5034
g2422 nand P1_U3086 P1_REG3_REG_9__SCAN_IN ; P1_U5035
g2423 nand P1_U3041 P1_U3484 ; P1_U5036
g2424 nand P1_R1162_U70 P1_U3039 ; P1_U5037
g2425 nand P1_U4932 P1_ADDR_REG_9__SCAN_IN ; P1_U5038
g2426 nand P1_R1105_U71 P1_U3042 ; P1_U5039
g2427 nand P1_U3040 P1_U3481 ; P1_U5040
g2428 nand P1_R1162_U71 P1_U3038 ; P1_U5041
g2429 nand P1_U5040 P1_U5039 P1_U5041 ; P1_U5042
g2430 nand P1_U3044 P1_U5042 ; P1_U5043
g2431 nand P1_R1105_U71 P1_U3043 ; P1_U5044
g2432 nand P1_U3086 P1_REG3_REG_8__SCAN_IN ; P1_U5045
g2433 nand P1_U3041 P1_U3481 ; P1_U5046
g2434 nand P1_R1162_U71 P1_U3039 ; P1_U5047
g2435 nand P1_U4932 P1_ADDR_REG_8__SCAN_IN ; P1_U5048
g2436 nand P1_R1105_U16 P1_U3042 ; P1_U5049
g2437 nand P1_U3040 P1_U3478 ; P1_U5050
g2438 nand P1_R1162_U16 P1_U3038 ; P1_U5051
g2439 nand P1_U5050 P1_U5049 P1_U5051 ; P1_U5052
g2440 nand P1_U3044 P1_U5052 ; P1_U5053
g2441 nand P1_R1105_U16 P1_U3043 ; P1_U5054
g2442 nand P1_U3086 P1_REG3_REG_7__SCAN_IN ; P1_U5055
g2443 nand P1_U3041 P1_U3478 ; P1_U5056
g2444 nand P1_R1162_U16 P1_U3039 ; P1_U5057
g2445 nand P1_U4932 P1_ADDR_REG_7__SCAN_IN ; P1_U5058
g2446 nand P1_R1105_U72 P1_U3042 ; P1_U5059
g2447 nand P1_U3040 P1_U3475 ; P1_U5060
g2448 nand P1_R1162_U72 P1_U3038 ; P1_U5061
g2449 nand P1_U5060 P1_U5059 P1_U5061 ; P1_U5062
g2450 nand P1_U3044 P1_U5062 ; P1_U5063
g2451 nand P1_R1105_U72 P1_U3043 ; P1_U5064
g2452 nand P1_U3086 P1_REG3_REG_6__SCAN_IN ; P1_U5065
g2453 nand P1_U3041 P1_U3475 ; P1_U5066
g2454 nand P1_R1162_U72 P1_U3039 ; P1_U5067
g2455 nand P1_U4932 P1_ADDR_REG_6__SCAN_IN ; P1_U5068
g2456 nand P1_R1105_U15 P1_U3042 ; P1_U5069
g2457 nand P1_U3040 P1_U3472 ; P1_U5070
g2458 nand P1_R1162_U15 P1_U3038 ; P1_U5071
g2459 nand P1_U5070 P1_U5069 P1_U5071 ; P1_U5072
g2460 nand P1_U3044 P1_U5072 ; P1_U5073
g2461 nand P1_R1105_U15 P1_U3043 ; P1_U5074
g2462 nand P1_U3086 P1_REG3_REG_5__SCAN_IN ; P1_U5075
g2463 nand P1_U3041 P1_U3472 ; P1_U5076
g2464 nand P1_R1162_U15 P1_U3039 ; P1_U5077
g2465 nand P1_U4932 P1_ADDR_REG_5__SCAN_IN ; P1_U5078
g2466 nand P1_R1105_U73 P1_U3042 ; P1_U5079
g2467 nand P1_U3040 P1_U3469 ; P1_U5080
g2468 nand P1_R1162_U73 P1_U3038 ; P1_U5081
g2469 nand P1_U5080 P1_U5079 P1_U5081 ; P1_U5082
g2470 nand P1_U3044 P1_U5082 ; P1_U5083
g2471 nand P1_R1105_U73 P1_U3043 ; P1_U5084
g2472 nand P1_U3086 P1_REG3_REG_4__SCAN_IN ; P1_U5085
g2473 nand P1_U3041 P1_U3469 ; P1_U5086
g2474 nand P1_R1162_U73 P1_U3039 ; P1_U5087
g2475 nand P1_U4932 P1_ADDR_REG_4__SCAN_IN ; P1_U5088
g2476 nand P1_R1105_U74 P1_U3042 ; P1_U5089
g2477 nand P1_U3040 P1_U3466 ; P1_U5090
g2478 nand P1_R1162_U74 P1_U3038 ; P1_U5091
g2479 nand P1_U5090 P1_U5089 P1_U5091 ; P1_U5092
g2480 nand P1_U3044 P1_U5092 ; P1_U5093
g2481 nand P1_R1105_U74 P1_U3043 ; P1_U5094
g2482 nand P1_U3086 P1_REG3_REG_3__SCAN_IN ; P1_U5095
g2483 nand P1_U3041 P1_U3466 ; P1_U5096
g2484 nand P1_R1162_U74 P1_U3039 ; P1_U5097
g2485 nand P1_U4932 P1_ADDR_REG_3__SCAN_IN ; P1_U5098
g2486 nand P1_R1105_U14 P1_U3042 ; P1_U5099
g2487 nand P1_U3040 P1_U3463 ; P1_U5100
g2488 nand P1_R1162_U14 P1_U3038 ; P1_U5101
g2489 nand P1_U5100 P1_U5099 P1_U5101 ; P1_U5102
g2490 nand P1_U3044 P1_U5102 ; P1_U5103
g2491 nand P1_R1105_U14 P1_U3043 ; P1_U5104
g2492 nand P1_U3086 P1_REG3_REG_2__SCAN_IN ; P1_U5105
g2493 nand P1_U3041 P1_U3463 ; P1_U5106
g2494 nand P1_R1162_U14 P1_U3039 ; P1_U5107
g2495 nand P1_U4932 P1_ADDR_REG_2__SCAN_IN ; P1_U5108
g2496 nand P1_R1105_U68 P1_U3042 ; P1_U5109
g2497 nand P1_U3040 P1_U3460 ; P1_U5110
g2498 nand P1_R1162_U68 P1_U3038 ; P1_U5111
g2499 nand P1_U5110 P1_U5109 P1_U5111 ; P1_U5112
g2500 nand P1_U3044 P1_U5112 ; P1_U5113
g2501 nand P1_R1105_U68 P1_U3043 ; P1_U5114
g2502 nand P1_U3086 P1_REG3_REG_1__SCAN_IN ; P1_U5115
g2503 nand P1_U3041 P1_U3460 ; P1_U5116
g2504 nand P1_R1162_U68 P1_U3039 ; P1_U5117
g2505 nand P1_U4932 P1_ADDR_REG_1__SCAN_IN ; P1_U5118
g2506 nand P1_R1105_U69 P1_U3042 ; P1_U5119
g2507 nand P1_U3040 P1_U3454 ; P1_U5120
g2508 nand P1_R1162_U69 P1_U3038 ; P1_U5121
g2509 nand P1_U5120 P1_U5119 P1_U5121 ; P1_U5122
g2510 nand P1_U3044 P1_U5122 ; P1_U5123
g2511 nand P1_R1105_U69 P1_U3043 ; P1_U5124
g2512 nand P1_U3086 P1_REG3_REG_0__SCAN_IN ; P1_U5125
g2513 nand P1_U3041 P1_U3454 ; P1_U5126
g2514 nand P1_R1162_U69 P1_U3039 ; P1_U5127
g2515 nand P1_U4932 P1_ADDR_REG_0__SCAN_IN ; P1_U5128
g2516 not P1_U3991 ; P1_U5129
g2517 nand P1_U6277 P1_U6276 P1_U3990 ; P1_U5130
g2518 nand P1_U3370 P1_U3373 ; P1_U5131
g2519 nand P1_U5802 P1_U3451 ; P1_U5132
g2520 nand P1_U3422 P1_U5132 ; P1_U5133
g2521 nand P1_U6279 P1_U6278 P1_U5772 ; P1_U5134
g2522 nand P1_U6281 P1_U6280 P1_U3845 ; P1_U5135
g2523 nand P1_U3022 P1_U4029 P1_U3432 ; P1_U5136
g2524 nand P1_U4043 P1_U5134 ; P1_U5137
g2525 nand P1_U5135 P1_B_REG_SCAN_IN ; P1_U5138
g2526 nand P1_U3037 P1_U3079 ; P1_U5139
g2527 nand P1_U3035 P1_U3073 ; P1_U5140
g2528 nand P1_ADD_99_U73 P1_U3434 ; P1_U5141
g2529 nand P1_U5141 P1_U5139 P1_U5140 ; P1_U5142
g2530 not P1_U3152 ; P1_U5143
g2531 nand P1_U3423 P1_U3999 ; P1_U5144
g2532 nand P1_U6283 P1_U6282 P1_U3849 P1_U3848 ; P1_U5145
g2533 nand P1_U5145 P1_U3434 ; P1_U5146
g2534 nand P1_U4012 P1_U5146 ; P1_U5147
g2535 nand P1_U3022 P1_U5147 ; P1_U5148
g2536 nand P1_U3503 P1_U5770 ; P1_U5149
g2537 nand P1_ADD_99_U73 P1_U5769 ; P1_U5150
g2538 nand P1_R1165_U105 P1_U3026 ; P1_U5151
g2539 nand P1_U4037 P1_U5142 ; P1_U5152
g2540 nand P1_U3086 P1_REG3_REG_15__SCAN_IN ; P1_U5153
g2541 nand P1_U3037 P1_U3058 ; P1_U5154
g2542 nand P1_U3035 P1_U3053 ; P1_U5155
g2543 nand P1_ADD_99_U62 P1_U3434 ; P1_U5156
g2544 nand P1_U5156 P1_U5154 P1_U5155 ; P1_U5157
g2545 nand P1_U4015 P1_U3426 ; P1_U5158
g2546 nand P1_U3421 P1_U5158 ; P1_U5159
g2547 nand P1_U3045 P1_U4019 ; P1_U5160
g2548 nand P1_ADD_99_U62 P1_U5769 ; P1_U5161
g2549 nand P1_R1165_U12 P1_U3026 ; P1_U5162
g2550 nand P1_U4037 P1_U5157 ; P1_U5163
g2551 nand P1_U3086 P1_REG3_REG_26__SCAN_IN ; P1_U5164
g2552 nand P1_U3037 P1_U3067 ; P1_U5165
g2553 nand P1_U3035 P1_U3070 ; P1_U5166
g2554 nand P1_ADD_99_U57 P1_U3434 ; P1_U5167
g2555 nand P1_U5166 P1_U5165 P1_U5167 ; P1_U5168
g2556 nand P1_U3476 P1_U5770 ; P1_U5169
g2557 nand P1_ADD_99_U57 P1_U5769 ; P1_U5170
g2558 nand P1_R1165_U90 P1_U3026 ; P1_U5171
g2559 nand P1_U4037 P1_U5168 ; P1_U5172
g2560 nand P1_U3086 P1_REG3_REG_6__SCAN_IN ; P1_U5173
g2561 nand P1_U3037 P1_U3069 ; P1_U5174
g2562 nand P1_U3035 P1_U3081 ; P1_U5175
g2563 nand P1_ADD_99_U70 P1_U3434 ; P1_U5176
g2564 nand P1_U5176 P1_U5174 P1_U5175 ; P1_U5177
g2565 nand P1_U3512 P1_U5770 ; P1_U5178
g2566 nand P1_ADD_99_U70 P1_U5769 ; P1_U5179
g2567 nand P1_R1165_U103 P1_U3026 ; P1_U5180
g2568 nand P1_U4037 P1_U5177 ; P1_U5181
g2569 nand P1_U3086 P1_REG3_REG_18__SCAN_IN ; P1_U5182
g2570 nand P1_U3037 P1_U3078 ; P1_U5183
g2571 nand P1_U3035 P1_U3064 ; P1_U5184
g2572 nand P1_U3434 P1_REG3_REG_2__SCAN_IN ; P1_U5185
g2573 nand P1_U5184 P1_U5183 P1_U5185 ; P1_U5186
g2574 nand P1_U3464 P1_U5770 ; P1_U5187
g2575 nand P1_U5769 P1_REG3_REG_2__SCAN_IN ; P1_U5188
g2576 nand P1_R1165_U93 P1_U3026 ; P1_U5189
g2577 nand P1_U4037 P1_U5186 ; P1_U5190
g2578 nand P1_U3086 P1_REG3_REG_2__SCAN_IN ; P1_U5191
g2579 nand P1_U3037 P1_U3062 ; P1_U5192
g2580 nand P1_U3035 P1_U3072 ; P1_U5193
g2581 nand P1_ADD_99_U77 P1_U3434 ; P1_U5194
g2582 nand P1_U5193 P1_U5192 P1_U5194 ; P1_U5195
g2583 nand P1_U3491 P1_U5770 ; P1_U5196
g2584 nand P1_ADD_99_U77 P1_U5769 ; P1_U5197
g2585 nand P1_R1165_U108 P1_U3026 ; P1_U5198
g2586 nand P1_U4037 P1_U5195 ; P1_U5199
g2587 nand P1_U3086 P1_REG3_REG_11__SCAN_IN ; P1_U5200
g2588 nand P1_U3037 P1_U3075 ; P1_U5201
g2589 nand P1_U3035 P1_U3066 ; P1_U5202
g2590 nand P1_ADD_99_U66 P1_U3434 ; P1_U5203
g2591 nand P1_U5203 P1_U5201 P1_U5202 ; P1_U5204
g2592 nand P1_U3045 P1_U4023 ; P1_U5205
g2593 nand P1_ADD_99_U66 P1_U5769 ; P1_U5206
g2594 nand P1_R1165_U99 P1_U3026 ; P1_U5207
g2595 nand P1_U4037 P1_U5204 ; P1_U5208
g2596 nand P1_U3086 P1_REG3_REG_22__SCAN_IN ; P1_U5209
g2597 nand P1_U3037 P1_U3072 ; P1_U5210
g2598 nand P1_U3035 P1_U3079 ; P1_U5211
g2599 nand P1_ADD_99_U75 P1_U3434 ; P1_U5212
g2600 nand P1_U5212 P1_U5210 P1_U5211 ; P1_U5213
g2601 nand P1_U3497 P1_U5770 ; P1_U5214
g2602 nand P1_ADD_99_U75 P1_U5769 ; P1_U5215
g2603 nand P1_R1165_U9 P1_U3026 ; P1_U5216
g2604 nand P1_U4037 P1_U5213 ; P1_U5217
g2605 nand P1_U3086 P1_REG3_REG_13__SCAN_IN ; P1_U5218
g2606 nand P1_U3037 P1_U3081 ; P1_U5219
g2607 nand P1_U3035 P1_U3075 ; P1_U5220
g2608 nand P1_ADD_99_U68 P1_U3434 ; P1_U5221
g2609 nand P1_U5221 P1_U5219 P1_U5220 ; P1_U5222
g2610 nand P1_U3045 P1_U4025 ; P1_U5223
g2611 nand P1_ADD_99_U68 P1_U5769 ; P1_U5224
g2612 nand P1_R1165_U100 P1_U3026 ; P1_U5225
g2613 nand P1_U4037 P1_U5222 ; P1_U5226
g2614 nand P1_U3086 P1_REG3_REG_20__SCAN_IN ; P1_U5227
g2615 nand P1_U3435 P1_U3433 ; P1_U5228
g2616 nand P1_U5228 P1_U3434 ; P1_U5229
g2617 nand P1_U3050 P1_U5229 ; P1_U5230
g2618 nand P1_U3858 P1_U3035 ; P1_U5231
g2619 nand P1_U3456 P1_U5770 ; P1_U5232
g2620 nand P1_U5230 P1_REG3_REG_0__SCAN_IN ; P1_U5233
g2621 nand P1_R1165_U87 P1_U3026 ; P1_U5234
g2622 nand P1_U3086 P1_REG3_REG_0__SCAN_IN ; P1_U5235
g2623 nand P1_U3037 P1_U3084 ; P1_U5236
g2624 nand P1_U3035 P1_U3062 ; P1_U5237
g2625 nand P1_ADD_99_U54 P1_U3434 ; P1_U5238
g2626 nand P1_U5237 P1_U5236 P1_U5238 ; P1_U5239
g2627 nand P1_U3485 P1_U5770 ; P1_U5240
g2628 nand P1_ADD_99_U54 P1_U5769 ; P1_U5241
g2629 nand P1_R1165_U88 P1_U3026 ; P1_U5242
g2630 nand P1_U4037 P1_U5239 ; P1_U5243
g2631 nand P1_U3086 P1_REG3_REG_9__SCAN_IN ; P1_U5244
g2632 nand P1_U3037 P1_U3064 ; P1_U5245
g2633 nand P1_U3035 P1_U3067 ; P1_U5246
g2634 nand P1_ADD_99_U59 P1_U3434 ; P1_U5247
g2635 nand P1_U5246 P1_U5245 P1_U5247 ; P1_U5248
g2636 nand P1_U3470 P1_U5770 ; P1_U5249
g2637 nand P1_ADD_99_U59 P1_U5769 ; P1_U5250
g2638 nand P1_R1165_U92 P1_U3026 ; P1_U5251
g2639 nand P1_U4037 P1_U5248 ; P1_U5252
g2640 nand P1_U3086 P1_REG3_REG_4__SCAN_IN ; P1_U5253
g2641 nand P1_U3037 P1_U3066 ; P1_U5254
g2642 nand P1_U3035 P1_U3058 ; P1_U5255
g2643 nand P1_ADD_99_U64 P1_U3434 ; P1_U5256
g2644 nand P1_U5256 P1_U5254 P1_U5255 ; P1_U5257
g2645 nand P1_U3045 P1_U4021 ; P1_U5258
g2646 nand P1_ADD_99_U64 P1_U5769 ; P1_U5259
g2647 nand P1_R1165_U97 P1_U3026 ; P1_U5260
g2648 nand P1_U4037 P1_U5257 ; P1_U5261
g2649 nand P1_U3086 P1_REG3_REG_24__SCAN_IN ; P1_U5262
g2650 nand P1_U3037 P1_U3073 ; P1_U5263
g2651 nand P1_U3035 P1_U3082 ; P1_U5264
g2652 nand P1_ADD_99_U71 P1_U3434 ; P1_U5265
g2653 nand P1_U5265 P1_U5263 P1_U5264 ; P1_U5266
g2654 nand P1_U3509 P1_U5770 ; P1_U5267
g2655 nand P1_ADD_99_U71 P1_U5769 ; P1_U5268
g2656 nand P1_R1165_U10 P1_U3026 ; P1_U5269
g2657 nand P1_U4037 P1_U5266 ; P1_U5270
g2658 nand P1_U3086 P1_REG3_REG_17__SCAN_IN ; P1_U5271
g2659 nand P1_U3037 P1_U3060 ; P1_U5272
g2660 nand P1_U3035 P1_U3071 ; P1_U5273
g2661 nand P1_ADD_99_U58 P1_U3434 ; P1_U5274
g2662 nand P1_U5273 P1_U5272 P1_U5274 ; P1_U5275
g2663 nand P1_U3473 P1_U5770 ; P1_U5276
g2664 nand P1_ADD_99_U58 P1_U5769 ; P1_U5277
g2665 nand P1_R1165_U91 P1_U3026 ; P1_U5278
g2666 nand P1_U4037 P1_U5275 ; P1_U5279
g2667 nand P1_U3086 P1_REG3_REG_5__SCAN_IN ; P1_U5280
g2668 nand P1_U3037 P1_U3074 ; P1_U5281
g2669 nand P1_U3035 P1_U3069 ; P1_U5282
g2670 nand P1_ADD_99_U72 P1_U3434 ; P1_U5283
g2671 nand P1_U5283 P1_U5281 P1_U5282 ; P1_U5284
g2672 nand P1_U3506 P1_U5770 ; P1_U5285
g2673 nand P1_ADD_99_U72 P1_U5769 ; P1_U5286
g2674 nand P1_R1165_U104 P1_U3026 ; P1_U5287
g2675 nand P1_U4037 P1_U5284 ; P1_U5288
g2676 nand P1_U3086 P1_REG3_REG_16__SCAN_IN ; P1_U5289
g2677 nand P1_U3037 P1_U3065 ; P1_U5290
g2678 nand P1_U3035 P1_U3057 ; P1_U5291
g2679 nand P1_ADD_99_U63 P1_U3434 ; P1_U5292
g2680 nand P1_U5292 P1_U5290 P1_U5291 ; P1_U5293
g2681 nand P1_U3045 P1_U4020 ; P1_U5294
g2682 nand P1_ADD_99_U63 P1_U5769 ; P1_U5295
g2683 nand P1_R1165_U96 P1_U3026 ; P1_U5296
g2684 nand P1_U4037 P1_U5293 ; P1_U5297
g2685 nand P1_U3086 P1_REG3_REG_25__SCAN_IN ; P1_U5298
g2686 nand P1_U3037 P1_U3063 ; P1_U5299
g2687 nand P1_U3035 P1_U3080 ; P1_U5300
g2688 nand P1_ADD_99_U76 P1_U3434 ; P1_U5301
g2689 nand P1_U5301 P1_U5299 P1_U5300 ; P1_U5302
g2690 nand P1_U3494 P1_U5770 ; P1_U5303
g2691 nand P1_ADD_99_U76 P1_U5769 ; P1_U5304
g2692 nand P1_R1165_U107 P1_U3026 ; P1_U5305
g2693 nand P1_U4037 P1_U5302 ; P1_U5306
g2694 nand P1_U3086 P1_REG3_REG_12__SCAN_IN ; P1_U5307
g2695 nand P1_U3037 P1_U3076 ; P1_U5308
g2696 nand P1_U3035 P1_U3061 ; P1_U5309
g2697 nand P1_ADD_99_U67 P1_U3434 ; P1_U5310
g2698 nand P1_U5310 P1_U5308 P1_U5309 ; P1_U5311
g2699 nand P1_U3045 P1_U4024 ; P1_U5312
g2700 nand P1_ADD_99_U67 P1_U5769 ; P1_U5313
g2701 nand P1_R1165_U11 P1_U3026 ; P1_U5314
g2702 nand P1_U4037 P1_U5311 ; P1_U5315
g2703 nand P1_U3086 P1_REG3_REG_21__SCAN_IN ; P1_U5316
g2704 nand P1_U3037 P1_U3077 ; P1_U5317
g2705 nand P1_U3035 P1_U3068 ; P1_U5318
g2706 nand P1_U3434 P1_REG3_REG_1__SCAN_IN ; P1_U5319
g2707 nand P1_U5318 P1_U5317 P1_U5319 ; P1_U5320
g2708 nand P1_U3461 P1_U5770 ; P1_U5321
g2709 nand P1_U5769 P1_REG3_REG_1__SCAN_IN ; P1_U5322
g2710 nand P1_R1165_U101 P1_U3026 ; P1_U5323
g2711 nand P1_U4037 P1_U5320 ; P1_U5324
g2712 nand P1_U3086 P1_REG3_REG_1__SCAN_IN ; P1_U5325
g2713 nand P1_U3037 P1_U3070 ; P1_U5326
g2714 nand P1_U3035 P1_U3083 ; P1_U5327
g2715 nand P1_ADD_99_U55 P1_U3434 ; P1_U5328
g2716 nand P1_U5327 P1_U5326 P1_U5328 ; P1_U5329
g2717 nand P1_U3482 P1_U5770 ; P1_U5330
g2718 nand P1_ADD_99_U55 P1_U5769 ; P1_U5331
g2719 nand P1_R1165_U89 P1_U3026 ; P1_U5332
g2720 nand P1_U4037 P1_U5329 ; P1_U5333
g2721 nand P1_U3086 P1_REG3_REG_8__SCAN_IN ; P1_U5334
g2722 nand P1_U3037 P1_U3053 ; P1_U5335
g2723 nand P1_U3035 P1_U3055 ; P1_U5336
g2724 nand P1_ADD_99_U60 P1_U3434 ; P1_U5337
g2725 nand P1_U5336 P1_U5335 P1_U5337 ; P1_U5338
g2726 nand P1_U3045 P1_U4017 ; P1_U5339
g2727 nand P1_ADD_99_U60 P1_U5769 ; P1_U5340
g2728 nand P1_R1165_U94 P1_U3026 ; P1_U5341
g2729 nand P1_U4037 P1_U5338 ; P1_U5342
g2730 nand P1_U3086 P1_REG3_REG_28__SCAN_IN ; P1_U5343
g2731 nand P1_U3037 P1_U3082 ; P1_U5344
g2732 nand P1_U3035 P1_U3076 ; P1_U5345
g2733 nand P1_ADD_99_U69 P1_U3434 ; P1_U5346
g2734 nand P1_U5346 P1_U5344 P1_U5345 ; P1_U5347
g2735 nand P1_U3514 P1_U5770 ; P1_U5348
g2736 nand P1_ADD_99_U69 P1_U5769 ; P1_U5349
g2737 nand P1_R1165_U102 P1_U3026 ; P1_U5350
g2738 nand P1_U4037 P1_U5347 ; P1_U5351
g2739 nand P1_U3086 P1_REG3_REG_19__SCAN_IN ; P1_U5352
g2740 nand P1_U3037 P1_U3068 ; P1_U5353
g2741 nand P1_U3035 P1_U3060 ; P1_U5354
g2742 nand P1_ADD_99_U4 P1_U3434 ; P1_U5355
g2743 nand P1_U5354 P1_U5353 P1_U5355 ; P1_U5356
g2744 nand P1_U3467 P1_U5770 ; P1_U5357
g2745 nand P1_ADD_99_U4 P1_U5769 ; P1_U5358
g2746 nand P1_R1165_U13 P1_U3026 ; P1_U5359
g2747 nand P1_U4037 P1_U5356 ; P1_U5360
g2748 nand P1_U3086 P1_REG3_REG_3__SCAN_IN ; P1_U5361
g2749 nand P1_U3037 P1_U3083 ; P1_U5362
g2750 nand P1_U3035 P1_U3063 ; P1_U5363
g2751 nand P1_ADD_99_U78 P1_U3434 ; P1_U5364
g2752 nand P1_U5363 P1_U5362 P1_U5364 ; P1_U5365
g2753 nand P1_U3488 P1_U5770 ; P1_U5366
g2754 nand P1_ADD_99_U78 P1_U5769 ; P1_U5367
g2755 nand P1_R1165_U109 P1_U3026 ; P1_U5368
g2756 nand P1_U4037 P1_U5365 ; P1_U5369
g2757 nand P1_U3086 P1_REG3_REG_10__SCAN_IN ; P1_U5370
g2758 nand P1_U3037 P1_U3061 ; P1_U5371
g2759 nand P1_U3035 P1_U3065 ; P1_U5372
g2760 nand P1_ADD_99_U65 P1_U3434 ; P1_U5373
g2761 nand P1_U5373 P1_U5371 P1_U5372 ; P1_U5374
g2762 nand P1_U3045 P1_U4022 ; P1_U5375
g2763 nand P1_ADD_99_U65 P1_U5769 ; P1_U5376
g2764 nand P1_R1165_U98 P1_U3026 ; P1_U5377
g2765 nand P1_U4037 P1_U5374 ; P1_U5378
g2766 nand P1_U3086 P1_REG3_REG_23__SCAN_IN ; P1_U5379
g2767 nand P1_U3037 P1_U3080 ; P1_U5380
g2768 nand P1_U3035 P1_U3074 ; P1_U5381
g2769 nand P1_ADD_99_U74 P1_U3434 ; P1_U5382
g2770 nand P1_U5382 P1_U5380 P1_U5381 ; P1_U5383
g2771 nand P1_U3500 P1_U5770 ; P1_U5384
g2772 nand P1_ADD_99_U74 P1_U5769 ; P1_U5385
g2773 nand P1_R1165_U106 P1_U3026 ; P1_U5386
g2774 nand P1_U4037 P1_U5383 ; P1_U5387
g2775 nand P1_U3086 P1_REG3_REG_14__SCAN_IN ; P1_U5388
g2776 nand P1_U3037 P1_U3057 ; P1_U5389
g2777 nand P1_U3035 P1_U3054 ; P1_U5390
g2778 nand P1_ADD_99_U61 P1_U3434 ; P1_U5391
g2779 nand P1_U5391 P1_U5389 P1_U5390 ; P1_U5392
g2780 nand P1_U3045 P1_U4018 ; P1_U5393
g2781 nand P1_ADD_99_U61 P1_U5769 ; P1_U5394
g2782 nand P1_R1165_U95 P1_U3026 ; P1_U5395
g2783 nand P1_U4037 P1_U5392 ; P1_U5396
g2784 nand P1_U3086 P1_REG3_REG_27__SCAN_IN ; P1_U5397
g2785 nand P1_U3037 P1_U3071 ; P1_U5398
g2786 nand P1_U3035 P1_U3084 ; P1_U5399
g2787 nand P1_ADD_99_U56 P1_U3434 ; P1_U5400
g2788 nand P1_U5399 P1_U5398 P1_U5400 ; P1_U5401
g2789 nand P1_U3479 P1_U5770 ; P1_U5402
g2790 nand P1_ADD_99_U56 P1_U5769 ; P1_U5403
g2791 nand P1_R1165_U14 P1_U3026 ; P1_U5404
g2792 nand P1_U4037 P1_U5401 ; P1_U5405
g2793 nand P1_U3086 P1_REG3_REG_7__SCAN_IN ; P1_U5406
g2794 nand P1_U3455 P1_U3377 ; P1_U5407
g2795 nand P1_U3449 P1_U5407 ; P1_U5408
g2796 nand P1_U5817 P1_U3449 P1_R1165_U87 ; P1_U5409
g2797 nand P1_U3450 P1_U3453 ; P1_U5410
g2798 nand P1_U3874 P1_U4013 ; P1_U5411
g2799 nand P1_U3370 P1_U3422 ; P1_U5412
g2800 nand P1_U4006 P1_U3363 P1_U3365 ; P1_U5413
g2801 nand P1_U4041 P1_U3425 ; P1_U5414
g2802 nand P1_U5413 P1_U3425 ; P1_U5415
g2803 not P1_U3436 ; P1_U5416
g2804 nand P1_U5416 P1_U4013 ; P1_U5417
g2805 nand P1_U3485 P1_U5417 ; P1_U5418
g2806 nand P1_U3021 P1_U3083 ; P1_U5419
g2807 nand P1_U3482 P1_U5417 ; P1_U5420
g2808 nand P1_U3021 P1_U3084 ; P1_U5421
g2809 nand P1_U3479 P1_U5417 ; P1_U5422
g2810 nand P1_U3021 P1_U3070 ; P1_U5423
g2811 nand P1_U3476 P1_U5417 ; P1_U5424
g2812 nand P1_U3021 P1_U3071 ; P1_U5425
g2813 nand P1_U3473 P1_U5417 ; P1_U5426
g2814 nand P1_U3021 P1_U3067 ; P1_U5427
g2815 nand P1_U3470 P1_U5417 ; P1_U5428
g2816 nand P1_U3021 P1_U3060 ; P1_U5429
g2817 nand P1_U3467 P1_U5417 ; P1_U5430
g2818 nand P1_U3021 P1_U3064 ; P1_U5431
g2819 nand P1_U4017 P1_U5417 ; P1_U5432
g2820 nand P1_U3021 P1_U3054 ; P1_U5433
g2821 nand P1_U4018 P1_U5417 ; P1_U5434
g2822 nand P1_U3021 P1_U3053 ; P1_U5435
g2823 nand P1_U4019 P1_U5417 ; P1_U5436
g2824 nand P1_U3021 P1_U3057 ; P1_U5437
g2825 nand P1_U4020 P1_U5417 ; P1_U5438
g2826 nand P1_U3021 P1_U3058 ; P1_U5439
g2827 nand P1_U4021 P1_U5417 ; P1_U5440
g2828 nand P1_U3021 P1_U3065 ; P1_U5441
g2829 nand P1_U4022 P1_U5417 ; P1_U5442
g2830 nand P1_U3021 P1_U3066 ; P1_U5443
g2831 nand P1_U4023 P1_U5417 ; P1_U5444
g2832 nand P1_U3021 P1_U3061 ; P1_U5445
g2833 nand P1_U4024 P1_U5417 ; P1_U5446
g2834 nand P1_U3021 P1_U3075 ; P1_U5447
g2835 nand P1_U4025 P1_U5417 ; P1_U5448
g2836 nand P1_U3021 P1_U3076 ; P1_U5449
g2837 nand P1_U3464 P1_U5417 ; P1_U5450
g2838 nand P1_U3021 P1_U3068 ; P1_U5451
g2839 nand P1_U3514 P1_U5417 ; P1_U5452
g2840 nand P1_U3021 P1_U3081 ; P1_U5453
g2841 nand P1_U3512 P1_U5417 ; P1_U5454
g2842 nand P1_U3021 P1_U3082 ; P1_U5455
g2843 nand P1_U3509 P1_U5417 ; P1_U5456
g2844 nand P1_U3021 P1_U3069 ; P1_U5457
g2845 nand P1_U3506 P1_U5417 ; P1_U5458
g2846 nand P1_U3021 P1_U3073 ; P1_U5459
g2847 nand P1_U3503 P1_U5417 ; P1_U5460
g2848 nand P1_U3021 P1_U3074 ; P1_U5461
g2849 nand P1_U3500 P1_U5417 ; P1_U5462
g2850 nand P1_U3021 P1_U3079 ; P1_U5463
g2851 nand P1_U3497 P1_U5417 ; P1_U5464
g2852 nand P1_U3021 P1_U3080 ; P1_U5465
g2853 nand P1_U3494 P1_U5417 ; P1_U5466
g2854 nand P1_U3021 P1_U3072 ; P1_U5467
g2855 nand P1_U3491 P1_U5417 ; P1_U5468
g2856 nand P1_U3021 P1_U3063 ; P1_U5469
g2857 nand P1_U3488 P1_U5417 ; P1_U5470
g2858 nand P1_U3021 P1_U3062 ; P1_U5471
g2859 nand P1_U3461 P1_U5417 ; P1_U5472
g2860 nand P1_U3021 P1_U3078 ; P1_U5473
g2861 nand P1_U3456 P1_U5417 ; P1_U5474
g2862 nand P1_U3021 P1_U3077 ; P1_U5475
g2863 nand P1_U4145 P1_REG1_REG_0__SCAN_IN ; P1_U5476
g2864 nand P1_U3021 P1_U3485 ; P1_U5477
g2865 nand P1_U3436 P1_U3083 ; P1_U5478
g2866 nand P1_U3021 P1_U3482 ; P1_U5479
g2867 nand P1_U3436 P1_U3084 ; P1_U5480
g2868 nand P1_U3021 P1_U3479 ; P1_U5481
g2869 nand P1_U3436 P1_U3070 ; P1_U5482
g2870 nand P1_U3021 P1_U3476 ; P1_U5483
g2871 nand P1_U3436 P1_U3071 ; P1_U5484
g2872 nand P1_U3021 P1_U3473 ; P1_U5485
g2873 nand P1_U3436 P1_U3067 ; P1_U5486
g2874 nand P1_U3021 P1_U3470 ; P1_U5487
g2875 nand P1_U3436 P1_U3060 ; P1_U5488
g2876 nand P1_U3021 P1_U3467 ; P1_U5489
g2877 nand P1_U3436 P1_U3064 ; P1_U5490
g2878 nand P1_U3021 P1_U4017 ; P1_U5491
g2879 nand P1_U3436 P1_U3054 ; P1_U5492
g2880 nand P1_U3021 P1_U4018 ; P1_U5493
g2881 nand P1_U3436 P1_U3053 ; P1_U5494
g2882 nand P1_U3021 P1_U4019 ; P1_U5495
g2883 nand P1_U3436 P1_U3057 ; P1_U5496
g2884 nand P1_U3021 P1_U4020 ; P1_U5497
g2885 nand P1_U3436 P1_U3058 ; P1_U5498
g2886 nand P1_U3021 P1_U4021 ; P1_U5499
g2887 nand P1_U3436 P1_U3065 ; P1_U5500
g2888 nand P1_U3021 P1_U4022 ; P1_U5501
g2889 nand P1_U3436 P1_U3066 ; P1_U5502
g2890 nand P1_U3021 P1_U4023 ; P1_U5503
g2891 nand P1_U3436 P1_U3061 ; P1_U5504
g2892 nand P1_U3021 P1_U4024 ; P1_U5505
g2893 nand P1_U3436 P1_U3075 ; P1_U5506
g2894 nand P1_U3021 P1_U4025 ; P1_U5507
g2895 nand P1_U3436 P1_U3076 ; P1_U5508
g2896 nand P1_U3021 P1_U3464 ; P1_U5509
g2897 nand P1_U3436 P1_U3068 ; P1_U5510
g2898 nand P1_U3021 P1_U3514 ; P1_U5511
g2899 nand P1_U3436 P1_U3081 ; P1_U5512
g2900 nand P1_U3021 P1_U3512 ; P1_U5513
g2901 nand P1_U3436 P1_U3082 ; P1_U5514
g2902 nand P1_U3021 P1_U3509 ; P1_U5515
g2903 nand P1_U3436 P1_U3069 ; P1_U5516
g2904 nand P1_U3021 P1_U3506 ; P1_U5517
g2905 nand P1_U3436 P1_U3073 ; P1_U5518
g2906 nand P1_U3021 P1_U3503 ; P1_U5519
g2907 nand P1_U3436 P1_U3074 ; P1_U5520
g2908 nand P1_U3021 P1_U3500 ; P1_U5521
g2909 nand P1_U3436 P1_U3079 ; P1_U5522
g2910 nand P1_U3021 P1_U3497 ; P1_U5523
g2911 nand P1_U3436 P1_U3080 ; P1_U5524
g2912 nand P1_U3021 P1_U3494 ; P1_U5525
g2913 nand P1_U3436 P1_U3072 ; P1_U5526
g2914 nand P1_U3021 P1_U3491 ; P1_U5527
g2915 nand P1_U3436 P1_U3063 ; P1_U5528
g2916 nand P1_U3021 P1_U3488 ; P1_U5529
g2917 nand P1_U3436 P1_U3062 ; P1_U5530
g2918 nand P1_U3021 P1_U3461 ; P1_U5531
g2919 nand P1_U3436 P1_U3078 ; P1_U5532
g2920 nand P1_U3021 P1_U3456 ; P1_U5533
g2921 nand P1_U3436 P1_U3077 ; P1_U5534
g2922 nand P1_U4145 P1_U3454 ; P1_U5535
g2923 not P1_U3437 ; P1_U5536
g2924 not P1_U3438 ; P1_U5537
g2925 nand P1_U5799 P1_U3450 ; P1_U5538
g2926 nand P1_U3437 P1_U3439 ; P1_U5539
g2927 nand P1_U3051 P1_U5539 ; P1_U5540
g2928 nand P1_U3014 P1_U3444 ; P1_U5541
g2929 not P1_U3440 ; P1_U5542
g2930 nand P1_U3052 P1_U5542 ; P1_U5543
g2931 nand P1_U3083 P1_U3027 ; P1_U5544
g2932 nand P1_U3485 P1_U5543 ; P1_U5545
g2933 nand P1_U5540 P1_U3083 ; P1_U5546
g2934 nand P1_U3084 P1_U3027 ; P1_U5547
g2935 nand P1_U3482 P1_U5543 ; P1_U5548
g2936 nand P1_U5540 P1_U3084 ; P1_U5549
g2937 nand P1_U3070 P1_U3027 ; P1_U5550
g2938 nand P1_U3479 P1_U5543 ; P1_U5551
g2939 nand P1_U5540 P1_U3070 ; P1_U5552
g2940 nand P1_U3071 P1_U3027 ; P1_U5553
g2941 nand P1_U3476 P1_U5543 ; P1_U5554
g2942 nand P1_U5540 P1_U3071 ; P1_U5555
g2943 nand P1_U3067 P1_U3027 ; P1_U5556
g2944 nand P1_U3473 P1_U5543 ; P1_U5557
g2945 nand P1_U5540 P1_U3067 ; P1_U5558
g2946 nand P1_U3060 P1_U3027 ; P1_U5559
g2947 nand P1_U3470 P1_U5543 ; P1_U5560
g2948 nand P1_U5540 P1_U3060 ; P1_U5561
g2949 nand P1_R1309_U8 P1_U3027 ; P1_U5562
g2950 nand P1_U4026 P1_U5543 ; P1_U5563
g2951 nand P1_U5540 P1_U3056 ; P1_U5564
g2952 nand P1_R1309_U6 P1_U3027 ; P1_U5565
g2953 nand P1_U4027 P1_U5543 ; P1_U5566
g2954 nand P1_U5540 P1_U3059 ; P1_U5567
g2955 nand P1_U3064 P1_U3027 ; P1_U5568
g2956 nand P1_U3467 P1_U5543 ; P1_U5569
g2957 nand P1_U5540 P1_U3064 ; P1_U5570
g2958 nand P1_U3055 P1_U3027 ; P1_U5571
g2959 nand P1_U4028 P1_U5543 ; P1_U5572
g2960 nand P1_U5540 P1_U3055 ; P1_U5573
g2961 nand P1_U3054 P1_U3027 ; P1_U5574
g2962 nand P1_U4017 P1_U5543 ; P1_U5575
g2963 nand P1_U5540 P1_U3054 ; P1_U5576
g2964 nand P1_U3053 P1_U3027 ; P1_U5577
g2965 nand P1_U4018 P1_U5543 ; P1_U5578
g2966 nand P1_U5540 P1_U3053 ; P1_U5579
g2967 nand P1_U3057 P1_U3027 ; P1_U5580
g2968 nand P1_U4019 P1_U5543 ; P1_U5581
g2969 nand P1_U5540 P1_U3057 ; P1_U5582
g2970 nand P1_U3058 P1_U3027 ; P1_U5583
g2971 nand P1_U4020 P1_U5543 ; P1_U5584
g2972 nand P1_U5540 P1_U3058 ; P1_U5585
g2973 nand P1_U3065 P1_U3027 ; P1_U5586
g2974 nand P1_U4021 P1_U5543 ; P1_U5587
g2975 nand P1_U5540 P1_U3065 ; P1_U5588
g2976 nand P1_U3066 P1_U3027 ; P1_U5589
g2977 nand P1_U4022 P1_U5543 ; P1_U5590
g2978 nand P1_U5540 P1_U3066 ; P1_U5591
g2979 nand P1_U3061 P1_U3027 ; P1_U5592
g2980 nand P1_U4023 P1_U5543 ; P1_U5593
g2981 nand P1_U5540 P1_U3061 ; P1_U5594
g2982 nand P1_U3075 P1_U3027 ; P1_U5595
g2983 nand P1_U4024 P1_U5543 ; P1_U5596
g2984 nand P1_U5540 P1_U3075 ; P1_U5597
g2985 nand P1_U3076 P1_U3027 ; P1_U5598
g2986 nand P1_U4025 P1_U5543 ; P1_U5599
g2987 nand P1_U5540 P1_U3076 ; P1_U5600
g2988 nand P1_U3068 P1_U3027 ; P1_U5601
g2989 nand P1_U3464 P1_U5543 ; P1_U5602
g2990 nand P1_U5540 P1_U3068 ; P1_U5603
g2991 nand P1_U3081 P1_U3027 ; P1_U5604
g2992 nand P1_U3514 P1_U5543 ; P1_U5605
g2993 nand P1_U5540 P1_U3081 ; P1_U5606
g2994 nand P1_U3082 P1_U3027 ; P1_U5607
g2995 nand P1_U3512 P1_U5543 ; P1_U5608
g2996 nand P1_U5540 P1_U3082 ; P1_U5609
g2997 nand P1_U3069 P1_U3027 ; P1_U5610
g2998 nand P1_U3509 P1_U5543 ; P1_U5611
g2999 nand P1_U5540 P1_U3069 ; P1_U5612
g3000 nand P1_U3073 P1_U3027 ; P1_U5613
g3001 nand P1_U3506 P1_U5543 ; P1_U5614
g3002 nand P1_U5540 P1_U3073 ; P1_U5615
g3003 nand P1_U3074 P1_U3027 ; P1_U5616
g3004 nand P1_U3503 P1_U5543 ; P1_U5617
g3005 nand P1_U5540 P1_U3074 ; P1_U5618
g3006 nand P1_U3079 P1_U3027 ; P1_U5619
g3007 nand P1_U3500 P1_U5543 ; P1_U5620
g3008 nand P1_U5540 P1_U3079 ; P1_U5621
g3009 nand P1_U3080 P1_U3027 ; P1_U5622
g3010 nand P1_U3497 P1_U5543 ; P1_U5623
g3011 nand P1_U5540 P1_U3080 ; P1_U5624
g3012 nand P1_U3072 P1_U3027 ; P1_U5625
g3013 nand P1_U3494 P1_U5543 ; P1_U5626
g3014 nand P1_U5540 P1_U3072 ; P1_U5627
g3015 nand P1_U3063 P1_U3027 ; P1_U5628
g3016 nand P1_U3491 P1_U5543 ; P1_U5629
g3017 nand P1_U5540 P1_U3063 ; P1_U5630
g3018 nand P1_U3062 P1_U3027 ; P1_U5631
g3019 nand P1_U3488 P1_U5543 ; P1_U5632
g3020 nand P1_U5540 P1_U3062 ; P1_U5633
g3021 nand P1_U3078 P1_U3027 ; P1_U5634
g3022 nand P1_U3461 P1_U5543 ; P1_U5635
g3023 nand P1_U5540 P1_U3078 ; P1_U5636
g3024 nand P1_U3077 P1_U3027 ; P1_U5637
g3025 nand P1_U3456 P1_U5543 ; P1_U5638
g3026 nand P1_U5540 P1_U3077 ; P1_U5639
g3027 nand P1_U3440 P1_U3439 ; P1_U5640
g3028 nand P1_U3052 P1_U5640 ; P1_U5641
g3029 nand P1_U3028 P1_U3083 ; P1_U5642
g3030 nand P1_U3485 P1_U3438 ; P1_U5643
g3031 nand P1_U5641 P1_U3083 ; P1_U5644
g3032 nand P1_U5786 P1_U3084 ; P1_U5645
g3033 nand P1_U3028 P1_U3084 ; P1_U5646
g3034 nand P1_U3482 P1_U3438 ; P1_U5647
g3035 nand P1_U5641 P1_U3084 ; P1_U5648
g3036 nand P1_U5786 P1_U3070 ; P1_U5649
g3037 nand P1_U3028 P1_U3070 ; P1_U5650
g3038 nand P1_U3479 P1_U3438 ; P1_U5651
g3039 nand P1_U5641 P1_U3070 ; P1_U5652
g3040 nand P1_U5786 P1_U3071 ; P1_U5653
g3041 nand P1_U3028 P1_U3071 ; P1_U5654
g3042 nand P1_U3476 P1_U3438 ; P1_U5655
g3043 nand P1_U5641 P1_U3071 ; P1_U5656
g3044 nand P1_U5786 P1_U3067 ; P1_U5657
g3045 nand P1_U3028 P1_U3067 ; P1_U5658
g3046 nand P1_U3473 P1_U3438 ; P1_U5659
g3047 nand P1_U5641 P1_U3067 ; P1_U5660
g3048 nand P1_U5786 P1_U3060 ; P1_U5661
g3049 nand P1_U3028 P1_U3060 ; P1_U5662
g3050 nand P1_U3470 P1_U3438 ; P1_U5663
g3051 nand P1_U5641 P1_U3060 ; P1_U5664
g3052 nand P1_U5786 P1_U3064 ; P1_U5665
g3053 nand P1_U3028 P1_R1309_U8 ; P1_U5666
g3054 nand P1_U4026 P1_U3438 ; P1_U5667
g3055 nand P1_U5641 P1_U3056 ; P1_U5668
g3056 nand P1_U3028 P1_R1309_U6 ; P1_U5669
g3057 nand P1_U4027 P1_U3438 ; P1_U5670
g3058 nand P1_U5641 P1_U3059 ; P1_U5671
g3059 nand P1_U3028 P1_U3064 ; P1_U5672
g3060 nand P1_U3467 P1_U3438 ; P1_U5673
g3061 nand P1_U5641 P1_U3064 ; P1_U5674
g3062 nand P1_U5786 P1_U3068 ; P1_U5675
g3063 nand P1_U3028 P1_U3055 ; P1_U5676
g3064 nand P1_U4028 P1_U3438 ; P1_U5677
g3065 nand P1_U5641 P1_U3055 ; P1_U5678
g3066 nand P1_U5786 P1_U3054 ; P1_U5679
g3067 nand P1_U3028 P1_U3054 ; P1_U5680
g3068 nand P1_U4017 P1_U3438 ; P1_U5681
g3069 nand P1_U5641 P1_U3054 ; P1_U5682
g3070 nand P1_U5786 P1_U3053 ; P1_U5683
g3071 nand P1_U3028 P1_U3053 ; P1_U5684
g3072 nand P1_U4018 P1_U3438 ; P1_U5685
g3073 nand P1_U5641 P1_U3053 ; P1_U5686
g3074 nand P1_U5786 P1_U3057 ; P1_U5687
g3075 nand P1_U3028 P1_U3057 ; P1_U5688
g3076 nand P1_U4019 P1_U3438 ; P1_U5689
g3077 nand P1_U5641 P1_U3057 ; P1_U5690
g3078 nand P1_U5786 P1_U3058 ; P1_U5691
g3079 nand P1_U3028 P1_U3058 ; P1_U5692
g3080 nand P1_U4020 P1_U3438 ; P1_U5693
g3081 nand P1_U5641 P1_U3058 ; P1_U5694
g3082 nand P1_U5786 P1_U3065 ; P1_U5695
g3083 nand P1_U3028 P1_U3065 ; P1_U5696
g3084 nand P1_U4021 P1_U3438 ; P1_U5697
g3085 nand P1_U5641 P1_U3065 ; P1_U5698
g3086 nand P1_U5786 P1_U3066 ; P1_U5699
g3087 nand P1_U3028 P1_U3066 ; P1_U5700
g3088 nand P1_U4022 P1_U3438 ; P1_U5701
g3089 nand P1_U5641 P1_U3066 ; P1_U5702
g3090 nand P1_U5786 P1_U3061 ; P1_U5703
g3091 nand P1_U3028 P1_U3061 ; P1_U5704
g3092 nand P1_U4023 P1_U3438 ; P1_U5705
g3093 nand P1_U5641 P1_U3061 ; P1_U5706
g3094 nand P1_U5786 P1_U3075 ; P1_U5707
g3095 nand P1_U3028 P1_U3075 ; P1_U5708
g3096 nand P1_U4024 P1_U3438 ; P1_U5709
g3097 nand P1_U5641 P1_U3075 ; P1_U5710
g3098 nand P1_U5786 P1_U3076 ; P1_U5711
g3099 nand P1_U3028 P1_U3076 ; P1_U5712
g3100 nand P1_U4025 P1_U3438 ; P1_U5713
g3101 nand P1_U5641 P1_U3076 ; P1_U5714
g3102 nand P1_U5786 P1_U3081 ; P1_U5715
g3103 nand P1_U3028 P1_U3068 ; P1_U5716
g3104 nand P1_U3464 P1_U3438 ; P1_U5717
g3105 nand P1_U5641 P1_U3068 ; P1_U5718
g3106 nand P1_U5786 P1_U3078 ; P1_U5719
g3107 nand P1_U3028 P1_U3081 ; P1_U5720
g3108 nand P1_U3514 P1_U3438 ; P1_U5721
g3109 nand P1_U5641 P1_U3081 ; P1_U5722
g3110 nand P1_U5786 P1_U3082 ; P1_U5723
g3111 nand P1_U3028 P1_U3082 ; P1_U5724
g3112 nand P1_U3512 P1_U3438 ; P1_U5725
g3113 nand P1_U5641 P1_U3082 ; P1_U5726
g3114 nand P1_U5786 P1_U3069 ; P1_U5727
g3115 nand P1_U3028 P1_U3069 ; P1_U5728
g3116 nand P1_U3509 P1_U3438 ; P1_U5729
g3117 nand P1_U5641 P1_U3069 ; P1_U5730
g3118 nand P1_U5786 P1_U3073 ; P1_U5731
g3119 nand P1_U3028 P1_U3073 ; P1_U5732
g3120 nand P1_U3506 P1_U3438 ; P1_U5733
g3121 nand P1_U5641 P1_U3073 ; P1_U5734
g3122 nand P1_U5786 P1_U3074 ; P1_U5735
g3123 nand P1_U3028 P1_U3074 ; P1_U5736
g3124 nand P1_U3503 P1_U3438 ; P1_U5737
g3125 nand P1_U5641 P1_U3074 ; P1_U5738
g3126 nand P1_U5786 P1_U3079 ; P1_U5739
g3127 nand P1_U3028 P1_U3079 ; P1_U5740
g3128 nand P1_U3500 P1_U3438 ; P1_U5741
g3129 nand P1_U5641 P1_U3079 ; P1_U5742
g3130 nand P1_U5786 P1_U3080 ; P1_U5743
g3131 nand P1_U3028 P1_U3080 ; P1_U5744
g3132 nand P1_U3497 P1_U3438 ; P1_U5745
g3133 nand P1_U5641 P1_U3080 ; P1_U5746
g3134 nand P1_U5786 P1_U3072 ; P1_U5747
g3135 nand P1_U3028 P1_U3072 ; P1_U5748
g3136 nand P1_U3494 P1_U3438 ; P1_U5749
g3137 nand P1_U5641 P1_U3072 ; P1_U5750
g3138 nand P1_U5786 P1_U3063 ; P1_U5751
g3139 nand P1_U3028 P1_U3063 ; P1_U5752
g3140 nand P1_U3491 P1_U3438 ; P1_U5753
g3141 nand P1_U5641 P1_U3063 ; P1_U5754
g3142 nand P1_U5786 P1_U3062 ; P1_U5755
g3143 nand P1_U3028 P1_U3062 ; P1_U5756
g3144 nand P1_U3488 P1_U3438 ; P1_U5757
g3145 nand P1_U5641 P1_U3062 ; P1_U5758
g3146 nand P1_U5786 P1_U3083 ; P1_U5759
g3147 nand P1_U3028 P1_U3078 ; P1_U5760
g3148 nand P1_U3461 P1_U3438 ; P1_U5761
g3149 nand P1_U5641 P1_U3078 ; P1_U5762
g3150 nand P1_U5786 P1_U3077 ; P1_U5763
g3151 nand P1_U3028 P1_U3077 ; P1_U5764
g3152 nand P1_U3456 P1_U3438 ; P1_U5765
g3153 nand P1_U5641 P1_U3077 ; P1_U5766
g3154 nand P1_U4038 P1_U3434 ; P1_U5767
g3155 nand P1_U4015 P1_U4038 ; P1_U5768
g3156 nand P1_U3050 P1_U5767 ; P1_U5769
g3157 nand P1_U5768 P1_U4039 ; P1_U5770
g3158 nand P1_U5775 P1_U5781 ; P1_U5771
g3159 nand P1_R1375_U9 P1_U5131 ; P1_U5772
g3160 nand P1_U3952 P1_IR_REG_24__SCAN_IN ; P1_U5773
g3161 nand P1_SUB_88_U17 P1_IR_REG_31__SCAN_IN ; P1_U5774
g3162 not P1_U3441 ; P1_U5775
g3163 nand P1_U3952 P1_IR_REG_25__SCAN_IN ; P1_U5776
g3164 nand P1_SUB_88_U170 P1_IR_REG_31__SCAN_IN ; P1_U5777
g3165 not P1_U3442 ; P1_U5778
g3166 nand P1_U3952 P1_IR_REG_26__SCAN_IN ; P1_U5779
g3167 nand P1_SUB_88_U18 P1_IR_REG_31__SCAN_IN ; P1_U5780
g3168 not P1_U3443 ; P1_U5781
g3169 nand P1_U3441 P1_U3359 ; P1_U5782
g3170 nand P1_U4046 P1_U5775 P1_B_REG_SCAN_IN ; P1_U5783
g3171 nand P1_U3952 P1_IR_REG_23__SCAN_IN ; P1_U5784
g3172 nand P1_SUB_88_U16 P1_IR_REG_31__SCAN_IN ; P1_U5785
g3173 not P1_U3444 ; P1_U5786
g3174 nand P1_U3953 P1_D_REG_0__SCAN_IN ; P1_U5787
g3175 nand P1_U4034 P1_U4146 ; P1_U5788
g3176 nand P1_U3953 P1_D_REG_1__SCAN_IN ; P1_U5789
g3177 nand P1_U4034 P1_U4147 ; P1_U5790
g3178 nand P1_U3952 P1_IR_REG_22__SCAN_IN ; P1_U5791
g3179 nand P1_SUB_88_U15 P1_IR_REG_31__SCAN_IN ; P1_U5792
g3180 not P1_U3451 ; P1_U5793
g3181 nand P1_U3952 P1_IR_REG_19__SCAN_IN ; P1_U5794
g3182 nand P1_SUB_88_U13 P1_IR_REG_31__SCAN_IN ; P1_U5795
g3183 not P1_U3452 ; P1_U5796
g3184 nand P1_U3952 P1_IR_REG_20__SCAN_IN ; P1_U5797
g3185 nand P1_SUB_88_U14 P1_IR_REG_31__SCAN_IN ; P1_U5798
g3186 not P1_U3453 ; P1_U5799
g3187 nand P1_U3952 P1_IR_REG_21__SCAN_IN ; P1_U5800
g3188 nand P1_SUB_88_U173 P1_IR_REG_31__SCAN_IN ; P1_U5801
g3189 not P1_U3450 ; P1_U5802
g3190 nand P1_U3952 P1_IR_REG_30__SCAN_IN ; P1_U5803
g3191 nand P1_SUB_88_U165 P1_IR_REG_31__SCAN_IN ; P1_U5804
g3192 not P1_U3447 ; P1_U5805
g3193 nand P1_U3952 P1_IR_REG_29__SCAN_IN ; P1_U5806
g3194 nand P1_SUB_88_U20 P1_IR_REG_31__SCAN_IN ; P1_U5807
g3195 not P1_U3448 ; P1_U5808
g3196 nand P1_U3952 P1_IR_REG_28__SCAN_IN ; P1_U5809
g3197 nand P1_SUB_88_U19 P1_IR_REG_31__SCAN_IN ; P1_U5810
g3198 not P1_U3449 ; P1_U5811
g3199 nand P1_U3952 P1_IR_REG_0__SCAN_IN ; P1_U5812
g3200 nand P1_IR_REG_0__SCAN_IN P1_IR_REG_31__SCAN_IN ; P1_U5813
g3201 not P1_U3454 ; P1_U5814
g3202 nand P1_U3952 P1_IR_REG_27__SCAN_IN ; P1_U5815
g3203 nand P1_SUB_88_U42 P1_IR_REG_31__SCAN_IN ; P1_U5816
g3204 not P1_U3455 ; P1_U5817
g3205 nand U125 P1_U3954 ; P1_U5818
g3206 nand P1_U4014 P1_U3454 ; P1_U5819
g3207 not P1_U3456 ; P1_U5820
g3208 nand P1_U3451 P1_U5802 ; P1_U5821
g3209 nand P1_U5793 P1_U4178 ; P1_U5822
g3210 nand P1_U4144 P1_D_REG_1__SCAN_IN ; P1_U5823
g3211 nand P1_U4147 P1_U3360 ; P1_U5824
g3212 not P1_U3458 ; P1_U5825
g3213 nand P1_U5771 P1_U3360 ; P1_U5826
g3214 nand P1_U4144 P1_D_REG_0__SCAN_IN ; P1_U5827
g3215 not P1_U3457 ; P1_U5828
g3216 nand P1_U3955 P1_REG0_REG_0__SCAN_IN ; P1_U5829
g3217 nand P1_U4033 P1_U4198 ; P1_U5830
g3218 nand P1_U3952 P1_IR_REG_1__SCAN_IN ; P1_U5831
g3219 nand P1_SUB_88_U40 P1_IR_REG_31__SCAN_IN ; P1_U5832
g3220 nand U114 P1_U3954 ; P1_U5833
g3221 nand P1_U3460 P1_U4014 ; P1_U5834
g3222 not P1_U3461 ; P1_U5835
g3223 nand P1_U3955 P1_REG0_REG_1__SCAN_IN ; P1_U5836
g3224 nand P1_U4033 P1_U4222 ; P1_U5837
g3225 nand P1_U3952 P1_IR_REG_2__SCAN_IN ; P1_U5838
g3226 nand P1_SUB_88_U21 P1_IR_REG_31__SCAN_IN ; P1_U5839
g3227 nand U103 P1_U3954 ; P1_U5840
g3228 nand P1_U3463 P1_U4014 ; P1_U5841
g3229 not P1_U3464 ; P1_U5842
g3230 nand P1_U3955 P1_REG0_REG_2__SCAN_IN ; P1_U5843
g3231 nand P1_U4033 P1_U4241 ; P1_U5844
g3232 nand P1_U3952 P1_IR_REG_3__SCAN_IN ; P1_U5845
g3233 nand P1_SUB_88_U22 P1_IR_REG_31__SCAN_IN ; P1_U5846
g3234 nand U100 P1_U3954 ; P1_U5847
g3235 nand P1_U3466 P1_U4014 ; P1_U5848
g3236 not P1_U3467 ; P1_U5849
g3237 nand P1_U3955 P1_REG0_REG_3__SCAN_IN ; P1_U5850
g3238 nand P1_U4033 P1_U4260 ; P1_U5851
g3239 nand P1_U3952 P1_IR_REG_4__SCAN_IN ; P1_U5852
g3240 nand P1_SUB_88_U23 P1_IR_REG_31__SCAN_IN ; P1_U5853
g3241 nand U99 P1_U3954 ; P1_U5854
g3242 nand P1_U3469 P1_U4014 ; P1_U5855
g3243 not P1_U3470 ; P1_U5856
g3244 nand P1_U3955 P1_REG0_REG_4__SCAN_IN ; P1_U5857
g3245 nand P1_U4033 P1_U4279 ; P1_U5858
g3246 nand P1_U3952 P1_IR_REG_5__SCAN_IN ; P1_U5859
g3247 nand P1_SUB_88_U162 P1_IR_REG_31__SCAN_IN ; P1_U5860
g3248 nand U98 P1_U3954 ; P1_U5861
g3249 nand P1_U3472 P1_U4014 ; P1_U5862
g3250 not P1_U3473 ; P1_U5863
g3251 nand P1_U3955 P1_REG0_REG_5__SCAN_IN ; P1_U5864
g3252 nand P1_U4033 P1_U4298 ; P1_U5865
g3253 nand P1_U3952 P1_IR_REG_6__SCAN_IN ; P1_U5866
g3254 nand P1_SUB_88_U24 P1_IR_REG_31__SCAN_IN ; P1_U5867
g3255 nand U97 P1_U3954 ; P1_U5868
g3256 nand P1_U3475 P1_U4014 ; P1_U5869
g3257 not P1_U3476 ; P1_U5870
g3258 nand P1_U3955 P1_REG0_REG_6__SCAN_IN ; P1_U5871
g3259 nand P1_U4033 P1_U4317 ; P1_U5872
g3260 nand P1_U3952 P1_IR_REG_7__SCAN_IN ; P1_U5873
g3261 nand P1_SUB_88_U25 P1_IR_REG_31__SCAN_IN ; P1_U5874
g3262 nand U96 P1_U3954 ; P1_U5875
g3263 nand P1_U3478 P1_U4014 ; P1_U5876
g3264 not P1_U3479 ; P1_U5877
g3265 nand P1_U3955 P1_REG0_REG_7__SCAN_IN ; P1_U5878
g3266 nand P1_U4033 P1_U4336 ; P1_U5879
g3267 nand P1_U3952 P1_IR_REG_8__SCAN_IN ; P1_U5880
g3268 nand P1_SUB_88_U26 P1_IR_REG_31__SCAN_IN ; P1_U5881
g3269 nand U95 P1_U3954 ; P1_U5882
g3270 nand P1_U3481 P1_U4014 ; P1_U5883
g3271 not P1_U3482 ; P1_U5884
g3272 nand P1_U3955 P1_REG0_REG_8__SCAN_IN ; P1_U5885
g3273 nand P1_U4033 P1_U4355 ; P1_U5886
g3274 nand P1_U3952 P1_IR_REG_9__SCAN_IN ; P1_U5887
g3275 nand P1_SUB_88_U160 P1_IR_REG_31__SCAN_IN ; P1_U5888
g3276 nand U94 P1_U3954 ; P1_U5889
g3277 nand P1_U3484 P1_U4014 ; P1_U5890
g3278 not P1_U3485 ; P1_U5891
g3279 nand P1_U3955 P1_REG0_REG_9__SCAN_IN ; P1_U5892
g3280 nand P1_U4033 P1_U4374 ; P1_U5893
g3281 nand P1_U3952 P1_IR_REG_10__SCAN_IN ; P1_U5894
g3282 nand P1_SUB_88_U6 P1_IR_REG_31__SCAN_IN ; P1_U5895
g3283 nand U124 P1_U3954 ; P1_U5896
g3284 nand P1_U3487 P1_U4014 ; P1_U5897
g3285 not P1_U3488 ; P1_U5898
g3286 nand P1_U3955 P1_REG0_REG_10__SCAN_IN ; P1_U5899
g3287 nand P1_U4033 P1_U4393 ; P1_U5900
g3288 nand P1_U3952 P1_IR_REG_11__SCAN_IN ; P1_U5901
g3289 nand P1_SUB_88_U7 P1_IR_REG_31__SCAN_IN ; P1_U5902
g3290 nand U123 P1_U3954 ; P1_U5903
g3291 nand P1_U3490 P1_U4014 ; P1_U5904
g3292 not P1_U3491 ; P1_U5905
g3293 nand P1_U3955 P1_REG0_REG_11__SCAN_IN ; P1_U5906
g3294 nand P1_U4033 P1_U4412 ; P1_U5907
g3295 nand P1_U3952 P1_IR_REG_12__SCAN_IN ; P1_U5908
g3296 nand P1_SUB_88_U8 P1_IR_REG_31__SCAN_IN ; P1_U5909
g3297 nand U122 P1_U3954 ; P1_U5910
g3298 nand P1_U3493 P1_U4014 ; P1_U5911
g3299 not P1_U3494 ; P1_U5912
g3300 nand P1_U3955 P1_REG0_REG_12__SCAN_IN ; P1_U5913
g3301 nand P1_U4033 P1_U4431 ; P1_U5914
g3302 nand P1_U3952 P1_IR_REG_13__SCAN_IN ; P1_U5915
g3303 nand P1_SUB_88_U179 P1_IR_REG_31__SCAN_IN ; P1_U5916
g3304 nand U121 P1_U3954 ; P1_U5917
g3305 nand P1_U3496 P1_U4014 ; P1_U5918
g3306 not P1_U3497 ; P1_U5919
g3307 nand P1_U3955 P1_REG0_REG_13__SCAN_IN ; P1_U5920
g3308 nand P1_U4033 P1_U4450 ; P1_U5921
g3309 nand P1_U3952 P1_IR_REG_14__SCAN_IN ; P1_U5922
g3310 nand P1_SUB_88_U9 P1_IR_REG_31__SCAN_IN ; P1_U5923
g3311 nand U120 P1_U3954 ; P1_U5924
g3312 nand P1_U3499 P1_U4014 ; P1_U5925
g3313 not P1_U3500 ; P1_U5926
g3314 nand P1_U3955 P1_REG0_REG_14__SCAN_IN ; P1_U5927
g3315 nand P1_U4033 P1_U4469 ; P1_U5928
g3316 nand P1_U3952 P1_IR_REG_15__SCAN_IN ; P1_U5929
g3317 nand P1_SUB_88_U10 P1_IR_REG_31__SCAN_IN ; P1_U5930
g3318 nand U119 P1_U3954 ; P1_U5931
g3319 nand P1_U3502 P1_U4014 ; P1_U5932
g3320 not P1_U3503 ; P1_U5933
g3321 nand P1_U3955 P1_REG0_REG_15__SCAN_IN ; P1_U5934
g3322 nand P1_U4033 P1_U4488 ; P1_U5935
g3323 nand P1_U3952 P1_IR_REG_16__SCAN_IN ; P1_U5936
g3324 nand P1_SUB_88_U11 P1_IR_REG_31__SCAN_IN ; P1_U5937
g3325 nand U118 P1_U3954 ; P1_U5938
g3326 nand P1_U3505 P1_U4014 ; P1_U5939
g3327 not P1_U3506 ; P1_U5940
g3328 nand P1_U3955 P1_REG0_REG_16__SCAN_IN ; P1_U5941
g3329 nand P1_U4033 P1_U4507 ; P1_U5942
g3330 nand P1_U3952 P1_IR_REG_17__SCAN_IN ; P1_U5943
g3331 nand P1_SUB_88_U177 P1_IR_REG_31__SCAN_IN ; P1_U5944
g3332 nand U117 P1_U3954 ; P1_U5945
g3333 nand P1_U3508 P1_U4014 ; P1_U5946
g3334 not P1_U3509 ; P1_U5947
g3335 nand P1_U3955 P1_REG0_REG_17__SCAN_IN ; P1_U5948
g3336 nand P1_U4033 P1_U4526 ; P1_U5949
g3337 nand P1_U3952 P1_IR_REG_18__SCAN_IN ; P1_U5950
g3338 nand P1_SUB_88_U12 P1_IR_REG_31__SCAN_IN ; P1_U5951
g3339 nand U116 P1_U3954 ; P1_U5952
g3340 nand P1_U3511 P1_U4014 ; P1_U5953
g3341 not P1_U3512 ; P1_U5954
g3342 nand P1_U3955 P1_REG0_REG_18__SCAN_IN ; P1_U5955
g3343 nand P1_U4033 P1_U4545 ; P1_U5956
g3344 nand U115 P1_U3954 ; P1_U5957
g3345 nand P1_U4014 P1_U3452 ; P1_U5958
g3346 not P1_U3514 ; P1_U5959
g3347 nand P1_U3955 P1_REG0_REG_19__SCAN_IN ; P1_U5960
g3348 nand P1_U4033 P1_U4564 ; P1_U5961
g3349 nand P1_U3955 P1_REG0_REG_20__SCAN_IN ; P1_U5962
g3350 nand P1_U4033 P1_U4583 ; P1_U5963
g3351 nand P1_U3955 P1_REG0_REG_21__SCAN_IN ; P1_U5964
g3352 nand P1_U4033 P1_U4602 ; P1_U5965
g3353 nand P1_U3955 P1_REG0_REG_22__SCAN_IN ; P1_U5966
g3354 nand P1_U4033 P1_U4621 ; P1_U5967
g3355 nand P1_U3955 P1_REG0_REG_23__SCAN_IN ; P1_U5968
g3356 nand P1_U4033 P1_U4640 ; P1_U5969
g3357 nand P1_U3955 P1_REG0_REG_24__SCAN_IN ; P1_U5970
g3358 nand P1_U4033 P1_U4659 ; P1_U5971
g3359 nand P1_U3955 P1_REG0_REG_25__SCAN_IN ; P1_U5972
g3360 nand P1_U4033 P1_U4678 ; P1_U5973
g3361 nand P1_U3955 P1_REG0_REG_26__SCAN_IN ; P1_U5974
g3362 nand P1_U4033 P1_U4697 ; P1_U5975
g3363 nand P1_U3955 P1_REG0_REG_27__SCAN_IN ; P1_U5976
g3364 nand P1_U4033 P1_U4716 ; P1_U5977
g3365 nand P1_U3955 P1_REG0_REG_28__SCAN_IN ; P1_U5978
g3366 nand P1_U4033 P1_U4735 ; P1_U5979
g3367 nand P1_U3955 P1_REG0_REG_29__SCAN_IN ; P1_U5980
g3368 nand P1_U4033 P1_U4755 ; P1_U5981
g3369 nand P1_U3955 P1_REG0_REG_30__SCAN_IN ; P1_U5982
g3370 nand P1_U4033 P1_U4762 ; P1_U5983
g3371 nand P1_U3955 P1_REG0_REG_31__SCAN_IN ; P1_U5984
g3372 nand P1_U4033 P1_U4765 ; P1_U5985
g3373 nand P1_U3956 P1_REG1_REG_0__SCAN_IN ; P1_U5986
g3374 nand P1_U4032 P1_U4198 ; P1_U5987
g3375 nand P1_U3956 P1_REG1_REG_1__SCAN_IN ; P1_U5988
g3376 nand P1_U4032 P1_U4222 ; P1_U5989
g3377 nand P1_U3956 P1_REG1_REG_2__SCAN_IN ; P1_U5990
g3378 nand P1_U4032 P1_U4241 ; P1_U5991
g3379 nand P1_U3956 P1_REG1_REG_3__SCAN_IN ; P1_U5992
g3380 nand P1_U4032 P1_U4260 ; P1_U5993
g3381 nand P1_U3956 P1_REG1_REG_4__SCAN_IN ; P1_U5994
g3382 nand P1_U4032 P1_U4279 ; P1_U5995
g3383 nand P1_U3956 P1_REG1_REG_5__SCAN_IN ; P1_U5996
g3384 nand P1_U4032 P1_U4298 ; P1_U5997
g3385 nand P1_U3956 P1_REG1_REG_6__SCAN_IN ; P1_U5998
g3386 nand P1_U4032 P1_U4317 ; P1_U5999
g3387 nand P1_U3956 P1_REG1_REG_7__SCAN_IN ; P1_U6000
g3388 nand P1_U4032 P1_U4336 ; P1_U6001
g3389 nand P1_U3956 P1_REG1_REG_8__SCAN_IN ; P1_U6002
g3390 nand P1_U4032 P1_U4355 ; P1_U6003
g3391 nand P1_U3956 P1_REG1_REG_9__SCAN_IN ; P1_U6004
g3392 nand P1_U4032 P1_U4374 ; P1_U6005
g3393 nand P1_U3956 P1_REG1_REG_10__SCAN_IN ; P1_U6006
g3394 nand P1_U4032 P1_U4393 ; P1_U6007
g3395 nand P1_U3956 P1_REG1_REG_11__SCAN_IN ; P1_U6008
g3396 nand P1_U4032 P1_U4412 ; P1_U6009
g3397 nand P1_U3956 P1_REG1_REG_12__SCAN_IN ; P1_U6010
g3398 nand P1_U4032 P1_U4431 ; P1_U6011
g3399 nand P1_U3956 P1_REG1_REG_13__SCAN_IN ; P1_U6012
g3400 nand P1_U4032 P1_U4450 ; P1_U6013
g3401 nand P1_U3956 P1_REG1_REG_14__SCAN_IN ; P1_U6014
g3402 nand P1_U4032 P1_U4469 ; P1_U6015
g3403 nand P1_U3956 P1_REG1_REG_15__SCAN_IN ; P1_U6016
g3404 nand P1_U4032 P1_U4488 ; P1_U6017
g3405 nand P1_U3956 P1_REG1_REG_16__SCAN_IN ; P1_U6018
g3406 nand P1_U4032 P1_U4507 ; P1_U6019
g3407 nand P1_U3956 P1_REG1_REG_17__SCAN_IN ; P1_U6020
g3408 nand P1_U4032 P1_U4526 ; P1_U6021
g3409 nand P1_U3956 P1_REG1_REG_18__SCAN_IN ; P1_U6022
g3410 nand P1_U4032 P1_U4545 ; P1_U6023
g3411 nand P1_U3956 P1_REG1_REG_19__SCAN_IN ; P1_U6024
g3412 nand P1_U4032 P1_U4564 ; P1_U6025
g3413 nand P1_U3956 P1_REG1_REG_20__SCAN_IN ; P1_U6026
g3414 nand P1_U4032 P1_U4583 ; P1_U6027
g3415 nand P1_U3956 P1_REG1_REG_21__SCAN_IN ; P1_U6028
g3416 nand P1_U4032 P1_U4602 ; P1_U6029
g3417 nand P1_U3956 P1_REG1_REG_22__SCAN_IN ; P1_U6030
g3418 nand P1_U4032 P1_U4621 ; P1_U6031
g3419 nand P1_U3956 P1_REG1_REG_23__SCAN_IN ; P1_U6032
g3420 nand P1_U4032 P1_U4640 ; P1_U6033
g3421 nand P1_U3956 P1_REG1_REG_24__SCAN_IN ; P1_U6034
g3422 nand P1_U4032 P1_U4659 ; P1_U6035
g3423 nand P1_U3956 P1_REG1_REG_25__SCAN_IN ; P1_U6036
g3424 nand P1_U4032 P1_U4678 ; P1_U6037
g3425 nand P1_U3956 P1_REG1_REG_26__SCAN_IN ; P1_U6038
g3426 nand P1_U4032 P1_U4697 ; P1_U6039
g3427 nand P1_U3956 P1_REG1_REG_27__SCAN_IN ; P1_U6040
g3428 nand P1_U4032 P1_U4716 ; P1_U6041
g3429 nand P1_U3956 P1_REG1_REG_28__SCAN_IN ; P1_U6042
g3430 nand P1_U4032 P1_U4735 ; P1_U6043
g3431 nand P1_U3956 P1_REG1_REG_29__SCAN_IN ; P1_U6044
g3432 nand P1_U4032 P1_U4755 ; P1_U6045
g3433 nand P1_U3956 P1_REG1_REG_30__SCAN_IN ; P1_U6046
g3434 nand P1_U4032 P1_U4762 ; P1_U6047
g3435 nand P1_U3956 P1_REG1_REG_31__SCAN_IN ; P1_U6048
g3436 nand P1_U4032 P1_U4765 ; P1_U6049
g3437 nand P1_U3420 P1_REG2_REG_0__SCAN_IN ; P1_U6050
g3438 nand P1_U4031 P1_U3376 ; P1_U6051
g3439 nand P1_U3420 P1_REG2_REG_1__SCAN_IN ; P1_U6052
g3440 nand P1_U4031 P1_U3378 ; P1_U6053
g3441 nand P1_U3420 P1_REG2_REG_2__SCAN_IN ; P1_U6054
g3442 nand P1_U4031 P1_U3379 ; P1_U6055
g3443 nand P1_U3420 P1_REG2_REG_3__SCAN_IN ; P1_U6056
g3444 nand P1_U4031 P1_U3380 ; P1_U6057
g3445 nand P1_U3420 P1_REG2_REG_4__SCAN_IN ; P1_U6058
g3446 nand P1_U4031 P1_U3381 ; P1_U6059
g3447 nand P1_U3420 P1_REG2_REG_5__SCAN_IN ; P1_U6060
g3448 nand P1_U4031 P1_U3382 ; P1_U6061
g3449 nand P1_U3420 P1_REG2_REG_6__SCAN_IN ; P1_U6062
g3450 nand P1_U4031 P1_U3383 ; P1_U6063
g3451 nand P1_U3420 P1_REG2_REG_7__SCAN_IN ; P1_U6064
g3452 nand P1_U4031 P1_U3384 ; P1_U6065
g3453 nand P1_U3420 P1_REG2_REG_8__SCAN_IN ; P1_U6066
g3454 nand P1_U4031 P1_U3385 ; P1_U6067
g3455 nand P1_U3420 P1_REG2_REG_9__SCAN_IN ; P1_U6068
g3456 nand P1_U4031 P1_U3386 ; P1_U6069
g3457 nand P1_U3420 P1_REG2_REG_10__SCAN_IN ; P1_U6070
g3458 nand P1_U4031 P1_U3387 ; P1_U6071
g3459 nand P1_U3420 P1_REG2_REG_11__SCAN_IN ; P1_U6072
g3460 nand P1_U4031 P1_U3388 ; P1_U6073
g3461 nand P1_U3420 P1_REG2_REG_12__SCAN_IN ; P1_U6074
g3462 nand P1_U4031 P1_U3389 ; P1_U6075
g3463 nand P1_U3420 P1_REG2_REG_13__SCAN_IN ; P1_U6076
g3464 nand P1_U4031 P1_U3390 ; P1_U6077
g3465 nand P1_U3420 P1_REG2_REG_14__SCAN_IN ; P1_U6078
g3466 nand P1_U4031 P1_U3391 ; P1_U6079
g3467 nand P1_U3420 P1_REG2_REG_15__SCAN_IN ; P1_U6080
g3468 nand P1_U4031 P1_U3392 ; P1_U6081
g3469 nand P1_U3420 P1_REG2_REG_16__SCAN_IN ; P1_U6082
g3470 nand P1_U4031 P1_U3393 ; P1_U6083
g3471 nand P1_U3420 P1_REG2_REG_17__SCAN_IN ; P1_U6084
g3472 nand P1_U4031 P1_U3394 ; P1_U6085
g3473 nand P1_U3420 P1_REG2_REG_18__SCAN_IN ; P1_U6086
g3474 nand P1_U4031 P1_U3395 ; P1_U6087
g3475 nand P1_U3420 P1_REG2_REG_19__SCAN_IN ; P1_U6088
g3476 nand P1_U4031 P1_U3396 ; P1_U6089
g3477 nand P1_U3420 P1_REG2_REG_20__SCAN_IN ; P1_U6090
g3478 nand P1_U4031 P1_U3398 ; P1_U6091
g3479 nand P1_U3420 P1_REG2_REG_21__SCAN_IN ; P1_U6092
g3480 nand P1_U4031 P1_U3400 ; P1_U6093
g3481 nand P1_U3420 P1_REG2_REG_22__SCAN_IN ; P1_U6094
g3482 nand P1_U4031 P1_U3402 ; P1_U6095
g3483 nand P1_U3420 P1_REG2_REG_23__SCAN_IN ; P1_U6096
g3484 nand P1_U4031 P1_U3404 ; P1_U6097
g3485 nand P1_U3420 P1_REG2_REG_24__SCAN_IN ; P1_U6098
g3486 nand P1_U4031 P1_U3406 ; P1_U6099
g3487 nand P1_U3420 P1_REG2_REG_25__SCAN_IN ; P1_U6100
g3488 nand P1_U4031 P1_U3408 ; P1_U6101
g3489 nand P1_U3420 P1_REG2_REG_26__SCAN_IN ; P1_U6102
g3490 nand P1_U4031 P1_U3410 ; P1_U6103
g3491 nand P1_U3420 P1_REG2_REG_27__SCAN_IN ; P1_U6104
g3492 nand P1_U4031 P1_U3412 ; P1_U6105
g3493 nand P1_U3420 P1_REG2_REG_28__SCAN_IN ; P1_U6106
g3494 nand P1_U4031 P1_U3414 ; P1_U6107
g3495 nand P1_U3420 P1_REG2_REG_29__SCAN_IN ; P1_U6108
g3496 nand P1_U4031 P1_U3416 ; P1_U6109
g3497 nand P1_U3420 P1_REG2_REG_30__SCAN_IN ; P1_U6110
g3498 nand P1_U4035 P1_U4031 ; P1_U6111
g3499 nand P1_U3420 P1_REG2_REG_31__SCAN_IN ; P1_U6112
g3500 nand P1_U4035 P1_U4031 ; P1_U6113
g3501 nand P1_U3430 P1_DATAO_REG_0__SCAN_IN ; P1_U6114
g3502 nand P1_U4016 P1_U3077 ; P1_U6115
g3503 nand P1_U3430 P1_DATAO_REG_1__SCAN_IN ; P1_U6116
g3504 nand P1_U4016 P1_U3078 ; P1_U6117
g3505 nand P1_U3430 P1_DATAO_REG_2__SCAN_IN ; P1_U6118
g3506 nand P1_U4016 P1_U3068 ; P1_U6119
g3507 nand P1_U3430 P1_DATAO_REG_3__SCAN_IN ; P1_U6120
g3508 nand P1_U4016 P1_U3064 ; P1_U6121
g3509 nand P1_U3430 P1_DATAO_REG_4__SCAN_IN ; P1_U6122
g3510 nand P1_U4016 P1_U3060 ; P1_U6123
g3511 nand P1_U3430 P1_DATAO_REG_5__SCAN_IN ; P1_U6124
g3512 nand P1_U4016 P1_U3067 ; P1_U6125
g3513 nand P1_U3430 P1_DATAO_REG_6__SCAN_IN ; P1_U6126
g3514 nand P1_U4016 P1_U3071 ; P1_U6127
g3515 nand P1_U3430 P1_DATAO_REG_7__SCAN_IN ; P1_U6128
g3516 nand P1_U4016 P1_U3070 ; P1_U6129
g3517 nand P1_U3430 P1_DATAO_REG_8__SCAN_IN ; P1_U6130
g3518 nand P1_U4016 P1_U3084 ; P1_U6131
g3519 nand P1_U3430 P1_DATAO_REG_9__SCAN_IN ; P1_U6132
g3520 nand P1_U4016 P1_U3083 ; P1_U6133
g3521 nand P1_U3430 P1_DATAO_REG_10__SCAN_IN ; P1_U6134
g3522 nand P1_U4016 P1_U3062 ; P1_U6135
g3523 nand P1_U3430 P1_DATAO_REG_11__SCAN_IN ; P1_U6136
g3524 nand P1_U4016 P1_U3063 ; P1_U6137
g3525 nand P1_U3430 P1_DATAO_REG_12__SCAN_IN ; P1_U6138
g3526 nand P1_U4016 P1_U3072 ; P1_U6139
g3527 nand P1_U3430 P1_DATAO_REG_13__SCAN_IN ; P1_U6140
g3528 nand P1_U4016 P1_U3080 ; P1_U6141
g3529 nand P1_U3430 P1_DATAO_REG_14__SCAN_IN ; P1_U6142
g3530 nand P1_U4016 P1_U3079 ; P1_U6143
g3531 nand P1_U3430 P1_DATAO_REG_15__SCAN_IN ; P1_U6144
g3532 nand P1_U4016 P1_U3074 ; P1_U6145
g3533 nand P1_U3430 P1_DATAO_REG_16__SCAN_IN ; P1_U6146
g3534 nand P1_U4016 P1_U3073 ; P1_U6147
g3535 nand P1_U3430 P1_DATAO_REG_17__SCAN_IN ; P1_U6148
g3536 nand P1_U4016 P1_U3069 ; P1_U6149
g3537 nand P1_U3430 P1_DATAO_REG_18__SCAN_IN ; P1_U6150
g3538 nand P1_U4016 P1_U3082 ; P1_U6151
g3539 nand P1_U3430 P1_DATAO_REG_19__SCAN_IN ; P1_U6152
g3540 nand P1_U4016 P1_U3081 ; P1_U6153
g3541 nand P1_U3430 P1_DATAO_REG_20__SCAN_IN ; P1_U6154
g3542 nand P1_U4016 P1_U3076 ; P1_U6155
g3543 nand P1_U3430 P1_DATAO_REG_21__SCAN_IN ; P1_U6156
g3544 nand P1_U4016 P1_U3075 ; P1_U6157
g3545 nand P1_U3430 P1_DATAO_REG_22__SCAN_IN ; P1_U6158
g3546 nand P1_U4016 P1_U3061 ; P1_U6159
g3547 nand P1_U3430 P1_DATAO_REG_23__SCAN_IN ; P1_U6160
g3548 nand P1_U4016 P1_U3066 ; P1_U6161
g3549 nand P1_U3430 P1_DATAO_REG_24__SCAN_IN ; P1_U6162
g3550 nand P1_U4016 P1_U3065 ; P1_U6163
g3551 nand P1_U3430 P1_DATAO_REG_25__SCAN_IN ; P1_U6164
g3552 nand P1_U4016 P1_U3058 ; P1_U6165
g3553 nand P1_U3430 P1_DATAO_REG_26__SCAN_IN ; P1_U6166
g3554 nand P1_U4016 P1_U3057 ; P1_U6167
g3555 nand P1_U3430 P1_DATAO_REG_27__SCAN_IN ; P1_U6168
g3556 nand P1_U4016 P1_U3053 ; P1_U6169
g3557 nand P1_U3430 P1_DATAO_REG_28__SCAN_IN ; P1_U6170
g3558 nand P1_U4016 P1_U3054 ; P1_U6171
g3559 nand P1_U3430 P1_DATAO_REG_29__SCAN_IN ; P1_U6172
g3560 nand P1_U4016 P1_U3055 ; P1_U6173
g3561 nand P1_U3430 P1_DATAO_REG_30__SCAN_IN ; P1_U6174
g3562 nand P1_U4016 P1_U3059 ; P1_U6175
g3563 nand P1_U3430 P1_DATAO_REG_31__SCAN_IN ; P1_U6176
g3564 nand P1_U4016 P1_U3056 ; P1_U6177
g3565 nand P1_U3450 P1_U5793 P1_U3432 ; P1_U6178
g3566 nand P1_R1375_U9 P1_U4030 ; P1_U6179
g3567 nand P1_U4017 P1_U3054 ; P1_U6180
g3568 nand P1_U3413 P1_U4702 ; P1_U6181
g3569 nand P1_U6181 P1_U6180 ; P1_U6182
g3570 nand P1_U4026 P1_U3056 ; P1_U6183
g3571 nand P1_U3418 P1_U4759 ; P1_U6184
g3572 nand P1_U6184 P1_U6183 ; P1_U6185
g3573 nand P1_U4025 P1_U3076 ; P1_U6186
g3574 nand P1_U3397 P1_U4550 ; P1_U6187
g3575 nand P1_U6187 P1_U6186 ; P1_U6188
g3576 nand P1_U4027 P1_U3059 ; P1_U6189
g3577 nand P1_U3417 P1_U4739 ; P1_U6190
g3578 nand P1_U6190 P1_U6189 ; P1_U6191
g3579 nand P1_U5959 P1_U4531 ; P1_U6192
g3580 nand P1_U3514 P1_U3081 ; P1_U6193
g3581 nand P1_U6193 P1_U6192 ; P1_U6194
g3582 nand P1_U5905 P1_U4379 ; P1_U6195
g3583 nand P1_U3491 P1_U3063 ; P1_U6196
g3584 nand P1_U6196 P1_U6195 ; P1_U6197
g3585 nand P1_U5856 P1_U4246 ; P1_U6198
g3586 nand P1_U3470 P1_U3060 ; P1_U6199
g3587 nand P1_U6199 P1_U6198 ; P1_U6200
g3588 nand P1_U5898 P1_U4360 ; P1_U6201
g3589 nand P1_U3488 P1_U3062 ; P1_U6202
g3590 nand P1_U6202 P1_U6201 ; P1_U6203
g3591 nand P1_U4028 P1_U3055 ; P1_U6204
g3592 nand P1_U3415 P1_U4721 ; P1_U6205
g3593 nand P1_U6205 P1_U6204 ; P1_U6206
g3594 nand P1_U4018 P1_U3053 ; P1_U6207
g3595 nand P1_U3411 P1_U4683 ; P1_U6208
g3596 nand P1_U6208 P1_U6207 ; P1_U6209
g3597 nand P1_U5947 P1_U4493 ; P1_U6210
g3598 nand P1_U3509 P1_U3069 ; P1_U6211
g3599 nand P1_U6211 P1_U6210 ; P1_U6212
g3600 nand P1_U5884 P1_U4322 ; P1_U6213
g3601 nand P1_U3482 P1_U3084 ; P1_U6214
g3602 nand P1_U6214 P1_U6213 ; P1_U6215
g3603 nand P1_U5891 P1_U4341 ; P1_U6216
g3604 nand P1_U3485 P1_U3083 ; P1_U6217
g3605 nand P1_U6217 P1_U6216 ; P1_U6218
g3606 nand P1_U5919 P1_U4417 ; P1_U6219
g3607 nand P1_U3497 P1_U3080 ; P1_U6220
g3608 nand P1_U6220 P1_U6219 ; P1_U6221
g3609 nand P1_U5926 P1_U4436 ; P1_U6222
g3610 nand P1_U3500 P1_U3079 ; P1_U6223
g3611 nand P1_U6223 P1_U6222 ; P1_U6224
g3612 nand P1_U5820 P1_U4208 ; P1_U6225
g3613 nand P1_U3456 P1_U3077 ; P1_U6226
g3614 nand P1_U6226 P1_U6225 ; P1_U6227
g3615 nand P1_U5835 P1_U4184 ; P1_U6228
g3616 nand P1_U3461 P1_U3078 ; P1_U6229
g3617 nand P1_U6229 P1_U6228 ; P1_U6230
g3618 nand P1_U5933 P1_U4455 ; P1_U6231
g3619 nand P1_U3503 P1_U3074 ; P1_U6232
g3620 nand P1_U6232 P1_U6231 ; P1_U6233
g3621 nand P1_U5940 P1_U4474 ; P1_U6234
g3622 nand P1_U3506 P1_U3073 ; P1_U6235
g3623 nand P1_U6235 P1_U6234 ; P1_U6236
g3624 nand P1_U5870 P1_U4284 ; P1_U6237
g3625 nand P1_U3476 P1_U3071 ; P1_U6238
g3626 nand P1_U6238 P1_U6237 ; P1_U6239
g3627 nand P1_U5877 P1_U4303 ; P1_U6240
g3628 nand P1_U3479 P1_U3070 ; P1_U6241
g3629 nand P1_U6241 P1_U6240 ; P1_U6242
g3630 nand P1_U5912 P1_U4398 ; P1_U6243
g3631 nand P1_U3494 P1_U3072 ; P1_U6244
g3632 nand P1_U6244 P1_U6243 ; P1_U6245
g3633 nand P1_U5842 P1_U4203 ; P1_U6246
g3634 nand P1_U3464 P1_U3068 ; P1_U6247
g3635 nand P1_U6247 P1_U6246 ; P1_U6248
g3636 nand P1_U5849 P1_U4227 ; P1_U6249
g3637 nand P1_U3467 P1_U3064 ; P1_U6250
g3638 nand P1_U6250 P1_U6249 ; P1_U6251
g3639 nand P1_U5863 P1_U4265 ; P1_U6252
g3640 nand P1_U3473 P1_U3067 ; P1_U6253
g3641 nand P1_U6253 P1_U6252 ; P1_U6254
g3642 nand P1_U5954 P1_U4512 ; P1_U6255
g3643 nand P1_U3512 P1_U3082 ; P1_U6256
g3644 nand P1_U6256 P1_U6255 ; P1_U6257
g3645 nand P1_U4021 P1_U3065 ; P1_U6258
g3646 nand P1_U3405 P1_U4626 ; P1_U6259
g3647 nand P1_U6259 P1_U6258 ; P1_U6260
g3648 nand P1_U4022 P1_U3066 ; P1_U6261
g3649 nand P1_U3403 P1_U4607 ; P1_U6262
g3650 nand P1_U6262 P1_U6261 ; P1_U6263
g3651 nand P1_U4024 P1_U3075 ; P1_U6264
g3652 nand P1_U3399 P1_U4569 ; P1_U6265
g3653 nand P1_U6265 P1_U6264 ; P1_U6266
g3654 nand P1_U4023 P1_U3061 ; P1_U6267
g3655 nand P1_U3401 P1_U4588 ; P1_U6268
g3656 nand P1_U6268 P1_U6267 ; P1_U6269
g3657 nand P1_U4020 P1_U3058 ; P1_U6270
g3658 nand P1_U3407 P1_U4645 ; P1_U6271
g3659 nand P1_U6271 P1_U6270 ; P1_U6272
g3660 nand P1_U4019 P1_U3057 ; P1_U6273
g3661 nand P1_U3409 P1_U4664 ; P1_U6274
g3662 nand P1_U6274 P1_U6273 ; P1_U6275
g3663 nand P1_U4041 P1_U3991 ; P1_U6276
g3664 nand P1_U5129 P1_U3049 ; P1_U6277
g3665 nand P1_U5133 P1_U3432 P1_U5799 ; P1_U6278
g3666 nand P1_U3453 P1_U5130 ; P1_U6279
g3667 nand P1_U5786 P1_U3431 ; P1_U6280
g3668 nand P1_U3451 P1_U3444 ; P1_U6281
g3669 nand P1_U3450 P1_U5144 ; P1_U6282
g3670 nand P1_U5802 P1_U3994 ; P1_U6283
g3671 nand P1_U3454 P1_U5408 ; P1_U6284
g3672 nand P1_U3015 P1_U5814 P1_REG2_REG_0__SCAN_IN ; P1_U6285
g3673 and P2_U3924 P2_U5671 ; P2_U3014
g3674 and P2_U3937 P2_U3419 ; P2_U3015
g3675 and P2_U3575 P2_U3570 ; P2_U3016
g3676 and P2_U5688 P2_U3423 ; P2_U3017
g3677 and P2_U3426 P2_U3423 ; P2_U3018
g3678 and P2_U3421 P2_U3422 ; P2_U3019
g3679 and P2_U5680 P2_U3421 ; P2_U3020
g3680 and P2_U5677 P2_U3422 ; P2_U3021
g3681 and P2_U5677 P2_U5680 ; P2_U3022
g3682 and P2_U3048 P2_STATE_REG_SCAN_IN ; P2_U3023
g3683 and P2_U3757 P2_U3401 ; P2_U3024
g3684 and P2_U3976 P2_U5671 ; P2_U3025
g3685 and P2_U3963 P2_U5683 ; P2_U3026
g3686 and P2_U3944 P2_U5671 ; P2_U3027
g3687 and P2_U3803 P2_U3946 ; P2_U3028
g3688 and P2_R1299_U6 P2_U3411 ; P2_U3029
g3689 and P2_U3329 P2_STATE_REG_SCAN_IN ; P2_U3030
g3690 and P2_U3932 P2_U3964 ; P2_U3031
g3691 and P2_U3964 P2_U3398 ; P2_U3032
g3692 and P2_U3933 P2_U3964 ; P2_U3033
g3693 and P2_U3938 P2_U3964 ; P2_U3034
g3694 and P2_U3963 P2_U3423 ; P2_U3035
g3695 and P2_U3946 P2_U5683 ; P2_U3036
g3696 and P2_U3964 P2_U3026 ; P2_U3037
g3697 and P2_U3946 P2_U3423 ; P2_U3038
g3698 and P2_U5688 P2_U4854 ; P2_U3039
g3699 and P2_U3024 P2_U5688 ; P2_U3040
g3700 and P2_U5683 P2_U4854 ; P2_U3041
g3701 and P2_U3024 P2_U5683 ; P2_U3042
g3702 and P2_U3018 P2_U4854 ; P2_U3043
g3703 and P2_U3024 P2_U3018 ; P2_U3044
g3704 and P2_U3023 P2_U3401 ; P2_U3045
g3705 and P2_U5184 P2_STATE_REG_SCAN_IN ; P2_U3046
g3706 and P2_U3023 P2_U5186 ; P2_U3047
g3707 and P2_U5658 P2_U3396 ; P2_U3048
g3708 and P2_U3418 P2_U5668 ; P2_U3049
g3709 and P2_U3576 P2_U3016 ; P2_U3050
g3710 and P2_U3341 P2_U3402 P2_U3392 P2_U3338 P2_U3337 ; P2_U3051
g3711 and P2_U3399 P2_STATE_REG_SCAN_IN ; P2_U3052
g3712 and P2_U3820 P2_U5439 P2_U3819 ; P2_U3053
g3713 and P2_U5461 P2_U5460 ; P2_U3054
g3714 nand P2_U4611 P2_U4612 P2_U4610 P2_U4613 ; P2_U3055
g3715 nand P2_U4630 P2_U4631 P2_U4629 P2_U4632 ; P2_U3056
g3716 nand P2_U4651 P2_U4650 P2_U4649 P2_U4648 ; P2_U3057
g3717 nand P2_U4688 P2_U4689 P2_U4687 ; P2_U3058
g3718 nand P2_U4592 P2_U4593 P2_U4591 P2_U4594 ; P2_U3059
g3719 nand P2_U4573 P2_U4574 P2_U4572 P2_U4575 ; P2_U3060
g3720 nand P2_U4668 P2_U4669 P2_U4667 ; P2_U3061
g3721 nand P2_U4176 P2_U4175 P2_U4174 P2_U4173 ; P2_U3062
g3722 nand P2_U4516 P2_U4517 P2_U4515 P2_U4518 ; P2_U3063
g3723 nand P2_U4290 P2_U4289 P2_U4288 P2_U4287 ; P2_U3064
g3724 nand P2_U4309 P2_U4308 P2_U4307 P2_U4306 ; P2_U3065
g3725 nand P2_U4157 P2_U4156 P2_U4155 P2_U4154 ; P2_U3066
g3726 nand P2_U4554 P2_U4555 P2_U4553 P2_U4556 ; P2_U3067
g3727 nand P2_U4535 P2_U4536 P2_U4534 P2_U4537 ; P2_U3068
g3728 nand P2_U4195 P2_U4194 P2_U4193 P2_U4192 ; P2_U3069
g3729 nand P2_U4133 P2_U4132 P2_U4131 P2_U4130 ; P2_U3070
g3730 nand P2_U4421 P2_U4422 P2_U4420 P2_U4423 ; P2_U3071
g3731 nand P2_U4233 P2_U4232 P2_U4231 P2_U4230 ; P2_U3072
g3732 nand P2_U4214 P2_U4213 P2_U4212 P2_U4211 ; P2_U3073
g3733 nand P2_U4328 P2_U4327 P2_U4326 P2_U4325 ; P2_U3074
g3734 nand P2_U4404 P2_U4403 P2_U4402 P2_U4401 ; P2_U3075
g3735 nand P2_U4385 P2_U4384 P2_U4383 P2_U4382 ; P2_U3076
g3736 nand P2_U4497 P2_U4498 P2_U4496 P2_U4499 ; P2_U3077
g3737 nand P2_U4478 P2_U4479 P2_U4477 P2_U4480 ; P2_U3078
g3738 nand P2_U4138 P2_U4137 P2_U4136 P2_U4135 ; P2_U3079
g3739 nand P2_U4114 P2_U4113 P2_U4112 P2_U4111 ; P2_U3080
g3740 nand P2_U4366 P2_U4365 P2_U4364 P2_U4363 ; P2_U3081
g3741 nand P2_U4347 P2_U4346 P2_U4345 P2_U4344 ; P2_U3082
g3742 nand P2_U4459 P2_U4460 P2_U4458 P2_U4461 ; P2_U3083
g3743 nand P2_U4440 P2_U4441 P2_U4439 P2_U4442 ; P2_U3084
g3744 nand P2_U4271 P2_U4270 P2_U4269 P2_U4268 ; P2_U3085
g3745 nand P2_U4252 P2_U4251 P2_U4250 P2_U4249 ; P2_U3086
g3746 nand P2_U3815 P2_U5434 ; P2_U3087
g3747 not P2_STATE_REG_SCAN_IN ; P2_U3088
g3748 nand P2_U5557 P2_U5556 ; P2_U3089
g3749 nand P2_U5559 P2_U5558 ; P2_U3090
g3750 nand P2_U3859 P2_U5563 ; P2_U3091
g3751 nand P2_U3860 P2_U5566 ; P2_U3092
g3752 nand P2_U3861 P2_U5569 ; P2_U3093
g3753 nand P2_U3862 P2_U5572 ; P2_U3094
g3754 nand P2_U3863 P2_U5575 ; P2_U3095
g3755 nand P2_U3864 P2_U5578 ; P2_U3096
g3756 nand P2_U3865 P2_U5581 ; P2_U3097
g3757 nand P2_U3866 P2_U5584 ; P2_U3098
g3758 nand P2_U3867 P2_U5587 ; P2_U3099
g3759 nand P2_U3868 P2_U5590 ; P2_U3100
g3760 nand P2_U3869 P2_U5596 ; P2_U3101
g3761 nand P2_U3870 P2_U5599 ; P2_U3102
g3762 nand P2_U3871 P2_U5602 ; P2_U3103
g3763 nand P2_U3872 P2_U5605 ; P2_U3104
g3764 nand P2_U3873 P2_U5608 ; P2_U3105
g3765 nand P2_U3874 P2_U5611 ; P2_U3106
g3766 nand P2_U3875 P2_U5614 ; P2_U3107
g3767 nand P2_U3876 P2_U5617 ; P2_U3108
g3768 nand P2_U3877 P2_U5620 ; P2_U3109
g3769 nand P2_U3878 P2_U5623 ; P2_U3110
g3770 nand P2_U3857 P2_U5538 ; P2_U3111
g3771 nand P2_U3858 P2_U5541 ; P2_U3112
g3772 nand P2_U5545 P2_U5544 P2_U5546 ; P2_U3113
g3773 nand P2_U5548 P2_U5547 P2_U5549 ; P2_U3114
g3774 nand P2_U5551 P2_U5550 P2_U5552 ; P2_U3115
g3775 nand P2_U5554 P2_U5553 P2_U5555 ; P2_U3116
g3776 nand P2_U5561 P2_U5560 P2_U5562 ; P2_U3117
g3777 nand P2_U5594 P2_U5593 P2_U5595 ; P2_U3118
g3778 nand P2_U5627 P2_U5626 P2_U5628 ; P2_U3119
g3779 nand P2_U5630 P2_U5629 ; P2_U3120
g3780 and P2_U5637 P2_U5632 P2_U5638 ; P2_U3121
g3781 nand P2_U5463 P2_U5462 P2_U5464 ; P2_U3122
g3782 nand P2_U5469 P2_U3831 P2_U5470 ; P2_U3123
g3783 nand P2_U5472 P2_U3832 P2_U5473 ; P2_U3124
g3784 nand P2_U5475 P2_U3833 P2_U5476 ; P2_U3125
g3785 nand P2_U5478 P2_U3834 P2_U5479 ; P2_U3126
g3786 nand P2_U5481 P2_U3835 P2_U5482 ; P2_U3127
g3787 nand P2_U5484 P2_U3836 P2_U5485 ; P2_U3128
g3788 nand P2_U5487 P2_U3837 P2_U5488 ; P2_U3129
g3789 nand P2_U5490 P2_U3838 P2_U5491 ; P2_U3130
g3790 nand P2_U5493 P2_U3839 P2_U5494 ; P2_U3131
g3791 nand P2_U5496 P2_U3840 P2_U5497 ; P2_U3132
g3792 nand P2_U5502 P2_U3843 P2_U5503 ; P2_U3133
g3793 nand P2_U5505 P2_U3844 P2_U5506 ; P2_U3134
g3794 nand P2_U5508 P2_U3845 P2_U5509 ; P2_U3135
g3795 nand P2_U5511 P2_U3846 P2_U5512 ; P2_U3136
g3796 nand P2_U5514 P2_U3847 P2_U5515 ; P2_U3137
g3797 nand P2_U5517 P2_U3848 P2_U5518 ; P2_U3138
g3798 nand P2_U5520 P2_U3849 P2_U5521 ; P2_U3139
g3799 nand P2_U5523 P2_U3850 P2_U5524 ; P2_U3140
g3800 nand P2_U5526 P2_U5525 P2_U3851 ; P2_U3141
g3801 nand P2_U5529 P2_U5528 P2_U3852 ; P2_U3142
g3802 nand P2_U5443 P2_U5442 P2_U3821 ; P2_U3143
g3803 nand P2_U5446 P2_U5445 P2_U3822 ; P2_U3144
g3804 nand P2_U5449 P2_U5448 P2_U3823 ; P2_U3145
g3805 nand P2_U5452 P2_U5451 P2_U3824 ; P2_U3146
g3806 nand P2_U5455 P2_U5454 P2_U3825 ; P2_U3147
g3807 nand P2_U5458 P2_U3826 ; P2_U3148
g3808 nand P2_U5466 P2_U3829 ; P2_U3149
g3809 nand P2_U5499 P2_U3841 ; P2_U3150
g3810 nand P2_U5532 P2_U3853 ; P2_U3151
g3811 nand P2_U5535 P2_U3855 ; P2_U3152
g3812 nand P2_U3817 P2_U3345 P2_U3415 ; P2_U3153
g3813 nand P2_U3015 P2_U5658 ; P2_U3154
g3814 and P2_U5437 P2_U3056 ; P2_U3155
g3815 and P2_U5437 P2_U3055 ; P2_U3156
g3816 and P2_U5437 P2_U3059 ; P2_U3157
g3817 and P2_U5437 P2_U3060 ; P2_U3158
g3818 and P2_U5437 P2_U3067 ; P2_U3159
g3819 and P2_U5437 P2_U3068 ; P2_U3160
g3820 and P2_U5437 P2_U3063 ; P2_U3161
g3821 and P2_U5437 P2_U3077 ; P2_U3162
g3822 and P2_U5437 P2_U3078 ; P2_U3163
g3823 and P2_U5437 P2_U3083 ; P2_U3164
g3824 and P2_U5437 P2_U3084 ; P2_U3165
g3825 and P2_U5437 P2_U3071 ; P2_U3166
g3826 and P2_U5437 P2_U3075 ; P2_U3167
g3827 and P2_U5437 P2_U3076 ; P2_U3168
g3828 and P2_U5437 P2_U3081 ; P2_U3169
g3829 and P2_U5437 P2_U3082 ; P2_U3170
g3830 and P2_U5437 P2_U3074 ; P2_U3171
g3831 and P2_U5437 P2_U3065 ; P2_U3172
g3832 and P2_U5437 P2_U3064 ; P2_U3173
g3833 and P2_U5437 P2_U3085 ; P2_U3174
g3834 and P2_U5437 P2_U3086 ; P2_U3175
g3835 and P2_U5437 P2_U3072 ; P2_U3176
g3836 and P2_U5437 P2_U3073 ; P2_U3177
g3837 and P2_U5437 P2_U3069 ; P2_U3178
g3838 and P2_U5437 P2_U3062 ; P2_U3179
g3839 and P2_U5437 P2_U3066 ; P2_U3180
g3840 and P2_U5437 P2_U3070 ; P2_U3181
g3841 and P2_U5437 P2_U3080 ; P2_U3182
g3842 and P2_U5437 P2_U3079 ; P2_U3183
g3843 nand P2_U3404 P2_U5436 P2_U3343 ; P2_U3184
g3844 nand P2_U5433 P2_U5432 P2_U3814 P2_U5430 ; P2_U3185
g3845 nand P2_U5424 P2_U5423 P2_U5421 P2_U5420 P2_U5422 ; P2_U3186
g3846 nand P2_U5412 P2_U5411 P2_U5415 P2_U5414 P2_U5413 ; P2_U3187
g3847 nand P2_U5406 P2_U5405 P2_U5403 P2_U5402 P2_U5404 ; P2_U3188
g3848 nand P2_U5394 P2_U5393 P2_U5395 P2_U5397 P2_U5396 ; P2_U3189
g3849 nand P2_U5388 P2_U5387 P2_U3813 P2_U5385 ; P2_U3190
g3850 nand P2_U5376 P2_U5375 P2_U5379 P2_U5378 P2_U5377 ; P2_U3191
g3851 nand P2_U5370 P2_U5369 P2_U5367 P2_U5366 P2_U5368 ; P2_U3192
g3852 nand P2_U5361 P2_U5360 P2_U3812 P2_U5358 ; P2_U3193
g3853 nand P2_U5352 P2_U5351 P2_U3811 P2_U5349 ; P2_U3194
g3854 nand P2_U5340 P2_U5339 P2_U5343 P2_U5342 P2_U5341 ; P2_U3195
g3855 nand P2_U5331 P2_U5330 P2_U5334 P2_U5333 P2_U5332 ; P2_U3196
g3856 nand P2_U5325 P2_U5324 P2_U5322 P2_U5321 P2_U5323 ; P2_U3197
g3857 nand P2_U5313 P2_U5312 P2_U5316 P2_U5315 P2_U5314 ; P2_U3198
g3858 nand P2_U5307 P2_U5306 P2_U3810 P2_U5304 ; P2_U3199
g3859 nand P2_U5295 P2_U5294 P2_U5298 P2_U5297 P2_U5296 ; P2_U3200
g3860 nand P2_U5289 P2_U5288 P2_U5286 P2_U5285 P2_U5287 ; P2_U3201
g3861 nand P2_U5280 P2_U5279 P2_U3809 P2_U5277 ; P2_U3202
g3862 nand P2_U5268 P2_U5267 P2_U5269 P2_U5271 P2_U5270 ; P2_U3203
g3863 nand P2_U3808 P2_U5260 P2_U3807 ; P2_U3204
g3864 nand P2_U5251 P2_U5250 P2_U5254 P2_U5253 P2_U5252 ; P2_U3205
g3865 nand P2_U5242 P2_U5241 P2_U5245 P2_U5244 P2_U5243 ; P2_U3206
g3866 nand P2_U5236 P2_U5235 P2_U5233 P2_U5232 P2_U5234 ; P2_U3207
g3867 nand P2_U5224 P2_U5223 P2_U5225 P2_U5227 P2_U5226 ; P2_U3208
g3868 nand P2_U5218 P2_U5217 P2_U3805 P2_U5215 ; P2_U3209
g3869 nand P2_U5206 P2_U5205 P2_U5209 P2_U5208 P2_U5207 ; P2_U3210
g3870 nand P2_U5200 P2_U5199 P2_U3804 P2_U5197 ; P2_U3211
g3871 nand P2_U5191 P2_U5190 P2_U5188 P2_U5187 P2_U5189 ; P2_U3212
g3872 nand P2_U5175 P2_U5174 P2_U5178 P2_U5177 P2_U5176 ; P2_U3213
g3873 nand P2_U5150 P2_U5149 P2_U3785 P2_U3786 ; P2_U3214
g3874 nand P2_U5135 P2_U5134 P2_U3783 P2_U3784 ; P2_U3215
g3875 nand P2_U5120 P2_U5119 P2_U3781 P2_U3782 ; P2_U3216
g3876 nand P2_U5105 P2_U5104 P2_U3779 P2_U3780 ; P2_U3217
g3877 nand P2_U5090 P2_U5089 P2_U3777 P2_U3778 ; P2_U3218
g3878 nand P2_U5075 P2_U5074 P2_U3775 P2_U3776 ; P2_U3219
g3879 nand P2_U5060 P2_U5059 P2_U3773 P2_U3774 ; P2_U3220
g3880 nand P2_U5045 P2_U5044 P2_U3771 P2_U3772 ; P2_U3221
g3881 nand P2_U5030 P2_U5029 P2_U3769 P2_U3770 ; P2_U3222
g3882 nand P2_U5015 P2_U5014 P2_U3768 ; P2_U3223
g3883 nand P2_U5000 P2_U4999 P2_U3767 ; P2_U3224
g3884 nand P2_U4985 P2_U4984 P2_U3766 ; P2_U3225
g3885 nand P2_U4970 P2_U4969 P2_U3765 ; P2_U3226
g3886 nand P2_U4955 P2_U4954 P2_U3764 ; P2_U3227
g3887 nand P2_U4940 P2_U4939 P2_U3763 ; P2_U3228
g3888 nand P2_U4925 P2_U4924 P2_U3762 ; P2_U3229
g3889 nand P2_U4910 P2_U4909 P2_U3761 ; P2_U3230
g3890 nand P2_U4895 P2_U4894 P2_U3760 ; P2_U3231
g3891 nand P2_U4880 P2_U4879 P2_U3759 ; P2_U3232
g3892 nand P2_U4865 P2_U4864 P2_U3758 ; P2_U3233
g3893 nand P2_U3915 P2_U4852 P2_U4853 ; P2_U3234
g3894 nand P2_U3914 P2_U4850 P2_U4851 ; P2_U3235
g3895 nand P2_U4847 P2_U4848 P2_U4849 P2_U4846 P2_U3912 ; P2_U3236
g3896 nand P2_U3753 P2_U3754 P2_U4842 P2_U3911 ; P2_U3237
g3897 nand P2_U3751 P2_U3752 P2_U4837 P2_U3910 ; P2_U3238
g3898 nand P2_U3749 P2_U3750 P2_U4832 P2_U3909 ; P2_U3239
g3899 nand P2_U3747 P2_U3748 P2_U4827 P2_U3908 ; P2_U3240
g3900 nand P2_U3745 P2_U3746 P2_U4822 P2_U3907 ; P2_U3241
g3901 nand P2_U3743 P2_U3744 P2_U4817 P2_U3906 ; P2_U3242
g3902 nand P2_U3741 P2_U3742 P2_U4812 P2_U3905 ; P2_U3243
g3903 nand P2_U3739 P2_U3740 P2_U4807 P2_U3904 ; P2_U3244
g3904 nand P2_U3737 P2_U3738 P2_U4802 P2_U3903 ; P2_U3245
g3905 nand P2_U3735 P2_U3736 P2_U4797 P2_U3902 ; P2_U3246
g3906 nand P2_U3733 P2_U3734 P2_U4792 P2_U3901 ; P2_U3247
g3907 nand P2_U3731 P2_U3732 P2_U4787 P2_U3900 ; P2_U3248
g3908 nand P2_U3729 P2_U3730 P2_U4782 P2_U3899 ; P2_U3249
g3909 nand P2_U3728 P2_U3727 P2_U3898 ; P2_U3250
g3910 nand P2_U3726 P2_U3725 P2_U3897 ; P2_U3251
g3911 nand P2_U3724 P2_U3723 P2_U3896 ; P2_U3252
g3912 nand P2_U3722 P2_U3721 P2_U3895 ; P2_U3253
g3913 nand P2_U3720 P2_U3719 P2_U3894 ; P2_U3254
g3914 nand P2_U3718 P2_U3717 P2_U3893 ; P2_U3255
g3915 nand P2_U3716 P2_U3715 ; P2_U3256
g3916 nand P2_U3714 P2_U3713 ; P2_U3257
g3917 nand P2_U3712 P2_U3711 ; P2_U3258
g3918 nand P2_U3710 P2_U3709 ; P2_U3259
g3919 nand P2_U3708 P2_U3707 ; P2_U3260
g3920 nand P2_U3706 P2_U3705 ; P2_U3261
g3921 nand P2_U3704 P2_U3703 ; P2_U3262
g3922 nand P2_U3702 P2_U3701 ; P2_U3263
g3923 nand P2_U3700 P2_U3699 ; P2_U3264
g3924 nand P2_U3698 P2_U3697 ; P2_U3265
g3925 and P2_U3880 P2_D_REG_31__SCAN_IN ; P2_U3266
g3926 and P2_U3880 P2_D_REG_30__SCAN_IN ; P2_U3267
g3927 and P2_U3880 P2_D_REG_29__SCAN_IN ; P2_U3268
g3928 and P2_U3880 P2_D_REG_28__SCAN_IN ; P2_U3269
g3929 and P2_U3880 P2_D_REG_27__SCAN_IN ; P2_U3270
g3930 and P2_U3880 P2_D_REG_26__SCAN_IN ; P2_U3271
g3931 and P2_U3880 P2_D_REG_25__SCAN_IN ; P2_U3272
g3932 and P2_U3880 P2_D_REG_24__SCAN_IN ; P2_U3273
g3933 and P2_U3880 P2_D_REG_23__SCAN_IN ; P2_U3274
g3934 and P2_U3880 P2_D_REG_22__SCAN_IN ; P2_U3275
g3935 and P2_U3880 P2_D_REG_21__SCAN_IN ; P2_U3276
g3936 and P2_U3880 P2_D_REG_20__SCAN_IN ; P2_U3277
g3937 and P2_U3880 P2_D_REG_19__SCAN_IN ; P2_U3278
g3938 and P2_U3880 P2_D_REG_18__SCAN_IN ; P2_U3279
g3939 and P2_U3880 P2_D_REG_17__SCAN_IN ; P2_U3280
g3940 and P2_U3880 P2_D_REG_16__SCAN_IN ; P2_U3281
g3941 and P2_U3880 P2_D_REG_15__SCAN_IN ; P2_U3282
g3942 and P2_U3880 P2_D_REG_14__SCAN_IN ; P2_U3283
g3943 and P2_U3880 P2_D_REG_13__SCAN_IN ; P2_U3284
g3944 and P2_U3880 P2_D_REG_12__SCAN_IN ; P2_U3285
g3945 and P2_U3880 P2_D_REG_11__SCAN_IN ; P2_U3286
g3946 and P2_U3880 P2_D_REG_10__SCAN_IN ; P2_U3287
g3947 and P2_U3880 P2_D_REG_9__SCAN_IN ; P2_U3288
g3948 and P2_U3880 P2_D_REG_8__SCAN_IN ; P2_U3289
g3949 and P2_U3880 P2_D_REG_7__SCAN_IN ; P2_U3290
g3950 and P2_U3880 P2_D_REG_6__SCAN_IN ; P2_U3291
g3951 and P2_U3880 P2_D_REG_5__SCAN_IN ; P2_U3292
g3952 and P2_U3880 P2_D_REG_4__SCAN_IN ; P2_U3293
g3953 and P2_U3880 P2_D_REG_3__SCAN_IN ; P2_U3294
g3954 and P2_U3880 P2_D_REG_2__SCAN_IN ; P2_U3295
g3955 nand P2_U4073 P2_U4074 P2_U4072 ; P2_U3296
g3956 nand P2_U4070 P2_U4071 P2_U4069 ; P2_U3297
g3957 nand P2_U4067 P2_U4068 P2_U4066 ; P2_U3298
g3958 nand P2_U4064 P2_U4065 P2_U4063 ; P2_U3299
g3959 nand P2_U4061 P2_U4062 P2_U4060 ; P2_U3300
g3960 nand P2_U4058 P2_U4059 P2_U4057 ; P2_U3301
g3961 nand P2_U4055 P2_U4056 P2_U4054 ; P2_U3302
g3962 nand P2_U4052 P2_U4053 P2_U4051 ; P2_U3303
g3963 nand P2_U4049 P2_U4050 P2_U4048 ; P2_U3304
g3964 nand P2_U4046 P2_U4047 P2_U4045 ; P2_U3305
g3965 nand P2_U4043 P2_U4044 P2_U4042 ; P2_U3306
g3966 nand P2_U4040 P2_U4041 P2_U4039 ; P2_U3307
g3967 nand P2_U4037 P2_U4038 P2_U4036 ; P2_U3308
g3968 nand P2_U4034 P2_U4035 P2_U4033 ; P2_U3309
g3969 nand P2_U4031 P2_U4032 P2_U4030 ; P2_U3310
g3970 nand P2_U4028 P2_U4029 P2_U4027 ; P2_U3311
g3971 nand P2_U4025 P2_U4026 P2_U4024 ; P2_U3312
g3972 nand P2_U4022 P2_U4023 P2_U4021 ; P2_U3313
g3973 nand P2_U4019 P2_U4020 P2_U4018 ; P2_U3314
g3974 nand P2_U4016 P2_U4017 P2_U4015 ; P2_U3315
g3975 nand P2_U4013 P2_U4014 P2_U4012 ; P2_U3316
g3976 nand P2_U4010 P2_U4011 P2_U4009 ; P2_U3317
g3977 nand P2_U4007 P2_U4008 P2_U4006 ; P2_U3318
g3978 nand P2_U4004 P2_U4005 P2_U4003 ; P2_U3319
g3979 nand P2_U4001 P2_U4002 P2_U4000 ; P2_U3320
g3980 nand P2_U3998 P2_U3999 P2_U3997 ; P2_U3321
g3981 nand P2_U3995 P2_U3996 P2_U3994 ; P2_U3322
g3982 nand P2_U3992 P2_U3993 P2_U3991 ; P2_U3323
g3983 nand P2_U3989 P2_U3990 P2_U3988 ; P2_U3324
g3984 nand P2_U3986 P2_U3987 P2_U3985 ; P2_U3325
g3985 nand P2_U3983 P2_U3984 P2_U3982 ; P2_U3326
g3986 nand P2_U3980 P2_U3981 P2_U3979 ; P2_U3327
g3987 and P2_U3797 P2_U5641 ; P2_U3328
g3988 nand P2_U3879 P2_STATE_REG_SCAN_IN ; P2_U3329
g3989 not U69 ; P2_U3330
g3990 not P2_B_REG_SCAN_IN ; P2_U3331
g3991 nand P2_U3414 P2_U5649 ; P2_U3332
g3992 nand P2_U3414 P2_U4075 ; P2_U3333
g3993 nand P2_U5671 P2_U3424 P2_U3420 ; P2_U3334
g3994 nand P2_U3418 P2_U3424 P2_U3420 ; P2_U3335
g3995 nand P2_U3049 P2_U3420 ; P2_U3336
g3996 nand P2_U3418 P2_U3424 P2_U3419 ; P2_U3337
g3997 nand P2_U3049 P2_U3419 ; P2_U3338
g3998 nand P2_U5668 P2_U5674 P2_U3420 ; P2_U3339
g3999 nand P2_U5671 P2_U5668 ; P2_U3340
g4000 nand P2_U3974 P2_U3419 ; P2_U3341
g4001 nand P2_U3939 P2_U5665 ; P2_U3342
g4002 nand P2_U5665 P2_U5674 ; P2_U3343
g4003 nand P2_U3420 P2_U3419 ; P2_U3344
g4004 nand P2_U5665 P2_U3424 ; P2_U3345
g4005 nand P2_U3049 P2_U5665 ; P2_U3346
g4006 nand P2_U5688 P2_U5683 ; P2_U3347
g4007 nand P2_U3564 P2_U4123 P2_U3563 ; P2_U3348
g4008 nand P2_U4141 P2_U4140 P2_U3578 P2_U3580 ; P2_U3349
g4009 nand P2_U4160 P2_U4159 P2_U3582 P2_U3584 ; P2_U3350
g4010 nand P2_U4179 P2_U4178 P2_U3586 P2_U3588 ; P2_U3351
g4011 nand P2_U4198 P2_U4197 P2_U3590 P2_U3592 ; P2_U3352
g4012 nand P2_U4217 P2_U4216 P2_U3594 P2_U3596 ; P2_U3353
g4013 nand P2_U4236 P2_U4235 P2_U3598 P2_U3600 ; P2_U3354
g4014 nand P2_U4255 P2_U4254 P2_U3602 P2_U3604 ; P2_U3355
g4015 nand P2_U4274 P2_U4273 P2_U3606 P2_U3608 ; P2_U3356
g4016 nand P2_U4293 P2_U4292 P2_U3610 P2_U3612 ; P2_U3357
g4017 nand P2_U4312 P2_U4311 P2_U3614 P2_U3616 ; P2_U3358
g4018 nand P2_U4331 P2_U4330 P2_U3618 P2_U3620 ; P2_U3359
g4019 nand P2_U4350 P2_U4349 P2_U3622 P2_U3624 ; P2_U3360
g4020 nand P2_U4369 P2_U4368 P2_U3626 P2_U3628 ; P2_U3361
g4021 nand P2_U4388 P2_U4387 P2_U3630 P2_U3632 ; P2_U3362
g4022 nand P2_U4407 P2_U4406 P2_U3634 P2_U3636 ; P2_U3363
g4023 nand P2_U4426 P2_U4425 P2_U3638 P2_U3640 ; P2_U3364
g4024 nand P2_U4445 P2_U4444 P2_U3642 P2_U3644 ; P2_U3365
g4025 nand P2_U4464 P2_U4463 P2_U3646 P2_U3648 ; P2_U3366
g4026 nand P2_U4483 P2_U4482 P2_U3650 P2_U3652 ; P2_U3367
g4027 nand U81 P2_U3347 ; P2_U3368
g4028 nand P2_U4502 P2_U4501 P2_U3654 P2_U3656 ; P2_U3369
g4029 nand U80 P2_U3347 ; P2_U3370
g4030 nand P2_U4521 P2_U4520 P2_U3658 P2_U3660 ; P2_U3371
g4031 nand U79 P2_U3347 ; P2_U3372
g4032 nand P2_U4540 P2_U4539 P2_U3662 P2_U3664 ; P2_U3373
g4033 nand U78 P2_U3347 ; P2_U3374
g4034 nand P2_U4559 P2_U4558 P2_U3666 P2_U3668 ; P2_U3375
g4035 nand U77 P2_U3347 ; P2_U3376
g4036 nand P2_U4578 P2_U4577 P2_U3670 P2_U3672 ; P2_U3377
g4037 nand U76 P2_U3347 ; P2_U3378
g4038 nand P2_U4597 P2_U4596 P2_U3674 P2_U3676 ; P2_U3379
g4039 nand U75 P2_U3347 ; P2_U3380
g4040 nand P2_U4616 P2_U4615 P2_U3678 P2_U3680 ; P2_U3381
g4041 nand U74 P2_U3347 ; P2_U3382
g4042 nand P2_U4635 P2_U4634 P2_U3682 P2_U3684 ; P2_U3383
g4043 nand U73 P2_U3347 ; P2_U3384
g4044 nand P2_U4654 P2_U4653 P2_U4655 P2_U4656 P2_U3687 ; P2_U3385
g4045 nand U72 P2_U3347 ; P2_U3386
g4046 nand P2_U4674 P2_U4673 P2_U4675 P2_U3690 P2_U3692 ; P2_U3387
g4047 nand U70 P2_U3347 ; P2_U3388
g4048 nand U69 P2_U3347 ; P2_U3389
g4049 nand P2_U3944 P2_U3424 ; P2_U3390
g4050 nand P2_U3023 P2_U4698 ; P2_U3391
g4051 nand P2_U5671 P2_U3424 P2_U3419 ; P2_U3392
g4052 nand P2_U3921 P2_U5671 ; P2_U3393
g4053 nand P2_U3944 P2_U5668 ; P2_U3394
g4054 nand P2_U3927 P2_U5671 ; P2_U3395
g4055 nand P2_U3413 P2_U3412 P2_U3414 ; P2_U3396
g4056 nand P2_U3344 P2_U3347 ; P2_U3397
g4057 nand P2_U3934 P2_U4699 ; P2_U3398
g4058 nand P2_U3962 P2_U5658 ; P2_U3399
g4059 nand P2_U3977 P2_STATE_REG_SCAN_IN ; P2_U3400
g4060 nand P2_U3756 P2_U3052 ; P2_U3401
g4061 nand P2_U3974 P2_U3420 ; P2_U3402
g4062 nand P2_U3015 P2_U3018 ; P2_U3403
g4063 nand P2_U5674 P2_U3424 ; P2_U3404
g4064 nand P2_U3023 P2_U3398 ; P2_U3405
g4065 nand P2_U3798 P2_U3016 ; P2_U3406
g4066 nand P2_U5168 P2_U3396 P2_STATE_REG_SCAN_IN ; P2_U3407
g4067 nand P2_U3802 P2_U5172 ; P2_U3408
g4068 not P2_R1299_U6 ; P2_U3409
g4069 nand P2_U3938 P2_U5665 ; P2_U3410
g4070 nand P2_U3335 P2_U3336 P2_U3346 P2_U3923 ; P2_U3411
g4071 nand P2_U5645 P2_U5644 ; P2_U3412
g4072 nand P2_U5648 P2_U5647 ; P2_U3413
g4073 nand P2_U5651 P2_U5650 ; P2_U3414
g4074 nand P2_U5657 P2_U5656 ; P2_U3415
g4075 nand P2_U5660 P2_U5659 ; P2_U3416
g4076 nand P2_U5662 P2_U5661 ; P2_U3417
g4077 nand P2_U5670 P2_U5669 ; P2_U3418
g4078 nand P2_U5673 P2_U5672 ; P2_U3419
g4079 nand P2_U5664 P2_U5663 ; P2_U3420
g4080 nand P2_U5676 P2_U5675 ; P2_U3421
g4081 nand P2_U5679 P2_U5678 ; P2_U3422
g4082 nand P2_U5682 P2_U5681 ; P2_U3423
g4083 nand P2_U5667 P2_U5666 ; P2_U3424
g4084 nand P2_U5685 P2_U5684 ; P2_U3425
g4085 nand P2_U5687 P2_U5686 ; P2_U3426
g4086 nand P2_U5690 P2_U5689 ; P2_U3427
g4087 nand P2_U5698 P2_U5697 ; P2_U3428
g4088 nand P2_U5695 P2_U5694 ; P2_U3429
g4089 nand P2_U5701 P2_U5700 ; P2_U3430
g4090 nand P2_U5703 P2_U5702 ; P2_U3431
g4091 nand P2_U5705 P2_U5704 ; P2_U3432
g4092 nand P2_U5708 P2_U5707 ; P2_U3433
g4093 nand P2_U5710 P2_U5709 ; P2_U3434
g4094 nand P2_U5712 P2_U5711 ; P2_U3435
g4095 nand P2_U5715 P2_U5714 ; P2_U3436
g4096 nand P2_U5717 P2_U5716 ; P2_U3437
g4097 nand P2_U5719 P2_U5718 ; P2_U3438
g4098 nand P2_U5722 P2_U5721 ; P2_U3439
g4099 nand P2_U5724 P2_U5723 ; P2_U3440
g4100 nand P2_U5726 P2_U5725 ; P2_U3441
g4101 nand P2_U5729 P2_U5728 ; P2_U3442
g4102 nand P2_U5731 P2_U5730 ; P2_U3443
g4103 nand P2_U5733 P2_U5732 ; P2_U3444
g4104 nand P2_U5736 P2_U5735 ; P2_U3445
g4105 nand P2_U5738 P2_U5737 ; P2_U3446
g4106 nand P2_U5740 P2_U5739 ; P2_U3447
g4107 nand P2_U5743 P2_U5742 ; P2_U3448
g4108 nand P2_U5745 P2_U5744 ; P2_U3449
g4109 nand P2_U5747 P2_U5746 ; P2_U3450
g4110 nand P2_U5750 P2_U5749 ; P2_U3451
g4111 nand P2_U5752 P2_U5751 ; P2_U3452
g4112 nand P2_U5754 P2_U5753 ; P2_U3453
g4113 nand P2_U5757 P2_U5756 ; P2_U3454
g4114 nand P2_U5759 P2_U5758 ; P2_U3455
g4115 nand P2_U5761 P2_U5760 ; P2_U3456
g4116 nand P2_U5764 P2_U5763 ; P2_U3457
g4117 nand P2_U5766 P2_U5765 ; P2_U3458
g4118 nand P2_U5768 P2_U5767 ; P2_U3459
g4119 nand P2_U5771 P2_U5770 ; P2_U3460
g4120 nand P2_U5773 P2_U5772 ; P2_U3461
g4121 nand P2_U5775 P2_U5774 ; P2_U3462
g4122 nand P2_U5778 P2_U5777 ; P2_U3463
g4123 nand P2_U5780 P2_U5779 ; P2_U3464
g4124 nand P2_U5782 P2_U5781 ; P2_U3465
g4125 nand P2_U5785 P2_U5784 ; P2_U3466
g4126 nand P2_U5787 P2_U5786 ; P2_U3467
g4127 nand P2_U5789 P2_U5788 ; P2_U3468
g4128 nand P2_U5792 P2_U5791 ; P2_U3469
g4129 nand P2_U5794 P2_U5793 ; P2_U3470
g4130 nand P2_U5796 P2_U5795 ; P2_U3471
g4131 nand P2_U5799 P2_U5798 ; P2_U3472
g4132 nand P2_U5801 P2_U5800 ; P2_U3473
g4133 nand P2_U5803 P2_U5802 ; P2_U3474
g4134 nand P2_U5806 P2_U5805 ; P2_U3475
g4135 nand P2_U5808 P2_U5807 ; P2_U3476
g4136 nand P2_U5810 P2_U5809 ; P2_U3477
g4137 nand P2_U5813 P2_U5812 ; P2_U3478
g4138 nand P2_U5815 P2_U5814 ; P2_U3479
g4139 nand P2_U5817 P2_U5816 ; P2_U3480
g4140 nand P2_U5820 P2_U5819 ; P2_U3481
g4141 nand P2_U5822 P2_U5821 ; P2_U3482
g4142 nand P2_U5824 P2_U5823 ; P2_U3483
g4143 nand P2_U5827 P2_U5826 ; P2_U3484
g4144 nand P2_U5829 P2_U5828 ; P2_U3485
g4145 nand P2_U5832 P2_U5831 ; P2_U3486
g4146 nand P2_U5834 P2_U5833 ; P2_U3487
g4147 nand P2_U5836 P2_U5835 ; P2_U3488
g4148 nand P2_U5838 P2_U5837 ; P2_U3489
g4149 nand P2_U5840 P2_U5839 ; P2_U3490
g4150 nand P2_U5842 P2_U5841 ; P2_U3491
g4151 nand P2_U5844 P2_U5843 ; P2_U3492
g4152 nand P2_U5846 P2_U5845 ; P2_U3493
g4153 nand P2_U5848 P2_U5847 ; P2_U3494
g4154 nand P2_U5850 P2_U5849 ; P2_U3495
g4155 nand P2_U5852 P2_U5851 ; P2_U3496
g4156 nand P2_U5854 P2_U5853 ; P2_U3497
g4157 nand P2_U5856 P2_U5855 ; P2_U3498
g4158 nand P2_U5858 P2_U5857 ; P2_U3499
g4159 nand P2_U5860 P2_U5859 ; P2_U3500
g4160 nand P2_U5862 P2_U5861 ; P2_U3501
g4161 nand P2_U5864 P2_U5863 ; P2_U3502
g4162 nand P2_U5866 P2_U5865 ; P2_U3503
g4163 nand P2_U5868 P2_U5867 ; P2_U3504
g4164 nand P2_U5870 P2_U5869 ; P2_U3505
g4165 nand P2_U5872 P2_U5871 ; P2_U3506
g4166 nand P2_U5874 P2_U5873 ; P2_U3507
g4167 nand P2_U5876 P2_U5875 ; P2_U3508
g4168 nand P2_U5878 P2_U5877 ; P2_U3509
g4169 nand P2_U5880 P2_U5879 ; P2_U3510
g4170 nand P2_U5882 P2_U5881 ; P2_U3511
g4171 nand P2_U5884 P2_U5883 ; P2_U3512
g4172 nand P2_U5886 P2_U5885 ; P2_U3513
g4173 nand P2_U5888 P2_U5887 ; P2_U3514
g4174 nand P2_U5890 P2_U5889 ; P2_U3515
g4175 nand P2_U5892 P2_U5891 ; P2_U3516
g4176 nand P2_U5894 P2_U5893 ; P2_U3517
g4177 nand P2_U5896 P2_U5895 ; P2_U3518
g4178 nand P2_U5898 P2_U5897 ; P2_U3519
g4179 nand P2_U5900 P2_U5899 ; P2_U3520
g4180 nand P2_U5902 P2_U5901 ; P2_U3521
g4181 nand P2_U5904 P2_U5903 ; P2_U3522
g4182 nand P2_U5906 P2_U5905 ; P2_U3523
g4183 nand P2_U5908 P2_U5907 ; P2_U3524
g4184 nand P2_U5910 P2_U5909 ; P2_U3525
g4185 nand P2_U5912 P2_U5911 ; P2_U3526
g4186 nand P2_U5914 P2_U5913 ; P2_U3527
g4187 nand P2_U5916 P2_U5915 ; P2_U3528
g4188 nand P2_U5918 P2_U5917 ; P2_U3529
g4189 nand P2_U5920 P2_U5919 ; P2_U3530
g4190 nand P2_U5986 P2_U5985 ; P2_U3531
g4191 nand P2_U5988 P2_U5987 ; P2_U3532
g4192 nand P2_U5990 P2_U5989 ; P2_U3533
g4193 nand P2_U5992 P2_U5991 ; P2_U3534
g4194 nand P2_U5994 P2_U5993 ; P2_U3535
g4195 nand P2_U5996 P2_U5995 ; P2_U3536
g4196 nand P2_U5998 P2_U5997 ; P2_U3537
g4197 nand P2_U6000 P2_U5999 ; P2_U3538
g4198 nand P2_U6002 P2_U6001 ; P2_U3539
g4199 nand P2_U6004 P2_U6003 ; P2_U3540
g4200 nand P2_U6006 P2_U6005 ; P2_U3541
g4201 nand P2_U6008 P2_U6007 ; P2_U3542
g4202 nand P2_U6010 P2_U6009 ; P2_U3543
g4203 nand P2_U6012 P2_U6011 ; P2_U3544
g4204 nand P2_U6014 P2_U6013 ; P2_U3545
g4205 nand P2_U6016 P2_U6015 ; P2_U3546
g4206 nand P2_U6018 P2_U6017 ; P2_U3547
g4207 nand P2_U6020 P2_U6019 ; P2_U3548
g4208 nand P2_U6022 P2_U6021 ; P2_U3549
g4209 nand P2_U6024 P2_U6023 ; P2_U3550
g4210 nand P2_U6026 P2_U6025 ; P2_U3551
g4211 nand P2_U6028 P2_U6027 ; P2_U3552
g4212 nand P2_U6030 P2_U6029 ; P2_U3553
g4213 nand P2_U6032 P2_U6031 ; P2_U3554
g4214 nand P2_U6034 P2_U6033 ; P2_U3555
g4215 nand P2_U6036 P2_U6035 ; P2_U3556
g4216 nand P2_U6038 P2_U6037 ; P2_U3557
g4217 nand P2_U6040 P2_U6039 ; P2_U3558
g4218 nand P2_U6042 P2_U6041 ; P2_U3559
g4219 nand P2_U6044 P2_U6043 ; P2_U3560
g4220 nand P2_U6046 P2_U6045 ; P2_U3561
g4221 nand P2_U6048 P2_U6047 ; P2_U3562
g4222 and P2_U4120 P2_U4119 P2_U4118 P2_U4117 ; P2_U3563
g4223 and P2_U4122 P2_U4121 ; P2_U3564
g4224 and P2_U4127 P2_U4125 ; P2_U3565
g4225 and P2_U4082 P2_U4081 P2_U4080 P2_U4079 ; P2_U3566
g4226 and P2_U4086 P2_U4085 P2_U4084 P2_U4083 ; P2_U3567
g4227 and P2_U4090 P2_U4089 P2_U4088 P2_U4087 ; P2_U3568
g4228 and P2_U4092 P2_U4091 P2_U4093 ; P2_U3569
g4229 and P2_U3569 P2_U3568 P2_U3567 P2_U3566 ; P2_U3570
g4230 and P2_U4097 P2_U4096 P2_U4095 P2_U4094 ; P2_U3571
g4231 and P2_U4101 P2_U4100 P2_U4099 P2_U4098 ; P2_U3572
g4232 and P2_U4105 P2_U4104 P2_U4103 P2_U4102 ; P2_U3573
g4233 and P2_U4107 P2_U4106 P2_U4108 ; P2_U3574
g4234 and P2_U3574 P2_U3573 P2_U3572 P2_U3571 ; P2_U3575
g4235 and P2_U5696 P2_U4110 ; P2_U3576
g4236 and P2_U5699 P2_U3023 ; P2_U3577
g4237 and P2_U4143 P2_U4142 ; P2_U3578
g4238 and P2_U4145 P2_U4144 ; P2_U3579
g4239 and P2_U4147 P2_U4146 P2_U3579 ; P2_U3580
g4240 and P2_U4150 P2_U4149 P2_U4152 P2_U4151 ; P2_U3581
g4241 and P2_U4162 P2_U4161 ; P2_U3582
g4242 and P2_U4164 P2_U4163 ; P2_U3583
g4243 and P2_U4166 P2_U4165 P2_U3583 ; P2_U3584
g4244 and P2_U4169 P2_U4168 P2_U4171 P2_U4170 ; P2_U3585
g4245 and P2_U4181 P2_U4180 ; P2_U3586
g4246 and P2_U4183 P2_U4182 ; P2_U3587
g4247 and P2_U4185 P2_U4184 P2_U3587 ; P2_U3588
g4248 and P2_U4188 P2_U4187 P2_U4190 P2_U4189 ; P2_U3589
g4249 and P2_U4200 P2_U4199 ; P2_U3590
g4250 and P2_U4202 P2_U4201 ; P2_U3591
g4251 and P2_U4204 P2_U4203 P2_U3591 ; P2_U3592
g4252 and P2_U4207 P2_U4206 P2_U4209 P2_U4208 ; P2_U3593
g4253 and P2_U4219 P2_U4218 ; P2_U3594
g4254 and P2_U4221 P2_U4220 ; P2_U3595
g4255 and P2_U4223 P2_U4222 P2_U3595 ; P2_U3596
g4256 and P2_U4226 P2_U4225 P2_U4228 P2_U4227 ; P2_U3597
g4257 and P2_U4238 P2_U4237 ; P2_U3598
g4258 and P2_U4240 P2_U4239 ; P2_U3599
g4259 and P2_U4242 P2_U4241 P2_U3599 ; P2_U3600
g4260 and P2_U4245 P2_U4244 P2_U4247 P2_U4246 ; P2_U3601
g4261 and P2_U4257 P2_U4256 ; P2_U3602
g4262 and P2_U4259 P2_U4258 ; P2_U3603
g4263 and P2_U4261 P2_U4260 P2_U3603 ; P2_U3604
g4264 and P2_U4264 P2_U4263 P2_U4266 P2_U4265 ; P2_U3605
g4265 and P2_U4276 P2_U4275 ; P2_U3606
g4266 and P2_U4278 P2_U4277 ; P2_U3607
g4267 and P2_U4280 P2_U4279 P2_U3607 ; P2_U3608
g4268 and P2_U4283 P2_U4282 P2_U4285 P2_U4284 ; P2_U3609
g4269 and P2_U4295 P2_U4294 ; P2_U3610
g4270 and P2_U4297 P2_U4296 ; P2_U3611
g4271 and P2_U4299 P2_U4298 P2_U3611 ; P2_U3612
g4272 and P2_U4302 P2_U4301 P2_U4304 P2_U4303 ; P2_U3613
g4273 and P2_U4314 P2_U4313 ; P2_U3614
g4274 and P2_U4316 P2_U4315 ; P2_U3615
g4275 and P2_U4318 P2_U4317 P2_U3615 ; P2_U3616
g4276 and P2_U4321 P2_U4320 P2_U4323 P2_U4322 ; P2_U3617
g4277 and P2_U4333 P2_U4332 ; P2_U3618
g4278 and P2_U4335 P2_U4334 ; P2_U3619
g4279 and P2_U4337 P2_U4336 P2_U3619 ; P2_U3620
g4280 and P2_U4340 P2_U4339 P2_U4342 P2_U4341 ; P2_U3621
g4281 and P2_U4352 P2_U4351 ; P2_U3622
g4282 and P2_U4354 P2_U4353 ; P2_U3623
g4283 and P2_U4356 P2_U4355 P2_U3623 ; P2_U3624
g4284 and P2_U4359 P2_U4358 P2_U4361 P2_U4360 ; P2_U3625
g4285 and P2_U4371 P2_U4370 ; P2_U3626
g4286 and P2_U4373 P2_U4372 ; P2_U3627
g4287 and P2_U4375 P2_U4374 P2_U3627 ; P2_U3628
g4288 and P2_U4378 P2_U4377 P2_U4380 P2_U4379 ; P2_U3629
g4289 and P2_U4390 P2_U4389 ; P2_U3630
g4290 and P2_U4392 P2_U4391 ; P2_U3631
g4291 and P2_U4394 P2_U4393 P2_U3631 ; P2_U3632
g4292 and P2_U4397 P2_U4396 P2_U4399 P2_U4398 ; P2_U3633
g4293 and P2_U4409 P2_U4408 ; P2_U3634
g4294 and P2_U4411 P2_U4410 ; P2_U3635
g4295 and P2_U4413 P2_U4412 P2_U3635 ; P2_U3636
g4296 and P2_U4416 P2_U4415 P2_U4418 P2_U4417 ; P2_U3637
g4297 and P2_U4428 P2_U4427 ; P2_U3638
g4298 and P2_U4430 P2_U4429 ; P2_U3639
g4299 and P2_U4432 P2_U4431 P2_U3639 ; P2_U3640
g4300 and P2_U4435 P2_U4434 P2_U4437 P2_U4436 ; P2_U3641
g4301 and P2_U4447 P2_U4446 ; P2_U3642
g4302 and P2_U4449 P2_U4448 ; P2_U3643
g4303 and P2_U4451 P2_U4450 P2_U3643 ; P2_U3644
g4304 and P2_U4454 P2_U4453 P2_U4456 P2_U4455 ; P2_U3645
g4305 and P2_U4466 P2_U4465 ; P2_U3646
g4306 and P2_U4468 P2_U4467 ; P2_U3647
g4307 and P2_U4470 P2_U4469 P2_U3647 ; P2_U3648
g4308 and P2_U4473 P2_U4472 P2_U4475 P2_U4474 ; P2_U3649
g4309 and P2_U4485 P2_U4484 ; P2_U3650
g4310 and P2_U4487 P2_U4486 ; P2_U3651
g4311 and P2_U4489 P2_U4488 P2_U3651 ; P2_U3652
g4312 and P2_U4492 P2_U4491 P2_U4494 P2_U4493 ; P2_U3653
g4313 and P2_U4504 P2_U4503 ; P2_U3654
g4314 and P2_U4506 P2_U4505 ; P2_U3655
g4315 and P2_U4508 P2_U4507 P2_U3655 ; P2_U3656
g4316 and P2_U4511 P2_U4510 P2_U4513 P2_U4512 ; P2_U3657
g4317 and P2_U4523 P2_U4522 ; P2_U3658
g4318 and P2_U4525 P2_U4524 ; P2_U3659
g4319 and P2_U4527 P2_U4526 P2_U3659 ; P2_U3660
g4320 and P2_U4530 P2_U4529 P2_U4532 P2_U4531 ; P2_U3661
g4321 and P2_U4542 P2_U4541 ; P2_U3662
g4322 and P2_U4544 P2_U4543 ; P2_U3663
g4323 and P2_U4546 P2_U4545 P2_U3663 ; P2_U3664
g4324 and P2_U4549 P2_U4548 P2_U4551 P2_U4550 ; P2_U3665
g4325 and P2_U4561 P2_U4560 ; P2_U3666
g4326 and P2_U4563 P2_U4562 ; P2_U3667
g4327 and P2_U4565 P2_U4564 P2_U3667 ; P2_U3668
g4328 and P2_U4568 P2_U4567 P2_U4570 P2_U4569 ; P2_U3669
g4329 and P2_U4580 P2_U4579 ; P2_U3670
g4330 and P2_U4582 P2_U4581 ; P2_U3671
g4331 and P2_U4584 P2_U4583 P2_U3671 ; P2_U3672
g4332 and P2_U4587 P2_U4586 P2_U4589 P2_U4588 ; P2_U3673
g4333 and P2_U4599 P2_U4598 ; P2_U3674
g4334 and P2_U4601 P2_U4600 ; P2_U3675
g4335 and P2_U4603 P2_U4602 P2_U3675 ; P2_U3676
g4336 and P2_U4606 P2_U4605 P2_U4608 P2_U4607 ; P2_U3677
g4337 and P2_U4618 P2_U4617 ; P2_U3678
g4338 and P2_U4620 P2_U4619 ; P2_U3679
g4339 and P2_U4622 P2_U4621 P2_U3679 ; P2_U3680
g4340 and P2_U4625 P2_U4624 P2_U4627 P2_U4626 ; P2_U3681
g4341 and P2_U4637 P2_U4636 ; P2_U3682
g4342 and P2_U4639 P2_U4638 ; P2_U3683
g4343 and P2_U4641 P2_U4640 P2_U3683 ; P2_U3684
g4344 and P2_U4644 P2_U4643 P2_U4646 P2_U4645 ; P2_U3685
g4345 and P2_U4658 P2_U4657 ; P2_U3686
g4346 and P2_U4660 P2_U4659 P2_U3686 ; P2_U3687
g4347 and P2_U4663 P2_U4662 P2_U4665 P2_U4664 ; P2_U3688
g4348 and P2_U4672 P2_U3963 ; P2_U3689
g4349 and P2_U4677 P2_U4676 ; P2_U3690
g4350 and P2_U4679 P2_U4678 ; P2_U3691
g4351 and P2_U4681 P2_U4680 P2_U3691 ; P2_U3692
g4352 and P2_U4685 P2_U4683 P2_U4684 ; P2_U3693
g4353 and P2_U3963 P2_U4672 ; P2_U3694
g4354 and P2_U3023 P2_U3428 ; P2_U3695
g4355 and P2_U5699 P2_U3935 P2_U3429 ; P2_U3696
g4356 and P2_U4702 P2_U4701 P2_U4703 ; P2_U3697
g4357 and P2_U4705 P2_U4704 P2_U3883 ; P2_U3698
g4358 and P2_U4707 P2_U4706 P2_U4708 ; P2_U3699
g4359 and P2_U4710 P2_U4709 P2_U3884 ; P2_U3700
g4360 and P2_U4712 P2_U4711 P2_U4713 ; P2_U3701
g4361 and P2_U4715 P2_U4714 P2_U3885 ; P2_U3702
g4362 and P2_U4717 P2_U4716 P2_U4718 ; P2_U3703
g4363 and P2_U4720 P2_U4719 P2_U3886 ; P2_U3704
g4364 and P2_U4722 P2_U4721 P2_U4723 ; P2_U3705
g4365 and P2_U4725 P2_U4724 P2_U3887 ; P2_U3706
g4366 and P2_U4727 P2_U4726 P2_U4728 ; P2_U3707
g4367 and P2_U4730 P2_U4729 P2_U3888 ; P2_U3708
g4368 and P2_U4732 P2_U4731 P2_U4733 ; P2_U3709
g4369 and P2_U4735 P2_U4734 P2_U3889 ; P2_U3710
g4370 and P2_U4737 P2_U4736 P2_U4738 ; P2_U3711
g4371 and P2_U4740 P2_U4739 P2_U3890 ; P2_U3712
g4372 and P2_U4742 P2_U4741 P2_U4743 ; P2_U3713
g4373 and P2_U4745 P2_U4744 P2_U3891 ; P2_U3714
g4374 and P2_U4747 P2_U4746 P2_U4748 ; P2_U3715
g4375 and P2_U4750 P2_U4749 P2_U3892 ; P2_U3716
g4376 and P2_U4752 P2_U4751 P2_U4753 ; P2_U3717
g4377 and P2_U4755 P2_U4754 ; P2_U3718
g4378 and P2_U4757 P2_U4756 P2_U4758 ; P2_U3719
g4379 and P2_U4760 P2_U4759 ; P2_U3720
g4380 and P2_U4762 P2_U4761 P2_U4763 ; P2_U3721
g4381 and P2_U4765 P2_U4764 ; P2_U3722
g4382 and P2_U4768 P2_U4766 P2_U4767 ; P2_U3723
g4383 and P2_U4770 P2_U4769 ; P2_U3724
g4384 and P2_U4772 P2_U4771 P2_U4773 ; P2_U3725
g4385 and P2_U4775 P2_U4774 ; P2_U3726
g4386 and P2_U4778 P2_U4776 P2_U4777 ; P2_U3727
g4387 and P2_U4780 P2_U4779 ; P2_U3728
g4388 and P2_U4783 P2_U4781 ; P2_U3729
g4389 and P2_U4785 P2_U4784 ; P2_U3730
g4390 and P2_U4788 P2_U4786 ; P2_U3731
g4391 and P2_U4790 P2_U4789 ; P2_U3732
g4392 and P2_U4793 P2_U4791 ; P2_U3733
g4393 and P2_U4795 P2_U4794 ; P2_U3734
g4394 and P2_U4798 P2_U4796 ; P2_U3735
g4395 and P2_U4800 P2_U4799 ; P2_U3736
g4396 and P2_U4803 P2_U4801 ; P2_U3737
g4397 and P2_U4805 P2_U4804 ; P2_U3738
g4398 and P2_U4808 P2_U4806 ; P2_U3739
g4399 and P2_U4810 P2_U4809 ; P2_U3740
g4400 and P2_U4813 P2_U4811 ; P2_U3741
g4401 and P2_U4815 P2_U4814 ; P2_U3742
g4402 and P2_U4818 P2_U4816 ; P2_U3743
g4403 and P2_U4820 P2_U4819 ; P2_U3744
g4404 and P2_U4823 P2_U4821 ; P2_U3745
g4405 and P2_U4825 P2_U4824 ; P2_U3746
g4406 and P2_U4828 P2_U4826 ; P2_U3747
g4407 and P2_U4830 P2_U4829 ; P2_U3748
g4408 and P2_U4833 P2_U4831 ; P2_U3749
g4409 and P2_U4835 P2_U4834 ; P2_U3750
g4410 and P2_U4838 P2_U4836 ; P2_U3751
g4411 and P2_U4840 P2_U4839 ; P2_U3752
g4412 and P2_U4843 P2_U4841 ; P2_U3753
g4413 and P2_U4845 P2_U4844 ; P2_U3754
g4414 and P2_U3335 P2_U3336 P2_U3334 ; P2_U3755
g4415 and P2_U5643 P2_U3397 ; P2_U3756
g4416 and P2_U3415 P2_STATE_REG_SCAN_IN ; P2_U3757
g4417 and P2_U4870 P2_U4868 P2_U4869 P2_U4867 P2_U4866 ; P2_U3758
g4418 and P2_U4885 P2_U4883 P2_U4884 P2_U4882 P2_U4881 ; P2_U3759
g4419 and P2_U4900 P2_U4898 P2_U4899 P2_U4897 P2_U4896 ; P2_U3760
g4420 and P2_U4915 P2_U4913 P2_U4914 P2_U4912 P2_U4911 ; P2_U3761
g4421 and P2_U4930 P2_U4928 P2_U4929 P2_U4927 P2_U4926 ; P2_U3762
g4422 and P2_U4945 P2_U4943 P2_U4944 P2_U4942 P2_U4941 ; P2_U3763
g4423 and P2_U4960 P2_U4958 P2_U4959 P2_U4957 P2_U4956 ; P2_U3764
g4424 and P2_U4975 P2_U4973 P2_U4974 P2_U4972 P2_U4971 ; P2_U3765
g4425 and P2_U4989 P2_U4988 P2_U4990 P2_U4987 P2_U4986 ; P2_U3766
g4426 and P2_U5005 P2_U5003 P2_U5004 P2_U5002 P2_U5001 ; P2_U3767
g4427 and P2_U5019 P2_U5018 P2_U5020 P2_U5017 P2_U5016 ; P2_U3768
g4428 and P2_U5032 P2_U5031 ; P2_U3769
g4429 and P2_U5034 P2_U5033 P2_U5035 ; P2_U3770
g4430 and P2_U5047 P2_U5046 ; P2_U3771
g4431 and P2_U5049 P2_U5048 P2_U5050 ; P2_U3772
g4432 and P2_U5062 P2_U5061 ; P2_U3773
g4433 and P2_U5064 P2_U5063 P2_U5065 ; P2_U3774
g4434 and P2_U5077 P2_U5076 ; P2_U3775
g4435 and P2_U5079 P2_U5078 P2_U5080 ; P2_U3776
g4436 and P2_U5092 P2_U5091 ; P2_U3777
g4437 and P2_U5094 P2_U5093 P2_U5095 ; P2_U3778
g4438 and P2_U5107 P2_U5106 ; P2_U3779
g4439 and P2_U5109 P2_U5108 P2_U5110 ; P2_U3780
g4440 and P2_U5122 P2_U5121 ; P2_U3781
g4441 and P2_U5124 P2_U5123 P2_U5125 ; P2_U3782
g4442 and P2_U5137 P2_U5136 ; P2_U3783
g4443 and P2_U5139 P2_U5138 P2_U5140 ; P2_U3784
g4444 and P2_U5152 P2_U5151 ; P2_U3785
g4445 and P2_U5154 P2_U5153 P2_U5155 ; P2_U3786
g4446 and P2_U5639 P2_U5658 ; P2_U3787
g4447 and P2_U6103 P2_U6100 P2_U6106 ; P2_U3788
g4448 and P2_U6097 P2_U6094 P2_U6091 P2_U6088 ; P2_U3789
g4449 and P2_U6121 P2_U6118 P2_U6115 P2_U6112 ; P2_U3790
g4450 and P2_U6127 P2_U6124 P2_U6130 P2_U6133 ; P2_U3791
g4451 and P2_U3788 P2_U3789 P2_U6109 P2_U3791 P2_U3790 ; P2_U3792
g4452 and P2_U3796 P2_U3795 P2_U6061 P2_U6058 P2_U6055 ; P2_U3793
g4453 and P2_U6145 P2_U6142 P2_U6139 P2_U6136 P2_U6148 ; P2_U3794
g4454 and P2_U6073 P2_U6070 P2_U6067 P2_U6064 ; P2_U3795
g4455 and P2_U6079 P2_U6076 ; P2_U3796
g4456 and P2_U5640 P2_U5631 ; P2_U3797
g4457 and P2_U3428 P2_U3429 ; P2_U3798
g4458 and P2_U3339 P2_U3928 ; P2_U3799
g4459 and P2_U3799 P2_U3342 ; P2_U3800
g4460 and P2_U3395 P2_U3410 ; P2_U3801
g4461 and P2_U5658 P2_U3935 P2_U3399 ; P2_U3802
g4462 and P2_U3023 P2_U5171 ; P2_U3803
g4463 and P2_U5198 P2_U5196 ; P2_U3804
g4464 and P2_U5216 P2_U5214 ; P2_U3805
g4465 and P2_U3969 P2_U3080 ; P2_U3806
g4466 and P2_U5259 P2_U5258 ; P2_U3807
g4467 and P2_U5262 P2_U5261 ; P2_U3808
g4468 and P2_U5278 P2_U5276 ; P2_U3809
g4469 and P2_U5305 P2_U5303 ; P2_U3810
g4470 and P2_U5350 P2_U5348 ; P2_U3811
g4471 and P2_U5359 P2_U5357 ; P2_U3812
g4472 and P2_U5386 P2_U5384 ; P2_U3813
g4473 and P2_U5431 P2_U5429 ; P2_U3814
g4474 and P2_U5435 P2_STATE_REG_SCAN_IN ; P2_U3815
g4475 and P2_U3919 P2_U3936 P2_U3920 ; P2_U3816
g4476 and P2_U5671 P2_U3419 ; P2_U3817
g4477 and P2_U3394 P2_U3339 ; P2_U3818
g4478 and P2_U3342 P2_U3390 P2_U3818 ; P2_U3819
g4479 and P2_U3334 P2_U3928 ; P2_U3820
g4480 and P2_U3415 P2_U5444 ; P2_U3821
g4481 and P2_U3415 P2_U5447 ; P2_U3822
g4482 and P2_U3415 P2_U5450 ; P2_U3823
g4483 and P2_U3415 P2_U5453 ; P2_U3824
g4484 and P2_U3415 P2_U5456 ; P2_U3825
g4485 and P2_U3827 P2_U5457 ; P2_U3826
g4486 and P2_U3415 P2_U5459 ; P2_U3827
g4487 and P2_U5460 P2_U3410 ; P2_U3828
g4488 and P2_U3830 P2_U5465 ; P2_U3829
g4489 and P2_U3415 P2_U5467 ; P2_U3830
g4490 and P2_U3415 P2_U5468 ; P2_U3831
g4491 and P2_U3415 P2_U5471 ; P2_U3832
g4492 and P2_U3415 P2_U5474 ; P2_U3833
g4493 and P2_U3415 P2_U5477 ; P2_U3834
g4494 and P2_U3415 P2_U5480 ; P2_U3835
g4495 and P2_U3415 P2_U5483 ; P2_U3836
g4496 and P2_U3415 P2_U5486 ; P2_U3837
g4497 and P2_U3415 P2_U5489 ; P2_U3838
g4498 and P2_U3415 P2_U5492 ; P2_U3839
g4499 and P2_U3415 P2_U5495 ; P2_U3840
g4500 and P2_U3842 P2_U5498 ; P2_U3841
g4501 and P2_U3415 P2_U5500 ; P2_U3842
g4502 and P2_U3415 P2_U5501 ; P2_U3843
g4503 and P2_U3415 P2_U5504 ; P2_U3844
g4504 and P2_U3415 P2_U5507 ; P2_U3845
g4505 and P2_U3415 P2_U5510 ; P2_U3846
g4506 and P2_U3415 P2_U5513 ; P2_U3847
g4507 and P2_U3415 P2_U5516 ; P2_U3848
g4508 and P2_U3415 P2_U5519 ; P2_U3849
g4509 and P2_U3415 P2_U5522 ; P2_U3850
g4510 and P2_U3415 P2_U5527 ; P2_U3851
g4511 and P2_U3415 P2_U5530 ; P2_U3852
g4512 and P2_U3854 P2_U5531 ; P2_U3853
g4513 and P2_U3415 P2_U5533 ; P2_U3854
g4514 and P2_U3856 P2_U5534 ; P2_U3855
g4515 and P2_U3415 P2_U5536 ; P2_U3856
g4516 and P2_U5539 P2_U5540 ; P2_U3857
g4517 and P2_U5542 P2_U5543 ; P2_U3858
g4518 and P2_U5564 P2_U5565 ; P2_U3859
g4519 and P2_U5567 P2_U5568 ; P2_U3860
g4520 and P2_U5570 P2_U5571 ; P2_U3861
g4521 and P2_U5573 P2_U5574 ; P2_U3862
g4522 and P2_U5576 P2_U5577 ; P2_U3863
g4523 and P2_U5579 P2_U5580 ; P2_U3864
g4524 and P2_U5582 P2_U5583 ; P2_U3865
g4525 and P2_U5585 P2_U5586 ; P2_U3866
g4526 and P2_U5588 P2_U5589 ; P2_U3867
g4527 and P2_U5591 P2_U5592 ; P2_U3868
g4528 and P2_U5597 P2_U5598 ; P2_U3869
g4529 and P2_U5600 P2_U5601 ; P2_U3870
g4530 and P2_U5603 P2_U5604 ; P2_U3871
g4531 and P2_U5606 P2_U5607 ; P2_U3872
g4532 and P2_U5609 P2_U5610 ; P2_U3873
g4533 and P2_U5612 P2_U5613 ; P2_U3874
g4534 and P2_U5615 P2_U5616 ; P2_U3875
g4535 and P2_U5618 P2_U5619 ; P2_U3876
g4536 and P2_U5621 P2_U5622 ; P2_U3877
g4537 and P2_U5624 P2_U5625 ; P2_U3878
g4538 not P2_IR_REG_31__SCAN_IN ; P2_U3879
g4539 nand P2_U3023 P2_U3333 ; P2_U3880
g4540 nand P2_U3577 P2_U3050 ; P2_U3881
g4541 nand P2_U3695 P2_U3050 ; P2_U3882
g4542 and P2_U5922 P2_U5921 ; P2_U3883
g4543 and P2_U5924 P2_U5923 ; P2_U3884
g4544 and P2_U5926 P2_U5925 ; P2_U3885
g4545 and P2_U5928 P2_U5927 ; P2_U3886
g4546 and P2_U5930 P2_U5929 ; P2_U3887
g4547 and P2_U5932 P2_U5931 ; P2_U3888
g4548 and P2_U5934 P2_U5933 ; P2_U3889
g4549 and P2_U5936 P2_U5935 ; P2_U3890
g4550 and P2_U5938 P2_U5937 ; P2_U3891
g4551 and P2_U5940 P2_U5939 ; P2_U3892
g4552 and P2_U5942 P2_U5941 ; P2_U3893
g4553 and P2_U5944 P2_U5943 ; P2_U3894
g4554 and P2_U5946 P2_U5945 ; P2_U3895
g4555 and P2_U5948 P2_U5947 ; P2_U3896
g4556 and P2_U5950 P2_U5949 ; P2_U3897
g4557 and P2_U5952 P2_U5951 ; P2_U3898
g4558 and P2_U5954 P2_U5953 ; P2_U3899
g4559 and P2_U5956 P2_U5955 ; P2_U3900
g4560 and P2_U5958 P2_U5957 ; P2_U3901
g4561 and P2_U5960 P2_U5959 ; P2_U3902
g4562 and P2_U5962 P2_U5961 ; P2_U3903
g4563 and P2_U5964 P2_U5963 ; P2_U3904
g4564 and P2_U5966 P2_U5965 ; P2_U3905
g4565 and P2_U5968 P2_U5967 ; P2_U3906
g4566 and P2_U5970 P2_U5969 ; P2_U3907
g4567 and P2_U5972 P2_U5971 ; P2_U3908
g4568 and P2_U5974 P2_U5973 ; P2_U3909
g4569 and P2_U5976 P2_U5975 ; P2_U3910
g4570 and P2_U5978 P2_U5977 ; P2_U3911
g4571 and P2_U5980 P2_U5979 ; P2_U3912
g4572 nand P2_U3694 P2_U3058 ; P2_U3913
g4573 and P2_U5982 P2_U5981 ; P2_U3914
g4574 and P2_U5984 P2_U5983 ; P2_U3915
g4575 not P2_R1312_U18 ; P2_U3916
g4576 and P2_U6050 P2_U6049 ; P2_U3917
g4577 nand P2_U3794 P2_U3792 P2_U6085 P2_U6082 P2_U3793 ; P2_U3918
g4578 nand P2_U3049 P2_U5674 ; P2_U3919
g4579 nand P2_U3973 P2_U3418 ; P2_U3920
g4580 not P2_U3390 ; P2_U3921
g4581 not P2_U3342 ; P2_U3922
g4582 nand P2_U3976 P2_U3418 ; P2_U3923
g4583 not P2_U3339 ; P2_U3924
g4584 not P2_U3346 ; P2_U3925
g4585 not P2_U3336 ; P2_U3926
g4586 not P2_U3394 ; P2_U3927
g4587 nand P2_U3973 P2_U3420 ; P2_U3928
g4588 not P2_U3410 ; P2_U3929
g4589 not P2_U3335 ; P2_U3930
g4590 not P2_U3334 ; P2_U3931
g4591 not P2_U3395 ; P2_U3932
g4592 not P2_U3393 ; P2_U3933
g4593 nand P2_U3925 P2_U5674 ; P2_U3934
g4594 nand P2_U3963 P2_U3340 ; P2_U3935
g4595 nand P2_U3973 P2_U5671 ; P2_U3936
g4596 not P2_U3402 ; P2_U3937
g4597 not P2_U3392 ; P2_U3938
g4598 not P2_U3341 ; P2_U3939
g4599 not P2_U3919 ; P2_U3940
g4600 not P2_U3337 ; P2_U3941
g4601 not P2_U3920 ; P2_U3942
g4602 not P2_U3338 ; P2_U3943
g4603 not P2_U3343 ; P2_U3944
g4604 not P2_U3347 ; P2_U3945
g4605 not P2_U3406 ; P2_U3946
g4606 not P2_U3400 ; P2_U3947
g4607 not P2_U3397 ; P2_U3948
g4608 not P2_U3384 ; P2_U3949
g4609 not P2_U3382 ; P2_U3950
g4610 not P2_U3380 ; P2_U3951
g4611 not P2_U3378 ; P2_U3952
g4612 not P2_U3376 ; P2_U3953
g4613 not P2_U3374 ; P2_U3954
g4614 not P2_U3372 ; P2_U3955
g4615 not P2_U3370 ; P2_U3956
g4616 not P2_U3368 ; P2_U3957
g4617 not P2_U3389 ; P2_U3958
g4618 not P2_U3388 ; P2_U3959
g4619 not P2_U3386 ; P2_U3960
g4620 not P2_U3403 ; P2_U3961
g4621 not P2_U3396 ; P2_U3962
g4622 not P2_U3344 ; P2_U3963
g4623 not P2_U3391 ; P2_U3964
g4624 not P2_U3882 ; P2_U3965
g4625 not P2_U3881 ; P2_U3966
g4626 not P2_U3880 ; P2_U3967
g4627 not P2_U3913 ; P2_U3968
g4628 not P2_U3407 ; P2_U3969
g4629 nand P2_U3408 P2_STATE_REG_SCAN_IN ; P2_U3970
g4630 nand P2_U3933 P2_U3023 ; P2_U3971
g4631 not P2_U3405 ; P2_U3972
g4632 not P2_U3404 ; P2_U3973
g4633 not P2_U3340 ; P2_U3974
g4634 not P2_U3332 ; P2_U3975
g4635 not P2_U3345 ; P2_U3976
g4636 not P2_U3399 ; P2_U3977
g4637 not P2_U3329 ; P2_U3978
g4638 nand U93 P2_U3088 ; P2_U3979
g4639 nand P2_U3030 P2_IR_REG_0__SCAN_IN ; P2_U3980
g4640 nand P2_U3978 P2_IR_REG_0__SCAN_IN ; P2_U3981
g4641 nand U82 P2_U3088 ; P2_U3982
g4642 nand P2_SUB_1108_U42 P2_U3030 ; P2_U3983
g4643 nand P2_U3978 P2_IR_REG_1__SCAN_IN ; P2_U3984
g4644 nand U71 P2_U3088 ; P2_U3985
g4645 nand P2_SUB_1108_U17 P2_U3030 ; P2_U3986
g4646 nand P2_U3978 P2_IR_REG_2__SCAN_IN ; P2_U3987
g4647 nand U68 P2_U3088 ; P2_U3988
g4648 nand P2_SUB_1108_U18 P2_U3030 ; P2_U3989
g4649 nand P2_U3978 P2_IR_REG_3__SCAN_IN ; P2_U3990
g4650 nand U67 P2_U3088 ; P2_U3991
g4651 nand P2_SUB_1108_U19 P2_U3030 ; P2_U3992
g4652 nand P2_U3978 P2_IR_REG_4__SCAN_IN ; P2_U3993
g4653 nand U66 P2_U3088 ; P2_U3994
g4654 nand P2_SUB_1108_U101 P2_U3030 ; P2_U3995
g4655 nand P2_U3978 P2_IR_REG_5__SCAN_IN ; P2_U3996
g4656 nand U65 P2_U3088 ; P2_U3997
g4657 nand P2_SUB_1108_U20 P2_U3030 ; P2_U3998
g4658 nand P2_U3978 P2_IR_REG_6__SCAN_IN ; P2_U3999
g4659 nand U64 P2_U3088 ; P2_U4000
g4660 nand P2_SUB_1108_U21 P2_U3030 ; P2_U4001
g4661 nand P2_U3978 P2_IR_REG_7__SCAN_IN ; P2_U4002
g4662 nand U63 P2_U3088 ; P2_U4003
g4663 nand P2_SUB_1108_U22 P2_U3030 ; P2_U4004
g4664 nand P2_U3978 P2_IR_REG_8__SCAN_IN ; P2_U4005
g4665 nand U62 P2_U3088 ; P2_U4006
g4666 nand P2_SUB_1108_U99 P2_U3030 ; P2_U4007
g4667 nand P2_U3978 P2_IR_REG_9__SCAN_IN ; P2_U4008
g4668 nand U92 P2_U3088 ; P2_U4009
g4669 nand P2_SUB_1108_U6 P2_U3030 ; P2_U4010
g4670 nand P2_U3978 P2_IR_REG_10__SCAN_IN ; P2_U4011
g4671 nand U91 P2_U3088 ; P2_U4012
g4672 nand P2_SUB_1108_U7 P2_U3030 ; P2_U4013
g4673 nand P2_U3978 P2_IR_REG_11__SCAN_IN ; P2_U4014
g4674 nand U90 P2_U3088 ; P2_U4015
g4675 nand P2_SUB_1108_U8 P2_U3030 ; P2_U4016
g4676 nand P2_U3978 P2_IR_REG_12__SCAN_IN ; P2_U4017
g4677 nand U89 P2_U3088 ; P2_U4018
g4678 nand P2_SUB_1108_U127 P2_U3030 ; P2_U4019
g4679 nand P2_U3978 P2_IR_REG_13__SCAN_IN ; P2_U4020
g4680 nand U88 P2_U3088 ; P2_U4021
g4681 nand P2_SUB_1108_U9 P2_U3030 ; P2_U4022
g4682 nand P2_U3978 P2_IR_REG_14__SCAN_IN ; P2_U4023
g4683 nand U87 P2_U3088 ; P2_U4024
g4684 nand P2_SUB_1108_U10 P2_U3030 ; P2_U4025
g4685 nand P2_U3978 P2_IR_REG_15__SCAN_IN ; P2_U4026
g4686 nand U86 P2_U3088 ; P2_U4027
g4687 nand P2_SUB_1108_U11 P2_U3030 ; P2_U4028
g4688 nand P2_U3978 P2_IR_REG_16__SCAN_IN ; P2_U4029
g4689 nand U85 P2_U3088 ; P2_U4030
g4690 nand P2_SUB_1108_U125 P2_U3030 ; P2_U4031
g4691 nand P2_U3978 P2_IR_REG_17__SCAN_IN ; P2_U4032
g4692 nand U84 P2_U3088 ; P2_U4033
g4693 nand P2_SUB_1108_U12 P2_U3030 ; P2_U4034
g4694 nand P2_U3978 P2_IR_REG_18__SCAN_IN ; P2_U4035
g4695 nand U83 P2_U3088 ; P2_U4036
g4696 nand P2_SUB_1108_U123 P2_U3030 ; P2_U4037
g4697 nand P2_U3978 P2_IR_REG_19__SCAN_IN ; P2_U4038
g4698 nand U81 P2_U3088 ; P2_U4039
g4699 nand P2_SUB_1108_U119 P2_U3030 ; P2_U4040
g4700 nand P2_U3978 P2_IR_REG_20__SCAN_IN ; P2_U4041
g4701 nand U80 P2_U3088 ; P2_U4042
g4702 nand P2_SUB_1108_U116 P2_U3030 ; P2_U4043
g4703 nand P2_U3978 P2_IR_REG_21__SCAN_IN ; P2_U4044
g4704 nand U79 P2_U3088 ; P2_U4045
g4705 nand P2_SUB_1108_U114 P2_U3030 ; P2_U4046
g4706 nand P2_U3978 P2_IR_REG_22__SCAN_IN ; P2_U4047
g4707 nand U78 P2_U3088 ; P2_U4048
g4708 nand P2_SUB_1108_U13 P2_U3030 ; P2_U4049
g4709 nand P2_U3978 P2_IR_REG_23__SCAN_IN ; P2_U4050
g4710 nand U77 P2_U3088 ; P2_U4051
g4711 nand P2_SUB_1108_U14 P2_U3030 ; P2_U4052
g4712 nand P2_U3978 P2_IR_REG_24__SCAN_IN ; P2_U4053
g4713 nand U76 P2_U3088 ; P2_U4054
g4714 nand P2_SUB_1108_U112 P2_U3030 ; P2_U4055
g4715 nand P2_U3978 P2_IR_REG_25__SCAN_IN ; P2_U4056
g4716 nand U75 P2_U3088 ; P2_U4057
g4717 nand P2_SUB_1108_U15 P2_U3030 ; P2_U4058
g4718 nand P2_U3978 P2_IR_REG_26__SCAN_IN ; P2_U4059
g4719 nand U74 P2_U3088 ; P2_U4060
g4720 nand P2_SUB_1108_U110 P2_U3030 ; P2_U4061
g4721 nand P2_U3978 P2_IR_REG_27__SCAN_IN ; P2_U4062
g4722 nand U73 P2_U3088 ; P2_U4063
g4723 nand P2_SUB_1108_U107 P2_U3030 ; P2_U4064
g4724 nand P2_U3978 P2_IR_REG_28__SCAN_IN ; P2_U4065
g4725 nand U72 P2_U3088 ; P2_U4066
g4726 nand P2_SUB_1108_U16 P2_U3030 ; P2_U4067
g4727 nand P2_U3978 P2_IR_REG_29__SCAN_IN ; P2_U4068
g4728 nand U70 P2_U3088 ; P2_U4069
g4729 nand P2_SUB_1108_U104 P2_U3030 ; P2_U4070
g4730 nand P2_U3978 P2_IR_REG_30__SCAN_IN ; P2_U4071
g4731 nand U69 P2_U3088 ; P2_U4072
g4732 nand P2_SUB_1108_U43 P2_U3030 ; P2_U4073
g4733 nand P2_U3978 P2_IR_REG_31__SCAN_IN ; P2_U4074
g4734 nand P2_U3975 P2_U5655 ; P2_U4075
g4735 not P2_U3333 ; P2_U4076
g4736 nand P2_U3332 P2_U5646 ; P2_U4077
g4737 nand P2_U3332 P2_U5649 ; P2_U4078
g4738 nand P2_U4076 P2_D_REG_10__SCAN_IN ; P2_U4079
g4739 nand P2_U4076 P2_D_REG_11__SCAN_IN ; P2_U4080
g4740 nand P2_U4076 P2_D_REG_12__SCAN_IN ; P2_U4081
g4741 nand P2_U4076 P2_D_REG_13__SCAN_IN ; P2_U4082
g4742 nand P2_U4076 P2_D_REG_14__SCAN_IN ; P2_U4083
g4743 nand P2_U4076 P2_D_REG_15__SCAN_IN ; P2_U4084
g4744 nand P2_U4076 P2_D_REG_16__SCAN_IN ; P2_U4085
g4745 nand P2_U4076 P2_D_REG_17__SCAN_IN ; P2_U4086
g4746 nand P2_U4076 P2_D_REG_18__SCAN_IN ; P2_U4087
g4747 nand P2_U4076 P2_D_REG_19__SCAN_IN ; P2_U4088
g4748 nand P2_U4076 P2_D_REG_20__SCAN_IN ; P2_U4089
g4749 nand P2_U4076 P2_D_REG_21__SCAN_IN ; P2_U4090
g4750 nand P2_U4076 P2_D_REG_22__SCAN_IN ; P2_U4091
g4751 nand P2_U4076 P2_D_REG_23__SCAN_IN ; P2_U4092
g4752 nand P2_U4076 P2_D_REG_24__SCAN_IN ; P2_U4093
g4753 nand P2_U4076 P2_D_REG_25__SCAN_IN ; P2_U4094
g4754 nand P2_U4076 P2_D_REG_26__SCAN_IN ; P2_U4095
g4755 nand P2_U4076 P2_D_REG_27__SCAN_IN ; P2_U4096
g4756 nand P2_U4076 P2_D_REG_28__SCAN_IN ; P2_U4097
g4757 nand P2_U4076 P2_D_REG_29__SCAN_IN ; P2_U4098
g4758 nand P2_U4076 P2_D_REG_2__SCAN_IN ; P2_U4099
g4759 nand P2_U4076 P2_D_REG_30__SCAN_IN ; P2_U4100
g4760 nand P2_U4076 P2_D_REG_31__SCAN_IN ; P2_U4101
g4761 nand P2_U4076 P2_D_REG_3__SCAN_IN ; P2_U4102
g4762 nand P2_U4076 P2_D_REG_4__SCAN_IN ; P2_U4103
g4763 nand P2_U4076 P2_D_REG_5__SCAN_IN ; P2_U4104
g4764 nand P2_U4076 P2_D_REG_6__SCAN_IN ; P2_U4105
g4765 nand P2_U4076 P2_D_REG_7__SCAN_IN ; P2_U4106
g4766 nand P2_U4076 P2_D_REG_8__SCAN_IN ; P2_U4107
g4767 nand P2_U4076 P2_D_REG_9__SCAN_IN ; P2_U4108
g4768 nand P2_U5674 P2_U5671 ; P2_U4109
g4769 nand P2_U5693 P2_U5692 P2_U3340 ; P2_U4110
g4770 nand P2_U3020 P2_REG2_REG_1__SCAN_IN ; P2_U4111
g4771 nand P2_U3021 P2_REG1_REG_1__SCAN_IN ; P2_U4112
g4772 nand P2_U3022 P2_REG0_REG_1__SCAN_IN ; P2_U4113
g4773 nand P2_U3019 P2_REG3_REG_1__SCAN_IN ; P2_U4114
g4774 not P2_U3080 ; P2_U4115
g4775 nand P2_U3390 P2_U3934 ; P2_U4116
g4776 nand P2_U3931 P2_R1146_U20 ; P2_U4117
g4777 nand P2_U3930 P2_R1113_U20 ; P2_U4118
g4778 nand P2_U3926 P2_R1131_U95 ; P2_U4119
g4779 nand P2_U3941 P2_R1179_U20 ; P2_U4120
g4780 nand P2_U3943 P2_R1203_U20 ; P2_U4121
g4781 nand P2_U3014 P2_R1164_U95 ; P2_U4122
g4782 nand P2_U3922 P2_R1233_U95 ; P2_U4123
g4783 not P2_U3348 ; P2_U4124
g4784 nand P2_U3427 P2_U3027 ; P2_U4125
g4785 nand P2_U3026 P2_U3080 ; P2_U4126
g4786 nand P2_R1215_U96 P2_U3025 ; P2_U4127
g4787 nand P2_U3427 P2_U4116 ; P2_U4128
g4788 nand P2_U4128 P2_U4126 P2_U3565 P2_U4124 ; P2_U4129
g4789 nand P2_U3020 P2_REG2_REG_2__SCAN_IN ; P2_U4130
g4790 nand P2_U3021 P2_REG1_REG_2__SCAN_IN ; P2_U4131
g4791 nand P2_U3022 P2_REG0_REG_2__SCAN_IN ; P2_U4132
g4792 nand P2_U3019 P2_REG3_REG_2__SCAN_IN ; P2_U4133
g4793 not P2_U3070 ; P2_U4134
g4794 nand P2_U3020 P2_REG2_REG_0__SCAN_IN ; P2_U4135
g4795 nand P2_U3021 P2_REG1_REG_0__SCAN_IN ; P2_U4136
g4796 nand P2_U3022 P2_REG0_REG_0__SCAN_IN ; P2_U4137
g4797 nand P2_U3019 P2_REG3_REG_0__SCAN_IN ; P2_U4138
g4798 not P2_U3079 ; P2_U4139
g4799 nand P2_U3035 P2_U3079 ; P2_U4140
g4800 nand P2_R1146_U97 P2_U3931 ; P2_U4141
g4801 nand P2_R1113_U97 P2_U3930 ; P2_U4142
g4802 nand P2_R1131_U94 P2_U3926 ; P2_U4143
g4803 nand P2_R1179_U97 P2_U3941 ; P2_U4144
g4804 nand P2_R1203_U97 P2_U3943 ; P2_U4145
g4805 nand P2_R1164_U94 P2_U3014 ; P2_U4146
g4806 nand P2_R1233_U94 P2_U3922 ; P2_U4147
g4807 not P2_U3349 ; P2_U4148
g4808 nand P2_R1275_U55 P2_U3027 ; P2_U4149
g4809 nand P2_U3026 P2_U3070 ; P2_U4150
g4810 nand P2_R1215_U95 P2_U3025 ; P2_U4151
g4811 nand P2_U3432 P2_U4116 ; P2_U4152
g4812 nand P2_U3581 P2_U4148 ; P2_U4153
g4813 nand P2_U3020 P2_REG2_REG_3__SCAN_IN ; P2_U4154
g4814 nand P2_U3021 P2_REG1_REG_3__SCAN_IN ; P2_U4155
g4815 nand P2_U3022 P2_REG0_REG_3__SCAN_IN ; P2_U4156
g4816 nand P2_ADD_1119_U4 P2_U3019 ; P2_U4157
g4817 not P2_U3066 ; P2_U4158
g4818 nand P2_U3035 P2_U3080 ; P2_U4159
g4819 nand P2_R1146_U107 P2_U3931 ; P2_U4160
g4820 nand P2_R1113_U107 P2_U3930 ; P2_U4161
g4821 nand P2_R1131_U16 P2_U3926 ; P2_U4162
g4822 nand P2_R1179_U107 P2_U3941 ; P2_U4163
g4823 nand P2_R1203_U107 P2_U3943 ; P2_U4164
g4824 nand P2_R1164_U16 P2_U3014 ; P2_U4165
g4825 nand P2_R1233_U16 P2_U3922 ; P2_U4166
g4826 not P2_U3350 ; P2_U4167
g4827 nand P2_R1275_U18 P2_U3027 ; P2_U4168
g4828 nand P2_U3026 P2_U3066 ; P2_U4169
g4829 nand P2_R1215_U17 P2_U3025 ; P2_U4170
g4830 nand P2_U3435 P2_U4116 ; P2_U4171
g4831 nand P2_U3585 P2_U4167 ; P2_U4172
g4832 nand P2_U3020 P2_REG2_REG_4__SCAN_IN ; P2_U4173
g4833 nand P2_U3021 P2_REG1_REG_4__SCAN_IN ; P2_U4174
g4834 nand P2_U3022 P2_REG0_REG_4__SCAN_IN ; P2_U4175
g4835 nand P2_ADD_1119_U55 P2_U3019 ; P2_U4176
g4836 not P2_U3062 ; P2_U4177
g4837 nand P2_U3035 P2_U3070 ; P2_U4178
g4838 nand P2_R1146_U17 P2_U3931 ; P2_U4179
g4839 nand P2_R1113_U17 P2_U3930 ; P2_U4180
g4840 nand P2_R1131_U100 P2_U3926 ; P2_U4181
g4841 nand P2_R1179_U17 P2_U3941 ; P2_U4182
g4842 nand P2_R1203_U17 P2_U3943 ; P2_U4183
g4843 nand P2_R1164_U100 P2_U3014 ; P2_U4184
g4844 nand P2_R1233_U100 P2_U3922 ; P2_U4185
g4845 not P2_U3351 ; P2_U4186
g4846 nand P2_R1275_U20 P2_U3027 ; P2_U4187
g4847 nand P2_U3026 P2_U3062 ; P2_U4188
g4848 nand P2_R1215_U101 P2_U3025 ; P2_U4189
g4849 nand P2_U3438 P2_U4116 ; P2_U4190
g4850 nand P2_U3589 P2_U4186 ; P2_U4191
g4851 nand P2_U3020 P2_REG2_REG_5__SCAN_IN ; P2_U4192
g4852 nand P2_U3021 P2_REG1_REG_5__SCAN_IN ; P2_U4193
g4853 nand P2_U3022 P2_REG0_REG_5__SCAN_IN ; P2_U4194
g4854 nand P2_ADD_1119_U54 P2_U3019 ; P2_U4195
g4855 not P2_U3069 ; P2_U4196
g4856 nand P2_U3035 P2_U3066 ; P2_U4197
g4857 nand P2_R1146_U106 P2_U3931 ; P2_U4198
g4858 nand P2_R1113_U106 P2_U3930 ; P2_U4199
g4859 nand P2_R1131_U99 P2_U3926 ; P2_U4200
g4860 nand P2_R1179_U106 P2_U3941 ; P2_U4201
g4861 nand P2_R1203_U106 P2_U3943 ; P2_U4202
g4862 nand P2_R1164_U99 P2_U3014 ; P2_U4203
g4863 nand P2_R1233_U99 P2_U3922 ; P2_U4204
g4864 not P2_U3352 ; P2_U4205
g4865 nand P2_R1275_U21 P2_U3027 ; P2_U4206
g4866 nand P2_U3026 P2_U3069 ; P2_U4207
g4867 nand P2_R1215_U100 P2_U3025 ; P2_U4208
g4868 nand P2_U3441 P2_U4116 ; P2_U4209
g4869 nand P2_U3593 P2_U4205 ; P2_U4210
g4870 nand P2_U3020 P2_REG2_REG_6__SCAN_IN ; P2_U4211
g4871 nand P2_U3021 P2_REG1_REG_6__SCAN_IN ; P2_U4212
g4872 nand P2_U3022 P2_REG0_REG_6__SCAN_IN ; P2_U4213
g4873 nand P2_ADD_1119_U53 P2_U3019 ; P2_U4214
g4874 not P2_U3073 ; P2_U4215
g4875 nand P2_U3035 P2_U3062 ; P2_U4216
g4876 nand P2_R1146_U105 P2_U3931 ; P2_U4217
g4877 nand P2_R1113_U105 P2_U3930 ; P2_U4218
g4878 nand P2_R1131_U17 P2_U3926 ; P2_U4219
g4879 nand P2_R1179_U105 P2_U3941 ; P2_U4220
g4880 nand P2_R1203_U105 P2_U3943 ; P2_U4221
g4881 nand P2_R1164_U17 P2_U3014 ; P2_U4222
g4882 nand P2_R1233_U17 P2_U3922 ; P2_U4223
g4883 not P2_U3353 ; P2_U4224
g4884 nand P2_R1275_U65 P2_U3027 ; P2_U4225
g4885 nand P2_U3026 P2_U3073 ; P2_U4226
g4886 nand P2_R1215_U18 P2_U3025 ; P2_U4227
g4887 nand P2_U3444 P2_U4116 ; P2_U4228
g4888 nand P2_U3597 P2_U4224 ; P2_U4229
g4889 nand P2_U3020 P2_REG2_REG_7__SCAN_IN ; P2_U4230
g4890 nand P2_U3021 P2_REG1_REG_7__SCAN_IN ; P2_U4231
g4891 nand P2_U3022 P2_REG0_REG_7__SCAN_IN ; P2_U4232
g4892 nand P2_ADD_1119_U52 P2_U3019 ; P2_U4233
g4893 not P2_U3072 ; P2_U4234
g4894 nand P2_U3035 P2_U3069 ; P2_U4235
g4895 nand P2_R1146_U18 P2_U3931 ; P2_U4236
g4896 nand P2_R1113_U18 P2_U3930 ; P2_U4237
g4897 nand P2_R1131_U98 P2_U3926 ; P2_U4238
g4898 nand P2_R1179_U18 P2_U3941 ; P2_U4239
g4899 nand P2_R1203_U18 P2_U3943 ; P2_U4240
g4900 nand P2_R1164_U98 P2_U3014 ; P2_U4241
g4901 nand P2_R1233_U98 P2_U3922 ; P2_U4242
g4902 not P2_U3354 ; P2_U4243
g4903 nand P2_R1275_U22 P2_U3027 ; P2_U4244
g4904 nand P2_U3026 P2_U3072 ; P2_U4245
g4905 nand P2_R1215_U99 P2_U3025 ; P2_U4246
g4906 nand P2_U3447 P2_U4116 ; P2_U4247
g4907 nand P2_U3601 P2_U4243 ; P2_U4248
g4908 nand P2_U3020 P2_REG2_REG_8__SCAN_IN ; P2_U4249
g4909 nand P2_U3021 P2_REG1_REG_8__SCAN_IN ; P2_U4250
g4910 nand P2_U3022 P2_REG0_REG_8__SCAN_IN ; P2_U4251
g4911 nand P2_ADD_1119_U51 P2_U3019 ; P2_U4252
g4912 not P2_U3086 ; P2_U4253
g4913 nand P2_U3035 P2_U3073 ; P2_U4254
g4914 nand P2_R1146_U104 P2_U3931 ; P2_U4255
g4915 nand P2_R1113_U104 P2_U3930 ; P2_U4256
g4916 nand P2_R1131_U18 P2_U3926 ; P2_U4257
g4917 nand P2_R1179_U104 P2_U3941 ; P2_U4258
g4918 nand P2_R1203_U104 P2_U3943 ; P2_U4259
g4919 nand P2_R1164_U18 P2_U3014 ; P2_U4260
g4920 nand P2_R1233_U18 P2_U3922 ; P2_U4261
g4921 not P2_U3355 ; P2_U4262
g4922 nand P2_R1275_U23 P2_U3027 ; P2_U4263
g4923 nand P2_U3026 P2_U3086 ; P2_U4264
g4924 nand P2_R1215_U19 P2_U3025 ; P2_U4265
g4925 nand P2_U3450 P2_U4116 ; P2_U4266
g4926 nand P2_U3605 P2_U4262 ; P2_U4267
g4927 nand P2_U3020 P2_REG2_REG_9__SCAN_IN ; P2_U4268
g4928 nand P2_U3021 P2_REG1_REG_9__SCAN_IN ; P2_U4269
g4929 nand P2_U3022 P2_REG0_REG_9__SCAN_IN ; P2_U4270
g4930 nand P2_ADD_1119_U50 P2_U3019 ; P2_U4271
g4931 not P2_U3085 ; P2_U4272
g4932 nand P2_U3035 P2_U3072 ; P2_U4273
g4933 nand P2_R1146_U19 P2_U3931 ; P2_U4274
g4934 nand P2_R1113_U19 P2_U3930 ; P2_U4275
g4935 nand P2_R1131_U97 P2_U3926 ; P2_U4276
g4936 nand P2_R1179_U19 P2_U3941 ; P2_U4277
g4937 nand P2_R1203_U19 P2_U3943 ; P2_U4278
g4938 nand P2_R1164_U97 P2_U3014 ; P2_U4279
g4939 nand P2_R1233_U97 P2_U3922 ; P2_U4280
g4940 not P2_U3356 ; P2_U4281
g4941 nand P2_R1275_U24 P2_U3027 ; P2_U4282
g4942 nand P2_U3026 P2_U3085 ; P2_U4283
g4943 nand P2_R1215_U98 P2_U3025 ; P2_U4284
g4944 nand P2_U3453 P2_U4116 ; P2_U4285
g4945 nand P2_U3609 P2_U4281 ; P2_U4286
g4946 nand P2_U3020 P2_REG2_REG_10__SCAN_IN ; P2_U4287
g4947 nand P2_U3021 P2_REG1_REG_10__SCAN_IN ; P2_U4288
g4948 nand P2_U3022 P2_REG0_REG_10__SCAN_IN ; P2_U4289
g4949 nand P2_ADD_1119_U74 P2_U3019 ; P2_U4290
g4950 not P2_U3064 ; P2_U4291
g4951 nand P2_U3035 P2_U3086 ; P2_U4292
g4952 nand P2_R1146_U103 P2_U3931 ; P2_U4293
g4953 nand P2_R1113_U103 P2_U3930 ; P2_U4294
g4954 nand P2_R1131_U96 P2_U3926 ; P2_U4295
g4955 nand P2_R1179_U103 P2_U3941 ; P2_U4296
g4956 nand P2_R1203_U103 P2_U3943 ; P2_U4297
g4957 nand P2_R1164_U96 P2_U3014 ; P2_U4298
g4958 nand P2_R1233_U96 P2_U3922 ; P2_U4299
g4959 not P2_U3357 ; P2_U4300
g4960 nand P2_R1275_U63 P2_U3027 ; P2_U4301
g4961 nand P2_U3026 P2_U3064 ; P2_U4302
g4962 nand P2_R1215_U97 P2_U3025 ; P2_U4303
g4963 nand P2_U3456 P2_U4116 ; P2_U4304
g4964 nand P2_U3613 P2_U4300 ; P2_U4305
g4965 nand P2_U3020 P2_REG2_REG_11__SCAN_IN ; P2_U4306
g4966 nand P2_U3021 P2_REG1_REG_11__SCAN_IN ; P2_U4307
g4967 nand P2_U3022 P2_REG0_REG_11__SCAN_IN ; P2_U4308
g4968 nand P2_ADD_1119_U73 P2_U3019 ; P2_U4309
g4969 not P2_U3065 ; P2_U4310
g4970 nand P2_U3035 P2_U3085 ; P2_U4311
g4971 nand P2_R1146_U113 P2_U3931 ; P2_U4312
g4972 nand P2_R1113_U113 P2_U3930 ; P2_U4313
g4973 nand P2_R1131_U10 P2_U3926 ; P2_U4314
g4974 nand P2_R1179_U113 P2_U3941 ; P2_U4315
g4975 nand P2_R1203_U113 P2_U3943 ; P2_U4316
g4976 nand P2_R1164_U10 P2_U3014 ; P2_U4317
g4977 nand P2_R1233_U10 P2_U3922 ; P2_U4318
g4978 not P2_U3358 ; P2_U4319
g4979 nand P2_R1275_U6 P2_U3027 ; P2_U4320
g4980 nand P2_U3026 P2_U3065 ; P2_U4321
g4981 nand P2_R1215_U11 P2_U3025 ; P2_U4322
g4982 nand P2_U3459 P2_U4116 ; P2_U4323
g4983 nand P2_U3617 P2_U4319 ; P2_U4324
g4984 nand P2_U3020 P2_REG2_REG_12__SCAN_IN ; P2_U4325
g4985 nand P2_U3021 P2_REG1_REG_12__SCAN_IN ; P2_U4326
g4986 nand P2_U3022 P2_REG0_REG_12__SCAN_IN ; P2_U4327
g4987 nand P2_ADD_1119_U72 P2_U3019 ; P2_U4328
g4988 not P2_U3074 ; P2_U4329
g4989 nand P2_U3035 P2_U3064 ; P2_U4330
g4990 nand P2_R1146_U12 P2_U3931 ; P2_U4331
g4991 nand P2_R1113_U12 P2_U3930 ; P2_U4332
g4992 nand P2_R1131_U114 P2_U3926 ; P2_U4333
g4993 nand P2_R1179_U12 P2_U3941 ; P2_U4334
g4994 nand P2_R1203_U12 P2_U3943 ; P2_U4335
g4995 nand P2_R1164_U114 P2_U3014 ; P2_U4336
g4996 nand P2_R1233_U114 P2_U3922 ; P2_U4337
g4997 not P2_U3359 ; P2_U4338
g4998 nand P2_R1275_U7 P2_U3027 ; P2_U4339
g4999 nand P2_U3026 P2_U3074 ; P2_U4340
g5000 nand P2_R1215_U115 P2_U3025 ; P2_U4341
g5001 nand P2_U3462 P2_U4116 ; P2_U4342
g5002 nand P2_U3621 P2_U4338 ; P2_U4343
g5003 nand P2_U3020 P2_REG2_REG_13__SCAN_IN ; P2_U4344
g5004 nand P2_U3021 P2_REG1_REG_13__SCAN_IN ; P2_U4345
g5005 nand P2_U3022 P2_REG0_REG_13__SCAN_IN ; P2_U4346
g5006 nand P2_ADD_1119_U71 P2_U3019 ; P2_U4347
g5007 not P2_U3082 ; P2_U4348
g5008 nand P2_U3035 P2_U3065 ; P2_U4349
g5009 nand P2_R1146_U102 P2_U3931 ; P2_U4350
g5010 nand P2_R1113_U102 P2_U3930 ; P2_U4351
g5011 nand P2_R1131_U113 P2_U3926 ; P2_U4352
g5012 nand P2_R1179_U102 P2_U3941 ; P2_U4353
g5013 nand P2_R1203_U102 P2_U3943 ; P2_U4354
g5014 nand P2_R1164_U113 P2_U3014 ; P2_U4355
g5015 nand P2_R1233_U113 P2_U3922 ; P2_U4356
g5016 not P2_U3360 ; P2_U4357
g5017 nand P2_R1275_U8 P2_U3027 ; P2_U4358
g5018 nand P2_U3026 P2_U3082 ; P2_U4359
g5019 nand P2_R1215_U114 P2_U3025 ; P2_U4360
g5020 nand P2_U3465 P2_U4116 ; P2_U4361
g5021 nand P2_U3625 P2_U4357 ; P2_U4362
g5022 nand P2_U3020 P2_REG2_REG_14__SCAN_IN ; P2_U4363
g5023 nand P2_U3021 P2_REG1_REG_14__SCAN_IN ; P2_U4364
g5024 nand P2_U3022 P2_REG0_REG_14__SCAN_IN ; P2_U4365
g5025 nand P2_ADD_1119_U70 P2_U3019 ; P2_U4366
g5026 not P2_U3081 ; P2_U4367
g5027 nand P2_U3035 P2_U3074 ; P2_U4368
g5028 nand P2_R1146_U101 P2_U3931 ; P2_U4369
g5029 nand P2_R1113_U101 P2_U3930 ; P2_U4370
g5030 nand P2_R1131_U11 P2_U3926 ; P2_U4371
g5031 nand P2_R1179_U101 P2_U3941 ; P2_U4372
g5032 nand P2_R1203_U101 P2_U3943 ; P2_U4373
g5033 nand P2_R1164_U11 P2_U3014 ; P2_U4374
g5034 nand P2_R1233_U11 P2_U3922 ; P2_U4375
g5035 not P2_U3361 ; P2_U4376
g5036 nand P2_R1275_U86 P2_U3027 ; P2_U4377
g5037 nand P2_U3026 P2_U3081 ; P2_U4378
g5038 nand P2_R1215_U12 P2_U3025 ; P2_U4379
g5039 nand P2_U3468 P2_U4116 ; P2_U4380
g5040 nand P2_U3629 P2_U4376 ; P2_U4381
g5041 nand P2_U3020 P2_REG2_REG_15__SCAN_IN ; P2_U4382
g5042 nand P2_U3021 P2_REG1_REG_15__SCAN_IN ; P2_U4383
g5043 nand P2_U3022 P2_REG0_REG_15__SCAN_IN ; P2_U4384
g5044 nand P2_ADD_1119_U69 P2_U3019 ; P2_U4385
g5045 not P2_U3076 ; P2_U4386
g5046 nand P2_U3035 P2_U3082 ; P2_U4387
g5047 nand P2_R1146_U112 P2_U3931 ; P2_U4388
g5048 nand P2_R1113_U112 P2_U3930 ; P2_U4389
g5049 nand P2_R1131_U112 P2_U3926 ; P2_U4390
g5050 nand P2_R1179_U112 P2_U3941 ; P2_U4391
g5051 nand P2_R1203_U112 P2_U3943 ; P2_U4392
g5052 nand P2_R1164_U112 P2_U3014 ; P2_U4393
g5053 nand P2_R1233_U112 P2_U3922 ; P2_U4394
g5054 not P2_U3362 ; P2_U4395
g5055 nand P2_R1275_U9 P2_U3027 ; P2_U4396
g5056 nand P2_U3026 P2_U3076 ; P2_U4397
g5057 nand P2_R1215_U113 P2_U3025 ; P2_U4398
g5058 nand P2_U3471 P2_U4116 ; P2_U4399
g5059 nand P2_U3633 P2_U4395 ; P2_U4400
g5060 nand P2_U3020 P2_REG2_REG_16__SCAN_IN ; P2_U4401
g5061 nand P2_U3021 P2_REG1_REG_16__SCAN_IN ; P2_U4402
g5062 nand P2_U3022 P2_REG0_REG_16__SCAN_IN ; P2_U4403
g5063 nand P2_ADD_1119_U68 P2_U3019 ; P2_U4404
g5064 not P2_U3075 ; P2_U4405
g5065 nand P2_U3035 P2_U3081 ; P2_U4406
g5066 nand P2_R1146_U111 P2_U3931 ; P2_U4407
g5067 nand P2_R1113_U111 P2_U3930 ; P2_U4408
g5068 nand P2_R1131_U111 P2_U3926 ; P2_U4409
g5069 nand P2_R1179_U111 P2_U3941 ; P2_U4410
g5070 nand P2_R1203_U111 P2_U3943 ; P2_U4411
g5071 nand P2_R1164_U111 P2_U3014 ; P2_U4412
g5072 nand P2_R1233_U111 P2_U3922 ; P2_U4413
g5073 not P2_U3363 ; P2_U4414
g5074 nand P2_R1275_U10 P2_U3027 ; P2_U4415
g5075 nand P2_U3026 P2_U3075 ; P2_U4416
g5076 nand P2_R1215_U112 P2_U3025 ; P2_U4417
g5077 nand P2_U3474 P2_U4116 ; P2_U4418
g5078 nand P2_U3637 P2_U4414 ; P2_U4419
g5079 nand P2_U3020 P2_REG2_REG_17__SCAN_IN ; P2_U4420
g5080 nand P2_U3021 P2_REG1_REG_17__SCAN_IN ; P2_U4421
g5081 nand P2_U3022 P2_REG0_REG_17__SCAN_IN ; P2_U4422
g5082 nand P2_ADD_1119_U67 P2_U3019 ; P2_U4423
g5083 not P2_U3071 ; P2_U4424
g5084 nand P2_U3035 P2_U3076 ; P2_U4425
g5085 nand P2_R1146_U13 P2_U3931 ; P2_U4426
g5086 nand P2_R1113_U13 P2_U3930 ; P2_U4427
g5087 nand P2_R1131_U110 P2_U3926 ; P2_U4428
g5088 nand P2_R1179_U13 P2_U3941 ; P2_U4429
g5089 nand P2_R1203_U13 P2_U3943 ; P2_U4430
g5090 nand P2_R1164_U110 P2_U3014 ; P2_U4431
g5091 nand P2_R1233_U110 P2_U3922 ; P2_U4432
g5092 not P2_U3364 ; P2_U4433
g5093 nand P2_R1275_U11 P2_U3027 ; P2_U4434
g5094 nand P2_U3026 P2_U3071 ; P2_U4435
g5095 nand P2_R1215_U111 P2_U3025 ; P2_U4436
g5096 nand P2_U3477 P2_U4116 ; P2_U4437
g5097 nand P2_U3641 P2_U4433 ; P2_U4438
g5098 nand P2_U3020 P2_REG2_REG_18__SCAN_IN ; P2_U4439
g5099 nand P2_U3021 P2_REG1_REG_18__SCAN_IN ; P2_U4440
g5100 nand P2_U3022 P2_REG0_REG_18__SCAN_IN ; P2_U4441
g5101 nand P2_ADD_1119_U66 P2_U3019 ; P2_U4442
g5102 not P2_U3084 ; P2_U4443
g5103 nand P2_U3035 P2_U3075 ; P2_U4444
g5104 nand P2_R1146_U100 P2_U3931 ; P2_U4445
g5105 nand P2_R1113_U100 P2_U3930 ; P2_U4446
g5106 nand P2_R1131_U12 P2_U3926 ; P2_U4447
g5107 nand P2_R1179_U100 P2_U3941 ; P2_U4448
g5108 nand P2_R1203_U100 P2_U3943 ; P2_U4449
g5109 nand P2_R1164_U12 P2_U3014 ; P2_U4450
g5110 nand P2_R1233_U12 P2_U3922 ; P2_U4451
g5111 not P2_U3365 ; P2_U4452
g5112 nand P2_R1275_U84 P2_U3027 ; P2_U4453
g5113 nand P2_U3026 P2_U3084 ; P2_U4454
g5114 nand P2_R1215_U13 P2_U3025 ; P2_U4455
g5115 nand P2_U3480 P2_U4116 ; P2_U4456
g5116 nand P2_U3645 P2_U4452 ; P2_U4457
g5117 nand P2_U3020 P2_REG2_REG_19__SCAN_IN ; P2_U4458
g5118 nand P2_U3021 P2_REG1_REG_19__SCAN_IN ; P2_U4459
g5119 nand P2_U3022 P2_REG0_REG_19__SCAN_IN ; P2_U4460
g5120 nand P2_ADD_1119_U65 P2_U3019 ; P2_U4461
g5121 not P2_U3083 ; P2_U4462
g5122 nand P2_U3035 P2_U3071 ; P2_U4463
g5123 nand P2_R1146_U99 P2_U3931 ; P2_U4464
g5124 nand P2_R1113_U99 P2_U3930 ; P2_U4465
g5125 nand P2_R1131_U109 P2_U3926 ; P2_U4466
g5126 nand P2_R1179_U99 P2_U3941 ; P2_U4467
g5127 nand P2_R1203_U99 P2_U3943 ; P2_U4468
g5128 nand P2_R1164_U109 P2_U3014 ; P2_U4469
g5129 nand P2_R1233_U109 P2_U3922 ; P2_U4470
g5130 not P2_U3366 ; P2_U4471
g5131 nand P2_R1275_U12 P2_U3027 ; P2_U4472
g5132 nand P2_U3026 P2_U3083 ; P2_U4473
g5133 nand P2_R1215_U110 P2_U3025 ; P2_U4474
g5134 nand P2_U3483 P2_U4116 ; P2_U4475
g5135 nand P2_U3649 P2_U4471 ; P2_U4476
g5136 nand P2_U3020 P2_REG2_REG_20__SCAN_IN ; P2_U4477
g5137 nand P2_U3021 P2_REG1_REG_20__SCAN_IN ; P2_U4478
g5138 nand P2_U3022 P2_REG0_REG_20__SCAN_IN ; P2_U4479
g5139 nand P2_ADD_1119_U64 P2_U3019 ; P2_U4480
g5140 not P2_U3078 ; P2_U4481
g5141 nand P2_U3035 P2_U3084 ; P2_U4482
g5142 nand P2_R1146_U98 P2_U3931 ; P2_U4483
g5143 nand P2_R1113_U98 P2_U3930 ; P2_U4484
g5144 nand P2_R1131_U108 P2_U3926 ; P2_U4485
g5145 nand P2_R1179_U98 P2_U3941 ; P2_U4486
g5146 nand P2_R1203_U98 P2_U3943 ; P2_U4487
g5147 nand P2_R1164_U108 P2_U3014 ; P2_U4488
g5148 nand P2_R1233_U108 P2_U3922 ; P2_U4489
g5149 not P2_U3367 ; P2_U4490
g5150 nand P2_R1275_U82 P2_U3027 ; P2_U4491
g5151 nand P2_U3026 P2_U3078 ; P2_U4492
g5152 nand P2_R1215_U109 P2_U3025 ; P2_U4493
g5153 nand P2_U3485 P2_U4116 ; P2_U4494
g5154 nand P2_U3653 P2_U4490 ; P2_U4495
g5155 nand P2_U3020 P2_REG2_REG_21__SCAN_IN ; P2_U4496
g5156 nand P2_U3021 P2_REG1_REG_21__SCAN_IN ; P2_U4497
g5157 nand P2_U3022 P2_REG0_REG_21__SCAN_IN ; P2_U4498
g5158 nand P2_ADD_1119_U63 P2_U3019 ; P2_U4499
g5159 not P2_U3077 ; P2_U4500
g5160 nand P2_U3035 P2_U3083 ; P2_U4501
g5161 nand P2_R1146_U96 P2_U3931 ; P2_U4502
g5162 nand P2_R1113_U96 P2_U3930 ; P2_U4503
g5163 nand P2_R1131_U13 P2_U3926 ; P2_U4504
g5164 nand P2_R1179_U96 P2_U3941 ; P2_U4505
g5165 nand P2_R1203_U96 P2_U3943 ; P2_U4506
g5166 nand P2_R1164_U13 P2_U3014 ; P2_U4507
g5167 nand P2_R1233_U13 P2_U3922 ; P2_U4508
g5168 not P2_U3369 ; P2_U4509
g5169 nand P2_R1275_U13 P2_U3027 ; P2_U4510
g5170 nand P2_U3026 P2_U3077 ; P2_U4511
g5171 nand P2_R1215_U14 P2_U3025 ; P2_U4512
g5172 nand P2_U3957 P2_U4116 ; P2_U4513
g5173 nand P2_U3657 P2_U4509 ; P2_U4514
g5174 nand P2_U3020 P2_REG2_REG_22__SCAN_IN ; P2_U4515
g5175 nand P2_U3021 P2_REG1_REG_22__SCAN_IN ; P2_U4516
g5176 nand P2_U3022 P2_REG0_REG_22__SCAN_IN ; P2_U4517
g5177 nand P2_ADD_1119_U62 P2_U3019 ; P2_U4518
g5178 not P2_U3063 ; P2_U4519
g5179 nand P2_U3035 P2_U3078 ; P2_U4520
g5180 nand P2_R1146_U110 P2_U3931 ; P2_U4521
g5181 nand P2_R1113_U110 P2_U3930 ; P2_U4522
g5182 nand P2_R1131_U14 P2_U3926 ; P2_U4523
g5183 nand P2_R1179_U110 P2_U3941 ; P2_U4524
g5184 nand P2_R1203_U110 P2_U3943 ; P2_U4525
g5185 nand P2_R1164_U14 P2_U3014 ; P2_U4526
g5186 nand P2_R1233_U14 P2_U3922 ; P2_U4527
g5187 not P2_U3371 ; P2_U4528
g5188 nand P2_R1275_U78 P2_U3027 ; P2_U4529
g5189 nand P2_U3026 P2_U3063 ; P2_U4530
g5190 nand P2_R1215_U15 P2_U3025 ; P2_U4531
g5191 nand P2_U3956 P2_U4116 ; P2_U4532
g5192 nand P2_U3661 P2_U4528 ; P2_U4533
g5193 nand P2_U3020 P2_REG2_REG_23__SCAN_IN ; P2_U4534
g5194 nand P2_U3021 P2_REG1_REG_23__SCAN_IN ; P2_U4535
g5195 nand P2_U3022 P2_REG0_REG_23__SCAN_IN ; P2_U4536
g5196 nand P2_ADD_1119_U61 P2_U3019 ; P2_U4537
g5197 not P2_U3068 ; P2_U4538
g5198 nand P2_U3035 P2_U3077 ; P2_U4539
g5199 nand P2_R1146_U109 P2_U3931 ; P2_U4540
g5200 nand P2_R1113_U109 P2_U3930 ; P2_U4541
g5201 nand P2_R1131_U107 P2_U3926 ; P2_U4542
g5202 nand P2_R1179_U109 P2_U3941 ; P2_U4543
g5203 nand P2_R1203_U109 P2_U3943 ; P2_U4544
g5204 nand P2_R1164_U107 P2_U3014 ; P2_U4545
g5205 nand P2_R1233_U107 P2_U3922 ; P2_U4546
g5206 not P2_U3373 ; P2_U4547
g5207 nand P2_R1275_U14 P2_U3027 ; P2_U4548
g5208 nand P2_U3026 P2_U3068 ; P2_U4549
g5209 nand P2_R1215_U108 P2_U3025 ; P2_U4550
g5210 nand P2_U3955 P2_U4116 ; P2_U4551
g5211 nand P2_U3665 P2_U4547 ; P2_U4552
g5212 nand P2_U3020 P2_REG2_REG_24__SCAN_IN ; P2_U4553
g5213 nand P2_U3021 P2_REG1_REG_24__SCAN_IN ; P2_U4554
g5214 nand P2_U3022 P2_REG0_REG_24__SCAN_IN ; P2_U4555
g5215 nand P2_ADD_1119_U60 P2_U3019 ; P2_U4556
g5216 not P2_U3067 ; P2_U4557
g5217 nand P2_U3035 P2_U3063 ; P2_U4558
g5218 nand P2_R1146_U14 P2_U3931 ; P2_U4559
g5219 nand P2_R1113_U14 P2_U3930 ; P2_U4560
g5220 nand P2_R1131_U106 P2_U3926 ; P2_U4561
g5221 nand P2_R1179_U14 P2_U3941 ; P2_U4562
g5222 nand P2_R1203_U14 P2_U3943 ; P2_U4563
g5223 nand P2_R1164_U106 P2_U3014 ; P2_U4564
g5224 nand P2_R1233_U106 P2_U3922 ; P2_U4565
g5225 not P2_U3375 ; P2_U4566
g5226 nand P2_R1275_U76 P2_U3027 ; P2_U4567
g5227 nand P2_U3026 P2_U3067 ; P2_U4568
g5228 nand P2_R1215_U107 P2_U3025 ; P2_U4569
g5229 nand P2_U3954 P2_U4116 ; P2_U4570
g5230 nand P2_U3669 P2_U4566 ; P2_U4571
g5231 nand P2_U3020 P2_REG2_REG_25__SCAN_IN ; P2_U4572
g5232 nand P2_U3021 P2_REG1_REG_25__SCAN_IN ; P2_U4573
g5233 nand P2_U3022 P2_REG0_REG_25__SCAN_IN ; P2_U4574
g5234 nand P2_ADD_1119_U59 P2_U3019 ; P2_U4575
g5235 not P2_U3060 ; P2_U4576
g5236 nand P2_U3035 P2_U3068 ; P2_U4577
g5237 nand P2_R1146_U95 P2_U3931 ; P2_U4578
g5238 nand P2_R1113_U95 P2_U3930 ; P2_U4579
g5239 nand P2_R1131_U105 P2_U3926 ; P2_U4580
g5240 nand P2_R1179_U95 P2_U3941 ; P2_U4581
g5241 nand P2_R1203_U95 P2_U3943 ; P2_U4582
g5242 nand P2_R1164_U105 P2_U3014 ; P2_U4583
g5243 nand P2_R1233_U105 P2_U3922 ; P2_U4584
g5244 not P2_U3377 ; P2_U4585
g5245 nand P2_R1275_U15 P2_U3027 ; P2_U4586
g5246 nand P2_U3026 P2_U3060 ; P2_U4587
g5247 nand P2_R1215_U106 P2_U3025 ; P2_U4588
g5248 nand P2_U3953 P2_U4116 ; P2_U4589
g5249 nand P2_U3673 P2_U4585 ; P2_U4590
g5250 nand P2_U3020 P2_REG2_REG_26__SCAN_IN ; P2_U4591
g5251 nand P2_U3021 P2_REG1_REG_26__SCAN_IN ; P2_U4592
g5252 nand P2_U3022 P2_REG0_REG_26__SCAN_IN ; P2_U4593
g5253 nand P2_ADD_1119_U58 P2_U3019 ; P2_U4594
g5254 not P2_U3059 ; P2_U4595
g5255 nand P2_U3035 P2_U3067 ; P2_U4596
g5256 nand P2_R1146_U94 P2_U3931 ; P2_U4597
g5257 nand P2_R1113_U94 P2_U3930 ; P2_U4598
g5258 nand P2_R1131_U104 P2_U3926 ; P2_U4599
g5259 nand P2_R1179_U94 P2_U3941 ; P2_U4600
g5260 nand P2_R1203_U94 P2_U3943 ; P2_U4601
g5261 nand P2_R1164_U104 P2_U3014 ; P2_U4602
g5262 nand P2_R1233_U104 P2_U3922 ; P2_U4603
g5263 not P2_U3379 ; P2_U4604
g5264 nand P2_R1275_U74 P2_U3027 ; P2_U4605
g5265 nand P2_U3026 P2_U3059 ; P2_U4606
g5266 nand P2_R1215_U105 P2_U3025 ; P2_U4607
g5267 nand P2_U3952 P2_U4116 ; P2_U4608
g5268 nand P2_U3677 P2_U4604 ; P2_U4609
g5269 nand P2_U3020 P2_REG2_REG_27__SCAN_IN ; P2_U4610
g5270 nand P2_U3021 P2_REG1_REG_27__SCAN_IN ; P2_U4611
g5271 nand P2_U3022 P2_REG0_REG_27__SCAN_IN ; P2_U4612
g5272 nand P2_ADD_1119_U57 P2_U3019 ; P2_U4613
g5273 not P2_U3055 ; P2_U4614
g5274 nand P2_U3035 P2_U3060 ; P2_U4615
g5275 nand P2_R1146_U108 P2_U3931 ; P2_U4616
g5276 nand P2_R1113_U108 P2_U3930 ; P2_U4617
g5277 nand P2_R1131_U15 P2_U3926 ; P2_U4618
g5278 nand P2_R1179_U108 P2_U3941 ; P2_U4619
g5279 nand P2_R1203_U108 P2_U3943 ; P2_U4620
g5280 nand P2_R1164_U15 P2_U3014 ; P2_U4621
g5281 nand P2_R1233_U15 P2_U3922 ; P2_U4622
g5282 not P2_U3381 ; P2_U4623
g5283 nand P2_R1275_U16 P2_U3027 ; P2_U4624
g5284 nand P2_U3026 P2_U3055 ; P2_U4625
g5285 nand P2_R1215_U16 P2_U3025 ; P2_U4626
g5286 nand P2_U3951 P2_U4116 ; P2_U4627
g5287 nand P2_U3681 P2_U4623 ; P2_U4628
g5288 nand P2_U3020 P2_REG2_REG_28__SCAN_IN ; P2_U4629
g5289 nand P2_U3021 P2_REG1_REG_28__SCAN_IN ; P2_U4630
g5290 nand P2_U3022 P2_REG0_REG_28__SCAN_IN ; P2_U4631
g5291 nand P2_ADD_1119_U56 P2_U3019 ; P2_U4632
g5292 not P2_U3056 ; P2_U4633
g5293 nand P2_U3035 P2_U3059 ; P2_U4634
g5294 nand P2_R1146_U15 P2_U3931 ; P2_U4635
g5295 nand P2_R1113_U15 P2_U3930 ; P2_U4636
g5296 nand P2_R1131_U103 P2_U3926 ; P2_U4637
g5297 nand P2_R1179_U15 P2_U3941 ; P2_U4638
g5298 nand P2_R1203_U15 P2_U3943 ; P2_U4639
g5299 nand P2_R1164_U103 P2_U3014 ; P2_U4640
g5300 nand P2_R1233_U103 P2_U3922 ; P2_U4641
g5301 not P2_U3383 ; P2_U4642
g5302 nand P2_R1275_U72 P2_U3027 ; P2_U4643
g5303 nand P2_U3026 P2_U3056 ; P2_U4644
g5304 nand P2_R1215_U104 P2_U3025 ; P2_U4645
g5305 nand P2_U3950 P2_U4116 ; P2_U4646
g5306 nand P2_U3685 P2_U4642 ; P2_U4647
g5307 nand P2_ADD_1119_U5 P2_U3019 ; P2_U4648
g5308 nand P2_U3020 P2_REG2_REG_29__SCAN_IN ; P2_U4649
g5309 nand P2_U3021 P2_REG1_REG_29__SCAN_IN ; P2_U4650
g5310 nand P2_U3022 P2_REG0_REG_29__SCAN_IN ; P2_U4651
g5311 not P2_U3057 ; P2_U4652
g5312 nand P2_U3035 P2_U3055 ; P2_U4653
g5313 nand P2_R1146_U93 P2_U3931 ; P2_U4654
g5314 nand P2_R1113_U93 P2_U3930 ; P2_U4655
g5315 nand P2_R1131_U102 P2_U3926 ; P2_U4656
g5316 nand P2_R1179_U93 P2_U3941 ; P2_U4657
g5317 nand P2_R1203_U93 P2_U3943 ; P2_U4658
g5318 nand P2_R1164_U102 P2_U3014 ; P2_U4659
g5319 nand P2_R1233_U102 P2_U3922 ; P2_U4660
g5320 not P2_U3385 ; P2_U4661
g5321 nand P2_R1275_U17 P2_U3027 ; P2_U4662
g5322 nand P2_U3026 P2_U3057 ; P2_U4663
g5323 nand P2_R1215_U103 P2_U3025 ; P2_U4664
g5324 nand P2_U3949 P2_U4116 ; P2_U4665
g5325 nand P2_U3688 P2_U4661 ; P2_U4666
g5326 nand P2_U3020 P2_REG2_REG_30__SCAN_IN ; P2_U4667
g5327 nand P2_U3021 P2_REG1_REG_30__SCAN_IN ; P2_U4668
g5328 nand P2_U3022 P2_REG0_REG_30__SCAN_IN ; P2_U4669
g5329 not P2_U3061 ; P2_U4670
g5330 nand P2_U5683 P2_U3331 ; P2_U4671
g5331 nand P2_U3347 P2_U4671 ; P2_U4672
g5332 nand P2_U3689 P2_U3061 ; P2_U4673
g5333 nand P2_U3035 P2_U3056 ; P2_U4674
g5334 nand P2_R1146_U16 P2_U3931 ; P2_U4675
g5335 nand P2_R1113_U16 P2_U3930 ; P2_U4676
g5336 nand P2_R1131_U101 P2_U3926 ; P2_U4677
g5337 nand P2_R1179_U16 P2_U3941 ; P2_U4678
g5338 nand P2_R1203_U16 P2_U3943 ; P2_U4679
g5339 nand P2_R1164_U101 P2_U3014 ; P2_U4680
g5340 nand P2_R1233_U101 P2_U3922 ; P2_U4681
g5341 not P2_U3387 ; P2_U4682
g5342 nand P2_R1275_U70 P2_U3027 ; P2_U4683
g5343 nand P2_R1215_U102 P2_U3025 ; P2_U4684
g5344 nand P2_U3960 P2_U4116 ; P2_U4685
g5345 nand P2_U3693 P2_U4682 ; P2_U4686
g5346 nand P2_U3020 P2_REG2_REG_31__SCAN_IN ; P2_U4687
g5347 nand P2_U3021 P2_REG1_REG_31__SCAN_IN ; P2_U4688
g5348 nand P2_U3022 P2_REG0_REG_31__SCAN_IN ; P2_U4689
g5349 not P2_U3058 ; P2_U4690
g5350 nand P2_R1275_U19 P2_U3027 ; P2_U4691
g5351 nand P2_U3959 P2_U4116 ; P2_U4692
g5352 nand P2_U4692 P2_U3913 P2_U4691 ; P2_U4693
g5353 nand P2_R1275_U68 P2_U3027 ; P2_U4694
g5354 nand P2_U3958 P2_U4116 ; P2_U4695
g5355 nand P2_U4695 P2_U3913 P2_U4694 ; P2_U4696
g5356 nand P2_U3696 P2_U3016 ; P2_U4697
g5357 nand P2_U3393 P2_U4697 ; P2_U4698
g5358 nand P2_U3921 P2_U3418 ; P2_U4699
g5359 not P2_U3398 ; P2_U4700
g5360 nand P2_U3037 P2_U3080 ; P2_U4701
g5361 nand P2_U3034 P2_R1215_U96 ; P2_U4702
g5362 nand P2_U3033 P2_REG3_REG_0__SCAN_IN ; P2_U4703
g5363 nand P2_U3032 P2_U3427 ; P2_U4704
g5364 nand P2_U3031 P2_U3427 ; P2_U4705
g5365 nand P2_U3037 P2_U3070 ; P2_U4706
g5366 nand P2_U3034 P2_R1215_U95 ; P2_U4707
g5367 nand P2_U3033 P2_REG3_REG_1__SCAN_IN ; P2_U4708
g5368 nand P2_U3032 P2_U3432 ; P2_U4709
g5369 nand P2_U3031 P2_R1275_U55 ; P2_U4710
g5370 nand P2_U3037 P2_U3066 ; P2_U4711
g5371 nand P2_U3034 P2_R1215_U17 ; P2_U4712
g5372 nand P2_U3033 P2_REG3_REG_2__SCAN_IN ; P2_U4713
g5373 nand P2_U3032 P2_U3435 ; P2_U4714
g5374 nand P2_U3031 P2_R1275_U18 ; P2_U4715
g5375 nand P2_U3037 P2_U3062 ; P2_U4716
g5376 nand P2_U3034 P2_R1215_U101 ; P2_U4717
g5377 nand P2_U3033 P2_ADD_1119_U4 ; P2_U4718
g5378 nand P2_U3032 P2_U3438 ; P2_U4719
g5379 nand P2_U3031 P2_R1275_U20 ; P2_U4720
g5380 nand P2_U3037 P2_U3069 ; P2_U4721
g5381 nand P2_U3034 P2_R1215_U100 ; P2_U4722
g5382 nand P2_U3033 P2_ADD_1119_U55 ; P2_U4723
g5383 nand P2_U3032 P2_U3441 ; P2_U4724
g5384 nand P2_U3031 P2_R1275_U21 ; P2_U4725
g5385 nand P2_U3037 P2_U3073 ; P2_U4726
g5386 nand P2_U3034 P2_R1215_U18 ; P2_U4727
g5387 nand P2_U3033 P2_ADD_1119_U54 ; P2_U4728
g5388 nand P2_U3032 P2_U3444 ; P2_U4729
g5389 nand P2_U3031 P2_R1275_U65 ; P2_U4730
g5390 nand P2_U3037 P2_U3072 ; P2_U4731
g5391 nand P2_U3034 P2_R1215_U99 ; P2_U4732
g5392 nand P2_U3033 P2_ADD_1119_U53 ; P2_U4733
g5393 nand P2_U3032 P2_U3447 ; P2_U4734
g5394 nand P2_U3031 P2_R1275_U22 ; P2_U4735
g5395 nand P2_U3037 P2_U3086 ; P2_U4736
g5396 nand P2_U3034 P2_R1215_U19 ; P2_U4737
g5397 nand P2_U3033 P2_ADD_1119_U52 ; P2_U4738
g5398 nand P2_U3032 P2_U3450 ; P2_U4739
g5399 nand P2_U3031 P2_R1275_U23 ; P2_U4740
g5400 nand P2_U3037 P2_U3085 ; P2_U4741
g5401 nand P2_U3034 P2_R1215_U98 ; P2_U4742
g5402 nand P2_U3033 P2_ADD_1119_U51 ; P2_U4743
g5403 nand P2_U3032 P2_U3453 ; P2_U4744
g5404 nand P2_U3031 P2_R1275_U24 ; P2_U4745
g5405 nand P2_U3037 P2_U3064 ; P2_U4746
g5406 nand P2_U3034 P2_R1215_U97 ; P2_U4747
g5407 nand P2_U3033 P2_ADD_1119_U50 ; P2_U4748
g5408 nand P2_U3032 P2_U3456 ; P2_U4749
g5409 nand P2_U3031 P2_R1275_U63 ; P2_U4750
g5410 nand P2_U3037 P2_U3065 ; P2_U4751
g5411 nand P2_U3034 P2_R1215_U11 ; P2_U4752
g5412 nand P2_U3033 P2_ADD_1119_U74 ; P2_U4753
g5413 nand P2_U3032 P2_U3459 ; P2_U4754
g5414 nand P2_U3031 P2_R1275_U6 ; P2_U4755
g5415 nand P2_U3037 P2_U3074 ; P2_U4756
g5416 nand P2_U3034 P2_R1215_U115 ; P2_U4757
g5417 nand P2_U3033 P2_ADD_1119_U73 ; P2_U4758
g5418 nand P2_U3032 P2_U3462 ; P2_U4759
g5419 nand P2_U3031 P2_R1275_U7 ; P2_U4760
g5420 nand P2_U3037 P2_U3082 ; P2_U4761
g5421 nand P2_U3034 P2_R1215_U114 ; P2_U4762
g5422 nand P2_U3033 P2_ADD_1119_U72 ; P2_U4763
g5423 nand P2_U3032 P2_U3465 ; P2_U4764
g5424 nand P2_U3031 P2_R1275_U8 ; P2_U4765
g5425 nand P2_U3037 P2_U3081 ; P2_U4766
g5426 nand P2_U3034 P2_R1215_U12 ; P2_U4767
g5427 nand P2_U3033 P2_ADD_1119_U71 ; P2_U4768
g5428 nand P2_U3032 P2_U3468 ; P2_U4769
g5429 nand P2_U3031 P2_R1275_U86 ; P2_U4770
g5430 nand P2_U3037 P2_U3076 ; P2_U4771
g5431 nand P2_U3034 P2_R1215_U113 ; P2_U4772
g5432 nand P2_U3033 P2_ADD_1119_U70 ; P2_U4773
g5433 nand P2_U3032 P2_U3471 ; P2_U4774
g5434 nand P2_U3031 P2_R1275_U9 ; P2_U4775
g5435 nand P2_U3037 P2_U3075 ; P2_U4776
g5436 nand P2_U3034 P2_R1215_U112 ; P2_U4777
g5437 nand P2_U3033 P2_ADD_1119_U69 ; P2_U4778
g5438 nand P2_U3032 P2_U3474 ; P2_U4779
g5439 nand P2_U3031 P2_R1275_U10 ; P2_U4780
g5440 nand P2_U3037 P2_U3071 ; P2_U4781
g5441 nand P2_U3034 P2_R1215_U111 ; P2_U4782
g5442 nand P2_U3033 P2_ADD_1119_U68 ; P2_U4783
g5443 nand P2_U3032 P2_U3477 ; P2_U4784
g5444 nand P2_U3031 P2_R1275_U11 ; P2_U4785
g5445 nand P2_U3037 P2_U3084 ; P2_U4786
g5446 nand P2_U3034 P2_R1215_U13 ; P2_U4787
g5447 nand P2_U3033 P2_ADD_1119_U67 ; P2_U4788
g5448 nand P2_U3032 P2_U3480 ; P2_U4789
g5449 nand P2_U3031 P2_R1275_U84 ; P2_U4790
g5450 nand P2_U3037 P2_U3083 ; P2_U4791
g5451 nand P2_U3034 P2_R1215_U110 ; P2_U4792
g5452 nand P2_U3033 P2_ADD_1119_U66 ; P2_U4793
g5453 nand P2_U3032 P2_U3483 ; P2_U4794
g5454 nand P2_U3031 P2_R1275_U12 ; P2_U4795
g5455 nand P2_U3037 P2_U3078 ; P2_U4796
g5456 nand P2_U3034 P2_R1215_U109 ; P2_U4797
g5457 nand P2_U3033 P2_ADD_1119_U65 ; P2_U4798
g5458 nand P2_U3032 P2_U3485 ; P2_U4799
g5459 nand P2_U3031 P2_R1275_U82 ; P2_U4800
g5460 nand P2_U3037 P2_U3077 ; P2_U4801
g5461 nand P2_U3034 P2_R1215_U14 ; P2_U4802
g5462 nand P2_U3033 P2_ADD_1119_U64 ; P2_U4803
g5463 nand P2_U3032 P2_U3957 ; P2_U4804
g5464 nand P2_U3031 P2_R1275_U13 ; P2_U4805
g5465 nand P2_U3037 P2_U3063 ; P2_U4806
g5466 nand P2_U3034 P2_R1215_U15 ; P2_U4807
g5467 nand P2_U3033 P2_ADD_1119_U63 ; P2_U4808
g5468 nand P2_U3032 P2_U3956 ; P2_U4809
g5469 nand P2_U3031 P2_R1275_U78 ; P2_U4810
g5470 nand P2_U3037 P2_U3068 ; P2_U4811
g5471 nand P2_U3034 P2_R1215_U108 ; P2_U4812
g5472 nand P2_U3033 P2_ADD_1119_U62 ; P2_U4813
g5473 nand P2_U3032 P2_U3955 ; P2_U4814
g5474 nand P2_U3031 P2_R1275_U14 ; P2_U4815
g5475 nand P2_U3037 P2_U3067 ; P2_U4816
g5476 nand P2_U3034 P2_R1215_U107 ; P2_U4817
g5477 nand P2_U3033 P2_ADD_1119_U61 ; P2_U4818
g5478 nand P2_U3032 P2_U3954 ; P2_U4819
g5479 nand P2_U3031 P2_R1275_U76 ; P2_U4820
g5480 nand P2_U3037 P2_U3060 ; P2_U4821
g5481 nand P2_U3034 P2_R1215_U106 ; P2_U4822
g5482 nand P2_U3033 P2_ADD_1119_U60 ; P2_U4823
g5483 nand P2_U3032 P2_U3953 ; P2_U4824
g5484 nand P2_U3031 P2_R1275_U15 ; P2_U4825
g5485 nand P2_U3037 P2_U3059 ; P2_U4826
g5486 nand P2_U3034 P2_R1215_U105 ; P2_U4827
g5487 nand P2_U3033 P2_ADD_1119_U59 ; P2_U4828
g5488 nand P2_U3032 P2_U3952 ; P2_U4829
g5489 nand P2_U3031 P2_R1275_U74 ; P2_U4830
g5490 nand P2_U3037 P2_U3055 ; P2_U4831
g5491 nand P2_U3034 P2_R1215_U16 ; P2_U4832
g5492 nand P2_U3033 P2_ADD_1119_U58 ; P2_U4833
g5493 nand P2_U3032 P2_U3951 ; P2_U4834
g5494 nand P2_U3031 P2_R1275_U16 ; P2_U4835
g5495 nand P2_U3037 P2_U3056 ; P2_U4836
g5496 nand P2_U3034 P2_R1215_U104 ; P2_U4837
g5497 nand P2_U3033 P2_ADD_1119_U57 ; P2_U4838
g5498 nand P2_U3032 P2_U3950 ; P2_U4839
g5499 nand P2_U3031 P2_R1275_U72 ; P2_U4840
g5500 nand P2_U3037 P2_U3057 ; P2_U4841
g5501 nand P2_U3034 P2_R1215_U103 ; P2_U4842
g5502 nand P2_U3033 P2_ADD_1119_U56 ; P2_U4843
g5503 nand P2_U3032 P2_U3949 ; P2_U4844
g5504 nand P2_U3031 P2_R1275_U17 ; P2_U4845
g5505 nand P2_U3034 P2_R1215_U102 ; P2_U4846
g5506 nand P2_U3033 P2_ADD_1119_U5 ; P2_U4847
g5507 nand P2_U3032 P2_U3960 ; P2_U4848
g5508 nand P2_U3031 P2_R1275_U70 ; P2_U4849
g5509 nand P2_U3032 P2_U3959 ; P2_U4850
g5510 nand P2_U3031 P2_R1275_U19 ; P2_U4851
g5511 nand P2_U3032 P2_U3958 ; P2_U4852
g5512 nand P2_U3031 P2_R1275_U68 ; P2_U4853
g5513 nand P2_U3755 P2_U3395 P2_U3051 P2_U4700 P2_U3393 ; P2_U4854
g5514 nand P2_R1170_U13 P2_U3043 ; P2_U4855
g5515 nand P2_U3041 P2_U3424 ; P2_U4856
g5516 nand P2_R1209_U13 P2_U3039 ; P2_U4857
g5517 nand P2_U4856 P2_U4855 P2_U4857 ; P2_U4858
g5518 nand P2_R1170_U13 P2_U3018 ; P2_U4859
g5519 nand P2_U3017 P2_R1209_U13 ; P2_U4860
g5520 nand P2_U5683 P2_U3424 ; P2_U4861
g5521 nand P2_U4860 P2_U4859 P2_U4861 ; P2_U4862
g5522 not P2_U3401 ; P2_U4863
g5523 nand P2_U3045 P2_U4858 ; P2_U4864
g5524 nand P2_U3947 P2_U4862 ; P2_U4865
g5525 nand P2_U3044 P2_R1170_U13 ; P2_U4866
g5526 nand P2_U3088 P2_REG3_REG_19__SCAN_IN ; P2_U4867
g5527 nand P2_U3042 P2_U3424 ; P2_U4868
g5528 nand P2_U3040 P2_R1209_U13 ; P2_U4869
g5529 nand P2_U4863 P2_ADDR_REG_19__SCAN_IN ; P2_U4870
g5530 nand P2_R1170_U75 P2_U3043 ; P2_U4871
g5531 nand P2_U3041 P2_U3482 ; P2_U4872
g5532 nand P2_R1209_U75 P2_U3039 ; P2_U4873
g5533 nand P2_U4872 P2_U4871 P2_U4873 ; P2_U4874
g5534 nand P2_R1170_U75 P2_U3018 ; P2_U4875
g5535 nand P2_R1209_U75 P2_U3017 ; P2_U4876
g5536 nand P2_U5683 P2_U3482 ; P2_U4877
g5537 nand P2_U4876 P2_U4875 P2_U4877 ; P2_U4878
g5538 nand P2_U3045 P2_U4874 ; P2_U4879
g5539 nand P2_U3947 P2_U4878 ; P2_U4880
g5540 nand P2_R1170_U75 P2_U3044 ; P2_U4881
g5541 nand P2_U3088 P2_REG3_REG_18__SCAN_IN ; P2_U4882
g5542 nand P2_U3042 P2_U3482 ; P2_U4883
g5543 nand P2_R1209_U75 P2_U3040 ; P2_U4884
g5544 nand P2_U4863 P2_ADDR_REG_18__SCAN_IN ; P2_U4885
g5545 nand P2_R1170_U12 P2_U3043 ; P2_U4886
g5546 nand P2_U3041 P2_U3479 ; P2_U4887
g5547 nand P2_R1209_U12 P2_U3039 ; P2_U4888
g5548 nand P2_U4887 P2_U4886 P2_U4888 ; P2_U4889
g5549 nand P2_R1170_U12 P2_U3018 ; P2_U4890
g5550 nand P2_R1209_U12 P2_U3017 ; P2_U4891
g5551 nand P2_U5683 P2_U3479 ; P2_U4892
g5552 nand P2_U4891 P2_U4890 P2_U4892 ; P2_U4893
g5553 nand P2_U3045 P2_U4889 ; P2_U4894
g5554 nand P2_U3947 P2_U4893 ; P2_U4895
g5555 nand P2_R1170_U12 P2_U3044 ; P2_U4896
g5556 nand P2_U3088 P2_REG3_REG_17__SCAN_IN ; P2_U4897
g5557 nand P2_U3042 P2_U3479 ; P2_U4898
g5558 nand P2_R1209_U12 P2_U3040 ; P2_U4899
g5559 nand P2_U4863 P2_ADDR_REG_17__SCAN_IN ; P2_U4900
g5560 nand P2_R1170_U76 P2_U3043 ; P2_U4901
g5561 nand P2_U3041 P2_U3476 ; P2_U4902
g5562 nand P2_R1209_U76 P2_U3039 ; P2_U4903
g5563 nand P2_U4902 P2_U4901 P2_U4903 ; P2_U4904
g5564 nand P2_R1170_U76 P2_U3018 ; P2_U4905
g5565 nand P2_R1209_U76 P2_U3017 ; P2_U4906
g5566 nand P2_U5683 P2_U3476 ; P2_U4907
g5567 nand P2_U4906 P2_U4905 P2_U4907 ; P2_U4908
g5568 nand P2_U3045 P2_U4904 ; P2_U4909
g5569 nand P2_U3947 P2_U4908 ; P2_U4910
g5570 nand P2_R1170_U76 P2_U3044 ; P2_U4911
g5571 nand P2_U3088 P2_REG3_REG_16__SCAN_IN ; P2_U4912
g5572 nand P2_U3042 P2_U3476 ; P2_U4913
g5573 nand P2_R1209_U76 P2_U3040 ; P2_U4914
g5574 nand P2_U4863 P2_ADDR_REG_16__SCAN_IN ; P2_U4915
g5575 nand P2_R1170_U77 P2_U3043 ; P2_U4916
g5576 nand P2_U3041 P2_U3473 ; P2_U4917
g5577 nand P2_R1209_U77 P2_U3039 ; P2_U4918
g5578 nand P2_U4917 P2_U4916 P2_U4918 ; P2_U4919
g5579 nand P2_R1170_U77 P2_U3018 ; P2_U4920
g5580 nand P2_R1209_U77 P2_U3017 ; P2_U4921
g5581 nand P2_U5683 P2_U3473 ; P2_U4922
g5582 nand P2_U4921 P2_U4920 P2_U4922 ; P2_U4923
g5583 nand P2_U3045 P2_U4919 ; P2_U4924
g5584 nand P2_U3947 P2_U4923 ; P2_U4925
g5585 nand P2_R1170_U77 P2_U3044 ; P2_U4926
g5586 nand P2_U3088 P2_REG3_REG_15__SCAN_IN ; P2_U4927
g5587 nand P2_U3042 P2_U3473 ; P2_U4928
g5588 nand P2_R1209_U77 P2_U3040 ; P2_U4929
g5589 nand P2_U4863 P2_ADDR_REG_15__SCAN_IN ; P2_U4930
g5590 nand P2_R1170_U78 P2_U3043 ; P2_U4931
g5591 nand P2_U3041 P2_U3470 ; P2_U4932
g5592 nand P2_R1209_U78 P2_U3039 ; P2_U4933
g5593 nand P2_U4932 P2_U4931 P2_U4933 ; P2_U4934
g5594 nand P2_R1170_U78 P2_U3018 ; P2_U4935
g5595 nand P2_R1209_U78 P2_U3017 ; P2_U4936
g5596 nand P2_U5683 P2_U3470 ; P2_U4937
g5597 nand P2_U4936 P2_U4935 P2_U4937 ; P2_U4938
g5598 nand P2_U3045 P2_U4934 ; P2_U4939
g5599 nand P2_U3947 P2_U4938 ; P2_U4940
g5600 nand P2_R1170_U78 P2_U3044 ; P2_U4941
g5601 nand P2_U3088 P2_REG3_REG_14__SCAN_IN ; P2_U4942
g5602 nand P2_U3042 P2_U3470 ; P2_U4943
g5603 nand P2_R1209_U78 P2_U3040 ; P2_U4944
g5604 nand P2_U4863 P2_ADDR_REG_14__SCAN_IN ; P2_U4945
g5605 nand P2_R1170_U11 P2_U3043 ; P2_U4946
g5606 nand P2_U3041 P2_U3467 ; P2_U4947
g5607 nand P2_R1209_U11 P2_U3039 ; P2_U4948
g5608 nand P2_U4947 P2_U4946 P2_U4948 ; P2_U4949
g5609 nand P2_R1170_U11 P2_U3018 ; P2_U4950
g5610 nand P2_R1209_U11 P2_U3017 ; P2_U4951
g5611 nand P2_U5683 P2_U3467 ; P2_U4952
g5612 nand P2_U4951 P2_U4950 P2_U4952 ; P2_U4953
g5613 nand P2_U3045 P2_U4949 ; P2_U4954
g5614 nand P2_U3947 P2_U4953 ; P2_U4955
g5615 nand P2_R1170_U11 P2_U3044 ; P2_U4956
g5616 nand P2_U3088 P2_REG3_REG_13__SCAN_IN ; P2_U4957
g5617 nand P2_U3042 P2_U3467 ; P2_U4958
g5618 nand P2_R1209_U11 P2_U3040 ; P2_U4959
g5619 nand P2_U4863 P2_ADDR_REG_13__SCAN_IN ; P2_U4960
g5620 nand P2_R1170_U79 P2_U3043 ; P2_U4961
g5621 nand P2_U3041 P2_U3464 ; P2_U4962
g5622 nand P2_R1209_U79 P2_U3039 ; P2_U4963
g5623 nand P2_U4962 P2_U4961 P2_U4963 ; P2_U4964
g5624 nand P2_R1170_U79 P2_U3018 ; P2_U4965
g5625 nand P2_R1209_U79 P2_U3017 ; P2_U4966
g5626 nand P2_U5683 P2_U3464 ; P2_U4967
g5627 nand P2_U4966 P2_U4965 P2_U4967 ; P2_U4968
g5628 nand P2_U3045 P2_U4964 ; P2_U4969
g5629 nand P2_U3947 P2_U4968 ; P2_U4970
g5630 nand P2_R1170_U79 P2_U3044 ; P2_U4971
g5631 nand P2_U3088 P2_REG3_REG_12__SCAN_IN ; P2_U4972
g5632 nand P2_U3042 P2_U3464 ; P2_U4973
g5633 nand P2_R1209_U79 P2_U3040 ; P2_U4974
g5634 nand P2_U4863 P2_ADDR_REG_12__SCAN_IN ; P2_U4975
g5635 nand P2_R1170_U80 P2_U3043 ; P2_U4976
g5636 nand P2_U3041 P2_U3461 ; P2_U4977
g5637 nand P2_R1209_U80 P2_U3039 ; P2_U4978
g5638 nand P2_U4977 P2_U4976 P2_U4978 ; P2_U4979
g5639 nand P2_R1170_U80 P2_U3018 ; P2_U4980
g5640 nand P2_R1209_U80 P2_U3017 ; P2_U4981
g5641 nand P2_U5683 P2_U3461 ; P2_U4982
g5642 nand P2_U4981 P2_U4980 P2_U4982 ; P2_U4983
g5643 nand P2_U3045 P2_U4979 ; P2_U4984
g5644 nand P2_U3947 P2_U4983 ; P2_U4985
g5645 nand P2_R1170_U80 P2_U3044 ; P2_U4986
g5646 nand P2_U3088 P2_REG3_REG_11__SCAN_IN ; P2_U4987
g5647 nand P2_U3042 P2_U3461 ; P2_U4988
g5648 nand P2_R1209_U80 P2_U3040 ; P2_U4989
g5649 nand P2_U4863 P2_ADDR_REG_11__SCAN_IN ; P2_U4990
g5650 nand P2_R1170_U10 P2_U3043 ; P2_U4991
g5651 nand P2_U3041 P2_U3458 ; P2_U4992
g5652 nand P2_R1209_U10 P2_U3039 ; P2_U4993
g5653 nand P2_U4992 P2_U4991 P2_U4993 ; P2_U4994
g5654 nand P2_R1170_U10 P2_U3018 ; P2_U4995
g5655 nand P2_R1209_U10 P2_U3017 ; P2_U4996
g5656 nand P2_U5683 P2_U3458 ; P2_U4997
g5657 nand P2_U4996 P2_U4995 P2_U4997 ; P2_U4998
g5658 nand P2_U3045 P2_U4994 ; P2_U4999
g5659 nand P2_U3947 P2_U4998 ; P2_U5000
g5660 nand P2_R1170_U10 P2_U3044 ; P2_U5001
g5661 nand P2_U3088 P2_REG3_REG_10__SCAN_IN ; P2_U5002
g5662 nand P2_U3042 P2_U3458 ; P2_U5003
g5663 nand P2_R1209_U10 P2_U3040 ; P2_U5004
g5664 nand P2_U4863 P2_ADDR_REG_10__SCAN_IN ; P2_U5005
g5665 nand P2_R1170_U70 P2_U3043 ; P2_U5006
g5666 nand P2_U3041 P2_U3455 ; P2_U5007
g5667 nand P2_R1209_U70 P2_U3039 ; P2_U5008
g5668 nand P2_U5007 P2_U5006 P2_U5008 ; P2_U5009
g5669 nand P2_R1170_U70 P2_U3018 ; P2_U5010
g5670 nand P2_R1209_U70 P2_U3017 ; P2_U5011
g5671 nand P2_U5683 P2_U3455 ; P2_U5012
g5672 nand P2_U5011 P2_U5010 P2_U5012 ; P2_U5013
g5673 nand P2_U3045 P2_U5009 ; P2_U5014
g5674 nand P2_U3947 P2_U5013 ; P2_U5015
g5675 nand P2_R1170_U70 P2_U3044 ; P2_U5016
g5676 nand P2_U3088 P2_REG3_REG_9__SCAN_IN ; P2_U5017
g5677 nand P2_U3042 P2_U3455 ; P2_U5018
g5678 nand P2_R1209_U70 P2_U3040 ; P2_U5019
g5679 nand P2_U4863 P2_ADDR_REG_9__SCAN_IN ; P2_U5020
g5680 nand P2_R1170_U71 P2_U3043 ; P2_U5021
g5681 nand P2_U3041 P2_U3452 ; P2_U5022
g5682 nand P2_R1209_U71 P2_U3039 ; P2_U5023
g5683 nand P2_U5022 P2_U5021 P2_U5023 ; P2_U5024
g5684 nand P2_R1170_U71 P2_U3018 ; P2_U5025
g5685 nand P2_R1209_U71 P2_U3017 ; P2_U5026
g5686 nand P2_U5683 P2_U3452 ; P2_U5027
g5687 nand P2_U5026 P2_U5025 P2_U5027 ; P2_U5028
g5688 nand P2_U3045 P2_U5024 ; P2_U5029
g5689 nand P2_U3947 P2_U5028 ; P2_U5030
g5690 nand P2_R1170_U71 P2_U3044 ; P2_U5031
g5691 nand P2_U3088 P2_REG3_REG_8__SCAN_IN ; P2_U5032
g5692 nand P2_U3042 P2_U3452 ; P2_U5033
g5693 nand P2_R1209_U71 P2_U3040 ; P2_U5034
g5694 nand P2_U4863 P2_ADDR_REG_8__SCAN_IN ; P2_U5035
g5695 nand P2_R1170_U16 P2_U3043 ; P2_U5036
g5696 nand P2_U3041 P2_U3449 ; P2_U5037
g5697 nand P2_R1209_U16 P2_U3039 ; P2_U5038
g5698 nand P2_U5037 P2_U5036 P2_U5038 ; P2_U5039
g5699 nand P2_R1170_U16 P2_U3018 ; P2_U5040
g5700 nand P2_R1209_U16 P2_U3017 ; P2_U5041
g5701 nand P2_U5683 P2_U3449 ; P2_U5042
g5702 nand P2_U5041 P2_U5040 P2_U5042 ; P2_U5043
g5703 nand P2_U3045 P2_U5039 ; P2_U5044
g5704 nand P2_U3947 P2_U5043 ; P2_U5045
g5705 nand P2_R1170_U16 P2_U3044 ; P2_U5046
g5706 nand P2_U3088 P2_REG3_REG_7__SCAN_IN ; P2_U5047
g5707 nand P2_U3042 P2_U3449 ; P2_U5048
g5708 nand P2_R1209_U16 P2_U3040 ; P2_U5049
g5709 nand P2_U4863 P2_ADDR_REG_7__SCAN_IN ; P2_U5050
g5710 nand P2_R1170_U72 P2_U3043 ; P2_U5051
g5711 nand P2_U3041 P2_U3446 ; P2_U5052
g5712 nand P2_R1209_U72 P2_U3039 ; P2_U5053
g5713 nand P2_U5052 P2_U5051 P2_U5053 ; P2_U5054
g5714 nand P2_R1170_U72 P2_U3018 ; P2_U5055
g5715 nand P2_R1209_U72 P2_U3017 ; P2_U5056
g5716 nand P2_U5683 P2_U3446 ; P2_U5057
g5717 nand P2_U5056 P2_U5055 P2_U5057 ; P2_U5058
g5718 nand P2_U3045 P2_U5054 ; P2_U5059
g5719 nand P2_U3947 P2_U5058 ; P2_U5060
g5720 nand P2_R1170_U72 P2_U3044 ; P2_U5061
g5721 nand P2_U3088 P2_REG3_REG_6__SCAN_IN ; P2_U5062
g5722 nand P2_U3042 P2_U3446 ; P2_U5063
g5723 nand P2_R1209_U72 P2_U3040 ; P2_U5064
g5724 nand P2_U4863 P2_ADDR_REG_6__SCAN_IN ; P2_U5065
g5725 nand P2_R1170_U15 P2_U3043 ; P2_U5066
g5726 nand P2_U3041 P2_U3443 ; P2_U5067
g5727 nand P2_R1209_U15 P2_U3039 ; P2_U5068
g5728 nand P2_U5067 P2_U5066 P2_U5068 ; P2_U5069
g5729 nand P2_R1170_U15 P2_U3018 ; P2_U5070
g5730 nand P2_R1209_U15 P2_U3017 ; P2_U5071
g5731 nand P2_U5683 P2_U3443 ; P2_U5072
g5732 nand P2_U5071 P2_U5070 P2_U5072 ; P2_U5073
g5733 nand P2_U3045 P2_U5069 ; P2_U5074
g5734 nand P2_U3947 P2_U5073 ; P2_U5075
g5735 nand P2_R1170_U15 P2_U3044 ; P2_U5076
g5736 nand P2_U3088 P2_REG3_REG_5__SCAN_IN ; P2_U5077
g5737 nand P2_U3042 P2_U3443 ; P2_U5078
g5738 nand P2_R1209_U15 P2_U3040 ; P2_U5079
g5739 nand P2_U4863 P2_ADDR_REG_5__SCAN_IN ; P2_U5080
g5740 nand P2_R1170_U73 P2_U3043 ; P2_U5081
g5741 nand P2_U3041 P2_U3440 ; P2_U5082
g5742 nand P2_R1209_U73 P2_U3039 ; P2_U5083
g5743 nand P2_U5082 P2_U5081 P2_U5083 ; P2_U5084
g5744 nand P2_R1170_U73 P2_U3018 ; P2_U5085
g5745 nand P2_R1209_U73 P2_U3017 ; P2_U5086
g5746 nand P2_U5683 P2_U3440 ; P2_U5087
g5747 nand P2_U5086 P2_U5085 P2_U5087 ; P2_U5088
g5748 nand P2_U3045 P2_U5084 ; P2_U5089
g5749 nand P2_U3947 P2_U5088 ; P2_U5090
g5750 nand P2_R1170_U73 P2_U3044 ; P2_U5091
g5751 nand P2_U3088 P2_REG3_REG_4__SCAN_IN ; P2_U5092
g5752 nand P2_U3042 P2_U3440 ; P2_U5093
g5753 nand P2_R1209_U73 P2_U3040 ; P2_U5094
g5754 nand P2_U4863 P2_ADDR_REG_4__SCAN_IN ; P2_U5095
g5755 nand P2_R1170_U74 P2_U3043 ; P2_U5096
g5756 nand P2_U3041 P2_U3437 ; P2_U5097
g5757 nand P2_R1209_U74 P2_U3039 ; P2_U5098
g5758 nand P2_U5097 P2_U5096 P2_U5098 ; P2_U5099
g5759 nand P2_R1170_U74 P2_U3018 ; P2_U5100
g5760 nand P2_R1209_U74 P2_U3017 ; P2_U5101
g5761 nand P2_U5683 P2_U3437 ; P2_U5102
g5762 nand P2_U5101 P2_U5100 P2_U5102 ; P2_U5103
g5763 nand P2_U3045 P2_U5099 ; P2_U5104
g5764 nand P2_U3947 P2_U5103 ; P2_U5105
g5765 nand P2_R1170_U74 P2_U3044 ; P2_U5106
g5766 nand P2_U3088 P2_REG3_REG_3__SCAN_IN ; P2_U5107
g5767 nand P2_U3042 P2_U3437 ; P2_U5108
g5768 nand P2_R1209_U74 P2_U3040 ; P2_U5109
g5769 nand P2_U4863 P2_ADDR_REG_3__SCAN_IN ; P2_U5110
g5770 nand P2_R1170_U14 P2_U3043 ; P2_U5111
g5771 nand P2_U3041 P2_U3434 ; P2_U5112
g5772 nand P2_R1209_U14 P2_U3039 ; P2_U5113
g5773 nand P2_U5112 P2_U5111 P2_U5113 ; P2_U5114
g5774 nand P2_R1170_U14 P2_U3018 ; P2_U5115
g5775 nand P2_R1209_U14 P2_U3017 ; P2_U5116
g5776 nand P2_U5683 P2_U3434 ; P2_U5117
g5777 nand P2_U5116 P2_U5115 P2_U5117 ; P2_U5118
g5778 nand P2_U3045 P2_U5114 ; P2_U5119
g5779 nand P2_U3947 P2_U5118 ; P2_U5120
g5780 nand P2_R1170_U14 P2_U3044 ; P2_U5121
g5781 nand P2_U3088 P2_REG3_REG_2__SCAN_IN ; P2_U5122
g5782 nand P2_U3042 P2_U3434 ; P2_U5123
g5783 nand P2_R1209_U14 P2_U3040 ; P2_U5124
g5784 nand P2_U4863 P2_ADDR_REG_2__SCAN_IN ; P2_U5125
g5785 nand P2_R1170_U68 P2_U3043 ; P2_U5126
g5786 nand P2_U3041 P2_U3431 ; P2_U5127
g5787 nand P2_R1209_U68 P2_U3039 ; P2_U5128
g5788 nand P2_U5127 P2_U5126 P2_U5128 ; P2_U5129
g5789 nand P2_R1170_U68 P2_U3018 ; P2_U5130
g5790 nand P2_R1209_U68 P2_U3017 ; P2_U5131
g5791 nand P2_U5683 P2_U3431 ; P2_U5132
g5792 nand P2_U5131 P2_U5130 P2_U5132 ; P2_U5133
g5793 nand P2_U3045 P2_U5129 ; P2_U5134
g5794 nand P2_U3947 P2_U5133 ; P2_U5135
g5795 nand P2_R1170_U68 P2_U3044 ; P2_U5136
g5796 nand P2_U3088 P2_REG3_REG_1__SCAN_IN ; P2_U5137
g5797 nand P2_U3042 P2_U3431 ; P2_U5138
g5798 nand P2_R1209_U68 P2_U3040 ; P2_U5139
g5799 nand P2_U4863 P2_ADDR_REG_1__SCAN_IN ; P2_U5140
g5800 nand P2_R1170_U69 P2_U3043 ; P2_U5141
g5801 nand P2_U3041 P2_U3425 ; P2_U5142
g5802 nand P2_R1209_U69 P2_U3039 ; P2_U5143
g5803 nand P2_U5142 P2_U5141 P2_U5143 ; P2_U5144
g5804 nand P2_R1170_U69 P2_U3018 ; P2_U5145
g5805 nand P2_R1209_U69 P2_U3017 ; P2_U5146
g5806 nand P2_U5683 P2_U3425 ; P2_U5147
g5807 nand P2_U5146 P2_U5145 P2_U5147 ; P2_U5148
g5808 nand P2_U3045 P2_U5144 ; P2_U5149
g5809 nand P2_U3947 P2_U5148 ; P2_U5150
g5810 nand P2_R1170_U69 P2_U3044 ; P2_U5151
g5811 nand P2_U3088 P2_REG3_REG_0__SCAN_IN ; P2_U5152
g5812 nand P2_U3042 P2_U3425 ; P2_U5153
g5813 nand P2_R1209_U69 P2_U3040 ; P2_U5154
g5814 nand P2_U4863 P2_ADDR_REG_0__SCAN_IN ; P2_U5155
g5815 not P2_U3918 ; P2_U5156
g5816 nand P2_U3936 P2_U3334 P2_U3337 ; P2_U5157
g5817 nand P2_U5665 P2_U5671 ; P2_U5158
g5818 nand P2_U3424 P2_U5158 ; P2_U5159
g5819 nand P2_U3419 P2_U5159 ; P2_U5160
g5820 nand P2_U3340 P2_U5160 ; P2_U5161
g5821 nand P2_U6052 P2_U6051 P2_U3052 ; P2_U5162
g5822 nand P2_U5162 P2_B_REG_SCAN_IN ; P2_U5163
g5823 nand P2_U3038 P2_U3081 ; P2_U5164
g5824 nand P2_U3036 P2_U3075 ; P2_U5165
g5825 nand P2_ADD_1119_U69 P2_U3406 ; P2_U5166
g5826 nand P2_U5165 P2_U5164 P2_U5166 ; P2_U5167
g5827 not P2_U3154 ; P2_U5168
g5828 nand P2_U3923 P2_U3346 ; P2_U5169
g5829 nand P2_U3419 P2_U5169 ; P2_U5170
g5830 nand P2_U3800 P2_U5170 P2_U3801 ; P2_U5171
g5831 nand P2_U5171 P2_U3406 ; P2_U5172
g5832 not P2_U3408 ; P2_U5173
g5833 nand P2_U3474 P2_U5636 ; P2_U5174
g5834 nand P2_ADD_1119_U69 P2_U5635 ; P2_U5175
g5835 nand P2_R1176_U111 P2_U3028 ; P2_U5176
g5836 nand P2_U3969 P2_U5167 ; P2_U5177
g5837 nand P2_U3088 P2_REG3_REG_15__SCAN_IN ; P2_U5178
g5838 nand P2_U3038 P2_U3060 ; P2_U5179
g5839 nand P2_U3036 P2_U3055 ; P2_U5180
g5840 nand P2_ADD_1119_U58 P2_U3406 ; P2_U5181
g5841 nand P2_U5181 P2_U5179 P2_U5180 ; P2_U5182
g5842 nand P2_U3398 P2_U3406 ; P2_U5183
g5843 nand P2_U5173 P2_U5183 ; P2_U5184
g5844 nand P2_U3946 P2_U3398 ; P2_U5185
g5845 nand P2_U3393 P2_U5185 ; P2_U5186
g5846 nand P2_U3047 P2_U3951 ; P2_U5187
g5847 nand P2_U3046 P2_ADD_1119_U58 ; P2_U5188
g5848 nand P2_R1176_U16 P2_U3028 ; P2_U5189
g5849 nand P2_U3969 P2_U5182 ; P2_U5190
g5850 nand P2_U3088 P2_REG3_REG_26__SCAN_IN ; P2_U5191
g5851 nand P2_U3038 P2_U3069 ; P2_U5192
g5852 nand P2_U3036 P2_U3072 ; P2_U5193
g5853 nand P2_ADD_1119_U53 P2_U3406 ; P2_U5194
g5854 nand P2_U5193 P2_U5192 P2_U5194 ; P2_U5195
g5855 nand P2_U3447 P2_U5636 ; P2_U5196
g5856 nand P2_ADD_1119_U53 P2_U5635 ; P2_U5197
g5857 nand P2_R1176_U96 P2_U3028 ; P2_U5198
g5858 nand P2_U3969 P2_U5195 ; P2_U5199
g5859 nand P2_U3088 P2_REG3_REG_6__SCAN_IN ; P2_U5200
g5860 nand P2_U3038 P2_U3071 ; P2_U5201
g5861 nand P2_U3036 P2_U3083 ; P2_U5202
g5862 nand P2_ADD_1119_U66 P2_U3406 ; P2_U5203
g5863 nand P2_U5202 P2_U5201 P2_U5203 ; P2_U5204
g5864 nand P2_U3483 P2_U5636 ; P2_U5205
g5865 nand P2_ADD_1119_U66 P2_U5635 ; P2_U5206
g5866 nand P2_R1176_U109 P2_U3028 ; P2_U5207
g5867 nand P2_U3969 P2_U5204 ; P2_U5208
g5868 nand P2_U3088 P2_REG3_REG_18__SCAN_IN ; P2_U5209
g5869 nand P2_U3038 P2_U3080 ; P2_U5210
g5870 nand P2_U3036 P2_U3066 ; P2_U5211
g5871 nand P2_U3406 P2_REG3_REG_2__SCAN_IN ; P2_U5212
g5872 nand P2_U5211 P2_U5210 P2_U5212 ; P2_U5213
g5873 nand P2_U3435 P2_U5636 ; P2_U5214
g5874 nand P2_U5635 P2_REG3_REG_2__SCAN_IN ; P2_U5215
g5875 nand P2_R1176_U99 P2_U3028 ; P2_U5216
g5876 nand P2_U3969 P2_U5213 ; P2_U5217
g5877 nand P2_U3088 P2_REG3_REG_2__SCAN_IN ; P2_U5218
g5878 nand P2_U3038 P2_U3064 ; P2_U5219
g5879 nand P2_U3036 P2_U3074 ; P2_U5220
g5880 nand P2_ADD_1119_U73 P2_U3406 ; P2_U5221
g5881 nand P2_U5220 P2_U5219 P2_U5221 ; P2_U5222
g5882 nand P2_U3462 P2_U5636 ; P2_U5223
g5883 nand P2_ADD_1119_U73 P2_U5635 ; P2_U5224
g5884 nand P2_R1176_U114 P2_U3028 ; P2_U5225
g5885 nand P2_U3969 P2_U5222 ; P2_U5226
g5886 nand P2_U3088 P2_REG3_REG_11__SCAN_IN ; P2_U5227
g5887 nand P2_U3038 P2_U3077 ; P2_U5228
g5888 nand P2_U3036 P2_U3068 ; P2_U5229
g5889 nand P2_ADD_1119_U62 P2_U3406 ; P2_U5230
g5890 nand P2_U5229 P2_U5228 P2_U5230 ; P2_U5231
g5891 nand P2_U3047 P2_U3955 ; P2_U5232
g5892 nand P2_U3046 P2_ADD_1119_U62 ; P2_U5233
g5893 nand P2_R1176_U105 P2_U3028 ; P2_U5234
g5894 nand P2_U3969 P2_U5231 ; P2_U5235
g5895 nand P2_U3088 P2_REG3_REG_22__SCAN_IN ; P2_U5236
g5896 nand P2_U3038 P2_U3074 ; P2_U5237
g5897 nand P2_U3036 P2_U3081 ; P2_U5238
g5898 nand P2_ADD_1119_U71 P2_U3406 ; P2_U5239
g5899 nand P2_U5238 P2_U5237 P2_U5239 ; P2_U5240
g5900 nand P2_U3468 P2_U5636 ; P2_U5241
g5901 nand P2_ADD_1119_U71 P2_U5635 ; P2_U5242
g5902 nand P2_R1176_U13 P2_U3028 ; P2_U5243
g5903 nand P2_U3969 P2_U5240 ; P2_U5244
g5904 nand P2_U3088 P2_REG3_REG_13__SCAN_IN ; P2_U5245
g5905 nand P2_U3038 P2_U3083 ; P2_U5246
g5906 nand P2_U3036 P2_U3077 ; P2_U5247
g5907 nand P2_ADD_1119_U64 P2_U3406 ; P2_U5248
g5908 nand P2_U5247 P2_U5246 P2_U5248 ; P2_U5249
g5909 nand P2_U3047 P2_U3957 ; P2_U5250
g5910 nand P2_U3046 P2_ADD_1119_U64 ; P2_U5251
g5911 nand P2_R1176_U106 P2_U3028 ; P2_U5252
g5912 nand P2_U3969 P2_U5249 ; P2_U5253
g5913 nand P2_U3088 P2_REG3_REG_20__SCAN_IN ; P2_U5254
g5914 nand P2_U3407 P2_U3405 ; P2_U5255
g5915 nand P2_U5255 P2_U3406 ; P2_U5256
g5916 nand P2_U3970 P2_U5256 ; P2_U5257
g5917 nand P2_U3806 P2_U3036 ; P2_U5258
g5918 nand P2_U3427 P2_U5636 ; P2_U5259
g5919 nand P2_U5257 P2_REG3_REG_0__SCAN_IN ; P2_U5260
g5920 nand P2_R1176_U93 P2_U3028 ; P2_U5261
g5921 nand P2_U3088 P2_REG3_REG_0__SCAN_IN ; P2_U5262
g5922 nand P2_U3038 P2_U3086 ; P2_U5263
g5923 nand P2_U3036 P2_U3064 ; P2_U5264
g5924 nand P2_ADD_1119_U50 P2_U3406 ; P2_U5265
g5925 nand P2_U5264 P2_U5263 P2_U5265 ; P2_U5266
g5926 nand P2_U3456 P2_U5636 ; P2_U5267
g5927 nand P2_ADD_1119_U50 P2_U5635 ; P2_U5268
g5928 nand P2_R1176_U94 P2_U3028 ; P2_U5269
g5929 nand P2_U3969 P2_U5266 ; P2_U5270
g5930 nand P2_U3088 P2_REG3_REG_9__SCAN_IN ; P2_U5271
g5931 nand P2_U3038 P2_U3066 ; P2_U5272
g5932 nand P2_U3036 P2_U3069 ; P2_U5273
g5933 nand P2_ADD_1119_U55 P2_U3406 ; P2_U5274
g5934 nand P2_U5273 P2_U5272 P2_U5274 ; P2_U5275
g5935 nand P2_U3441 P2_U5636 ; P2_U5276
g5936 nand P2_ADD_1119_U55 P2_U5635 ; P2_U5277
g5937 nand P2_R1176_U98 P2_U3028 ; P2_U5278
g5938 nand P2_U3969 P2_U5275 ; P2_U5279
g5939 nand P2_U3088 P2_REG3_REG_4__SCAN_IN ; P2_U5280
g5940 nand P2_U3038 P2_U3068 ; P2_U5281
g5941 nand P2_U3036 P2_U3060 ; P2_U5282
g5942 nand P2_ADD_1119_U60 P2_U3406 ; P2_U5283
g5943 nand P2_U5282 P2_U5281 P2_U5283 ; P2_U5284
g5944 nand P2_U3047 P2_U3953 ; P2_U5285
g5945 nand P2_U3046 P2_ADD_1119_U60 ; P2_U5286
g5946 nand P2_R1176_U103 P2_U3028 ; P2_U5287
g5947 nand P2_U3969 P2_U5284 ; P2_U5288
g5948 nand P2_U3088 P2_REG3_REG_24__SCAN_IN ; P2_U5289
g5949 nand P2_U3038 P2_U3075 ; P2_U5290
g5950 nand P2_U3036 P2_U3084 ; P2_U5291
g5951 nand P2_ADD_1119_U67 P2_U3406 ; P2_U5292
g5952 nand P2_U5291 P2_U5290 P2_U5292 ; P2_U5293
g5953 nand P2_U3480 P2_U5636 ; P2_U5294
g5954 nand P2_ADD_1119_U67 P2_U5635 ; P2_U5295
g5955 nand P2_R1176_U14 P2_U3028 ; P2_U5296
g5956 nand P2_U3969 P2_U5293 ; P2_U5297
g5957 nand P2_U3088 P2_REG3_REG_17__SCAN_IN ; P2_U5298
g5958 nand P2_U3038 P2_U3062 ; P2_U5299
g5959 nand P2_U3036 P2_U3073 ; P2_U5300
g5960 nand P2_ADD_1119_U54 P2_U3406 ; P2_U5301
g5961 nand P2_U5300 P2_U5299 P2_U5301 ; P2_U5302
g5962 nand P2_U3444 P2_U5636 ; P2_U5303
g5963 nand P2_ADD_1119_U54 P2_U5635 ; P2_U5304
g5964 nand P2_R1176_U97 P2_U3028 ; P2_U5305
g5965 nand P2_U3969 P2_U5302 ; P2_U5306
g5966 nand P2_U3088 P2_REG3_REG_5__SCAN_IN ; P2_U5307
g5967 nand P2_U3038 P2_U3076 ; P2_U5308
g5968 nand P2_U3036 P2_U3071 ; P2_U5309
g5969 nand P2_ADD_1119_U68 P2_U3406 ; P2_U5310
g5970 nand P2_U5309 P2_U5308 P2_U5310 ; P2_U5311
g5971 nand P2_U3477 P2_U5636 ; P2_U5312
g5972 nand P2_ADD_1119_U68 P2_U5635 ; P2_U5313
g5973 nand P2_R1176_U110 P2_U3028 ; P2_U5314
g5974 nand P2_U3969 P2_U5311 ; P2_U5315
g5975 nand P2_U3088 P2_REG3_REG_16__SCAN_IN ; P2_U5316
g5976 nand P2_U3038 P2_U3067 ; P2_U5317
g5977 nand P2_U3036 P2_U3059 ; P2_U5318
g5978 nand P2_ADD_1119_U59 P2_U3406 ; P2_U5319
g5979 nand P2_U5318 P2_U5317 P2_U5319 ; P2_U5320
g5980 nand P2_U3047 P2_U3952 ; P2_U5321
g5981 nand P2_U3046 P2_ADD_1119_U59 ; P2_U5322
g5982 nand P2_R1176_U102 P2_U3028 ; P2_U5323
g5983 nand P2_U3969 P2_U5320 ; P2_U5324
g5984 nand P2_U3088 P2_REG3_REG_25__SCAN_IN ; P2_U5325
g5985 nand P2_U3038 P2_U3065 ; P2_U5326
g5986 nand P2_U3036 P2_U3082 ; P2_U5327
g5987 nand P2_ADD_1119_U72 P2_U3406 ; P2_U5328
g5988 nand P2_U5327 P2_U5326 P2_U5328 ; P2_U5329
g5989 nand P2_U3465 P2_U5636 ; P2_U5330
g5990 nand P2_ADD_1119_U72 P2_U5635 ; P2_U5331
g5991 nand P2_R1176_U113 P2_U3028 ; P2_U5332
g5992 nand P2_U3969 P2_U5329 ; P2_U5333
g5993 nand P2_U3088 P2_REG3_REG_12__SCAN_IN ; P2_U5334
g5994 nand P2_U3038 P2_U3078 ; P2_U5335
g5995 nand P2_U3036 P2_U3063 ; P2_U5336
g5996 nand P2_ADD_1119_U63 P2_U3406 ; P2_U5337
g5997 nand P2_U5336 P2_U5335 P2_U5337 ; P2_U5338
g5998 nand P2_U3047 P2_U3956 ; P2_U5339
g5999 nand P2_U3046 P2_ADD_1119_U63 ; P2_U5340
g6000 nand P2_R1176_U15 P2_U3028 ; P2_U5341
g6001 nand P2_U3969 P2_U5338 ; P2_U5342
g6002 nand P2_U3088 P2_REG3_REG_21__SCAN_IN ; P2_U5343
g6003 nand P2_U3038 P2_U3079 ; P2_U5344
g6004 nand P2_U3036 P2_U3070 ; P2_U5345
g6005 nand P2_U3406 P2_REG3_REG_1__SCAN_IN ; P2_U5346
g6006 nand P2_U5345 P2_U5344 P2_U5346 ; P2_U5347
g6007 nand P2_U3432 P2_U5636 ; P2_U5348
g6008 nand P2_U5635 P2_REG3_REG_1__SCAN_IN ; P2_U5349
g6009 nand P2_R1176_U107 P2_U3028 ; P2_U5350
g6010 nand P2_U3969 P2_U5347 ; P2_U5351
g6011 nand P2_U3088 P2_REG3_REG_1__SCAN_IN ; P2_U5352
g6012 nand P2_U3038 P2_U3072 ; P2_U5353
g6013 nand P2_U3036 P2_U3085 ; P2_U5354
g6014 nand P2_ADD_1119_U51 P2_U3406 ; P2_U5355
g6015 nand P2_U5354 P2_U5353 P2_U5355 ; P2_U5356
g6016 nand P2_U3453 P2_U5636 ; P2_U5357
g6017 nand P2_ADD_1119_U51 P2_U5635 ; P2_U5358
g6018 nand P2_R1176_U95 P2_U3028 ; P2_U5359
g6019 nand P2_U3969 P2_U5356 ; P2_U5360
g6020 nand P2_U3088 P2_REG3_REG_8__SCAN_IN ; P2_U5361
g6021 nand P2_U3038 P2_U3055 ; P2_U5362
g6022 nand P2_U3036 P2_U3057 ; P2_U5363
g6023 nand P2_ADD_1119_U56 P2_U3406 ; P2_U5364
g6024 nand P2_U5363 P2_U5364 P2_U5362 ; P2_U5365
g6025 nand P2_U3047 P2_U3949 ; P2_U5366
g6026 nand P2_U3046 P2_ADD_1119_U56 ; P2_U5367
g6027 nand P2_R1176_U100 P2_U3028 ; P2_U5368
g6028 nand P2_U3969 P2_U5365 ; P2_U5369
g6029 nand P2_U3088 P2_REG3_REG_28__SCAN_IN ; P2_U5370
g6030 nand P2_U3038 P2_U3084 ; P2_U5371
g6031 nand P2_U3036 P2_U3078 ; P2_U5372
g6032 nand P2_ADD_1119_U65 P2_U3406 ; P2_U5373
g6033 nand P2_U5372 P2_U5371 P2_U5373 ; P2_U5374
g6034 nand P2_U3485 P2_U5636 ; P2_U5375
g6035 nand P2_ADD_1119_U65 P2_U5635 ; P2_U5376
g6036 nand P2_R1176_U108 P2_U3028 ; P2_U5377
g6037 nand P2_U3969 P2_U5374 ; P2_U5378
g6038 nand P2_U3088 P2_REG3_REG_19__SCAN_IN ; P2_U5379
g6039 nand P2_U3038 P2_U3070 ; P2_U5380
g6040 nand P2_U3036 P2_U3062 ; P2_U5381
g6041 nand P2_ADD_1119_U4 P2_U3406 ; P2_U5382
g6042 nand P2_U5381 P2_U5380 P2_U5382 ; P2_U5383
g6043 nand P2_U3438 P2_U5636 ; P2_U5384
g6044 nand P2_ADD_1119_U4 P2_U5635 ; P2_U5385
g6045 nand P2_R1176_U17 P2_U3028 ; P2_U5386
g6046 nand P2_U3969 P2_U5383 ; P2_U5387
g6047 nand P2_U3088 P2_REG3_REG_3__SCAN_IN ; P2_U5388
g6048 nand P2_U3038 P2_U3085 ; P2_U5389
g6049 nand P2_U3036 P2_U3065 ; P2_U5390
g6050 nand P2_ADD_1119_U74 P2_U3406 ; P2_U5391
g6051 nand P2_U5390 P2_U5389 P2_U5391 ; P2_U5392
g6052 nand P2_U3459 P2_U5636 ; P2_U5393
g6053 nand P2_ADD_1119_U74 P2_U5635 ; P2_U5394
g6054 nand P2_R1176_U115 P2_U3028 ; P2_U5395
g6055 nand P2_U3969 P2_U5392 ; P2_U5396
g6056 nand P2_U3088 P2_REG3_REG_10__SCAN_IN ; P2_U5397
g6057 nand P2_U3038 P2_U3063 ; P2_U5398
g6058 nand P2_U3036 P2_U3067 ; P2_U5399
g6059 nand P2_ADD_1119_U61 P2_U3406 ; P2_U5400
g6060 nand P2_U5399 P2_U5398 P2_U5400 ; P2_U5401
g6061 nand P2_U3047 P2_U3954 ; P2_U5402
g6062 nand P2_U3046 P2_ADD_1119_U61 ; P2_U5403
g6063 nand P2_R1176_U104 P2_U3028 ; P2_U5404
g6064 nand P2_U3969 P2_U5401 ; P2_U5405
g6065 nand P2_U3088 P2_REG3_REG_23__SCAN_IN ; P2_U5406
g6066 nand P2_U3038 P2_U3082 ; P2_U5407
g6067 nand P2_U3036 P2_U3076 ; P2_U5408
g6068 nand P2_ADD_1119_U70 P2_U3406 ; P2_U5409
g6069 nand P2_U5408 P2_U5407 P2_U5409 ; P2_U5410
g6070 nand P2_U3471 P2_U5636 ; P2_U5411
g6071 nand P2_ADD_1119_U70 P2_U5635 ; P2_U5412
g6072 nand P2_R1176_U112 P2_U3028 ; P2_U5413
g6073 nand P2_U3969 P2_U5410 ; P2_U5414
g6074 nand P2_U3088 P2_REG3_REG_14__SCAN_IN ; P2_U5415
g6075 nand P2_U3038 P2_U3059 ; P2_U5416
g6076 nand P2_U3036 P2_U3056 ; P2_U5417
g6077 nand P2_ADD_1119_U57 P2_U3406 ; P2_U5418
g6078 nand P2_U5418 P2_U5416 P2_U5417 ; P2_U5419
g6079 nand P2_U3047 P2_U3950 ; P2_U5420
g6080 nand P2_U3046 P2_ADD_1119_U57 ; P2_U5421
g6081 nand P2_R1176_U101 P2_U3028 ; P2_U5422
g6082 nand P2_U3969 P2_U5419 ; P2_U5423
g6083 nand P2_U3088 P2_REG3_REG_27__SCAN_IN ; P2_U5424
g6084 nand P2_U3038 P2_U3073 ; P2_U5425
g6085 nand P2_U3036 P2_U3086 ; P2_U5426
g6086 nand P2_ADD_1119_U52 P2_U3406 ; P2_U5427
g6087 nand P2_U5426 P2_U5425 P2_U5427 ; P2_U5428
g6088 nand P2_U3450 P2_U5636 ; P2_U5429
g6089 nand P2_ADD_1119_U52 P2_U5635 ; P2_U5430
g6090 nand P2_R1176_U18 P2_U3028 ; P2_U5431
g6091 nand P2_U3969 P2_U5428 ; P2_U5432
g6092 nand P2_U3088 P2_REG3_REG_7__SCAN_IN ; P2_U5433
g6093 nand P2_U3948 P2_U3048 ; P2_U5434
g6094 nand P2_U3415 P2_U3347 ; P2_U5435
g6095 nand P2_U3419 P2_U3418 ; P2_U5436
g6096 nand P2_U3816 P2_U3051 ; P2_U5437
g6097 not P2_U3411 ; P2_U5438
g6098 nand P2_U3015 P2_U3415 ; P2_U5439
g6099 nand P2_U3411 P2_U3409 ; P2_U5440
g6100 nand P2_U3053 P2_U5440 ; P2_U5441
g6101 nand P2_U3085 P2_U3029 ; P2_U5442
g6102 nand P2_U5441 P2_U3085 ; P2_U5443
g6103 nand P2_U3929 P2_U3456 ; P2_U5444
g6104 nand P2_U3086 P2_U3029 ; P2_U5445
g6105 nand P2_U5441 P2_U3086 ; P2_U5446
g6106 nand P2_U3929 P2_U3453 ; P2_U5447
g6107 nand P2_U3072 P2_U3029 ; P2_U5448
g6108 nand P2_U5441 P2_U3072 ; P2_U5449
g6109 nand P2_U3929 P2_U3450 ; P2_U5450
g6110 nand P2_U3073 P2_U3029 ; P2_U5451
g6111 nand P2_U5441 P2_U3073 ; P2_U5452
g6112 nand P2_U3929 P2_U3447 ; P2_U5453
g6113 nand P2_U3069 P2_U3029 ; P2_U5454
g6114 nand P2_U5441 P2_U3069 ; P2_U5455
g6115 nand P2_U3929 P2_U3444 ; P2_U5456
g6116 nand P2_U3062 P2_U3029 ; P2_U5457
g6117 nand P2_U5441 P2_U3062 ; P2_U5458
g6118 nand P2_U3929 P2_U3441 ; P2_U5459
g6119 nand P2_R1335_U8 P2_U3029 ; P2_U5460
g6120 nand P2_U5441 P2_U3058 ; P2_U5461
g6121 nand P2_R1335_U6 P2_U3029 ; P2_U5462
g6122 nand P2_U5441 P2_U3061 ; P2_U5463
g6123 nand P2_U3929 P2_U3347 U70 ; P2_U5464
g6124 nand P2_U3066 P2_U3029 ; P2_U5465
g6125 nand P2_U5441 P2_U3066 ; P2_U5466
g6126 nand P2_U3929 P2_U3438 ; P2_U5467
g6127 nand P2_U3057 P2_U3029 ; P2_U5468
g6128 nand P2_U5441 P2_U3057 ; P2_U5469
g6129 nand P2_U3929 P2_U3960 ; P2_U5470
g6130 nand P2_U3056 P2_U3029 ; P2_U5471
g6131 nand P2_U5441 P2_U3056 ; P2_U5472
g6132 nand P2_U3929 P2_U3949 ; P2_U5473
g6133 nand P2_U3055 P2_U3029 ; P2_U5474
g6134 nand P2_U5441 P2_U3055 ; P2_U5475
g6135 nand P2_U3929 P2_U3950 ; P2_U5476
g6136 nand P2_U3059 P2_U3029 ; P2_U5477
g6137 nand P2_U5441 P2_U3059 ; P2_U5478
g6138 nand P2_U3929 P2_U3951 ; P2_U5479
g6139 nand P2_U3060 P2_U3029 ; P2_U5480
g6140 nand P2_U5441 P2_U3060 ; P2_U5481
g6141 nand P2_U3929 P2_U3952 ; P2_U5482
g6142 nand P2_U3067 P2_U3029 ; P2_U5483
g6143 nand P2_U5441 P2_U3067 ; P2_U5484
g6144 nand P2_U3929 P2_U3953 ; P2_U5485
g6145 nand P2_U3068 P2_U3029 ; P2_U5486
g6146 nand P2_U5441 P2_U3068 ; P2_U5487
g6147 nand P2_U3929 P2_U3954 ; P2_U5488
g6148 nand P2_U3063 P2_U3029 ; P2_U5489
g6149 nand P2_U5441 P2_U3063 ; P2_U5490
g6150 nand P2_U3929 P2_U3955 ; P2_U5491
g6151 nand P2_U3077 P2_U3029 ; P2_U5492
g6152 nand P2_U5441 P2_U3077 ; P2_U5493
g6153 nand P2_U3929 P2_U3956 ; P2_U5494
g6154 nand P2_U3078 P2_U3029 ; P2_U5495
g6155 nand P2_U5441 P2_U3078 ; P2_U5496
g6156 nand P2_U3929 P2_U3957 ; P2_U5497
g6157 nand P2_U3070 P2_U3029 ; P2_U5498
g6158 nand P2_U5441 P2_U3070 ; P2_U5499
g6159 nand P2_U3929 P2_U3435 ; P2_U5500
g6160 nand P2_U3083 P2_U3029 ; P2_U5501
g6161 nand P2_U5441 P2_U3083 ; P2_U5502
g6162 nand P2_U3929 P2_U3485 ; P2_U5503
g6163 nand P2_U3084 P2_U3029 ; P2_U5504
g6164 nand P2_U5441 P2_U3084 ; P2_U5505
g6165 nand P2_U3929 P2_U3483 ; P2_U5506
g6166 nand P2_U3071 P2_U3029 ; P2_U5507
g6167 nand P2_U5441 P2_U3071 ; P2_U5508
g6168 nand P2_U3929 P2_U3480 ; P2_U5509
g6169 nand P2_U3075 P2_U3029 ; P2_U5510
g6170 nand P2_U5441 P2_U3075 ; P2_U5511
g6171 nand P2_U3929 P2_U3477 ; P2_U5512
g6172 nand P2_U3076 P2_U3029 ; P2_U5513
g6173 nand P2_U5441 P2_U3076 ; P2_U5514
g6174 nand P2_U3929 P2_U3474 ; P2_U5515
g6175 nand P2_U3081 P2_U3029 ; P2_U5516
g6176 nand P2_U5441 P2_U3081 ; P2_U5517
g6177 nand P2_U3929 P2_U3471 ; P2_U5518
g6178 nand P2_U3082 P2_U3029 ; P2_U5519
g6179 nand P2_U5441 P2_U3082 ; P2_U5520
g6180 nand P2_U3929 P2_U3468 ; P2_U5521
g6181 nand P2_U3074 P2_U3029 ; P2_U5522
g6182 nand P2_U5441 P2_U3074 ; P2_U5523
g6183 nand P2_U3929 P2_U3465 ; P2_U5524
g6184 nand P2_U3065 P2_U3029 ; P2_U5525
g6185 nand P2_U5441 P2_U3065 ; P2_U5526
g6186 nand P2_U3929 P2_U3462 ; P2_U5527
g6187 nand P2_U3064 P2_U3029 ; P2_U5528
g6188 nand P2_U5441 P2_U3064 ; P2_U5529
g6189 nand P2_U3929 P2_U3459 ; P2_U5530
g6190 nand P2_U3080 P2_U3029 ; P2_U5531
g6191 nand P2_U5441 P2_U3080 ; P2_U5532
g6192 nand P2_U3929 P2_U3432 ; P2_U5533
g6193 nand P2_U3079 P2_U3029 ; P2_U5534
g6194 nand P2_U5441 P2_U3079 ; P2_U5535
g6195 nand P2_U3929 P2_U3427 ; P2_U5536
g6196 nand P2_U5438 P2_U3053 ; P2_U5537
g6197 nand P2_U3456 P2_U5537 ; P2_U5538
g6198 nand P2_U3929 P2_U3085 ; P2_U5539
g6199 nand P2_U5658 P2_U3086 ; P2_U5540
g6200 nand P2_U3453 P2_U5537 ; P2_U5541
g6201 nand P2_U3929 P2_U3086 ; P2_U5542
g6202 nand P2_U5658 P2_U3072 ; P2_U5543
g6203 nand P2_U3450 P2_U5537 ; P2_U5544
g6204 nand P2_U3929 P2_U3072 ; P2_U5545
g6205 nand P2_U5658 P2_U3073 ; P2_U5546
g6206 nand P2_U3447 P2_U5537 ; P2_U5547
g6207 nand P2_U3929 P2_U3073 ; P2_U5548
g6208 nand P2_U5658 P2_U3069 ; P2_U5549
g6209 nand P2_U3444 P2_U5537 ; P2_U5550
g6210 nand P2_U3929 P2_U3069 ; P2_U5551
g6211 nand P2_U5658 P2_U3062 ; P2_U5552
g6212 nand P2_U3441 P2_U5537 ; P2_U5553
g6213 nand P2_U3929 P2_U3062 ; P2_U5554
g6214 nand P2_U5658 P2_U3066 ; P2_U5555
g6215 nand P2_U5537 P2_U3347 U69 ; P2_U5556
g6216 nand P2_U3929 P2_U3058 ; P2_U5557
g6217 nand P2_U3959 P2_U5537 ; P2_U5558
g6218 nand P2_U3929 P2_U3061 ; P2_U5559
g6219 nand P2_U3438 P2_U5537 ; P2_U5560
g6220 nand P2_U3929 P2_U3066 ; P2_U5561
g6221 nand P2_U5658 P2_U3070 ; P2_U5562
g6222 nand P2_U3960 P2_U5537 ; P2_U5563
g6223 nand P2_U3929 P2_U3057 ; P2_U5564
g6224 nand P2_U5658 P2_U3056 ; P2_U5565
g6225 nand P2_U3949 P2_U5537 ; P2_U5566
g6226 nand P2_U3929 P2_U3056 ; P2_U5567
g6227 nand P2_U5658 P2_U3055 ; P2_U5568
g6228 nand P2_U3950 P2_U5537 ; P2_U5569
g6229 nand P2_U3929 P2_U3055 ; P2_U5570
g6230 nand P2_U5658 P2_U3059 ; P2_U5571
g6231 nand P2_U3951 P2_U5537 ; P2_U5572
g6232 nand P2_U3929 P2_U3059 ; P2_U5573
g6233 nand P2_U5658 P2_U3060 ; P2_U5574
g6234 nand P2_U3952 P2_U5537 ; P2_U5575
g6235 nand P2_U3929 P2_U3060 ; P2_U5576
g6236 nand P2_U5658 P2_U3067 ; P2_U5577
g6237 nand P2_U3953 P2_U5537 ; P2_U5578
g6238 nand P2_U3929 P2_U3067 ; P2_U5579
g6239 nand P2_U5658 P2_U3068 ; P2_U5580
g6240 nand P2_U3954 P2_U5537 ; P2_U5581
g6241 nand P2_U3929 P2_U3068 ; P2_U5582
g6242 nand P2_U5658 P2_U3063 ; P2_U5583
g6243 nand P2_U3955 P2_U5537 ; P2_U5584
g6244 nand P2_U3929 P2_U3063 ; P2_U5585
g6245 nand P2_U5658 P2_U3077 ; P2_U5586
g6246 nand P2_U3956 P2_U5537 ; P2_U5587
g6247 nand P2_U3929 P2_U3077 ; P2_U5588
g6248 nand P2_U5658 P2_U3078 ; P2_U5589
g6249 nand P2_U3957 P2_U5537 ; P2_U5590
g6250 nand P2_U3929 P2_U3078 ; P2_U5591
g6251 nand P2_U5658 P2_U3083 ; P2_U5592
g6252 nand P2_U3435 P2_U5537 ; P2_U5593
g6253 nand P2_U3929 P2_U3070 ; P2_U5594
g6254 nand P2_U5658 P2_U3080 ; P2_U5595
g6255 nand P2_U3485 P2_U5537 ; P2_U5596
g6256 nand P2_U3929 P2_U3083 ; P2_U5597
g6257 nand P2_U5658 P2_U3084 ; P2_U5598
g6258 nand P2_U3483 P2_U5537 ; P2_U5599
g6259 nand P2_U3929 P2_U3084 ; P2_U5600
g6260 nand P2_U5658 P2_U3071 ; P2_U5601
g6261 nand P2_U3480 P2_U5537 ; P2_U5602
g6262 nand P2_U3929 P2_U3071 ; P2_U5603
g6263 nand P2_U5658 P2_U3075 ; P2_U5604
g6264 nand P2_U3477 P2_U5537 ; P2_U5605
g6265 nand P2_U3929 P2_U3075 ; P2_U5606
g6266 nand P2_U5658 P2_U3076 ; P2_U5607
g6267 nand P2_U3474 P2_U5537 ; P2_U5608
g6268 nand P2_U3929 P2_U3076 ; P2_U5609
g6269 nand P2_U5658 P2_U3081 ; P2_U5610
g6270 nand P2_U3471 P2_U5537 ; P2_U5611
g6271 nand P2_U3929 P2_U3081 ; P2_U5612
g6272 nand P2_U5658 P2_U3082 ; P2_U5613
g6273 nand P2_U3468 P2_U5537 ; P2_U5614
g6274 nand P2_U3929 P2_U3082 ; P2_U5615
g6275 nand P2_U5658 P2_U3074 ; P2_U5616
g6276 nand P2_U3465 P2_U5537 ; P2_U5617
g6277 nand P2_U3929 P2_U3074 ; P2_U5618
g6278 nand P2_U5658 P2_U3065 ; P2_U5619
g6279 nand P2_U3462 P2_U5537 ; P2_U5620
g6280 nand P2_U3929 P2_U3065 ; P2_U5621
g6281 nand P2_U5658 P2_U3064 ; P2_U5622
g6282 nand P2_U3459 P2_U5537 ; P2_U5623
g6283 nand P2_U3929 P2_U3064 ; P2_U5624
g6284 nand P2_U5658 P2_U3085 ; P2_U5625
g6285 nand P2_U3432 P2_U5537 ; P2_U5626
g6286 nand P2_U3929 P2_U3080 ; P2_U5627
g6287 nand P2_U5658 P2_U3079 ; P2_U5628
g6288 nand P2_U3427 P2_U5537 ; P2_U5629
g6289 nand P2_U3929 P2_U3079 ; P2_U5630
g6290 nand P2_U5163 P2_U3088 ; P2_U5631
g6291 nand P2_U3828 P2_U5461 ; P2_U5632
g6292 nand P2_U3972 P2_U3406 ; P2_U5633
g6293 nand P2_U3946 P2_U3972 ; P2_U5634
g6294 nand P2_U5633 P2_U3970 ; P2_U5635
g6295 nand P2_U5634 P2_U3971 ; P2_U5636
g6296 nand P2_U3054 P2_U3945 ; P2_U5637
g6297 nand P2_U3054 P2_U3330 ; P2_U5638
g6298 nand P2_U3961 P2_U3023 ; P2_U5639
g6299 nand P2_U3787 P2_U5163 ; P2_U5640
g6300 nand P2_U6150 P2_U6149 P2_U5163 P2_U3917 ; P2_U5641
g6301 nand P2_U5652 P2_U5646 ; P2_U5642
g6302 nand P2_U3415 P2_U3347 ; P2_U5643
g6303 nand P2_U3879 P2_IR_REG_24__SCAN_IN ; P2_U5644
g6304 nand P2_SUB_1108_U14 P2_IR_REG_31__SCAN_IN ; P2_U5645
g6305 not P2_U3412 ; P2_U5646
g6306 nand P2_U3879 P2_IR_REG_25__SCAN_IN ; P2_U5647
g6307 nand P2_SUB_1108_U112 P2_IR_REG_31__SCAN_IN ; P2_U5648
g6308 not P2_U3413 ; P2_U5649
g6309 nand P2_U3879 P2_IR_REG_26__SCAN_IN ; P2_U5650
g6310 nand P2_SUB_1108_U15 P2_IR_REG_31__SCAN_IN ; P2_U5651
g6311 not P2_U3414 ; P2_U5652
g6312 nand P2_U5646 P2_B_REG_SCAN_IN ; P2_U5653
g6313 nand P2_U3412 P2_U3331 ; P2_U5654
g6314 nand P2_U5654 P2_U5653 ; P2_U5655
g6315 nand P2_U3879 P2_IR_REG_23__SCAN_IN ; P2_U5656
g6316 nand P2_SUB_1108_U13 P2_IR_REG_31__SCAN_IN ; P2_U5657
g6317 not P2_U3415 ; P2_U5658
g6318 nand P2_U3880 P2_D_REG_0__SCAN_IN ; P2_U5659
g6319 nand P2_U3967 P2_U4077 ; P2_U5660
g6320 nand P2_U3880 P2_D_REG_1__SCAN_IN ; P2_U5661
g6321 nand P2_U3967 P2_U4078 ; P2_U5662
g6322 nand P2_U3879 P2_IR_REG_22__SCAN_IN ; P2_U5663
g6323 nand P2_SUB_1108_U114 P2_IR_REG_31__SCAN_IN ; P2_U5664
g6324 not P2_U3420 ; P2_U5665
g6325 nand P2_U3879 P2_IR_REG_19__SCAN_IN ; P2_U5666
g6326 nand P2_SUB_1108_U123 P2_IR_REG_31__SCAN_IN ; P2_U5667
g6327 not P2_U3424 ; P2_U5668
g6328 nand P2_U3879 P2_IR_REG_20__SCAN_IN ; P2_U5669
g6329 nand P2_SUB_1108_U119 P2_IR_REG_31__SCAN_IN ; P2_U5670
g6330 not P2_U3418 ; P2_U5671
g6331 nand P2_U3879 P2_IR_REG_21__SCAN_IN ; P2_U5672
g6332 nand P2_SUB_1108_U116 P2_IR_REG_31__SCAN_IN ; P2_U5673
g6333 not P2_U3419 ; P2_U5674
g6334 nand P2_U3879 P2_IR_REG_30__SCAN_IN ; P2_U5675
g6335 nand P2_SUB_1108_U104 P2_IR_REG_31__SCAN_IN ; P2_U5676
g6336 not P2_U3421 ; P2_U5677
g6337 nand P2_U3879 P2_IR_REG_29__SCAN_IN ; P2_U5678
g6338 nand P2_SUB_1108_U16 P2_IR_REG_31__SCAN_IN ; P2_U5679
g6339 not P2_U3422 ; P2_U5680
g6340 nand P2_U3879 P2_IR_REG_28__SCAN_IN ; P2_U5681
g6341 nand P2_SUB_1108_U107 P2_IR_REG_31__SCAN_IN ; P2_U5682
g6342 not P2_U3423 ; P2_U5683
g6343 nand P2_U3879 P2_IR_REG_0__SCAN_IN ; P2_U5684
g6344 nand P2_IR_REG_0__SCAN_IN P2_IR_REG_31__SCAN_IN ; P2_U5685
g6345 nand P2_U3879 P2_IR_REG_27__SCAN_IN ; P2_U5686
g6346 nand P2_SUB_1108_U110 P2_IR_REG_31__SCAN_IN ; P2_U5687
g6347 not P2_U3426 ; P2_U5688
g6348 nand U93 P2_U3347 ; P2_U5689
g6349 nand P2_U3425 P2_U3945 ; P2_U5690
g6350 not P2_U3427 ; P2_U5691
g6351 nand P2_U3420 P2_U5674 ; P2_U5692
g6352 nand P2_U5665 P2_U4109 ; P2_U5693
g6353 nand P2_U4076 P2_D_REG_1__SCAN_IN ; P2_U5694
g6354 nand P2_U4078 P2_U3333 ; P2_U5695
g6355 not P2_U3429 ; P2_U5696
g6356 nand P2_U5642 P2_U3333 ; P2_U5697
g6357 nand P2_U4076 P2_D_REG_0__SCAN_IN ; P2_U5698
g6358 not P2_U3428 ; P2_U5699
g6359 nand P2_U3881 P2_REG0_REG_0__SCAN_IN ; P2_U5700
g6360 nand P2_U3966 P2_U4129 ; P2_U5701
g6361 nand P2_U3879 P2_IR_REG_1__SCAN_IN ; P2_U5702
g6362 nand P2_SUB_1108_U42 P2_IR_REG_31__SCAN_IN ; P2_U5703
g6363 nand U82 P2_U3347 ; P2_U5704
g6364 nand P2_U3431 P2_U3945 ; P2_U5705
g6365 not P2_U3432 ; P2_U5706
g6366 nand P2_U3881 P2_REG0_REG_1__SCAN_IN ; P2_U5707
g6367 nand P2_U3966 P2_U4153 ; P2_U5708
g6368 nand P2_U3879 P2_IR_REG_2__SCAN_IN ; P2_U5709
g6369 nand P2_SUB_1108_U17 P2_IR_REG_31__SCAN_IN ; P2_U5710
g6370 nand U71 P2_U3347 ; P2_U5711
g6371 nand P2_U3434 P2_U3945 ; P2_U5712
g6372 not P2_U3435 ; P2_U5713
g6373 nand P2_U3881 P2_REG0_REG_2__SCAN_IN ; P2_U5714
g6374 nand P2_U3966 P2_U4172 ; P2_U5715
g6375 nand P2_U3879 P2_IR_REG_3__SCAN_IN ; P2_U5716
g6376 nand P2_SUB_1108_U18 P2_IR_REG_31__SCAN_IN ; P2_U5717
g6377 nand U68 P2_U3347 ; P2_U5718
g6378 nand P2_U3437 P2_U3945 ; P2_U5719
g6379 not P2_U3438 ; P2_U5720
g6380 nand P2_U3881 P2_REG0_REG_3__SCAN_IN ; P2_U5721
g6381 nand P2_U3966 P2_U4191 ; P2_U5722
g6382 nand P2_U3879 P2_IR_REG_4__SCAN_IN ; P2_U5723
g6383 nand P2_SUB_1108_U19 P2_IR_REG_31__SCAN_IN ; P2_U5724
g6384 nand U67 P2_U3347 ; P2_U5725
g6385 nand P2_U3440 P2_U3945 ; P2_U5726
g6386 not P2_U3441 ; P2_U5727
g6387 nand P2_U3881 P2_REG0_REG_4__SCAN_IN ; P2_U5728
g6388 nand P2_U3966 P2_U4210 ; P2_U5729
g6389 nand P2_U3879 P2_IR_REG_5__SCAN_IN ; P2_U5730
g6390 nand P2_SUB_1108_U101 P2_IR_REG_31__SCAN_IN ; P2_U5731
g6391 nand U66 P2_U3347 ; P2_U5732
g6392 nand P2_U3443 P2_U3945 ; P2_U5733
g6393 not P2_U3444 ; P2_U5734
g6394 nand P2_U3881 P2_REG0_REG_5__SCAN_IN ; P2_U5735
g6395 nand P2_U3966 P2_U4229 ; P2_U5736
g6396 nand P2_U3879 P2_IR_REG_6__SCAN_IN ; P2_U5737
g6397 nand P2_SUB_1108_U20 P2_IR_REG_31__SCAN_IN ; P2_U5738
g6398 nand U65 P2_U3347 ; P2_U5739
g6399 nand P2_U3446 P2_U3945 ; P2_U5740
g6400 not P2_U3447 ; P2_U5741
g6401 nand P2_U3881 P2_REG0_REG_6__SCAN_IN ; P2_U5742
g6402 nand P2_U3966 P2_U4248 ; P2_U5743
g6403 nand P2_U3879 P2_IR_REG_7__SCAN_IN ; P2_U5744
g6404 nand P2_SUB_1108_U21 P2_IR_REG_31__SCAN_IN ; P2_U5745
g6405 nand U64 P2_U3347 ; P2_U5746
g6406 nand P2_U3449 P2_U3945 ; P2_U5747
g6407 not P2_U3450 ; P2_U5748
g6408 nand P2_U3881 P2_REG0_REG_7__SCAN_IN ; P2_U5749
g6409 nand P2_U3966 P2_U4267 ; P2_U5750
g6410 nand P2_U3879 P2_IR_REG_8__SCAN_IN ; P2_U5751
g6411 nand P2_SUB_1108_U22 P2_IR_REG_31__SCAN_IN ; P2_U5752
g6412 nand U63 P2_U3347 ; P2_U5753
g6413 nand P2_U3452 P2_U3945 ; P2_U5754
g6414 not P2_U3453 ; P2_U5755
g6415 nand P2_U3881 P2_REG0_REG_8__SCAN_IN ; P2_U5756
g6416 nand P2_U3966 P2_U4286 ; P2_U5757
g6417 nand P2_U3879 P2_IR_REG_9__SCAN_IN ; P2_U5758
g6418 nand P2_SUB_1108_U99 P2_IR_REG_31__SCAN_IN ; P2_U5759
g6419 nand U62 P2_U3347 ; P2_U5760
g6420 nand P2_U3455 P2_U3945 ; P2_U5761
g6421 not P2_U3456 ; P2_U5762
g6422 nand P2_U3881 P2_REG0_REG_9__SCAN_IN ; P2_U5763
g6423 nand P2_U3966 P2_U4305 ; P2_U5764
g6424 nand P2_U3879 P2_IR_REG_10__SCAN_IN ; P2_U5765
g6425 nand P2_SUB_1108_U6 P2_IR_REG_31__SCAN_IN ; P2_U5766
g6426 nand U92 P2_U3347 ; P2_U5767
g6427 nand P2_U3458 P2_U3945 ; P2_U5768
g6428 not P2_U3459 ; P2_U5769
g6429 nand P2_U3881 P2_REG0_REG_10__SCAN_IN ; P2_U5770
g6430 nand P2_U3966 P2_U4324 ; P2_U5771
g6431 nand P2_U3879 P2_IR_REG_11__SCAN_IN ; P2_U5772
g6432 nand P2_SUB_1108_U7 P2_IR_REG_31__SCAN_IN ; P2_U5773
g6433 nand U91 P2_U3347 ; P2_U5774
g6434 nand P2_U3461 P2_U3945 ; P2_U5775
g6435 not P2_U3462 ; P2_U5776
g6436 nand P2_U3881 P2_REG0_REG_11__SCAN_IN ; P2_U5777
g6437 nand P2_U3966 P2_U4343 ; P2_U5778
g6438 nand P2_U3879 P2_IR_REG_12__SCAN_IN ; P2_U5779
g6439 nand P2_SUB_1108_U8 P2_IR_REG_31__SCAN_IN ; P2_U5780
g6440 nand U90 P2_U3347 ; P2_U5781
g6441 nand P2_U3464 P2_U3945 ; P2_U5782
g6442 not P2_U3465 ; P2_U5783
g6443 nand P2_U3881 P2_REG0_REG_12__SCAN_IN ; P2_U5784
g6444 nand P2_U3966 P2_U4362 ; P2_U5785
g6445 nand P2_U3879 P2_IR_REG_13__SCAN_IN ; P2_U5786
g6446 nand P2_SUB_1108_U127 P2_IR_REG_31__SCAN_IN ; P2_U5787
g6447 nand U89 P2_U3347 ; P2_U5788
g6448 nand P2_U3467 P2_U3945 ; P2_U5789
g6449 not P2_U3468 ; P2_U5790
g6450 nand P2_U3881 P2_REG0_REG_13__SCAN_IN ; P2_U5791
g6451 nand P2_U3966 P2_U4381 ; P2_U5792
g6452 nand P2_U3879 P2_IR_REG_14__SCAN_IN ; P2_U5793
g6453 nand P2_SUB_1108_U9 P2_IR_REG_31__SCAN_IN ; P2_U5794
g6454 nand U88 P2_U3347 ; P2_U5795
g6455 nand P2_U3470 P2_U3945 ; P2_U5796
g6456 not P2_U3471 ; P2_U5797
g6457 nand P2_U3881 P2_REG0_REG_14__SCAN_IN ; P2_U5798
g6458 nand P2_U3966 P2_U4400 ; P2_U5799
g6459 nand P2_U3879 P2_IR_REG_15__SCAN_IN ; P2_U5800
g6460 nand P2_SUB_1108_U10 P2_IR_REG_31__SCAN_IN ; P2_U5801
g6461 nand U87 P2_U3347 ; P2_U5802
g6462 nand P2_U3473 P2_U3945 ; P2_U5803
g6463 not P2_U3474 ; P2_U5804
g6464 nand P2_U3881 P2_REG0_REG_15__SCAN_IN ; P2_U5805
g6465 nand P2_U3966 P2_U4419 ; P2_U5806
g6466 nand P2_U3879 P2_IR_REG_16__SCAN_IN ; P2_U5807
g6467 nand P2_SUB_1108_U11 P2_IR_REG_31__SCAN_IN ; P2_U5808
g6468 nand U86 P2_U3347 ; P2_U5809
g6469 nand P2_U3476 P2_U3945 ; P2_U5810
g6470 not P2_U3477 ; P2_U5811
g6471 nand P2_U3881 P2_REG0_REG_16__SCAN_IN ; P2_U5812
g6472 nand P2_U3966 P2_U4438 ; P2_U5813
g6473 nand P2_U3879 P2_IR_REG_17__SCAN_IN ; P2_U5814
g6474 nand P2_SUB_1108_U125 P2_IR_REG_31__SCAN_IN ; P2_U5815
g6475 nand U85 P2_U3347 ; P2_U5816
g6476 nand P2_U3479 P2_U3945 ; P2_U5817
g6477 not P2_U3480 ; P2_U5818
g6478 nand P2_U3881 P2_REG0_REG_17__SCAN_IN ; P2_U5819
g6479 nand P2_U3966 P2_U4457 ; P2_U5820
g6480 nand P2_U3879 P2_IR_REG_18__SCAN_IN ; P2_U5821
g6481 nand P2_SUB_1108_U12 P2_IR_REG_31__SCAN_IN ; P2_U5822
g6482 nand U84 P2_U3347 ; P2_U5823
g6483 nand P2_U3482 P2_U3945 ; P2_U5824
g6484 not P2_U3483 ; P2_U5825
g6485 nand P2_U3881 P2_REG0_REG_18__SCAN_IN ; P2_U5826
g6486 nand P2_U3966 P2_U4476 ; P2_U5827
g6487 nand U83 P2_U3347 ; P2_U5828
g6488 nand P2_U3424 P2_U3945 ; P2_U5829
g6489 not P2_U3485 ; P2_U5830
g6490 nand P2_U3881 P2_REG0_REG_19__SCAN_IN ; P2_U5831
g6491 nand P2_U3966 P2_U4495 ; P2_U5832
g6492 nand P2_U3881 P2_REG0_REG_20__SCAN_IN ; P2_U5833
g6493 nand P2_U3966 P2_U4514 ; P2_U5834
g6494 nand P2_U3881 P2_REG0_REG_21__SCAN_IN ; P2_U5835
g6495 nand P2_U3966 P2_U4533 ; P2_U5836
g6496 nand P2_U3881 P2_REG0_REG_22__SCAN_IN ; P2_U5837
g6497 nand P2_U3966 P2_U4552 ; P2_U5838
g6498 nand P2_U3881 P2_REG0_REG_23__SCAN_IN ; P2_U5839
g6499 nand P2_U3966 P2_U4571 ; P2_U5840
g6500 nand P2_U3881 P2_REG0_REG_24__SCAN_IN ; P2_U5841
g6501 nand P2_U3966 P2_U4590 ; P2_U5842
g6502 nand P2_U3881 P2_REG0_REG_25__SCAN_IN ; P2_U5843
g6503 nand P2_U3966 P2_U4609 ; P2_U5844
g6504 nand P2_U3881 P2_REG0_REG_26__SCAN_IN ; P2_U5845
g6505 nand P2_U3966 P2_U4628 ; P2_U5846
g6506 nand P2_U3881 P2_REG0_REG_27__SCAN_IN ; P2_U5847
g6507 nand P2_U3966 P2_U4647 ; P2_U5848
g6508 nand P2_U3881 P2_REG0_REG_28__SCAN_IN ; P2_U5849
g6509 nand P2_U3966 P2_U4666 ; P2_U5850
g6510 nand P2_U3881 P2_REG0_REG_29__SCAN_IN ; P2_U5851
g6511 nand P2_U3966 P2_U4686 ; P2_U5852
g6512 nand P2_U3881 P2_REG0_REG_30__SCAN_IN ; P2_U5853
g6513 nand P2_U3966 P2_U4693 ; P2_U5854
g6514 nand P2_U3881 P2_REG0_REG_31__SCAN_IN ; P2_U5855
g6515 nand P2_U3966 P2_U4696 ; P2_U5856
g6516 nand P2_U3882 P2_REG1_REG_0__SCAN_IN ; P2_U5857
g6517 nand P2_U3965 P2_U4129 ; P2_U5858
g6518 nand P2_U3882 P2_REG1_REG_1__SCAN_IN ; P2_U5859
g6519 nand P2_U3965 P2_U4153 ; P2_U5860
g6520 nand P2_U3882 P2_REG1_REG_2__SCAN_IN ; P2_U5861
g6521 nand P2_U3965 P2_U4172 ; P2_U5862
g6522 nand P2_U3882 P2_REG1_REG_3__SCAN_IN ; P2_U5863
g6523 nand P2_U3965 P2_U4191 ; P2_U5864
g6524 nand P2_U3882 P2_REG1_REG_4__SCAN_IN ; P2_U5865
g6525 nand P2_U3965 P2_U4210 ; P2_U5866
g6526 nand P2_U3882 P2_REG1_REG_5__SCAN_IN ; P2_U5867
g6527 nand P2_U3965 P2_U4229 ; P2_U5868
g6528 nand P2_U3882 P2_REG1_REG_6__SCAN_IN ; P2_U5869
g6529 nand P2_U3965 P2_U4248 ; P2_U5870
g6530 nand P2_U3882 P2_REG1_REG_7__SCAN_IN ; P2_U5871
g6531 nand P2_U3965 P2_U4267 ; P2_U5872
g6532 nand P2_U3882 P2_REG1_REG_8__SCAN_IN ; P2_U5873
g6533 nand P2_U3965 P2_U4286 ; P2_U5874
g6534 nand P2_U3882 P2_REG1_REG_9__SCAN_IN ; P2_U5875
g6535 nand P2_U3965 P2_U4305 ; P2_U5876
g6536 nand P2_U3882 P2_REG1_REG_10__SCAN_IN ; P2_U5877
g6537 nand P2_U3965 P2_U4324 ; P2_U5878
g6538 nand P2_U3882 P2_REG1_REG_11__SCAN_IN ; P2_U5879
g6539 nand P2_U3965 P2_U4343 ; P2_U5880
g6540 nand P2_U3882 P2_REG1_REG_12__SCAN_IN ; P2_U5881
g6541 nand P2_U3965 P2_U4362 ; P2_U5882
g6542 nand P2_U3882 P2_REG1_REG_13__SCAN_IN ; P2_U5883
g6543 nand P2_U3965 P2_U4381 ; P2_U5884
g6544 nand P2_U3882 P2_REG1_REG_14__SCAN_IN ; P2_U5885
g6545 nand P2_U3965 P2_U4400 ; P2_U5886
g6546 nand P2_U3882 P2_REG1_REG_15__SCAN_IN ; P2_U5887
g6547 nand P2_U3965 P2_U4419 ; P2_U5888
g6548 nand P2_U3882 P2_REG1_REG_16__SCAN_IN ; P2_U5889
g6549 nand P2_U3965 P2_U4438 ; P2_U5890
g6550 nand P2_U3882 P2_REG1_REG_17__SCAN_IN ; P2_U5891
g6551 nand P2_U3965 P2_U4457 ; P2_U5892
g6552 nand P2_U3882 P2_REG1_REG_18__SCAN_IN ; P2_U5893
g6553 nand P2_U3965 P2_U4476 ; P2_U5894
g6554 nand P2_U3882 P2_REG1_REG_19__SCAN_IN ; P2_U5895
g6555 nand P2_U3965 P2_U4495 ; P2_U5896
g6556 nand P2_U3882 P2_REG1_REG_20__SCAN_IN ; P2_U5897
g6557 nand P2_U3965 P2_U4514 ; P2_U5898
g6558 nand P2_U3882 P2_REG1_REG_21__SCAN_IN ; P2_U5899
g6559 nand P2_U3965 P2_U4533 ; P2_U5900
g6560 nand P2_U3882 P2_REG1_REG_22__SCAN_IN ; P2_U5901
g6561 nand P2_U3965 P2_U4552 ; P2_U5902
g6562 nand P2_U3882 P2_REG1_REG_23__SCAN_IN ; P2_U5903
g6563 nand P2_U3965 P2_U4571 ; P2_U5904
g6564 nand P2_U3882 P2_REG1_REG_24__SCAN_IN ; P2_U5905
g6565 nand P2_U3965 P2_U4590 ; P2_U5906
g6566 nand P2_U3882 P2_REG1_REG_25__SCAN_IN ; P2_U5907
g6567 nand P2_U3965 P2_U4609 ; P2_U5908
g6568 nand P2_U3882 P2_REG1_REG_26__SCAN_IN ; P2_U5909
g6569 nand P2_U3965 P2_U4628 ; P2_U5910
g6570 nand P2_U3882 P2_REG1_REG_27__SCAN_IN ; P2_U5911
g6571 nand P2_U3965 P2_U4647 ; P2_U5912
g6572 nand P2_U3882 P2_REG1_REG_28__SCAN_IN ; P2_U5913
g6573 nand P2_U3965 P2_U4666 ; P2_U5914
g6574 nand P2_U3882 P2_REG1_REG_29__SCAN_IN ; P2_U5915
g6575 nand P2_U3965 P2_U4686 ; P2_U5916
g6576 nand P2_U3882 P2_REG1_REG_30__SCAN_IN ; P2_U5917
g6577 nand P2_U3965 P2_U4693 ; P2_U5918
g6578 nand P2_U3882 P2_REG1_REG_31__SCAN_IN ; P2_U5919
g6579 nand P2_U3965 P2_U4696 ; P2_U5920
g6580 nand P2_U3391 P2_REG2_REG_0__SCAN_IN ; P2_U5921
g6581 nand P2_U3964 P2_U3348 ; P2_U5922
g6582 nand P2_U3391 P2_REG2_REG_1__SCAN_IN ; P2_U5923
g6583 nand P2_U3964 P2_U3349 ; P2_U5924
g6584 nand P2_U3391 P2_REG2_REG_2__SCAN_IN ; P2_U5925
g6585 nand P2_U3964 P2_U3350 ; P2_U5926
g6586 nand P2_U3391 P2_REG2_REG_3__SCAN_IN ; P2_U5927
g6587 nand P2_U3964 P2_U3351 ; P2_U5928
g6588 nand P2_U3391 P2_REG2_REG_4__SCAN_IN ; P2_U5929
g6589 nand P2_U3964 P2_U3352 ; P2_U5930
g6590 nand P2_U3391 P2_REG2_REG_5__SCAN_IN ; P2_U5931
g6591 nand P2_U3964 P2_U3353 ; P2_U5932
g6592 nand P2_U3391 P2_REG2_REG_6__SCAN_IN ; P2_U5933
g6593 nand P2_U3964 P2_U3354 ; P2_U5934
g6594 nand P2_U3391 P2_REG2_REG_7__SCAN_IN ; P2_U5935
g6595 nand P2_U3964 P2_U3355 ; P2_U5936
g6596 nand P2_U3391 P2_REG2_REG_8__SCAN_IN ; P2_U5937
g6597 nand P2_U3964 P2_U3356 ; P2_U5938
g6598 nand P2_U3391 P2_REG2_REG_9__SCAN_IN ; P2_U5939
g6599 nand P2_U3964 P2_U3357 ; P2_U5940
g6600 nand P2_U3391 P2_REG2_REG_10__SCAN_IN ; P2_U5941
g6601 nand P2_U3964 P2_U3358 ; P2_U5942
g6602 nand P2_U3391 P2_REG2_REG_11__SCAN_IN ; P2_U5943
g6603 nand P2_U3964 P2_U3359 ; P2_U5944
g6604 nand P2_U3391 P2_REG2_REG_12__SCAN_IN ; P2_U5945
g6605 nand P2_U3964 P2_U3360 ; P2_U5946
g6606 nand P2_U3391 P2_REG2_REG_13__SCAN_IN ; P2_U5947
g6607 nand P2_U3964 P2_U3361 ; P2_U5948
g6608 nand P2_U3391 P2_REG2_REG_14__SCAN_IN ; P2_U5949
g6609 nand P2_U3964 P2_U3362 ; P2_U5950
g6610 nand P2_U3391 P2_REG2_REG_15__SCAN_IN ; P2_U5951
g6611 nand P2_U3964 P2_U3363 ; P2_U5952
g6612 nand P2_U3391 P2_REG2_REG_16__SCAN_IN ; P2_U5953
g6613 nand P2_U3964 P2_U3364 ; P2_U5954
g6614 nand P2_U3391 P2_REG2_REG_17__SCAN_IN ; P2_U5955
g6615 nand P2_U3964 P2_U3365 ; P2_U5956
g6616 nand P2_U3391 P2_REG2_REG_18__SCAN_IN ; P2_U5957
g6617 nand P2_U3964 P2_U3366 ; P2_U5958
g6618 nand P2_U3391 P2_REG2_REG_19__SCAN_IN ; P2_U5959
g6619 nand P2_U3964 P2_U3367 ; P2_U5960
g6620 nand P2_U3391 P2_REG2_REG_20__SCAN_IN ; P2_U5961
g6621 nand P2_U3964 P2_U3369 ; P2_U5962
g6622 nand P2_U3391 P2_REG2_REG_21__SCAN_IN ; P2_U5963
g6623 nand P2_U3964 P2_U3371 ; P2_U5964
g6624 nand P2_U3391 P2_REG2_REG_22__SCAN_IN ; P2_U5965
g6625 nand P2_U3964 P2_U3373 ; P2_U5966
g6626 nand P2_U3391 P2_REG2_REG_23__SCAN_IN ; P2_U5967
g6627 nand P2_U3964 P2_U3375 ; P2_U5968
g6628 nand P2_U3391 P2_REG2_REG_24__SCAN_IN ; P2_U5969
g6629 nand P2_U3964 P2_U3377 ; P2_U5970
g6630 nand P2_U3391 P2_REG2_REG_25__SCAN_IN ; P2_U5971
g6631 nand P2_U3964 P2_U3379 ; P2_U5972
g6632 nand P2_U3391 P2_REG2_REG_26__SCAN_IN ; P2_U5973
g6633 nand P2_U3964 P2_U3381 ; P2_U5974
g6634 nand P2_U3391 P2_REG2_REG_27__SCAN_IN ; P2_U5975
g6635 nand P2_U3964 P2_U3383 ; P2_U5976
g6636 nand P2_U3391 P2_REG2_REG_28__SCAN_IN ; P2_U5977
g6637 nand P2_U3964 P2_U3385 ; P2_U5978
g6638 nand P2_U3391 P2_REG2_REG_29__SCAN_IN ; P2_U5979
g6639 nand P2_U3964 P2_U3387 ; P2_U5980
g6640 nand P2_U3391 P2_REG2_REG_30__SCAN_IN ; P2_U5981
g6641 nand P2_U3968 P2_U3964 ; P2_U5982
g6642 nand P2_U3391 P2_REG2_REG_31__SCAN_IN ; P2_U5983
g6643 nand P2_U3968 P2_U3964 ; P2_U5984
g6644 nand P2_U3400 P2_DATAO_REG_0__SCAN_IN ; P2_U5985
g6645 nand P2_U3947 P2_U3079 ; P2_U5986
g6646 nand P2_U3400 P2_DATAO_REG_1__SCAN_IN ; P2_U5987
g6647 nand P2_U3947 P2_U3080 ; P2_U5988
g6648 nand P2_U3400 P2_DATAO_REG_2__SCAN_IN ; P2_U5989
g6649 nand P2_U3947 P2_U3070 ; P2_U5990
g6650 nand P2_U3400 P2_DATAO_REG_3__SCAN_IN ; P2_U5991
g6651 nand P2_U3947 P2_U3066 ; P2_U5992
g6652 nand P2_U3400 P2_DATAO_REG_4__SCAN_IN ; P2_U5993
g6653 nand P2_U3947 P2_U3062 ; P2_U5994
g6654 nand P2_U3400 P2_DATAO_REG_5__SCAN_IN ; P2_U5995
g6655 nand P2_U3947 P2_U3069 ; P2_U5996
g6656 nand P2_U3400 P2_DATAO_REG_6__SCAN_IN ; P2_U5997
g6657 nand P2_U3947 P2_U3073 ; P2_U5998
g6658 nand P2_U3400 P2_DATAO_REG_7__SCAN_IN ; P2_U5999
g6659 nand P2_U3947 P2_U3072 ; P2_U6000
g6660 nand P2_U3400 P2_DATAO_REG_8__SCAN_IN ; P2_U6001
g6661 nand P2_U3947 P2_U3086 ; P2_U6002
g6662 nand P2_U3400 P2_DATAO_REG_9__SCAN_IN ; P2_U6003
g6663 nand P2_U3947 P2_U3085 ; P2_U6004
g6664 nand P2_U3400 P2_DATAO_REG_10__SCAN_IN ; P2_U6005
g6665 nand P2_U3947 P2_U3064 ; P2_U6006
g6666 nand P2_U3400 P2_DATAO_REG_11__SCAN_IN ; P2_U6007
g6667 nand P2_U3947 P2_U3065 ; P2_U6008
g6668 nand P2_U3400 P2_DATAO_REG_12__SCAN_IN ; P2_U6009
g6669 nand P2_U3947 P2_U3074 ; P2_U6010
g6670 nand P2_U3400 P2_DATAO_REG_13__SCAN_IN ; P2_U6011
g6671 nand P2_U3947 P2_U3082 ; P2_U6012
g6672 nand P2_U3400 P2_DATAO_REG_14__SCAN_IN ; P2_U6013
g6673 nand P2_U3947 P2_U3081 ; P2_U6014
g6674 nand P2_U3400 P2_DATAO_REG_15__SCAN_IN ; P2_U6015
g6675 nand P2_U3947 P2_U3076 ; P2_U6016
g6676 nand P2_U3400 P2_DATAO_REG_16__SCAN_IN ; P2_U6017
g6677 nand P2_U3947 P2_U3075 ; P2_U6018
g6678 nand P2_U3400 P2_DATAO_REG_17__SCAN_IN ; P2_U6019
g6679 nand P2_U3947 P2_U3071 ; P2_U6020
g6680 nand P2_U3400 P2_DATAO_REG_18__SCAN_IN ; P2_U6021
g6681 nand P2_U3947 P2_U3084 ; P2_U6022
g6682 nand P2_U3400 P2_DATAO_REG_19__SCAN_IN ; P2_U6023
g6683 nand P2_U3947 P2_U3083 ; P2_U6024
g6684 nand P2_U3400 P2_DATAO_REG_20__SCAN_IN ; P2_U6025
g6685 nand P2_U3947 P2_U3078 ; P2_U6026
g6686 nand P2_U3400 P2_DATAO_REG_21__SCAN_IN ; P2_U6027
g6687 nand P2_U3947 P2_U3077 ; P2_U6028
g6688 nand P2_U3400 P2_DATAO_REG_22__SCAN_IN ; P2_U6029
g6689 nand P2_U3947 P2_U3063 ; P2_U6030
g6690 nand P2_U3400 P2_DATAO_REG_23__SCAN_IN ; P2_U6031
g6691 nand P2_U3947 P2_U3068 ; P2_U6032
g6692 nand P2_U3400 P2_DATAO_REG_24__SCAN_IN ; P2_U6033
g6693 nand P2_U3947 P2_U3067 ; P2_U6034
g6694 nand P2_U3400 P2_DATAO_REG_25__SCAN_IN ; P2_U6035
g6695 nand P2_U3947 P2_U3060 ; P2_U6036
g6696 nand P2_U3400 P2_DATAO_REG_26__SCAN_IN ; P2_U6037
g6697 nand P2_U3947 P2_U3059 ; P2_U6038
g6698 nand P2_U3400 P2_DATAO_REG_27__SCAN_IN ; P2_U6039
g6699 nand P2_U3947 P2_U3055 ; P2_U6040
g6700 nand P2_U3400 P2_DATAO_REG_28__SCAN_IN ; P2_U6041
g6701 nand P2_U3947 P2_U3056 ; P2_U6042
g6702 nand P2_U3400 P2_DATAO_REG_29__SCAN_IN ; P2_U6043
g6703 nand P2_U3947 P2_U3057 ; P2_U6044
g6704 nand P2_U3400 P2_DATAO_REG_30__SCAN_IN ; P2_U6045
g6705 nand P2_U3947 P2_U3061 ; P2_U6046
g6706 nand P2_U3400 P2_DATAO_REG_31__SCAN_IN ; P2_U6047
g6707 nand P2_U3947 P2_U3058 ; P2_U6048
g6708 nand P2_R1312_U18 P2_U5157 ; P2_U6049
g6709 nand P2_U5161 P2_U3916 ; P2_U6050
g6710 nand P2_U5658 P2_U3403 ; P2_U6051
g6711 nand P2_U3420 P2_U3415 ; P2_U6052
g6712 nand P2_U3960 P2_U3057 ; P2_U6053
g6713 nand P2_U3386 P2_U4652 ; P2_U6054
g6714 nand P2_U6054 P2_U6053 ; P2_U6055
g6715 nand P2_U3949 P2_U3056 ; P2_U6056
g6716 nand P2_U3384 P2_U4633 ; P2_U6057
g6717 nand P2_U6057 P2_U6056 ; P2_U6058
g6718 nand P2_U3950 P2_U3055 ; P2_U6059
g6719 nand P2_U3382 P2_U4614 ; P2_U6060
g6720 nand P2_U6060 P2_U6059 ; P2_U6061
g6721 nand P2_U3953 P2_U3067 ; P2_U6062
g6722 nand P2_U3376 P2_U4557 ; P2_U6063
g6723 nand P2_U6063 P2_U6062 ; P2_U6064
g6724 nand P2_U3954 P2_U3068 ; P2_U6065
g6725 nand P2_U3374 P2_U4538 ; P2_U6066
g6726 nand P2_U6066 P2_U6065 ; P2_U6067
g6727 nand P2_U3956 P2_U3077 ; P2_U6068
g6728 nand P2_U3370 P2_U4500 ; P2_U6069
g6729 nand P2_U6069 P2_U6068 ; P2_U6070
g6730 nand P2_U3955 P2_U3063 ; P2_U6071
g6731 nand P2_U3372 P2_U4519 ; P2_U6072
g6732 nand P2_U6072 P2_U6071 ; P2_U6073
g6733 nand P2_U3952 P2_U3060 ; P2_U6074
g6734 nand P2_U3378 P2_U4576 ; P2_U6075
g6735 nand P2_U6075 P2_U6074 ; P2_U6076
g6736 nand P2_U3951 P2_U3059 ; P2_U6077
g6737 nand P2_U3380 P2_U4595 ; P2_U6078
g6738 nand P2_U6078 P2_U6077 ; P2_U6079
g6739 nand P2_U3959 P2_U3061 ; P2_U6080
g6740 nand P2_U3388 P2_U4670 ; P2_U6081
g6741 nand P2_U6081 P2_U6080 ; P2_U6082
g6742 nand P2_U3958 P2_U3058 ; P2_U6083
g6743 nand P2_U3389 P2_U4690 ; P2_U6084
g6744 nand P2_U6084 P2_U6083 ; P2_U6085
g6745 nand P2_U5797 P2_U4367 ; P2_U6086
g6746 nand P2_U3471 P2_U3081 ; P2_U6087
g6747 nand P2_U6087 P2_U6086 ; P2_U6088
g6748 nand P2_U5706 P2_U4115 ; P2_U6089
g6749 nand P2_U3432 P2_U3080 ; P2_U6090
g6750 nand P2_U6090 P2_U6089 ; P2_U6091
g6751 nand P2_U5691 P2_U4139 ; P2_U6092
g6752 nand P2_U3427 P2_U3079 ; P2_U6093
g6753 nand P2_U6093 P2_U6092 ; P2_U6094
g6754 nand P2_U5804 P2_U4386 ; P2_U6095
g6755 nand P2_U3474 P2_U3076 ; P2_U6096
g6756 nand P2_U6096 P2_U6095 ; P2_U6097
g6757 nand P2_U5755 P2_U4253 ; P2_U6098
g6758 nand P2_U3453 P2_U3086 ; P2_U6099
g6759 nand P2_U6099 P2_U6098 ; P2_U6100
g6760 nand P2_U5762 P2_U4272 ; P2_U6101
g6761 nand P2_U3456 P2_U3085 ; P2_U6102
g6762 nand P2_U6102 P2_U6101 ; P2_U6103
g6763 nand P2_U5790 P2_U4348 ; P2_U6104
g6764 nand P2_U3468 P2_U3082 ; P2_U6105
g6765 nand P2_U6105 P2_U6104 ; P2_U6106
g6766 nand P2_U5825 P2_U4443 ; P2_U6107
g6767 nand P2_U3483 P2_U3084 ; P2_U6108
g6768 nand P2_U6108 P2_U6107 ; P2_U6109
g6769 nand P2_U5811 P2_U4405 ; P2_U6110
g6770 nand P2_U3477 P2_U3075 ; P2_U6111
g6771 nand P2_U6111 P2_U6110 ; P2_U6112
g6772 nand P2_U5783 P2_U4329 ; P2_U6113
g6773 nand P2_U3465 P2_U3074 ; P2_U6114
g6774 nand P2_U6114 P2_U6113 ; P2_U6115
g6775 nand P2_U5741 P2_U4215 ; P2_U6116
g6776 nand P2_U3447 P2_U3073 ; P2_U6117
g6777 nand P2_U6117 P2_U6116 ; P2_U6118
g6778 nand P2_U5748 P2_U4234 ; P2_U6119
g6779 nand P2_U3450 P2_U3072 ; P2_U6120
g6780 nand P2_U6120 P2_U6119 ; P2_U6121
g6781 nand P2_U5734 P2_U4196 ; P2_U6122
g6782 nand P2_U3444 P2_U3069 ; P2_U6123
g6783 nand P2_U6123 P2_U6122 ; P2_U6124
g6784 nand P2_U5720 P2_U4158 ; P2_U6125
g6785 nand P2_U3438 P2_U3066 ; P2_U6126
g6786 nand P2_U6126 P2_U6125 ; P2_U6127
g6787 nand P2_U5713 P2_U4134 ; P2_U6128
g6788 nand P2_U3435 P2_U3070 ; P2_U6129
g6789 nand P2_U6129 P2_U6128 ; P2_U6130
g6790 nand P2_U5818 P2_U4424 ; P2_U6131
g6791 nand P2_U3480 P2_U3071 ; P2_U6132
g6792 nand P2_U6132 P2_U6131 ; P2_U6133
g6793 nand P2_U5830 P2_U4462 ; P2_U6134
g6794 nand P2_U3485 P2_U3083 ; P2_U6135
g6795 nand P2_U6135 P2_U6134 ; P2_U6136
g6796 nand P2_U5727 P2_U4177 ; P2_U6137
g6797 nand P2_U3441 P2_U3062 ; P2_U6138
g6798 nand P2_U6138 P2_U6137 ; P2_U6139
g6799 nand P2_U5776 P2_U4310 ; P2_U6140
g6800 nand P2_U3462 P2_U3065 ; P2_U6141
g6801 nand P2_U6141 P2_U6140 ; P2_U6142
g6802 nand P2_U5769 P2_U4291 ; P2_U6143
g6803 nand P2_U3459 P2_U3064 ; P2_U6144
g6804 nand P2_U6144 P2_U6143 ; P2_U6145
g6805 nand P2_U3957 P2_U3078 ; P2_U6146
g6806 nand P2_U3368 P2_U4481 ; P2_U6147
g6807 nand P2_U6147 P2_U6146 ; P2_U6148
g6808 nand P2_U3940 P2_U5156 ; P2_U6149
g6809 nand P2_U3942 P2_U3918 ; P2_U6150
g6810 and P3_U3380 P3_U5450 ; P3_U3013
g6811 and P3_U3380 P3_U3379 ; P3_U3014
g6812 and P3_U5453 P3_U3379 ; P3_U3015
g6813 and P3_U5453 P3_U5450 ; P3_U3016
g6814 and P3_U3874 P3_U5447 ; P3_U3017
g6815 and P3_U3587 P3_U3582 ; P3_U3018
g6816 and P3_U3381 P3_U3382 ; P3_U3019
g6817 and P3_U5462 P3_U3381 ; P3_U3020
g6818 and P3_U5459 P3_U3382 ; P3_U3021
g6819 and P3_U5462 P3_U5459 ; P3_U3022
g6820 and P3_U3046 P3_STATE_REG_SCAN_IN ; P3_U3023
g6821 and P3_U3696 P3_U3366 ; P3_U3024
g6822 and P3_U3911 P3_U4073 ; P3_U3025
g6823 and P3_U3015 P3_U5447 ; P3_U3026
g6824 and P3_U3297 P3_STATE_REG_SCAN_IN ; P3_U3027
g6825 and P3_U3886 P3_U3912 ; P3_U3028
g6826 and P3_U3912 P3_U3365 ; P3_U3029
g6827 and P3_U3693 P3_U3912 ; P3_U3030
g6828 and P3_U3890 P3_U3023 ; P3_U3031
g6829 and P3_U3895 P3_U4073 ; P3_U3032
g6830 and P3_U3911 P3_U4089 ; P3_U3033
g6831 and P3_U3912 P3_U3025 ; P3_U3034
g6832 and P3_U3023 P3_U4989 ; P3_U3035
g6833 and P3_U3895 P3_U4089 ; P3_U3036
g6834 and P3_U5468 P3_U4754 ; P3_U3037
g6835 and P3_U3024 P3_U5468 ; P3_U3038
g6836 and P3_U5465 P3_U4754 ; P3_U3039
g6837 and P3_U3892 P3_U4754 ; P3_U3040
g6838 and P3_U3024 P3_U3892 ; P3_U3041
g6839 and P3_U3023 P3_U3366 ; P3_U3042
g6840 and P3_U3023 P3_U3365 ; P3_U3043
g6841 and P3_U5004 P3_STATE_REG_SCAN_IN ; P3_U3044
g6842 and P3_U3023 P3_U5006 ; P3_U3045
g6843 and P3_U5440 P3_U3362 ; P3_U3046
g6844 and P3_U3692 P3_U3018 ; P3_U3047
g6845 and P3_U3691 P3_U3018 ; P3_U3048
g6846 and P3_U4749 P3_U4748 ; P3_U3049
g6847 and P3_U4759 P3_STATE_REG_SCAN_IN ; P3_U3050
g6848 and P3_U3897 P3_U4761 ; P3_U3051
g6849 nand P3_U4536 P3_U4537 P3_U4535 P3_U4538 ; P3_U3052
g6850 nand P3_U4556 P3_U4555 P3_U4554 P3_U4553 ; P3_U3053
g6851 nand P3_U4574 P3_U4573 P3_U4572 P3_U4571 ; P3_U3054
g6852 nand P3_U4612 P3_U4611 P3_U4610 P3_U4609 ; P3_U3055
g6853 nand P3_U4520 P3_U4519 P3_U4518 P3_U4517 ; P3_U3056
g6854 nand P3_U4502 P3_U4501 P3_U4500 P3_U4499 ; P3_U3057
g6855 nand P3_U4592 P3_U4591 P3_U4590 P3_U4589 ; P3_U3058
g6856 nand P3_U4124 P3_U4123 P3_U4122 P3_U4121 ; P3_U3059
g6857 nand P3_U4448 P3_U4447 P3_U4446 P3_U4445 ; P3_U3060
g6858 nand P3_U4232 P3_U4231 P3_U4230 P3_U4229 ; P3_U3061
g6859 nand P3_U4250 P3_U4249 P3_U4248 P3_U4247 ; P3_U3062
g6860 nand P3_U4106 P3_U4105 P3_U4104 P3_U4103 ; P3_U3063
g6861 nand P3_U4484 P3_U4483 P3_U4482 P3_U4481 ; P3_U3064
g6862 nand P3_U4466 P3_U4465 P3_U4464 P3_U4463 ; P3_U3065
g6863 nand P3_U4142 P3_U4141 P3_U4140 P3_U4139 ; P3_U3066
g6864 nand P3_U4081 P3_U4080 P3_U4079 P3_U4078 ; P3_U3067
g6865 nand P3_U4358 P3_U4357 P3_U4356 P3_U4355 ; P3_U3068
g6866 nand P3_U4178 P3_U4177 P3_U4176 P3_U4175 ; P3_U3069
g6867 nand P3_U4160 P3_U4159 P3_U4158 P3_U4157 ; P3_U3070
g6868 nand P3_U4268 P3_U4267 P3_U4266 P3_U4265 ; P3_U3071
g6869 nand P3_U4340 P3_U4339 P3_U4338 P3_U4337 ; P3_U3072
g6870 nand P3_U4322 P3_U4321 P3_U4320 P3_U4319 ; P3_U3073
g6871 nand P3_U4430 P3_U4429 P3_U4428 P3_U4427 ; P3_U3074
g6872 nand P3_U4412 P3_U4411 P3_U4410 P3_U4409 ; P3_U3075
g6873 nand P3_U4086 P3_U4085 P3_U4084 P3_U4083 ; P3_U3076
g6874 nand P3_U4062 P3_U4061 P3_U4060 P3_U4059 ; P3_U3077
g6875 nand P3_U4304 P3_U4303 P3_U4302 P3_U4301 ; P3_U3078
g6876 nand P3_U4286 P3_U4285 P3_U4284 P3_U4283 ; P3_U3079
g6877 nand P3_U4394 P3_U4393 P3_U4392 P3_U4391 ; P3_U3080
g6878 nand P3_U4376 P3_U4375 P3_U4374 P3_U4373 ; P3_U3081
g6879 nand P3_U4214 P3_U4213 P3_U4212 P3_U4211 ; P3_U3082
g6880 nand P3_U4196 P3_U4195 P3_U4194 P3_U4193 ; P3_U3083
g6881 nand P3_U5341 P3_U5340 ; P3_U3084
g6882 nand P3_U5343 P3_U5342 ; P3_U3085
g6883 nand P3_U5349 P3_U5347 P3_U5348 ; P3_U3086
g6884 nand P3_U5352 P3_U5350 P3_U5351 ; P3_U3087
g6885 nand P3_U5355 P3_U5353 P3_U5354 ; P3_U3088
g6886 nand P3_U5358 P3_U5356 P3_U5357 ; P3_U3089
g6887 nand P3_U5361 P3_U5359 P3_U5360 ; P3_U3090
g6888 nand P3_U5364 P3_U5362 P3_U5363 ; P3_U3091
g6889 nand P3_U5367 P3_U5365 P3_U5366 ; P3_U3092
g6890 nand P3_U5370 P3_U5368 P3_U5369 ; P3_U3093
g6891 nand P3_U5373 P3_U5371 P3_U5372 ; P3_U3094
g6892 nand P3_U5376 P3_U5374 P3_U5375 ; P3_U3095
g6893 nand P3_U5381 P3_U5382 P3_U5380 ; P3_U3096
g6894 nand P3_U5384 P3_U5385 P3_U5383 ; P3_U3097
g6895 nand P3_U5387 P3_U5388 P3_U5386 ; P3_U3098
g6896 nand P3_U5390 P3_U5391 P3_U5389 ; P3_U3099
g6897 nand P3_U5393 P3_U5394 P3_U5392 ; P3_U3100
g6898 nand P3_U5396 P3_U5397 P3_U5395 ; P3_U3101
g6899 nand P3_U5399 P3_U5398 P3_U5400 ; P3_U3102
g6900 nand P3_U5402 P3_U5401 P3_U5403 ; P3_U3103
g6901 nand P3_U5405 P3_U5404 P3_U5406 ; P3_U3104
g6902 nand P3_U5408 P3_U5407 P3_U5409 ; P3_U3105
g6903 nand P3_U5323 P3_U5322 P3_U5324 ; P3_U3106
g6904 nand P3_U5326 P3_U5325 P3_U5327 ; P3_U3107
g6905 nand P3_U5329 P3_U5328 P3_U5330 ; P3_U3108
g6906 nand P3_U5332 P3_U5331 P3_U5333 ; P3_U3109
g6907 nand P3_U5335 P3_U5334 P3_U5336 ; P3_U3110
g6908 nand P3_U5338 P3_U5337 P3_U5339 ; P3_U3111
g6909 nand P3_U5345 P3_U5344 P3_U5346 ; P3_U3112
g6910 nand P3_U5378 P3_U5377 P3_U5379 ; P3_U3113
g6911 nand P3_U5411 P3_U5410 P3_U5412 ; P3_U3114
g6912 nand P3_U5414 P3_U5413 ; P3_U3115
g6913 nand P3_U5271 P3_U5270 ; P3_U3116
g6914 nand P3_U5273 P3_U5272 ; P3_U3117
g6915 nand P3_U5277 P3_U3375 P3_U5276 ; P3_U3118
g6916 nand P3_U5279 P3_U3375 P3_U5278 ; P3_U3119
g6917 nand P3_U5281 P3_U3375 P3_U5280 ; P3_U3120
g6918 nand P3_U5283 P3_U3375 P3_U5282 ; P3_U3121
g6919 nand P3_U5285 P3_U3375 P3_U5284 ; P3_U3122
g6920 nand P3_U5287 P3_U3375 P3_U5286 ; P3_U3123
g6921 nand P3_U5289 P3_U3375 P3_U5288 ; P3_U3124
g6922 nand P3_U5291 P3_U3375 P3_U5290 ; P3_U3125
g6923 nand P3_U5293 P3_U3375 P3_U5292 ; P3_U3126
g6924 nand P3_U5295 P3_U3375 P3_U5294 ; P3_U3127
g6925 nand P3_U5299 P3_U3375 P3_U5298 ; P3_U3128
g6926 nand P3_U5301 P3_U3375 P3_U5300 ; P3_U3129
g6927 nand P3_U5303 P3_U3375 P3_U5302 ; P3_U3130
g6928 nand P3_U5305 P3_U3375 P3_U5304 ; P3_U3131
g6929 nand P3_U5307 P3_U3375 P3_U5306 ; P3_U3132
g6930 nand P3_U5309 P3_U3375 P3_U5308 ; P3_U3133
g6931 nand P3_U3825 P3_U5311 ; P3_U3134
g6932 nand P3_U3826 P3_U5313 ; P3_U3135
g6933 nand P3_U3827 P3_U5315 ; P3_U3136
g6934 nand P3_U3828 P3_U5317 ; P3_U3137
g6935 nand P3_U3817 P3_U5259 ; P3_U3138
g6936 nand P3_U3818 P3_U5261 ; P3_U3139
g6937 nand P3_U3819 P3_U5263 ; P3_U3140
g6938 nand P3_U3820 P3_U5265 ; P3_U3141
g6939 nand P3_U3821 P3_U5267 ; P3_U3142
g6940 nand P3_U3822 P3_U5269 ; P3_U3143
g6941 nand P3_U3823 P3_U5275 ; P3_U3144
g6942 nand P3_U3824 P3_U5297 ; P3_U3145
g6943 nand P3_U3829 P3_U5319 ; P3_U3146
g6944 nand P3_U3830 P3_U5321 ; P3_U3147
g6945 nand P3_U3385 P3_U5453 P3_U3375 ; P3_U3148
g6946 nand P3_U3813 P3_U3013 ; P3_U3149
g6947 nand P3_U3812 P3_U5253 ; P3_U3150
g6948 not P3_STATE_REG_SCAN_IN ; P3_U3151
g6949 nand P3_U5944 P3_U5943 P3_U3359 ; P3_U3152
g6950 nand P3_U5249 P3_U5248 P3_U3811 P3_U5250 ; P3_U3153
g6951 nand P3_U5240 P3_U3810 P3_U5239 P3_U5241 ; P3_U3154
g6952 nand P3_U5231 P3_U5230 P3_U3809 P3_U5232 ; P3_U3155
g6953 nand P3_U5222 P3_U3808 P3_U5221 P3_U5223 ; P3_U3156
g6954 nand P3_U5213 P3_U5212 P3_U3807 P3_U5214 ; P3_U3157
g6955 nand P3_U3805 P3_U5204 P3_U3806 ; P3_U3158
g6956 nand P3_U5195 P3_U3804 P3_U5194 P3_U5196 ; P3_U3159
g6957 nand P3_U5186 P3_U3803 P3_U5185 P3_U5187 ; P3_U3160
g6958 nand P3_U5177 P3_U5176 P3_U3802 P3_U5178 ; P3_U3161
g6959 nand P3_U3800 P3_U5168 P3_U3801 ; P3_U3162
g6960 nand P3_U5159 P3_U3799 P3_U5158 P3_U5160 ; P3_U3163
g6961 nand P3_U5150 P3_U5149 P3_U3798 P3_U5151 ; P3_U3164
g6962 nand P3_U5141 P3_U3797 P3_U5140 P3_U5142 ; P3_U3165
g6963 nand P3_U5132 P3_U5131 P3_U3796 P3_U5133 ; P3_U3166
g6964 nand P3_U5123 P3_U5122 P3_U3795 P3_U5124 ; P3_U3167
g6965 nand P3_U5114 P3_U5113 P3_U3794 P3_U5115 ; P3_U3168
g6966 nand P3_U5105 P3_U3793 P3_U5104 P3_U5106 ; P3_U3169
g6967 nand P3_U3791 P3_U5096 P3_U3792 ; P3_U3170
g6968 nand P3_U5087 P3_U5086 P3_U3790 P3_U5088 ; P3_U3171
g6969 nand P3_U5079 P3_U3789 ; P3_U3172
g6970 nand P3_U5071 P3_U3786 P3_U5070 P3_U5072 ; P3_U3173
g6971 nand P3_U5062 P3_U5061 P3_U3785 P3_U5063 ; P3_U3174
g6972 nand P3_U5053 P3_U3784 P3_U5052 P3_U5054 ; P3_U3175
g6973 nand P3_U5044 P3_U5043 P3_U3783 P3_U5045 ; P3_U3176
g6974 nand P3_U3781 P3_U5035 P3_U3782 ; P3_U3177
g6975 nand P3_U5026 P3_U5025 P3_U3780 P3_U5027 ; P3_U3178
g6976 nand P3_U5017 P3_U5016 P3_U3779 P3_U5018 ; P3_U3179
g6977 nand P3_U5008 P3_U3778 P3_U5007 P3_U5009 ; P3_U3180
g6978 nand P3_U4995 P3_U4994 P3_U3777 P3_U4996 ; P3_U3181
g6979 nand P3_U4973 P3_U3756 ; P3_U3182
g6980 nand P3_U4962 P3_U3753 ; P3_U3183
g6981 nand P3_U4951 P3_U3750 ; P3_U3184
g6982 nand P3_U4941 P3_U4940 P3_U3747 ; P3_U3185
g6983 nand P3_U4930 P3_U4929 P3_U3744 ; P3_U3186
g6984 nand P3_U4918 P3_U3741 P3_U3743 P3_U4916 ; P3_U3187
g6985 nand P3_U4907 P3_U3738 P3_U4905 ; P3_U3188
g6986 nand P3_U4896 P3_U3735 ; P3_U3189
g6987 nand P3_U4885 P3_U3732 ; P3_U3190
g6988 nand P3_U4874 P3_U3729 ; P3_U3191
g6989 nand P3_U4863 P3_U3726 ; P3_U3192
g6990 nand P3_U4852 P3_U3723 ; P3_U3193
g6991 nand P3_U4841 P3_U3720 ; P3_U3194
g6992 nand P3_U4830 P3_U3717 ; P3_U3195
g6993 nand P3_U4819 P3_U3714 ; P3_U3196
g6994 nand P3_U4808 P3_U3711 ; P3_U3197
g6995 nand P3_U4797 P3_U3708 ; P3_U3198
g6996 nand P3_U4786 P3_U3705 ; P3_U3199
g6997 nand P3_U4775 P3_U3702 ; P3_U3200
g6998 nand P3_U4764 P3_U3699 ; P3_U3201
g6999 nand P3_U4753 P3_U3049 P3_U4752 ; P3_U3202
g7000 nand P3_U4751 P3_U3049 P3_U4750 ; P3_U3203
g7001 nand P3_U4746 P3_U4747 P3_U4745 P3_U3866 ; P3_U3204
g7002 nand P3_U4743 P3_U4741 P3_U4744 P3_U4742 P3_U3865 ; P3_U3205
g7003 nand P3_U4739 P3_U4737 P3_U4740 P3_U4738 P3_U3864 ; P3_U3206
g7004 nand P3_U4735 P3_U4733 P3_U4736 P3_U4734 P3_U3863 ; P3_U3207
g7005 nand P3_U4731 P3_U4729 P3_U4732 P3_U4730 P3_U3862 ; P3_U3208
g7006 nand P3_U4727 P3_U4725 P3_U4728 P3_U4726 P3_U3861 ; P3_U3209
g7007 nand P3_U4723 P3_U4721 P3_U4724 P3_U4722 P3_U3860 ; P3_U3210
g7008 nand P3_U4719 P3_U4717 P3_U4720 P3_U4718 P3_U3859 ; P3_U3211
g7009 nand P3_U4715 P3_U4713 P3_U4716 P3_U4714 P3_U3858 ; P3_U3212
g7010 nand P3_U4711 P3_U4709 P3_U4712 P3_U4710 P3_U3857 ; P3_U3213
g7011 nand P3_U4707 P3_U4705 P3_U4708 P3_U4706 P3_U3856 ; P3_U3214
g7012 nand P3_U4703 P3_U4701 P3_U4704 P3_U4702 P3_U3855 ; P3_U3215
g7013 nand P3_U4699 P3_U4697 P3_U4700 P3_U4698 P3_U3854 ; P3_U3216
g7014 nand P3_U4695 P3_U4693 P3_U4696 P3_U4694 P3_U3853 ; P3_U3217
g7015 nand P3_U4691 P3_U4689 P3_U4692 P3_U4690 P3_U3852 ; P3_U3218
g7016 nand P3_U4687 P3_U4685 P3_U4688 P3_U4686 P3_U3851 ; P3_U3219
g7017 nand P3_U4684 P3_U4682 P3_U4683 P3_U4681 P3_U3850 ; P3_U3220
g7018 nand P3_U4680 P3_U4679 P3_U4678 P3_U4677 P3_U3849 ; P3_U3221
g7019 nand P3_U4676 P3_U4674 P3_U4675 P3_U4673 P3_U3848 ; P3_U3222
g7020 nand P3_U4672 P3_U4671 P3_U4670 P3_U4669 P3_U3847 ; P3_U3223
g7021 nand P3_U4666 P3_U4665 P3_U4667 P3_U3846 P3_U4668 ; P3_U3224
g7022 nand P3_U4662 P3_U4661 P3_U4663 P3_U3845 P3_U4664 ; P3_U3225
g7023 nand P3_U4658 P3_U4657 P3_U4659 P3_U3844 P3_U4660 ; P3_U3226
g7024 nand P3_U4654 P3_U4653 P3_U4655 P3_U3843 P3_U4656 ; P3_U3227
g7025 nand P3_U4650 P3_U4649 P3_U4651 P3_U3842 P3_U4652 ; P3_U3228
g7026 nand P3_U4646 P3_U4645 P3_U4647 P3_U3841 P3_U4648 ; P3_U3229
g7027 nand P3_U4642 P3_U4641 P3_U4643 P3_U3840 P3_U4644 ; P3_U3230
g7028 nand P3_U4638 P3_U4637 P3_U4639 P3_U3839 P3_U4640 ; P3_U3231
g7029 nand P3_U4634 P3_U4633 P3_U4635 P3_U3838 P3_U4636 ; P3_U3232
g7030 nand P3_U4630 P3_U4629 P3_U4631 P3_U3837 P3_U4632 ; P3_U3233
g7031 and P3_U3832 P3_D_REG_31__SCAN_IN ; P3_U3234
g7032 and P3_U3832 P3_D_REG_30__SCAN_IN ; P3_U3235
g7033 and P3_U3832 P3_D_REG_29__SCAN_IN ; P3_U3236
g7034 and P3_U3832 P3_D_REG_28__SCAN_IN ; P3_U3237
g7035 and P3_U3832 P3_D_REG_27__SCAN_IN ; P3_U3238
g7036 and P3_U3832 P3_D_REG_26__SCAN_IN ; P3_U3239
g7037 and P3_U3832 P3_D_REG_25__SCAN_IN ; P3_U3240
g7038 and P3_U3832 P3_D_REG_24__SCAN_IN ; P3_U3241
g7039 and P3_U3832 P3_D_REG_23__SCAN_IN ; P3_U3242
g7040 and P3_U3832 P3_D_REG_22__SCAN_IN ; P3_U3243
g7041 and P3_U3832 P3_D_REG_21__SCAN_IN ; P3_U3244
g7042 and P3_U3832 P3_D_REG_20__SCAN_IN ; P3_U3245
g7043 and P3_U3832 P3_D_REG_19__SCAN_IN ; P3_U3246
g7044 and P3_U3832 P3_D_REG_18__SCAN_IN ; P3_U3247
g7045 and P3_U3832 P3_D_REG_17__SCAN_IN ; P3_U3248
g7046 and P3_U3832 P3_D_REG_16__SCAN_IN ; P3_U3249
g7047 and P3_U3832 P3_D_REG_15__SCAN_IN ; P3_U3250
g7048 and P3_U3832 P3_D_REG_14__SCAN_IN ; P3_U3251
g7049 and P3_U3832 P3_D_REG_13__SCAN_IN ; P3_U3252
g7050 and P3_U3832 P3_D_REG_12__SCAN_IN ; P3_U3253
g7051 and P3_U3832 P3_D_REG_11__SCAN_IN ; P3_U3254
g7052 and P3_U3832 P3_D_REG_10__SCAN_IN ; P3_U3255
g7053 and P3_U3832 P3_D_REG_9__SCAN_IN ; P3_U3256
g7054 and P3_U3832 P3_D_REG_8__SCAN_IN ; P3_U3257
g7055 and P3_U3832 P3_D_REG_7__SCAN_IN ; P3_U3258
g7056 and P3_U3832 P3_D_REG_6__SCAN_IN ; P3_U3259
g7057 and P3_U3832 P3_D_REG_5__SCAN_IN ; P3_U3260
g7058 and P3_U3832 P3_D_REG_4__SCAN_IN ; P3_U3261
g7059 and P3_U3832 P3_D_REG_3__SCAN_IN ; P3_U3262
g7060 and P3_U3832 P3_D_REG_2__SCAN_IN ; P3_U3263
g7061 nand P3_U4016 P3_U4017 P3_U4015 ; P3_U3264
g7062 nand P3_U4013 P3_U4014 P3_U4012 ; P3_U3265
g7063 nand P3_U4010 P3_U4011 P3_U4009 ; P3_U3266
g7064 nand P3_U4007 P3_U4008 P3_U4006 ; P3_U3267
g7065 nand P3_U4004 P3_U4005 P3_U4003 ; P3_U3268
g7066 nand P3_U4001 P3_U4002 P3_U4000 ; P3_U3269
g7067 nand P3_U3998 P3_U3999 P3_U3997 ; P3_U3270
g7068 nand P3_U3995 P3_U3996 P3_U3994 ; P3_U3271
g7069 nand P3_U3992 P3_U3993 P3_U3991 ; P3_U3272
g7070 nand P3_U3989 P3_U3990 P3_U3988 ; P3_U3273
g7071 nand P3_U3986 P3_U3987 P3_U3985 ; P3_U3274
g7072 nand P3_U3983 P3_U3984 P3_U3982 ; P3_U3275
g7073 nand P3_U3980 P3_U3981 P3_U3979 ; P3_U3276
g7074 nand P3_U3977 P3_U3978 P3_U3976 ; P3_U3277
g7075 nand P3_U3974 P3_U3975 P3_U3973 ; P3_U3278
g7076 nand P3_U3971 P3_U3972 P3_U3970 ; P3_U3279
g7077 nand P3_U3968 P3_U3969 P3_U3967 ; P3_U3280
g7078 nand P3_U3965 P3_U3966 P3_U3964 ; P3_U3281
g7079 nand P3_U3962 P3_U3963 P3_U3961 ; P3_U3282
g7080 nand P3_U3959 P3_U3960 P3_U3958 ; P3_U3283
g7081 nand P3_U3956 P3_U3957 P3_U3955 ; P3_U3284
g7082 nand P3_U3953 P3_U3954 P3_U3952 ; P3_U3285
g7083 nand P3_U3950 P3_U3951 P3_U3949 ; P3_U3286
g7084 nand P3_U3947 P3_U3948 P3_U3946 ; P3_U3287
g7085 nand P3_U3944 P3_U3945 P3_U3943 ; P3_U3288
g7086 nand P3_U3941 P3_U3942 P3_U3940 ; P3_U3289
g7087 nand P3_U3938 P3_U3939 P3_U3937 ; P3_U3290
g7088 nand P3_U3935 P3_U3936 P3_U3934 ; P3_U3291
g7089 nand P3_U3932 P3_U3933 P3_U3931 ; P3_U3292
g7090 nand P3_U3929 P3_U3930 P3_U3928 ; P3_U3293
g7091 nand P3_U3926 P3_U3927 P3_U3925 ; P3_U3294
g7092 nand P3_U3923 P3_U3924 P3_U3922 ; P3_U3295
g7093 and P3_U3775 P3_U5421 ; P3_U3296
g7094 nand P3_U3831 P3_STATE_REG_SCAN_IN ; P3_U3297
g7095 not P3_B_REG_SCAN_IN ; P3_U3298
g7096 nand P3_U3374 P3_U5431 ; P3_U3299
g7097 nand P3_U3374 P3_U4018 ; P3_U3300
g7098 nand P3_U3013 P3_U5447 ; P3_U3301
g7099 nand P3_U3014 P3_U5456 ; P3_U3302
g7100 nand P3_U3588 P3_U3018 ; P3_U3303
g7101 nand P3_U3589 P3_U3018 ; P3_U3304
g7102 nand P3_U3014 P3_U5447 ; P3_U3305
g7103 nand P3_U3014 P3_U3378 ; P3_U3306
g7104 nand P3_U3013 P3_U3378 ; P3_U3307
g7105 nand P3_U3385 P3_U3379 P3_U3378 ; P3_U3308
g7106 nand P3_U5450 P3_U3385 P3_U3378 ; P3_U3309
g7107 nand P3_U5456 P3_U3013 ; P3_U3310
g7108 nand P3_U3878 P3_U5447 ; P3_U3311
g7109 nand P3_U3016 P3_U3385 ; P3_U3312
g7110 nand P3_U3385 P3_U3380 ; P3_U3313
g7111 nand P3_U4070 P3_U4069 P3_U4071 P3_U3576 P3_U3575 ; P3_U3314
g7112 nand P3_U4091 P3_U4090 P3_U3590 P3_U3592 ; P3_U3315
g7113 nand P3_U4109 P3_U4108 P3_U3594 P3_U3596 ; P3_U3316
g7114 nand P3_U4127 P3_U4126 P3_U3598 P3_U3600 ; P3_U3317
g7115 nand P3_U4145 P3_U4144 P3_U4146 P3_U4147 P3_U3603 ; P3_U3318
g7116 nand P3_U4163 P3_U4162 P3_U4164 P3_U4165 P3_U3606 ; P3_U3319
g7117 nand P3_U4181 P3_U4180 P3_U4182 P3_U4183 P3_U3609 ; P3_U3320
g7118 nand P3_U4199 P3_U4198 P3_U4200 P3_U4201 P3_U3612 ; P3_U3321
g7119 nand P3_U4217 P3_U4216 P3_U4218 P3_U4219 P3_U3615 ; P3_U3322
g7120 nand P3_U4235 P3_U4234 P3_U3617 P3_U3619 ; P3_U3323
g7121 nand P3_U4253 P3_U4252 P3_U3621 P3_U3623 ; P3_U3324
g7122 nand P3_U4271 P3_U4270 P3_U4272 P3_U4273 P3_U3626 ; P3_U3325
g7123 nand P3_U4289 P3_U4288 P3_U3628 P3_U3630 ; P3_U3326
g7124 nand P3_U4307 P3_U4306 P3_U3632 P3_U3634 ; P3_U3327
g7125 nand P3_U4325 P3_U4324 P3_U4326 P3_U4327 P3_U3637 ; P3_U3328
g7126 nand P3_U4343 P3_U4342 P3_U4344 P3_U4345 P3_U3640 ; P3_U3329
g7127 nand P3_U4361 P3_U4360 P3_U4362 P3_U4363 P3_U3643 ; P3_U3330
g7128 nand P3_U4379 P3_U4378 P3_U3645 P3_U3647 ; P3_U3331
g7129 nand P3_U4397 P3_U4396 P3_U4398 P3_U4399 P3_U3650 ; P3_U3332
g7130 nand P3_U4415 P3_U4414 P3_U4416 P3_U4417 P3_U3653 ; P3_U3333
g7131 nand U49 P3_U3833 ; P3_U3334
g7132 nand P3_U4433 P3_U4432 P3_U4434 P3_U4435 P3_U3656 ; P3_U3335
g7133 nand U48 P3_U3833 ; P3_U3336
g7134 nand P3_U4451 P3_U4450 P3_U4452 P3_U4453 P3_U3659 ; P3_U3337
g7135 nand U47 P3_U3833 ; P3_U3338
g7136 nand P3_U4469 P3_U4468 P3_U4470 P3_U4471 P3_U3662 ; P3_U3339
g7137 nand U46 P3_U3833 ; P3_U3340
g7138 nand P3_U4487 P3_U4486 P3_U4488 P3_U4489 P3_U3665 ; P3_U3341
g7139 nand U45 P3_U3833 ; P3_U3342
g7140 nand P3_U4505 P3_U4504 P3_U3667 P3_U3669 ; P3_U3343
g7141 nand U44 P3_U3833 ; P3_U3344
g7142 nand P3_U4523 P3_U4522 P3_U3671 P3_U3673 ; P3_U3345
g7143 nand U43 P3_U3833 ; P3_U3346
g7144 nand P3_U4541 P3_U4540 P3_U3675 P3_U3677 ; P3_U3347
g7145 nand U42 P3_U3833 ; P3_U3348
g7146 nand P3_U4559 P3_U4558 P3_U3679 P3_U3681 ; P3_U3349
g7147 nand U41 P3_U3833 ; P3_U3350
g7148 nand P3_U4577 P3_U4576 P3_U3683 P3_U3685 ; P3_U3351
g7149 nand P3_U3383 P3_U3384 ; P3_U3352
g7150 nand U40 P3_U3833 ; P3_U3353
g7151 nand P3_U4597 P3_U4596 P3_U4598 P3_U3687 P3_U3689 ; P3_U3354
g7152 nand U38 P3_U3833 ; P3_U3355
g7153 nand U37 P3_U3833 ; P3_U3356
g7154 nand P3_U3015 P3_U5456 ; P3_U3357
g7155 nand P3_U3023 P3_U4627 ; P3_U3358
g7156 nand P3_U5447 P3_U3385 ; P3_U3359
g7157 nand P3_U3879 P3_U5447 ; P3_U3360
g7158 nand P3_U3911 P3_U4595 P3_U3055 ; P3_U3361
g7159 nand P3_U3373 P3_U3374 P3_U3372 ; P3_U3362
g7160 nand P3_U3694 P3_U3910 ; P3_U3363
g7161 nand P3_U3313 P3_U3833 ; P3_U3364
g7162 nand P3_U3877 P3_U5423 ; P3_U3365
g7163 nand P3_U3695 P3_U3050 ; P3_U3366
g7164 nand P3_U3882 P3_U3385 ; P3_U3367
g7165 nand P3_U3759 P3_U3890 ; P3_U3368
g7166 nand P3_U3876 P3_U3378 ; P3_U3369
g7167 nand P3_U4992 P3_U4991 P3_U3776 ; P3_U3370
g7168 nand P3_U5417 P3_U3917 ; P3_U3371
g7169 nand P3_U5427 P3_U5426 ; P3_U3372
g7170 nand P3_U5430 P3_U5429 ; P3_U3373
g7171 nand P3_U5433 P3_U5432 ; P3_U3374
g7172 nand P3_U5439 P3_U5438 ; P3_U3375
g7173 nand P3_U5442 P3_U5441 ; P3_U3376
g7174 nand P3_U5444 P3_U5443 ; P3_U3377
g7175 nand P3_U5446 P3_U5445 ; P3_U3378
g7176 nand P3_U5449 P3_U5448 ; P3_U3379
g7177 nand P3_U5452 P3_U5451 ; P3_U3380
g7178 nand P3_U5458 P3_U5457 ; P3_U3381
g7179 nand P3_U5461 P3_U5460 ; P3_U3382
g7180 nand P3_U5464 P3_U5463 ; P3_U3383
g7181 nand P3_U5467 P3_U5466 ; P3_U3384
g7182 nand P3_U5455 P3_U5454 ; P3_U3385
g7183 nand P3_U5470 P3_U5469 ; P3_U3386
g7184 nand P3_U5472 P3_U5471 ; P3_U3387
g7185 nand P3_U5475 P3_U5474 ; P3_U3388
g7186 nand P3_U5478 P3_U5477 ; P3_U3389
g7187 nand P3_U5484 P3_U5483 ; P3_U3390
g7188 nand P3_U5486 P3_U5485 ; P3_U3391
g7189 nand P3_U5488 P3_U5487 ; P3_U3392
g7190 nand P3_U5491 P3_U5490 ; P3_U3393
g7191 nand P3_U5493 P3_U5492 ; P3_U3394
g7192 nand P3_U5495 P3_U5494 ; P3_U3395
g7193 nand P3_U5498 P3_U5497 ; P3_U3396
g7194 nand P3_U5500 P3_U5499 ; P3_U3397
g7195 nand P3_U5502 P3_U5501 ; P3_U3398
g7196 nand P3_U5505 P3_U5504 ; P3_U3399
g7197 nand P3_U5507 P3_U5506 ; P3_U3400
g7198 nand P3_U5509 P3_U5508 ; P3_U3401
g7199 nand P3_U5512 P3_U5511 ; P3_U3402
g7200 nand P3_U5514 P3_U5513 ; P3_U3403
g7201 nand P3_U5516 P3_U5515 ; P3_U3404
g7202 nand P3_U5519 P3_U5518 ; P3_U3405
g7203 nand P3_U5521 P3_U5520 ; P3_U3406
g7204 nand P3_U5523 P3_U5522 ; P3_U3407
g7205 nand P3_U5526 P3_U5525 ; P3_U3408
g7206 nand P3_U5528 P3_U5527 ; P3_U3409
g7207 nand P3_U5530 P3_U5529 ; P3_U3410
g7208 nand P3_U5533 P3_U5532 ; P3_U3411
g7209 nand P3_U5535 P3_U5534 ; P3_U3412
g7210 nand P3_U5537 P3_U5536 ; P3_U3413
g7211 nand P3_U5540 P3_U5539 ; P3_U3414
g7212 nand P3_U5542 P3_U5541 ; P3_U3415
g7213 nand P3_U5544 P3_U5543 ; P3_U3416
g7214 nand P3_U5547 P3_U5546 ; P3_U3417
g7215 nand P3_U5549 P3_U5548 ; P3_U3418
g7216 nand P3_U5551 P3_U5550 ; P3_U3419
g7217 nand P3_U5554 P3_U5553 ; P3_U3420
g7218 nand P3_U5556 P3_U5555 ; P3_U3421
g7219 nand P3_U5558 P3_U5557 ; P3_U3422
g7220 nand P3_U5561 P3_U5560 ; P3_U3423
g7221 nand P3_U5563 P3_U5562 ; P3_U3424
g7222 nand P3_U5565 P3_U5564 ; P3_U3425
g7223 nand P3_U5568 P3_U5567 ; P3_U3426
g7224 nand P3_U5570 P3_U5569 ; P3_U3427
g7225 nand P3_U5572 P3_U5571 ; P3_U3428
g7226 nand P3_U5575 P3_U5574 ; P3_U3429
g7227 nand P3_U5577 P3_U5576 ; P3_U3430
g7228 nand P3_U5579 P3_U5578 ; P3_U3431
g7229 nand P3_U5582 P3_U5581 ; P3_U3432
g7230 nand P3_U5584 P3_U5583 ; P3_U3433
g7231 nand P3_U5586 P3_U5585 ; P3_U3434
g7232 nand P3_U5589 P3_U5588 ; P3_U3435
g7233 nand P3_U5591 P3_U5590 ; P3_U3436
g7234 nand P3_U5593 P3_U5592 ; P3_U3437
g7235 nand P3_U5596 P3_U5595 ; P3_U3438
g7236 nand P3_U5598 P3_U5597 ; P3_U3439
g7237 nand P3_U5600 P3_U5599 ; P3_U3440
g7238 nand P3_U5603 P3_U5602 ; P3_U3441
g7239 nand P3_U5605 P3_U5604 ; P3_U3442
g7240 nand P3_U5607 P3_U5606 ; P3_U3443
g7241 nand P3_U5610 P3_U5609 ; P3_U3444
g7242 nand P3_U5612 P3_U5611 ; P3_U3445
g7243 nand P3_U5615 P3_U5614 ; P3_U3446
g7244 nand P3_U5617 P3_U5616 ; P3_U3447
g7245 nand P3_U5619 P3_U5618 ; P3_U3448
g7246 nand P3_U5621 P3_U5620 ; P3_U3449
g7247 nand P3_U5623 P3_U5622 ; P3_U3450
g7248 nand P3_U5625 P3_U5624 ; P3_U3451
g7249 nand P3_U5627 P3_U5626 ; P3_U3452
g7250 nand P3_U5629 P3_U5628 ; P3_U3453
g7251 nand P3_U5631 P3_U5630 ; P3_U3454
g7252 nand P3_U5633 P3_U5632 ; P3_U3455
g7253 nand P3_U5635 P3_U5634 ; P3_U3456
g7254 nand P3_U5637 P3_U5636 ; P3_U3457
g7255 nand P3_U5639 P3_U5638 ; P3_U3458
g7256 nand P3_U5643 P3_U5642 ; P3_U3459
g7257 nand P3_U5645 P3_U5644 ; P3_U3460
g7258 nand P3_U5647 P3_U5646 ; P3_U3461
g7259 nand P3_U5649 P3_U5648 ; P3_U3462
g7260 nand P3_U5651 P3_U5650 ; P3_U3463
g7261 nand P3_U5653 P3_U5652 ; P3_U3464
g7262 nand P3_U5655 P3_U5654 ; P3_U3465
g7263 nand P3_U5657 P3_U5656 ; P3_U3466
g7264 nand P3_U5659 P3_U5658 ; P3_U3467
g7265 nand P3_U5661 P3_U5660 ; P3_U3468
g7266 nand P3_U5663 P3_U5662 ; P3_U3469
g7267 nand P3_U5665 P3_U5664 ; P3_U3470
g7268 nand P3_U5667 P3_U5666 ; P3_U3471
g7269 nand P3_U5669 P3_U5668 ; P3_U3472
g7270 nand P3_U5671 P3_U5670 ; P3_U3473
g7271 nand P3_U5673 P3_U5672 ; P3_U3474
g7272 nand P3_U5675 P3_U5674 ; P3_U3475
g7273 nand P3_U5677 P3_U5676 ; P3_U3476
g7274 nand P3_U5679 P3_U5678 ; P3_U3477
g7275 nand P3_U5681 P3_U5680 ; P3_U3478
g7276 nand P3_U5683 P3_U5682 ; P3_U3479
g7277 nand P3_U5685 P3_U5684 ; P3_U3480
g7278 nand P3_U5687 P3_U5686 ; P3_U3481
g7279 nand P3_U5689 P3_U5688 ; P3_U3482
g7280 nand P3_U5691 P3_U5690 ; P3_U3483
g7281 nand P3_U5693 P3_U5692 ; P3_U3484
g7282 nand P3_U5695 P3_U5694 ; P3_U3485
g7283 nand P3_U5697 P3_U5696 ; P3_U3486
g7284 nand P3_U5699 P3_U5698 ; P3_U3487
g7285 nand P3_U5701 P3_U5700 ; P3_U3488
g7286 nand P3_U5703 P3_U5702 ; P3_U3489
g7287 nand P3_U5705 P3_U5704 ; P3_U3490
g7288 nand P3_U5770 P3_U5769 ; P3_U3491
g7289 nand P3_U5772 P3_U5771 ; P3_U3492
g7290 nand P3_U5774 P3_U5773 ; P3_U3493
g7291 nand P3_U5776 P3_U5775 ; P3_U3494
g7292 nand P3_U5778 P3_U5777 ; P3_U3495
g7293 nand P3_U5780 P3_U5779 ; P3_U3496
g7294 nand P3_U5782 P3_U5781 ; P3_U3497
g7295 nand P3_U5784 P3_U5783 ; P3_U3498
g7296 nand P3_U5786 P3_U5785 ; P3_U3499
g7297 nand P3_U5788 P3_U5787 ; P3_U3500
g7298 nand P3_U5790 P3_U5789 ; P3_U3501
g7299 nand P3_U5792 P3_U5791 ; P3_U3502
g7300 nand P3_U5794 P3_U5793 ; P3_U3503
g7301 nand P3_U5796 P3_U5795 ; P3_U3504
g7302 nand P3_U5798 P3_U5797 ; P3_U3505
g7303 nand P3_U5800 P3_U5799 ; P3_U3506
g7304 nand P3_U5802 P3_U5801 ; P3_U3507
g7305 nand P3_U5804 P3_U5803 ; P3_U3508
g7306 nand P3_U5806 P3_U5805 ; P3_U3509
g7307 nand P3_U5808 P3_U5807 ; P3_U3510
g7308 nand P3_U5810 P3_U5809 ; P3_U3511
g7309 nand P3_U5812 P3_U5811 ; P3_U3512
g7310 nand P3_U5814 P3_U5813 ; P3_U3513
g7311 nand P3_U5816 P3_U5815 ; P3_U3514
g7312 nand P3_U5818 P3_U5817 ; P3_U3515
g7313 nand P3_U5820 P3_U5819 ; P3_U3516
g7314 nand P3_U5822 P3_U5821 ; P3_U3517
g7315 nand P3_U5824 P3_U5823 ; P3_U3518
g7316 nand P3_U5826 P3_U5825 ; P3_U3519
g7317 nand P3_U5828 P3_U5827 ; P3_U3520
g7318 nand P3_U5830 P3_U5829 ; P3_U3521
g7319 nand P3_U5832 P3_U5831 ; P3_U3522
g7320 nand P3_U5946 P3_U5945 ; P3_U3523
g7321 nand P3_U5948 P3_U5947 ; P3_U3524
g7322 nand P3_U5950 P3_U5949 ; P3_U3525
g7323 nand P3_U5952 P3_U5951 ; P3_U3526
g7324 nand P3_U5954 P3_U5953 ; P3_U3527
g7325 nand P3_U5956 P3_U5955 ; P3_U3528
g7326 nand P3_U5958 P3_U5957 ; P3_U3529
g7327 nand P3_U5960 P3_U5959 ; P3_U3530
g7328 nand P3_U5962 P3_U5961 ; P3_U3531
g7329 nand P3_U5964 P3_U5963 ; P3_U3532
g7330 nand P3_U5966 P3_U5965 ; P3_U3533
g7331 nand P3_U5968 P3_U5967 ; P3_U3534
g7332 nand P3_U5970 P3_U5969 ; P3_U3535
g7333 nand P3_U5972 P3_U5971 ; P3_U3536
g7334 nand P3_U5974 P3_U5973 ; P3_U3537
g7335 nand P3_U5976 P3_U5975 ; P3_U3538
g7336 nand P3_U5978 P3_U5977 ; P3_U3539
g7337 nand P3_U5980 P3_U5979 ; P3_U3540
g7338 nand P3_U5982 P3_U5981 ; P3_U3541
g7339 nand P3_U5984 P3_U5983 ; P3_U3542
g7340 nand P3_U5986 P3_U5985 ; P3_U3543
g7341 nand P3_U5988 P3_U5987 ; P3_U3544
g7342 nand P3_U5990 P3_U5989 ; P3_U3545
g7343 nand P3_U5992 P3_U5991 ; P3_U3546
g7344 nand P3_U5994 P3_U5993 ; P3_U3547
g7345 nand P3_U5996 P3_U5995 ; P3_U3548
g7346 nand P3_U5998 P3_U5997 ; P3_U3549
g7347 nand P3_U6000 P3_U5999 ; P3_U3550
g7348 nand P3_U6002 P3_U6001 ; P3_U3551
g7349 nand P3_U6004 P3_U6003 ; P3_U3552
g7350 nand P3_U6006 P3_U6005 ; P3_U3553
g7351 nand P3_U6008 P3_U6007 ; P3_U3554
g7352 nand P3_U6010 P3_U6009 ; P3_U3555
g7353 nand P3_U6012 P3_U6011 ; P3_U3556
g7354 nand P3_U6014 P3_U6013 ; P3_U3557
g7355 nand P3_U6016 P3_U6015 ; P3_U3558
g7356 nand P3_U6018 P3_U6017 ; P3_U3559
g7357 nand P3_U6020 P3_U6019 ; P3_U3560
g7358 nand P3_U6022 P3_U6021 ; P3_U3561
g7359 nand P3_U6024 P3_U6023 ; P3_U3562
g7360 nand P3_U6026 P3_U6025 ; P3_U3563
g7361 nand P3_U6028 P3_U6027 ; P3_U3564
g7362 nand P3_U6030 P3_U6029 ; P3_U3565
g7363 nand P3_U6032 P3_U6031 ; P3_U3566
g7364 nand P3_U6034 P3_U6033 ; P3_U3567
g7365 nand P3_U6036 P3_U6035 ; P3_U3568
g7366 nand P3_U6038 P3_U6037 ; P3_U3569
g7367 nand P3_U6040 P3_U6039 ; P3_U3570
g7368 nand P3_U6042 P3_U6041 ; P3_U3571
g7369 nand P3_U6044 P3_U6043 ; P3_U3572
g7370 nand P3_U6046 P3_U6045 ; P3_U3573
g7371 nand P3_U6048 P3_U6047 ; P3_U3574
g7372 and P3_U4066 P3_U4065 ; P3_U3575
g7373 and P3_U4068 P3_U4067 ; P3_U3576
g7374 and P3_U4076 P3_U4074 P3_U4075 ; P3_U3577
g7375 and P3_U4025 P3_U4024 P3_U4023 P3_U4022 ; P3_U3578
g7376 and P3_U4029 P3_U4028 P3_U4027 P3_U4026 ; P3_U3579
g7377 and P3_U4033 P3_U4032 P3_U4031 P3_U4030 ; P3_U3580
g7378 and P3_U4035 P3_U4034 P3_U4036 ; P3_U3581
g7379 and P3_U3581 P3_U3580 P3_U3579 P3_U3578 ; P3_U3582
g7380 and P3_U4040 P3_U4039 P3_U4038 P3_U4037 ; P3_U3583
g7381 and P3_U4044 P3_U4043 P3_U4042 P3_U4041 ; P3_U3584
g7382 and P3_U4048 P3_U4047 P3_U4046 P3_U4045 ; P3_U3585
g7383 and P3_U4050 P3_U4049 P3_U4051 ; P3_U3586
g7384 and P3_U3586 P3_U3585 P3_U3584 P3_U3583 ; P3_U3587
g7385 and P3_U3389 P3_U3388 ; P3_U3588
g7386 and P3_U5479 P3_U5476 ; P3_U3589
g7387 and P3_U4093 P3_U4092 ; P3_U3590
g7388 and P3_U4095 P3_U4094 ; P3_U3591
g7389 and P3_U4097 P3_U4096 P3_U3591 ; P3_U3592
g7390 and P3_U4100 P3_U4101 P3_U4099 ; P3_U3593
g7391 and P3_U4111 P3_U4110 ; P3_U3594
g7392 and P3_U4113 P3_U4112 ; P3_U3595
g7393 and P3_U4115 P3_U4114 P3_U3595 ; P3_U3596
g7394 and P3_U4118 P3_U4119 P3_U4117 ; P3_U3597
g7395 and P3_U4129 P3_U4128 ; P3_U3598
g7396 and P3_U4131 P3_U4130 ; P3_U3599
g7397 and P3_U4133 P3_U4132 P3_U3599 ; P3_U3600
g7398 and P3_U4136 P3_U4137 P3_U4135 ; P3_U3601
g7399 and P3_U4149 P3_U4148 ; P3_U3602
g7400 and P3_U4151 P3_U4150 P3_U3602 ; P3_U3603
g7401 and P3_U4154 P3_U4155 P3_U4153 ; P3_U3604
g7402 and P3_U4167 P3_U4166 ; P3_U3605
g7403 and P3_U4169 P3_U4168 P3_U3605 ; P3_U3606
g7404 and P3_U4172 P3_U4173 P3_U4171 ; P3_U3607
g7405 and P3_U4185 P3_U4184 ; P3_U3608
g7406 and P3_U4187 P3_U4186 P3_U3608 ; P3_U3609
g7407 and P3_U4190 P3_U4191 P3_U4189 ; P3_U3610
g7408 and P3_U4203 P3_U4202 ; P3_U3611
g7409 and P3_U4205 P3_U4204 P3_U3611 ; P3_U3612
g7410 and P3_U4208 P3_U4209 P3_U4207 ; P3_U3613
g7411 and P3_U4221 P3_U4220 ; P3_U3614
g7412 and P3_U4223 P3_U4222 P3_U3614 ; P3_U3615
g7413 and P3_U4226 P3_U4227 P3_U4225 ; P3_U3616
g7414 and P3_U4237 P3_U4236 ; P3_U3617
g7415 and P3_U4239 P3_U4238 ; P3_U3618
g7416 and P3_U4241 P3_U4240 P3_U3618 ; P3_U3619
g7417 and P3_U4244 P3_U4245 P3_U4243 ; P3_U3620
g7418 and P3_U4255 P3_U4254 ; P3_U3621
g7419 and P3_U4257 P3_U4256 ; P3_U3622
g7420 and P3_U4259 P3_U4258 P3_U3622 ; P3_U3623
g7421 and P3_U4262 P3_U4263 P3_U4261 ; P3_U3624
g7422 and P3_U4275 P3_U4274 ; P3_U3625
g7423 and P3_U4277 P3_U4276 P3_U3625 ; P3_U3626
g7424 and P3_U4280 P3_U4281 P3_U4279 ; P3_U3627
g7425 and P3_U4291 P3_U4290 ; P3_U3628
g7426 and P3_U4293 P3_U4292 ; P3_U3629
g7427 and P3_U4295 P3_U4294 P3_U3629 ; P3_U3630
g7428 and P3_U4298 P3_U4299 P3_U4297 ; P3_U3631
g7429 and P3_U4309 P3_U4308 ; P3_U3632
g7430 and P3_U4311 P3_U4310 ; P3_U3633
g7431 and P3_U4313 P3_U4312 P3_U3633 ; P3_U3634
g7432 and P3_U4316 P3_U4317 P3_U4315 ; P3_U3635
g7433 and P3_U4329 P3_U4328 ; P3_U3636
g7434 and P3_U4331 P3_U4330 P3_U3636 ; P3_U3637
g7435 and P3_U4334 P3_U4335 P3_U4333 ; P3_U3638
g7436 and P3_U4347 P3_U4346 ; P3_U3639
g7437 and P3_U4349 P3_U4348 P3_U3639 ; P3_U3640
g7438 and P3_U4352 P3_U4353 P3_U4351 ; P3_U3641
g7439 and P3_U4365 P3_U4364 ; P3_U3642
g7440 and P3_U4367 P3_U4366 P3_U3642 ; P3_U3643
g7441 and P3_U4370 P3_U4371 P3_U4369 ; P3_U3644
g7442 and P3_U4381 P3_U4380 ; P3_U3645
g7443 and P3_U4383 P3_U4382 ; P3_U3646
g7444 and P3_U4385 P3_U4384 P3_U3646 ; P3_U3647
g7445 and P3_U4388 P3_U4389 P3_U4387 ; P3_U3648
g7446 and P3_U4401 P3_U4400 ; P3_U3649
g7447 and P3_U4403 P3_U4402 P3_U3649 ; P3_U3650
g7448 and P3_U4406 P3_U4407 P3_U4405 ; P3_U3651
g7449 and P3_U4419 P3_U4418 ; P3_U3652
g7450 and P3_U4421 P3_U4420 P3_U3652 ; P3_U3653
g7451 and P3_U4424 P3_U4425 P3_U4423 ; P3_U3654
g7452 and P3_U4437 P3_U4436 ; P3_U3655
g7453 and P3_U4439 P3_U4438 P3_U3655 ; P3_U3656
g7454 and P3_U4442 P3_U4443 P3_U4441 ; P3_U3657
g7455 and P3_U4455 P3_U4454 ; P3_U3658
g7456 and P3_U4457 P3_U4456 P3_U3658 ; P3_U3659
g7457 and P3_U4460 P3_U4461 P3_U4459 ; P3_U3660
g7458 and P3_U4473 P3_U4472 ; P3_U3661
g7459 and P3_U4475 P3_U4474 P3_U3661 ; P3_U3662
g7460 and P3_U4478 P3_U4479 P3_U4477 ; P3_U3663
g7461 and P3_U4491 P3_U4490 ; P3_U3664
g7462 and P3_U4493 P3_U4492 P3_U3664 ; P3_U3665
g7463 and P3_U4496 P3_U4497 P3_U4495 ; P3_U3666
g7464 and P3_U4507 P3_U4506 ; P3_U3667
g7465 and P3_U4509 P3_U4508 ; P3_U3668
g7466 and P3_U4511 P3_U4510 P3_U3668 ; P3_U3669
g7467 and P3_U4514 P3_U4515 P3_U4513 ; P3_U3670
g7468 and P3_U4525 P3_U4524 ; P3_U3671
g7469 and P3_U4527 P3_U4526 ; P3_U3672
g7470 and P3_U4529 P3_U4528 P3_U3672 ; P3_U3673
g7471 and P3_U4532 P3_U4533 P3_U4531 ; P3_U3674
g7472 and P3_U4543 P3_U4542 ; P3_U3675
g7473 and P3_U4545 P3_U4544 ; P3_U3676
g7474 and P3_U4547 P3_U4546 P3_U3676 ; P3_U3677
g7475 and P3_U4550 P3_U4551 P3_U4549 ; P3_U3678
g7476 and P3_U4561 P3_U4560 ; P3_U3679
g7477 and P3_U4563 P3_U4562 ; P3_U3680
g7478 and P3_U4565 P3_U4564 P3_U3680 ; P3_U3681
g7479 and P3_U4568 P3_U4569 P3_U4567 ; P3_U3682
g7480 and P3_U4579 P3_U4578 ; P3_U3683
g7481 and P3_U4581 P3_U4580 ; P3_U3684
g7482 and P3_U4583 P3_U4582 P3_U3684 ; P3_U3685
g7483 and P3_U4586 P3_U4587 P3_U4585 ; P3_U3686
g7484 and P3_U4600 P3_U4599 ; P3_U3687
g7485 and P3_U4602 P3_U4601 ; P3_U3688
g7486 and P3_U4604 P3_U4603 P3_U3688 ; P3_U3689
g7487 and P3_U4607 P3_U4606 ; P3_U3690
g7488 and P3_U5476 P3_U3389 ; P3_U3691
g7489 and P3_U5479 P3_U3388 ; P3_U3692
g7490 and P3_U3920 P3_U3379 ; P3_U3693
g7491 and P3_U5440 P3_STATE_REG_SCAN_IN ; P3_U3694
g7492 and P3_U5424 P3_U3364 ; P3_U3695
g7493 and P3_U3375 P3_STATE_REG_SCAN_IN ; P3_U3696
g7494 and P3_U3301 P3_U3308 P3_U3305 P3_U3306 P3_U3307 ; P3_U3697
g7495 and P3_U3309 P3_U3360 ; P3_U3698
g7496 and P3_U4763 P3_U4762 P3_U4765 P3_U3701 ; P3_U3699
g7497 and P3_U4768 P3_U4766 ; P3_U3700
g7498 and P3_U3700 P3_U4767 ; P3_U3701
g7499 and P3_U4774 P3_U4773 P3_U4776 P3_U3704 ; P3_U3702
g7500 and P3_U4779 P3_U4777 ; P3_U3703
g7501 and P3_U3703 P3_U4778 ; P3_U3704
g7502 and P3_U4785 P3_U4784 P3_U4787 P3_U3707 ; P3_U3705
g7503 and P3_U4790 P3_U4788 ; P3_U3706
g7504 and P3_U3706 P3_U4789 ; P3_U3707
g7505 and P3_U4796 P3_U4795 P3_U4798 P3_U3710 ; P3_U3708
g7506 and P3_U4801 P3_U4799 ; P3_U3709
g7507 and P3_U3709 P3_U4800 ; P3_U3710
g7508 and P3_U4807 P3_U4806 P3_U4809 P3_U3713 ; P3_U3711
g7509 and P3_U4812 P3_U4810 ; P3_U3712
g7510 and P3_U3712 P3_U4811 ; P3_U3713
g7511 and P3_U4818 P3_U4817 P3_U4820 P3_U3716 ; P3_U3714
g7512 and P3_U4823 P3_U4821 ; P3_U3715
g7513 and P3_U3715 P3_U4822 ; P3_U3716
g7514 and P3_U4829 P3_U4828 P3_U4831 P3_U3719 ; P3_U3717
g7515 and P3_U4834 P3_U4832 ; P3_U3718
g7516 and P3_U3718 P3_U4833 ; P3_U3719
g7517 and P3_U4840 P3_U4839 P3_U4842 P3_U3722 ; P3_U3720
g7518 and P3_U4845 P3_U4843 ; P3_U3721
g7519 and P3_U3721 P3_U4844 ; P3_U3722
g7520 and P3_U4851 P3_U4850 P3_U4853 P3_U3725 ; P3_U3723
g7521 and P3_U4856 P3_U4854 ; P3_U3724
g7522 and P3_U3724 P3_U4855 ; P3_U3725
g7523 and P3_U4862 P3_U4861 P3_U4864 P3_U3728 ; P3_U3726
g7524 and P3_U4867 P3_U4865 ; P3_U3727
g7525 and P3_U3727 P3_U4866 ; P3_U3728
g7526 and P3_U4873 P3_U4872 P3_U4875 P3_U3731 ; P3_U3729
g7527 and P3_U4878 P3_U4876 ; P3_U3730
g7528 and P3_U3730 P3_U4877 ; P3_U3731
g7529 and P3_U4884 P3_U4886 P3_U4883 P3_U3734 ; P3_U3732
g7530 and P3_U4889 P3_U4887 ; P3_U3733
g7531 and P3_U3733 P3_U4888 ; P3_U3734
g7532 and P3_U4895 P3_U4897 P3_U4894 P3_U3737 ; P3_U3735
g7533 and P3_U4900 P3_U4898 ; P3_U3736
g7534 and P3_U3736 P3_U4899 ; P3_U3737
g7535 and P3_U4908 P3_U4906 P3_U3740 ; P3_U3738
g7536 and P3_U4911 P3_U4909 ; P3_U3739
g7537 and P3_U3739 P3_U4910 ; P3_U3740
g7538 and P3_U4919 P3_U4917 ; P3_U3741
g7539 and P3_U4922 P3_U4920 ; P3_U3742
g7540 and P3_U3742 P3_U4921 ; P3_U3743
g7541 and P3_U4928 P3_U3746 P3_U4927 ; P3_U3744
g7542 and P3_U4933 P3_U4931 ; P3_U3745
g7543 and P3_U3745 P3_U4932 ; P3_U3746
g7544 and P3_U4939 P3_U3749 P3_U4938 ; P3_U3747
g7545 and P3_U4944 P3_U4942 ; P3_U3748
g7546 and P3_U3748 P3_U4943 ; P3_U3749
g7547 and P3_U4950 P3_U4952 P3_U4949 P3_U3752 ; P3_U3750
g7548 and P3_U4955 P3_U4953 ; P3_U3751
g7549 and P3_U3751 P3_U4954 ; P3_U3752
g7550 and P3_U4961 P3_U4960 P3_U4963 P3_U3755 ; P3_U3753
g7551 and P3_U4966 P3_U4964 ; P3_U3754
g7552 and P3_U3754 P3_U4965 ; P3_U3755
g7553 and P3_U4972 P3_U4971 P3_U4974 P3_U3758 ; P3_U3756
g7554 and P3_U4977 P3_U4975 ; P3_U3757
g7555 and P3_U3757 P3_U4976 ; P3_U3758
g7556 and P3_U5468 P3_U3383 ; P3_U3759
g7557 nand P3_U5834 P3_U5833 ; P3_U3760
g7558 and P3_U5915 P3_U5912 ; P3_U3761
g7559 and P3_U3764 P3_U3763 P3_U3761 P3_U5897 ; P3_U3762
g7560 and P3_U5903 P3_U5900 ; P3_U3763
g7561 and P3_U5909 P3_U5906 ; P3_U3764
g7562 and P3_U5885 P3_U5882 P3_U5879 ; P3_U3765
g7563 and P3_U5894 P3_U5891 P3_U5888 ; P3_U3766
g7564 and P3_U3766 P3_U3765 P3_U5876 P3_U5873 ; P3_U3767
g7565 and P3_U5867 P3_U5864 P3_U5861 P3_U5858 ; P3_U3768
g7566 and P3_U5855 P3_U5852 ; P3_U3769
g7567 and P3_U5930 P3_U5927 P3_U5924 P3_U5921 ; P3_U3770
g7568 and P3_U5843 P3_U5840 P3_U5846 ; P3_U3771
g7569 and P3_U3768 P3_U3769 P3_U5870 P3_U5849 P3_U3771 ; P3_U3772
g7570 and P3_U3762 P3_U3767 P3_U5918 P3_U3770 P3_U5933 ; P3_U3773
g7571 and P3_U4981 P3_U3870 P3_U4980 ; P3_U3774
g7572 and P3_U5416 P3_U5415 ; P3_U3775
g7573 and P3_U5440 P3_U3362 P3_U4990 P3_U3880 ; P3_U3776
g7574 and P3_U4998 P3_U4997 ; P3_U3777
g7575 and P3_U5011 P3_U5010 ; P3_U3778
g7576 and P3_U5020 P3_U5019 ; P3_U3779
g7577 and P3_U5029 P3_U5028 ; P3_U3780
g7578 and P3_U5036 P3_U5034 ; P3_U3781
g7579 and P3_U5038 P3_U5037 ; P3_U3782
g7580 and P3_U5047 P3_U5046 ; P3_U3783
g7581 and P3_U5056 P3_U5055 ; P3_U3784
g7582 and P3_U5065 P3_U5064 ; P3_U3785
g7583 and P3_U5074 P3_U5073 ; P3_U3786
g7584 and P3_U3031 P3_U3077 ; P3_U3787
g7585 and P3_U5078 P3_U5077 ; P3_U3788
g7586 and P3_U5081 P3_U5080 P3_U3788 ; P3_U3789
g7587 and P3_U5090 P3_U5089 ; P3_U3790
g7588 and P3_U5097 P3_U5095 ; P3_U3791
g7589 and P3_U5099 P3_U5098 ; P3_U3792
g7590 and P3_U5108 P3_U5107 ; P3_U3793
g7591 and P3_U5117 P3_U5116 ; P3_U3794
g7592 and P3_U5126 P3_U5125 ; P3_U3795
g7593 and P3_U5135 P3_U5134 ; P3_U3796
g7594 and P3_U5144 P3_U5143 ; P3_U3797
g7595 and P3_U5153 P3_U5152 ; P3_U3798
g7596 and P3_U5162 P3_U5161 ; P3_U3799
g7597 and P3_U5169 P3_U5167 ; P3_U3800
g7598 and P3_U5171 P3_U5170 ; P3_U3801
g7599 and P3_U5180 P3_U5179 ; P3_U3802
g7600 and P3_U5189 P3_U5188 ; P3_U3803
g7601 and P3_U5198 P3_U5197 ; P3_U3804
g7602 and P3_U5205 P3_U5203 ; P3_U3805
g7603 and P3_U5207 P3_U5206 ; P3_U3806
g7604 and P3_U5216 P3_U5215 ; P3_U3807
g7605 and P3_U5225 P3_U5224 ; P3_U3808
g7606 and P3_U5234 P3_U5233 ; P3_U3809
g7607 and P3_U5243 P3_U5242 ; P3_U3810
g7608 and P3_U5252 P3_U5251 ; P3_U3811
g7609 and P3_U5254 P3_STATE_REG_SCAN_IN ; P3_U3812
g7610 and P3_U5440 P3_U3385 ; P3_U3813
g7611 and P3_U3385 P3_U3375 ; P3_U3814
g7612 and P3_U3875 P3_U3312 P3_U3302 ; P3_U3815
g7613 and P3_U3357 P3_U3877 P3_U3310 ; P3_U3816
g7614 and P3_U3375 P3_U5258 ; P3_U3817
g7615 and P3_U3375 P3_U5260 ; P3_U3818
g7616 and P3_U3375 P3_U5262 ; P3_U3819
g7617 and P3_U3375 P3_U5264 ; P3_U3820
g7618 and P3_U3375 P3_U5266 ; P3_U3821
g7619 and P3_U3375 P3_U5268 ; P3_U3822
g7620 and P3_U3375 P3_U5274 ; P3_U3823
g7621 and P3_U3375 P3_U5296 ; P3_U3824
g7622 and P3_U3375 P3_U5310 ; P3_U3825
g7623 and P3_U3375 P3_U5312 ; P3_U3826
g7624 and P3_U3375 P3_U5314 ; P3_U3827
g7625 and P3_U3375 P3_U5316 ; P3_U3828
g7626 and P3_U3375 P3_U5318 ; P3_U3829
g7627 and P3_U3375 P3_U5320 ; P3_U3830
g7628 not P3_IR_REG_31__SCAN_IN ; P3_U3831
g7629 nand P3_U3023 P3_U3300 ; P3_U3832
g7630 nand P3_U5468 P3_U5465 ; P3_U3833
g7631 nand P3_U5456 P3_U5447 ; P3_U3834
g7632 nand P3_U3023 P3_U4058 ; P3_U3835
g7633 nand P3_U3023 P3_U4622 ; P3_U3836
g7634 and P3_U5707 P3_U5706 ; P3_U3837
g7635 and P3_U5709 P3_U5708 ; P3_U3838
g7636 and P3_U5711 P3_U5710 ; P3_U3839
g7637 and P3_U5713 P3_U5712 ; P3_U3840
g7638 and P3_U5715 P3_U5714 ; P3_U3841
g7639 and P3_U5717 P3_U5716 ; P3_U3842
g7640 and P3_U5719 P3_U5718 ; P3_U3843
g7641 and P3_U5721 P3_U5720 ; P3_U3844
g7642 and P3_U5723 P3_U5722 ; P3_U3845
g7643 and P3_U5725 P3_U5724 ; P3_U3846
g7644 and P3_U5727 P3_U5726 ; P3_U3847
g7645 and P3_U5729 P3_U5728 ; P3_U3848
g7646 and P3_U5731 P3_U5730 ; P3_U3849
g7647 and P3_U5733 P3_U5732 ; P3_U3850
g7648 and P3_U5735 P3_U5734 ; P3_U3851
g7649 and P3_U5737 P3_U5736 ; P3_U3852
g7650 and P3_U5739 P3_U5738 ; P3_U3853
g7651 and P3_U5741 P3_U5740 ; P3_U3854
g7652 and P3_U5743 P3_U5742 ; P3_U3855
g7653 and P3_U5745 P3_U5744 ; P3_U3856
g7654 and P3_U5747 P3_U5746 ; P3_U3857
g7655 and P3_U5749 P3_U5748 ; P3_U3858
g7656 and P3_U5751 P3_U5750 ; P3_U3859
g7657 and P3_U5753 P3_U5752 ; P3_U3860
g7658 and P3_U5755 P3_U5754 ; P3_U3861
g7659 and P3_U5757 P3_U5756 ; P3_U3862
g7660 and P3_U5759 P3_U5758 ; P3_U3863
g7661 and P3_U5761 P3_U5760 ; P3_U3864
g7662 and P3_U5763 P3_U5762 ; P3_U3865
g7663 and P3_U5765 P3_U5764 ; P3_U3866
g7664 not P3_R1269_U11 ; P3_U3867
g7665 nand P3_U3773 P3_U3772 ; P3_U3868
g7666 not P3_R693_U14 ; P3_U3869
g7667 and P3_U5940 P3_U5939 ; P3_U3870
g7668 not P3_R1297_U6 ; P3_U3871
g7669 not P3_U3356 ; P3_U3872
g7670 not P3_U3355 ; P3_U3873
g7671 not P3_U3312 ; P3_U3874
g7672 nand P3_U3015 P3_U3385 ; P3_U3875
g7673 not P3_U3302 ; P3_U3876
g7674 nand P3_U3016 P3_U5456 ; P3_U3877
g7675 not P3_U3310 ; P3_U3878
g7676 not P3_U3357 ; P3_U3879
g7677 nand P3_U3014 P3_U3385 ; P3_U3880
g7678 not P3_U3308 ; P3_U3881
g7679 not P3_U3301 ; P3_U3882
g7680 not P3_U3305 ; P3_U3883
g7681 not P3_U3307 ; P3_U3884
g7682 not P3_U3306 ; P3_U3885
g7683 not P3_U3360 ; P3_U3886
g7684 not P3_U3311 ; P3_U3887
g7685 nand P3_U3878 P3_U3378 ; P3_U3888
g7686 not P3_U3369 ; P3_U3889
g7687 not P3_U3367 ; P3_U3890
g7688 not P3_U3309 ; P3_U3891
g7689 not P3_U3352 ; P3_U3892
g7690 not P3_U3833 ; P3_U3893
g7691 not P3_U3303 ; P3_U3894
g7692 not P3_U3304 ; P3_U3895
g7693 nand P3_U5465 P3_U3384 ; P3_U3896
g7694 not P3_U3363 ; P3_U3897
g7695 not P3_U3364 ; P3_U3898
g7696 not P3_U3350 ; P3_U3899
g7697 not P3_U3348 ; P3_U3900
g7698 not P3_U3346 ; P3_U3901
g7699 not P3_U3344 ; P3_U3902
g7700 not P3_U3342 ; P3_U3903
g7701 not P3_U3340 ; P3_U3904
g7702 not P3_U3338 ; P3_U3905
g7703 not P3_U3336 ; P3_U3906
g7704 not P3_U3334 ; P3_U3907
g7705 not P3_U3353 ; P3_U3908
g7706 not P3_U3368 ; P3_U3909
g7707 not P3_U3362 ; P3_U3910
g7708 not P3_U3313 ; P3_U3911
g7709 not P3_U3358 ; P3_U3912
g7710 not P3_U3836 ; P3_U3913
g7711 not P3_U3835 ; P3_U3914
g7712 not P3_U3832 ; P3_U3915
g7713 not P3_U3361 ; P3_U3916
g7714 nand P3_U3370 P3_STATE_REG_SCAN_IN ; P3_U3917
g7715 nand P3_U3886 P3_U3023 ; P3_U3918
g7716 not P3_U3299 ; P3_U3919
g7717 not P3_U3359 ; P3_U3920
g7718 not P3_U3297 ; P3_U3921
g7719 nand U61 P3_U3151 ; P3_U3922
g7720 nand P3_U3027 P3_IR_REG_0__SCAN_IN ; P3_U3923
g7721 nand P3_U3921 P3_IR_REG_0__SCAN_IN ; P3_U3924
g7722 nand U50 P3_U3151 ; P3_U3925
g7723 nand P3_SUB_598_U51 P3_U3027 ; P3_U3926
g7724 nand P3_U3921 P3_IR_REG_1__SCAN_IN ; P3_U3927
g7725 nand U39 P3_U3151 ; P3_U3928
g7726 nand P3_SUB_598_U22 P3_U3027 ; P3_U3929
g7727 nand P3_U3921 P3_IR_REG_2__SCAN_IN ; P3_U3930
g7728 nand U36 P3_U3151 ; P3_U3931
g7729 nand P3_SUB_598_U23 P3_U3027 ; P3_U3932
g7730 nand P3_U3921 P3_IR_REG_3__SCAN_IN ; P3_U3933
g7731 nand U35 P3_U3151 ; P3_U3934
g7732 nand P3_SUB_598_U24 P3_U3027 ; P3_U3935
g7733 nand P3_U3921 P3_IR_REG_4__SCAN_IN ; P3_U3936
g7734 nand U34 P3_U3151 ; P3_U3937
g7735 nand P3_SUB_598_U74 P3_U3027 ; P3_U3938
g7736 nand P3_U3921 P3_IR_REG_5__SCAN_IN ; P3_U3939
g7737 nand U33 P3_U3151 ; P3_U3940
g7738 nand P3_SUB_598_U25 P3_U3027 ; P3_U3941
g7739 nand P3_U3921 P3_IR_REG_6__SCAN_IN ; P3_U3942
g7740 nand U32 P3_U3151 ; P3_U3943
g7741 nand P3_SUB_598_U26 P3_U3027 ; P3_U3944
g7742 nand P3_U3921 P3_IR_REG_7__SCAN_IN ; P3_U3945
g7743 nand U31 P3_U3151 ; P3_U3946
g7744 nand P3_SUB_598_U27 P3_U3027 ; P3_U3947
g7745 nand P3_U3921 P3_IR_REG_8__SCAN_IN ; P3_U3948
g7746 nand U30 P3_U3151 ; P3_U3949
g7747 nand P3_SUB_598_U72 P3_U3027 ; P3_U3950
g7748 nand P3_U3921 P3_IR_REG_9__SCAN_IN ; P3_U3951
g7749 nand U60 P3_U3151 ; P3_U3952
g7750 nand P3_SUB_598_U7 P3_U3027 ; P3_U3953
g7751 nand P3_U3921 P3_IR_REG_10__SCAN_IN ; P3_U3954
g7752 nand U59 P3_U3151 ; P3_U3955
g7753 nand P3_SUB_598_U8 P3_U3027 ; P3_U3956
g7754 nand P3_U3921 P3_IR_REG_11__SCAN_IN ; P3_U3957
g7755 nand U58 P3_U3151 ; P3_U3958
g7756 nand P3_SUB_598_U9 P3_U3027 ; P3_U3959
g7757 nand P3_U3921 P3_IR_REG_12__SCAN_IN ; P3_U3960
g7758 nand U57 P3_U3151 ; P3_U3961
g7759 nand P3_SUB_598_U89 P3_U3027 ; P3_U3962
g7760 nand P3_U3921 P3_IR_REG_13__SCAN_IN ; P3_U3963
g7761 nand U56 P3_U3151 ; P3_U3964
g7762 nand P3_SUB_598_U10 P3_U3027 ; P3_U3965
g7763 nand P3_U3921 P3_IR_REG_14__SCAN_IN ; P3_U3966
g7764 nand U55 P3_U3151 ; P3_U3967
g7765 nand P3_SUB_598_U11 P3_U3027 ; P3_U3968
g7766 nand P3_U3921 P3_IR_REG_15__SCAN_IN ; P3_U3969
g7767 nand U54 P3_U3151 ; P3_U3970
g7768 nand P3_SUB_598_U12 P3_U3027 ; P3_U3971
g7769 nand P3_U3921 P3_IR_REG_16__SCAN_IN ; P3_U3972
g7770 nand U53 P3_U3151 ; P3_U3973
g7771 nand P3_SUB_598_U87 P3_U3027 ; P3_U3974
g7772 nand P3_U3921 P3_IR_REG_17__SCAN_IN ; P3_U3975
g7773 nand U52 P3_U3151 ; P3_U3976
g7774 nand P3_SUB_598_U13 P3_U3027 ; P3_U3977
g7775 nand P3_U3921 P3_IR_REG_18__SCAN_IN ; P3_U3978
g7776 nand U51 P3_U3151 ; P3_U3979
g7777 nand P3_SUB_598_U14 P3_U3027 ; P3_U3980
g7778 nand P3_U3921 P3_IR_REG_19__SCAN_IN ; P3_U3981
g7779 nand U49 P3_U3151 ; P3_U3982
g7780 nand P3_SUB_598_U15 P3_U3027 ; P3_U3983
g7781 nand P3_U3921 P3_IR_REG_20__SCAN_IN ; P3_U3984
g7782 nand U48 P3_U3151 ; P3_U3985
g7783 nand P3_SUB_598_U83 P3_U3027 ; P3_U3986
g7784 nand P3_U3921 P3_IR_REG_21__SCAN_IN ; P3_U3987
g7785 nand U47 P3_U3151 ; P3_U3988
g7786 nand P3_SUB_598_U16 P3_U3027 ; P3_U3989
g7787 nand P3_U3921 P3_IR_REG_22__SCAN_IN ; P3_U3990
g7788 nand U46 P3_U3151 ; P3_U3991
g7789 nand P3_SUB_598_U17 P3_U3027 ; P3_U3992
g7790 nand P3_U3921 P3_IR_REG_23__SCAN_IN ; P3_U3993
g7791 nand U45 P3_U3151 ; P3_U3994
g7792 nand P3_SUB_598_U18 P3_U3027 ; P3_U3995
g7793 nand P3_U3921 P3_IR_REG_24__SCAN_IN ; P3_U3996
g7794 nand U44 P3_U3151 ; P3_U3997
g7795 nand P3_SUB_598_U81 P3_U3027 ; P3_U3998
g7796 nand P3_U3921 P3_IR_REG_25__SCAN_IN ; P3_U3999
g7797 nand U43 P3_U3151 ; P3_U4000
g7798 nand P3_SUB_598_U19 P3_U3027 ; P3_U4001
g7799 nand P3_U3921 P3_IR_REG_26__SCAN_IN ; P3_U4002
g7800 nand U42 P3_U3151 ; P3_U4003
g7801 nand P3_SUB_598_U79 P3_U3027 ; P3_U4004
g7802 nand P3_U3921 P3_IR_REG_27__SCAN_IN ; P3_U4005
g7803 nand U41 P3_U3151 ; P3_U4006
g7804 nand P3_SUB_598_U20 P3_U3027 ; P3_U4007
g7805 nand P3_U3921 P3_IR_REG_28__SCAN_IN ; P3_U4008
g7806 nand U40 P3_U3151 ; P3_U4009
g7807 nand P3_SUB_598_U21 P3_U3027 ; P3_U4010
g7808 nand P3_U3921 P3_IR_REG_29__SCAN_IN ; P3_U4011
g7809 nand U38 P3_U3151 ; P3_U4012
g7810 nand P3_SUB_598_U77 P3_U3027 ; P3_U4013
g7811 nand P3_U3921 P3_IR_REG_30__SCAN_IN ; P3_U4014
g7812 nand U37 P3_U3151 ; P3_U4015
g7813 nand P3_SUB_598_U52 P3_U3027 ; P3_U4016
g7814 nand P3_U3921 P3_IR_REG_31__SCAN_IN ; P3_U4017
g7815 nand P3_U3919 P3_U5437 ; P3_U4018
g7816 not P3_U3300 ; P3_U4019
g7817 nand P3_U3299 P3_U5428 ; P3_U4020
g7818 nand P3_U3299 P3_U5431 ; P3_U4021
g7819 nand P3_U4019 P3_D_REG_10__SCAN_IN ; P3_U4022
g7820 nand P3_U4019 P3_D_REG_11__SCAN_IN ; P3_U4023
g7821 nand P3_U4019 P3_D_REG_12__SCAN_IN ; P3_U4024
g7822 nand P3_U4019 P3_D_REG_13__SCAN_IN ; P3_U4025
g7823 nand P3_U4019 P3_D_REG_14__SCAN_IN ; P3_U4026
g7824 nand P3_U4019 P3_D_REG_15__SCAN_IN ; P3_U4027
g7825 nand P3_U4019 P3_D_REG_16__SCAN_IN ; P3_U4028
g7826 nand P3_U4019 P3_D_REG_17__SCAN_IN ; P3_U4029
g7827 nand P3_U4019 P3_D_REG_18__SCAN_IN ; P3_U4030
g7828 nand P3_U4019 P3_D_REG_19__SCAN_IN ; P3_U4031
g7829 nand P3_U4019 P3_D_REG_20__SCAN_IN ; P3_U4032
g7830 nand P3_U4019 P3_D_REG_21__SCAN_IN ; P3_U4033
g7831 nand P3_U4019 P3_D_REG_22__SCAN_IN ; P3_U4034
g7832 nand P3_U4019 P3_D_REG_23__SCAN_IN ; P3_U4035
g7833 nand P3_U4019 P3_D_REG_24__SCAN_IN ; P3_U4036
g7834 nand P3_U4019 P3_D_REG_25__SCAN_IN ; P3_U4037
g7835 nand P3_U4019 P3_D_REG_26__SCAN_IN ; P3_U4038
g7836 nand P3_U4019 P3_D_REG_27__SCAN_IN ; P3_U4039
g7837 nand P3_U4019 P3_D_REG_28__SCAN_IN ; P3_U4040
g7838 nand P3_U4019 P3_D_REG_29__SCAN_IN ; P3_U4041
g7839 nand P3_U4019 P3_D_REG_2__SCAN_IN ; P3_U4042
g7840 nand P3_U4019 P3_D_REG_30__SCAN_IN ; P3_U4043
g7841 nand P3_U4019 P3_D_REG_31__SCAN_IN ; P3_U4044
g7842 nand P3_U4019 P3_D_REG_3__SCAN_IN ; P3_U4045
g7843 nand P3_U4019 P3_D_REG_4__SCAN_IN ; P3_U4046
g7844 nand P3_U4019 P3_D_REG_5__SCAN_IN ; P3_U4047
g7845 nand P3_U4019 P3_D_REG_6__SCAN_IN ; P3_U4048
g7846 nand P3_U4019 P3_D_REG_7__SCAN_IN ; P3_U4049
g7847 nand P3_U4019 P3_D_REG_8__SCAN_IN ; P3_U4050
g7848 nand P3_U4019 P3_D_REG_9__SCAN_IN ; P3_U4051
g7849 not P3_U3834 ; P3_U4052
g7850 nand P3_U5456 P3_U5450 ; P3_U4053
g7851 nand P3_U5482 P3_U4053 ; P3_U4054
g7852 nand P3_U3369 P3_U3367 ; P3_U4055
g7853 nand P3_U3894 P3_U4055 ; P3_U4056
g7854 nand P3_U3895 P3_U4054 ; P3_U4057
g7855 nand P3_U4057 P3_U4056 ; P3_U4058
g7856 nand P3_U3022 P3_REG0_REG_1__SCAN_IN ; P3_U4059
g7857 nand P3_U3021 P3_REG1_REG_1__SCAN_IN ; P3_U4060
g7858 nand P3_U3020 P3_REG2_REG_1__SCAN_IN ; P3_U4061
g7859 nand P3_U3019 P3_REG3_REG_1__SCAN_IN ; P3_U4062
g7860 not P3_U3077 ; P3_U4063
g7861 nand P3_U3877 P3_U3357 ; P3_U4064
g7862 nand P3_U3883 P3_R1110_U95 ; P3_U4065
g7863 nand P3_U3885 P3_R1077_U95 ; P3_U4066
g7864 nand P3_U3884 P3_R1095_U24 ; P3_U4067
g7865 nand P3_U3881 P3_R1143_U95 ; P3_U4068
g7866 nand P3_U3891 P3_R1161_U95 ; P3_U4069
g7867 nand P3_U3887 P3_R1131_U24 ; P3_U4070
g7868 nand P3_U3017 P3_R1200_U24 ; P3_U4071
g7869 not P3_U3314 ; P3_U4072
g7870 nand P3_U3352 P3_U3833 ; P3_U4073
g7871 nand P3_R1179_U24 P3_U3026 ; P3_U4074
g7872 nand P3_U3025 P3_U3077 ; P3_U4075
g7873 nand P3_U3387 P3_U4064 ; P3_U4076
g7874 nand P3_U3577 P3_U4072 ; P3_U4077
g7875 nand P3_U3022 P3_REG0_REG_2__SCAN_IN ; P3_U4078
g7876 nand P3_U3021 P3_REG1_REG_2__SCAN_IN ; P3_U4079
g7877 nand P3_U3020 P3_REG2_REG_2__SCAN_IN ; P3_U4080
g7878 nand P3_U3019 P3_REG3_REG_2__SCAN_IN ; P3_U4081
g7879 not P3_U3067 ; P3_U4082
g7880 nand P3_U3022 P3_REG0_REG_0__SCAN_IN ; P3_U4083
g7881 nand P3_U3021 P3_REG1_REG_0__SCAN_IN ; P3_U4084
g7882 nand P3_U3020 P3_REG2_REG_0__SCAN_IN ; P3_U4085
g7883 nand P3_U3019 P3_REG3_REG_0__SCAN_IN ; P3_U4086
g7884 not P3_U3076 ; P3_U4087
g7885 nand P3_U5468 P3_U3383 ; P3_U4088
g7886 nand P3_U3896 P3_U4088 ; P3_U4089
g7887 nand P3_U3033 P3_U3076 ; P3_U4090
g7888 nand P3_R1110_U94 P3_U3883 ; P3_U4091
g7889 nand P3_R1077_U94 P3_U3885 ; P3_U4092
g7890 nand P3_R1095_U100 P3_U3884 ; P3_U4093
g7891 nand P3_R1143_U94 P3_U3881 ; P3_U4094
g7892 nand P3_R1161_U94 P3_U3891 ; P3_U4095
g7893 nand P3_R1131_U100 P3_U3887 ; P3_U4096
g7894 nand P3_R1200_U100 P3_U3017 ; P3_U4097
g7895 not P3_U3315 ; P3_U4098
g7896 nand P3_R1179_U100 P3_U3026 ; P3_U4099
g7897 nand P3_U3025 P3_U3067 ; P3_U4100
g7898 nand P3_U3392 P3_U4064 ; P3_U4101
g7899 nand P3_U3593 P3_U4098 ; P3_U4102
g7900 nand P3_U3022 P3_REG0_REG_3__SCAN_IN ; P3_U4103
g7901 nand P3_U3021 P3_REG1_REG_3__SCAN_IN ; P3_U4104
g7902 nand P3_U3020 P3_REG2_REG_3__SCAN_IN ; P3_U4105
g7903 nand P3_SUB_609_U25 P3_U3019 ; P3_U4106
g7904 not P3_U3063 ; P3_U4107
g7905 nand P3_U3033 P3_U3077 ; P3_U4108
g7906 nand P3_R1110_U16 P3_U3883 ; P3_U4109
g7907 nand P3_R1077_U16 P3_U3885 ; P3_U4110
g7908 nand P3_R1095_U110 P3_U3884 ; P3_U4111
g7909 nand P3_R1143_U16 P3_U3881 ; P3_U4112
g7910 nand P3_R1161_U16 P3_U3891 ; P3_U4113
g7911 nand P3_R1131_U110 P3_U3887 ; P3_U4114
g7912 nand P3_R1200_U110 P3_U3017 ; P3_U4115
g7913 not P3_U3316 ; P3_U4116
g7914 nand P3_R1179_U110 P3_U3026 ; P3_U4117
g7915 nand P3_U3025 P3_U3063 ; P3_U4118
g7916 nand P3_U3395 P3_U4064 ; P3_U4119
g7917 nand P3_U3597 P3_U4116 ; P3_U4120
g7918 nand P3_U3022 P3_REG0_REG_4__SCAN_IN ; P3_U4121
g7919 nand P3_U3021 P3_REG1_REG_4__SCAN_IN ; P3_U4122
g7920 nand P3_U3020 P3_REG2_REG_4__SCAN_IN ; P3_U4123
g7921 nand P3_SUB_609_U29 P3_U3019 ; P3_U4124
g7922 not P3_U3059 ; P3_U4125
g7923 nand P3_U3033 P3_U3067 ; P3_U4126
g7924 nand P3_R1110_U100 P3_U3883 ; P3_U4127
g7925 nand P3_R1077_U100 P3_U3885 ; P3_U4128
g7926 nand P3_R1095_U21 P3_U3884 ; P3_U4129
g7927 nand P3_R1143_U100 P3_U3881 ; P3_U4130
g7928 nand P3_R1161_U100 P3_U3891 ; P3_U4131
g7929 nand P3_R1131_U21 P3_U3887 ; P3_U4132
g7930 nand P3_R1200_U21 P3_U3017 ; P3_U4133
g7931 not P3_U3317 ; P3_U4134
g7932 nand P3_R1179_U21 P3_U3026 ; P3_U4135
g7933 nand P3_U3025 P3_U3059 ; P3_U4136
g7934 nand P3_U3398 P3_U4064 ; P3_U4137
g7935 nand P3_U3601 P3_U4134 ; P3_U4138
g7936 nand P3_U3022 P3_REG0_REG_5__SCAN_IN ; P3_U4139
g7937 nand P3_U3021 P3_REG1_REG_5__SCAN_IN ; P3_U4140
g7938 nand P3_U3020 P3_REG2_REG_5__SCAN_IN ; P3_U4141
g7939 nand P3_SUB_609_U53 P3_U3019 ; P3_U4142
g7940 not P3_U3066 ; P3_U4143
g7941 nand P3_U3033 P3_U3063 ; P3_U4144
g7942 nand P3_R1110_U99 P3_U3883 ; P3_U4145
g7943 nand P3_R1077_U99 P3_U3885 ; P3_U4146
g7944 nand P3_R1095_U109 P3_U3884 ; P3_U4147
g7945 nand P3_R1143_U99 P3_U3881 ; P3_U4148
g7946 nand P3_R1161_U99 P3_U3891 ; P3_U4149
g7947 nand P3_R1131_U109 P3_U3887 ; P3_U4150
g7948 nand P3_R1200_U109 P3_U3017 ; P3_U4151
g7949 not P3_U3318 ; P3_U4152
g7950 nand P3_R1179_U109 P3_U3026 ; P3_U4153
g7951 nand P3_U3025 P3_U3066 ; P3_U4154
g7952 nand P3_U3401 P3_U4064 ; P3_U4155
g7953 nand P3_U3604 P3_U4152 ; P3_U4156
g7954 nand P3_U3022 P3_REG0_REG_6__SCAN_IN ; P3_U4157
g7955 nand P3_U3021 P3_REG1_REG_6__SCAN_IN ; P3_U4158
g7956 nand P3_U3020 P3_REG2_REG_6__SCAN_IN ; P3_U4159
g7957 nand P3_SUB_609_U8 P3_U3019 ; P3_U4160
g7958 not P3_U3070 ; P3_U4161
g7959 nand P3_U3033 P3_U3059 ; P3_U4162
g7960 nand P3_R1110_U17 P3_U3883 ; P3_U4163
g7961 nand P3_R1077_U17 P3_U3885 ; P3_U4164
g7962 nand P3_R1095_U108 P3_U3884 ; P3_U4165
g7963 nand P3_R1143_U17 P3_U3881 ; P3_U4166
g7964 nand P3_R1161_U17 P3_U3891 ; P3_U4167
g7965 nand P3_R1131_U108 P3_U3887 ; P3_U4168
g7966 nand P3_R1200_U108 P3_U3017 ; P3_U4169
g7967 not P3_U3319 ; P3_U4170
g7968 nand P3_R1179_U108 P3_U3026 ; P3_U4171
g7969 nand P3_U3025 P3_U3070 ; P3_U4172
g7970 nand P3_U3404 P3_U4064 ; P3_U4173
g7971 nand P3_U3607 P3_U4170 ; P3_U4174
g7972 nand P3_U3022 P3_REG0_REG_7__SCAN_IN ; P3_U4175
g7973 nand P3_U3021 P3_REG1_REG_7__SCAN_IN ; P3_U4176
g7974 nand P3_U3020 P3_REG2_REG_7__SCAN_IN ; P3_U4177
g7975 nand P3_SUB_609_U18 P3_U3019 ; P3_U4178
g7976 not P3_U3069 ; P3_U4179
g7977 nand P3_U3033 P3_U3066 ; P3_U4180
g7978 nand P3_R1110_U98 P3_U3883 ; P3_U4181
g7979 nand P3_R1077_U98 P3_U3885 ; P3_U4182
g7980 nand P3_R1095_U22 P3_U3884 ; P3_U4183
g7981 nand P3_R1143_U98 P3_U3881 ; P3_U4184
g7982 nand P3_R1161_U98 P3_U3891 ; P3_U4185
g7983 nand P3_R1131_U22 P3_U3887 ; P3_U4186
g7984 nand P3_R1200_U22 P3_U3017 ; P3_U4187
g7985 not P3_U3320 ; P3_U4188
g7986 nand P3_R1179_U22 P3_U3026 ; P3_U4189
g7987 nand P3_U3025 P3_U3069 ; P3_U4190
g7988 nand P3_U3407 P3_U4064 ; P3_U4191
g7989 nand P3_U3610 P3_U4188 ; P3_U4192
g7990 nand P3_U3022 P3_REG0_REG_8__SCAN_IN ; P3_U4193
g7991 nand P3_U3021 P3_REG1_REG_8__SCAN_IN ; P3_U4194
g7992 nand P3_U3020 P3_REG2_REG_8__SCAN_IN ; P3_U4195
g7993 nand P3_SUB_609_U12 P3_U3019 ; P3_U4196
g7994 not P3_U3083 ; P3_U4197
g7995 nand P3_U3033 P3_U3070 ; P3_U4198
g7996 nand P3_R1110_U18 P3_U3883 ; P3_U4199
g7997 nand P3_R1077_U18 P3_U3885 ; P3_U4200
g7998 nand P3_R1095_U107 P3_U3884 ; P3_U4201
g7999 nand P3_R1143_U18 P3_U3881 ; P3_U4202
g8000 nand P3_R1161_U18 P3_U3891 ; P3_U4203
g8001 nand P3_R1131_U107 P3_U3887 ; P3_U4204
g8002 nand P3_R1200_U107 P3_U3017 ; P3_U4205
g8003 not P3_U3321 ; P3_U4206
g8004 nand P3_R1179_U107 P3_U3026 ; P3_U4207
g8005 nand P3_U3025 P3_U3083 ; P3_U4208
g8006 nand P3_U3410 P3_U4064 ; P3_U4209
g8007 nand P3_U3613 P3_U4206 ; P3_U4210
g8008 nand P3_U3022 P3_REG0_REG_9__SCAN_IN ; P3_U4211
g8009 nand P3_U3021 P3_REG1_REG_9__SCAN_IN ; P3_U4212
g8010 nand P3_U3020 P3_REG2_REG_9__SCAN_IN ; P3_U4213
g8011 nand P3_SUB_609_U14 P3_U3019 ; P3_U4214
g8012 not P3_U3082 ; P3_U4215
g8013 nand P3_U3033 P3_U3069 ; P3_U4216
g8014 nand P3_R1110_U97 P3_U3883 ; P3_U4217
g8015 nand P3_R1077_U97 P3_U3885 ; P3_U4218
g8016 nand P3_R1095_U23 P3_U3884 ; P3_U4219
g8017 nand P3_R1143_U97 P3_U3881 ; P3_U4220
g8018 nand P3_R1161_U97 P3_U3891 ; P3_U4221
g8019 nand P3_R1131_U23 P3_U3887 ; P3_U4222
g8020 nand P3_R1200_U23 P3_U3017 ; P3_U4223
g8021 not P3_U3322 ; P3_U4224
g8022 nand P3_R1179_U23 P3_U3026 ; P3_U4225
g8023 nand P3_U3025 P3_U3082 ; P3_U4226
g8024 nand P3_U3413 P3_U4064 ; P3_U4227
g8025 nand P3_U3616 P3_U4224 ; P3_U4228
g8026 nand P3_U3022 P3_REG0_REG_10__SCAN_IN ; P3_U4229
g8027 nand P3_U3021 P3_REG1_REG_10__SCAN_IN ; P3_U4230
g8028 nand P3_U3020 P3_REG2_REG_10__SCAN_IN ; P3_U4231
g8029 nand P3_SUB_609_U13 P3_U3019 ; P3_U4232
g8030 not P3_U3061 ; P3_U4233
g8031 nand P3_U3033 P3_U3083 ; P3_U4234
g8032 nand P3_R1110_U96 P3_U3883 ; P3_U4235
g8033 nand P3_R1077_U96 P3_U3885 ; P3_U4236
g8034 nand P3_R1095_U106 P3_U3884 ; P3_U4237
g8035 nand P3_R1143_U96 P3_U3881 ; P3_U4238
g8036 nand P3_R1161_U96 P3_U3891 ; P3_U4239
g8037 nand P3_R1131_U106 P3_U3887 ; P3_U4240
g8038 nand P3_R1200_U106 P3_U3017 ; P3_U4241
g8039 not P3_U3323 ; P3_U4242
g8040 nand P3_R1179_U106 P3_U3026 ; P3_U4243
g8041 nand P3_U3025 P3_U3061 ; P3_U4244
g8042 nand P3_U3416 P3_U4064 ; P3_U4245
g8043 nand P3_U3620 P3_U4242 ; P3_U4246
g8044 nand P3_U3022 P3_REG0_REG_11__SCAN_IN ; P3_U4247
g8045 nand P3_U3021 P3_REG1_REG_11__SCAN_IN ; P3_U4248
g8046 nand P3_U3020 P3_REG2_REG_11__SCAN_IN ; P3_U4249
g8047 nand P3_SUB_609_U9 P3_U3019 ; P3_U4250
g8048 not P3_U3062 ; P3_U4251
g8049 nand P3_U3033 P3_U3082 ; P3_U4252
g8050 nand P3_R1110_U10 P3_U3883 ; P3_U4253
g8051 nand P3_R1077_U10 P3_U3885 ; P3_U4254
g8052 nand P3_R1095_U116 P3_U3884 ; P3_U4255
g8053 nand P3_R1143_U10 P3_U3881 ; P3_U4256
g8054 nand P3_R1161_U10 P3_U3891 ; P3_U4257
g8055 nand P3_R1131_U116 P3_U3887 ; P3_U4258
g8056 nand P3_R1200_U116 P3_U3017 ; P3_U4259
g8057 not P3_U3324 ; P3_U4260
g8058 nand P3_R1179_U116 P3_U3026 ; P3_U4261
g8059 nand P3_U3025 P3_U3062 ; P3_U4262
g8060 nand P3_U3419 P3_U4064 ; P3_U4263
g8061 nand P3_U3624 P3_U4260 ; P3_U4264
g8062 nand P3_U3022 P3_REG0_REG_12__SCAN_IN ; P3_U4265
g8063 nand P3_U3021 P3_REG1_REG_12__SCAN_IN ; P3_U4266
g8064 nand P3_U3020 P3_REG2_REG_12__SCAN_IN ; P3_U4267
g8065 nand P3_SUB_609_U23 P3_U3019 ; P3_U4268
g8066 not P3_U3071 ; P3_U4269
g8067 nand P3_U3033 P3_U3061 ; P3_U4270
g8068 nand P3_R1110_U114 P3_U3883 ; P3_U4271
g8069 nand P3_R1077_U114 P3_U3885 ; P3_U4272
g8070 nand P3_R1095_U16 P3_U3884 ; P3_U4273
g8071 nand P3_R1143_U114 P3_U3881 ; P3_U4274
g8072 nand P3_R1161_U114 P3_U3891 ; P3_U4275
g8073 nand P3_R1131_U16 P3_U3887 ; P3_U4276
g8074 nand P3_R1200_U16 P3_U3017 ; P3_U4277
g8075 not P3_U3325 ; P3_U4278
g8076 nand P3_R1179_U16 P3_U3026 ; P3_U4279
g8077 nand P3_U3025 P3_U3071 ; P3_U4280
g8078 nand P3_U3422 P3_U4064 ; P3_U4281
g8079 nand P3_U3627 P3_U4278 ; P3_U4282
g8080 nand P3_U3022 P3_REG0_REG_13__SCAN_IN ; P3_U4283
g8081 nand P3_U3021 P3_REG1_REG_13__SCAN_IN ; P3_U4284
g8082 nand P3_U3020 P3_REG2_REG_13__SCAN_IN ; P3_U4285
g8083 nand P3_SUB_609_U24 P3_U3019 ; P3_U4286
g8084 not P3_U3079 ; P3_U4287
g8085 nand P3_U3033 P3_U3062 ; P3_U4288
g8086 nand P3_R1110_U113 P3_U3883 ; P3_U4289
g8087 nand P3_R1077_U113 P3_U3885 ; P3_U4290
g8088 nand P3_R1095_U105 P3_U3884 ; P3_U4291
g8089 nand P3_R1143_U113 P3_U3881 ; P3_U4292
g8090 nand P3_R1161_U113 P3_U3891 ; P3_U4293
g8091 nand P3_R1131_U105 P3_U3887 ; P3_U4294
g8092 nand P3_R1200_U105 P3_U3017 ; P3_U4295
g8093 not P3_U3326 ; P3_U4296
g8094 nand P3_R1179_U105 P3_U3026 ; P3_U4297
g8095 nand P3_U3025 P3_U3079 ; P3_U4298
g8096 nand P3_U3425 P3_U4064 ; P3_U4299
g8097 nand P3_U3631 P3_U4296 ; P3_U4300
g8098 nand P3_U3022 P3_REG0_REG_14__SCAN_IN ; P3_U4301
g8099 nand P3_U3021 P3_REG1_REG_14__SCAN_IN ; P3_U4302
g8100 nand P3_U3020 P3_REG2_REG_14__SCAN_IN ; P3_U4303
g8101 nand P3_SUB_609_U30 P3_U3019 ; P3_U4304
g8102 not P3_U3078 ; P3_U4305
g8103 nand P3_U3033 P3_U3071 ; P3_U4306
g8104 nand P3_R1110_U11 P3_U3883 ; P3_U4307
g8105 nand P3_R1077_U11 P3_U3885 ; P3_U4308
g8106 nand P3_R1095_U104 P3_U3884 ; P3_U4309
g8107 nand P3_R1143_U11 P3_U3881 ; P3_U4310
g8108 nand P3_R1161_U11 P3_U3891 ; P3_U4311
g8109 nand P3_R1131_U104 P3_U3887 ; P3_U4312
g8110 nand P3_R1200_U104 P3_U3017 ; P3_U4313
g8111 not P3_U3327 ; P3_U4314
g8112 nand P3_R1179_U104 P3_U3026 ; P3_U4315
g8113 nand P3_U3025 P3_U3078 ; P3_U4316
g8114 nand P3_U3428 P3_U4064 ; P3_U4317
g8115 nand P3_U3635 P3_U4314 ; P3_U4318
g8116 nand P3_U3022 P3_REG0_REG_15__SCAN_IN ; P3_U4319
g8117 nand P3_U3021 P3_REG1_REG_15__SCAN_IN ; P3_U4320
g8118 nand P3_U3020 P3_REG2_REG_15__SCAN_IN ; P3_U4321
g8119 nand P3_SUB_609_U21 P3_U3019 ; P3_U4322
g8120 not P3_U3073 ; P3_U4323
g8121 nand P3_U3033 P3_U3079 ; P3_U4324
g8122 nand P3_R1110_U112 P3_U3883 ; P3_U4325
g8123 nand P3_R1077_U112 P3_U3885 ; P3_U4326
g8124 nand P3_R1095_U115 P3_U3884 ; P3_U4327
g8125 nand P3_R1143_U112 P3_U3881 ; P3_U4328
g8126 nand P3_R1161_U112 P3_U3891 ; P3_U4329
g8127 nand P3_R1131_U115 P3_U3887 ; P3_U4330
g8128 nand P3_R1200_U115 P3_U3017 ; P3_U4331
g8129 not P3_U3328 ; P3_U4332
g8130 nand P3_R1179_U115 P3_U3026 ; P3_U4333
g8131 nand P3_U3025 P3_U3073 ; P3_U4334
g8132 nand P3_U3431 P3_U4064 ; P3_U4335
g8133 nand P3_U3638 P3_U4332 ; P3_U4336
g8134 nand P3_U3022 P3_REG0_REG_16__SCAN_IN ; P3_U4337
g8135 nand P3_U3021 P3_REG1_REG_16__SCAN_IN ; P3_U4338
g8136 nand P3_U3020 P3_REG2_REG_16__SCAN_IN ; P3_U4339
g8137 nand P3_SUB_609_U7 P3_U3019 ; P3_U4340
g8138 not P3_U3072 ; P3_U4341
g8139 nand P3_U3033 P3_U3078 ; P3_U4342
g8140 nand P3_R1110_U111 P3_U3883 ; P3_U4343
g8141 nand P3_R1077_U111 P3_U3885 ; P3_U4344
g8142 nand P3_R1095_U114 P3_U3884 ; P3_U4345
g8143 nand P3_R1143_U111 P3_U3881 ; P3_U4346
g8144 nand P3_R1161_U111 P3_U3891 ; P3_U4347
g8145 nand P3_R1131_U114 P3_U3887 ; P3_U4348
g8146 nand P3_R1200_U114 P3_U3017 ; P3_U4349
g8147 not P3_U3329 ; P3_U4350
g8148 nand P3_R1179_U114 P3_U3026 ; P3_U4351
g8149 nand P3_U3025 P3_U3072 ; P3_U4352
g8150 nand P3_U3434 P3_U4064 ; P3_U4353
g8151 nand P3_U3641 P3_U4350 ; P3_U4354
g8152 nand P3_U3022 P3_REG0_REG_17__SCAN_IN ; P3_U4355
g8153 nand P3_U3021 P3_REG1_REG_17__SCAN_IN ; P3_U4356
g8154 nand P3_U3020 P3_REG2_REG_17__SCAN_IN ; P3_U4357
g8155 nand P3_SUB_609_U19 P3_U3019 ; P3_U4358
g8156 not P3_U3068 ; P3_U4359
g8157 nand P3_U3033 P3_U3073 ; P3_U4360
g8158 nand P3_R1110_U110 P3_U3883 ; P3_U4361
g8159 nand P3_R1077_U110 P3_U3885 ; P3_U4362
g8160 nand P3_R1095_U17 P3_U3884 ; P3_U4363
g8161 nand P3_R1143_U110 P3_U3881 ; P3_U4364
g8162 nand P3_R1161_U110 P3_U3891 ; P3_U4365
g8163 nand P3_R1131_U17 P3_U3887 ; P3_U4366
g8164 nand P3_R1200_U17 P3_U3017 ; P3_U4367
g8165 not P3_U3330 ; P3_U4368
g8166 nand P3_R1179_U17 P3_U3026 ; P3_U4369
g8167 nand P3_U3025 P3_U3068 ; P3_U4370
g8168 nand P3_U3437 P3_U4064 ; P3_U4371
g8169 nand P3_U3644 P3_U4368 ; P3_U4372
g8170 nand P3_U3022 P3_REG0_REG_18__SCAN_IN ; P3_U4373
g8171 nand P3_U3021 P3_REG1_REG_18__SCAN_IN ; P3_U4374
g8172 nand P3_U3020 P3_REG2_REG_18__SCAN_IN ; P3_U4375
g8173 nand P3_SUB_609_U11 P3_U3019 ; P3_U4376
g8174 not P3_U3081 ; P3_U4377
g8175 nand P3_U3033 P3_U3072 ; P3_U4378
g8176 nand P3_R1110_U12 P3_U3883 ; P3_U4379
g8177 nand P3_R1077_U12 P3_U3885 ; P3_U4380
g8178 nand P3_R1095_U103 P3_U3884 ; P3_U4381
g8179 nand P3_R1143_U12 P3_U3881 ; P3_U4382
g8180 nand P3_R1161_U12 P3_U3891 ; P3_U4383
g8181 nand P3_R1131_U103 P3_U3887 ; P3_U4384
g8182 nand P3_R1200_U103 P3_U3017 ; P3_U4385
g8183 not P3_U3331 ; P3_U4386
g8184 nand P3_R1179_U103 P3_U3026 ; P3_U4387
g8185 nand P3_U3025 P3_U3081 ; P3_U4388
g8186 nand P3_U3440 P3_U4064 ; P3_U4389
g8187 nand P3_U3648 P3_U4386 ; P3_U4390
g8188 nand P3_U3022 P3_REG0_REG_19__SCAN_IN ; P3_U4391
g8189 nand P3_U3021 P3_REG1_REG_19__SCAN_IN ; P3_U4392
g8190 nand P3_U3020 P3_REG2_REG_19__SCAN_IN ; P3_U4393
g8191 nand P3_SUB_609_U15 P3_U3019 ; P3_U4394
g8192 not P3_U3080 ; P3_U4395
g8193 nand P3_U3033 P3_U3068 ; P3_U4396
g8194 nand P3_R1110_U109 P3_U3883 ; P3_U4397
g8195 nand P3_R1077_U109 P3_U3885 ; P3_U4398
g8196 nand P3_R1095_U102 P3_U3884 ; P3_U4399
g8197 nand P3_R1143_U109 P3_U3881 ; P3_U4400
g8198 nand P3_R1161_U109 P3_U3891 ; P3_U4401
g8199 nand P3_R1131_U102 P3_U3887 ; P3_U4402
g8200 nand P3_R1200_U102 P3_U3017 ; P3_U4403
g8201 not P3_U3332 ; P3_U4404
g8202 nand P3_R1179_U102 P3_U3026 ; P3_U4405
g8203 nand P3_U3025 P3_U3080 ; P3_U4406
g8204 nand P3_U3443 P3_U4064 ; P3_U4407
g8205 nand P3_U3651 P3_U4404 ; P3_U4408
g8206 nand P3_U3020 P3_REG2_REG_20__SCAN_IN ; P3_U4409
g8207 nand P3_U3021 P3_REG1_REG_20__SCAN_IN ; P3_U4410
g8208 nand P3_U3022 P3_REG0_REG_20__SCAN_IN ; P3_U4411
g8209 nand P3_SUB_609_U20 P3_U3019 ; P3_U4412
g8210 not P3_U3075 ; P3_U4413
g8211 nand P3_U3033 P3_U3081 ; P3_U4414
g8212 nand P3_R1110_U108 P3_U3883 ; P3_U4415
g8213 nand P3_R1077_U108 P3_U3885 ; P3_U4416
g8214 nand P3_R1095_U101 P3_U3884 ; P3_U4417
g8215 nand P3_R1143_U108 P3_U3881 ; P3_U4418
g8216 nand P3_R1161_U108 P3_U3891 ; P3_U4419
g8217 nand P3_R1131_U101 P3_U3887 ; P3_U4420
g8218 nand P3_R1200_U101 P3_U3017 ; P3_U4421
g8219 not P3_U3333 ; P3_U4422
g8220 nand P3_R1179_U101 P3_U3026 ; P3_U4423
g8221 nand P3_U3025 P3_U3075 ; P3_U4424
g8222 nand P3_U3445 P3_U4064 ; P3_U4425
g8223 nand P3_U3654 P3_U4422 ; P3_U4426
g8224 nand P3_U3020 P3_REG2_REG_21__SCAN_IN ; P3_U4427
g8225 nand P3_U3021 P3_REG1_REG_21__SCAN_IN ; P3_U4428
g8226 nand P3_U3022 P3_REG0_REG_21__SCAN_IN ; P3_U4429
g8227 nand P3_SUB_609_U27 P3_U3019 ; P3_U4430
g8228 not P3_U3074 ; P3_U4431
g8229 nand P3_U3033 P3_U3080 ; P3_U4432
g8230 nand P3_R1110_U13 P3_U3883 ; P3_U4433
g8231 nand P3_R1077_U13 P3_U3885 ; P3_U4434
g8232 nand P3_R1095_U99 P3_U3884 ; P3_U4435
g8233 nand P3_R1143_U13 P3_U3881 ; P3_U4436
g8234 nand P3_R1161_U13 P3_U3891 ; P3_U4437
g8235 nand P3_R1131_U99 P3_U3887 ; P3_U4438
g8236 nand P3_R1200_U99 P3_U3017 ; P3_U4439
g8237 not P3_U3335 ; P3_U4440
g8238 nand P3_R1179_U99 P3_U3026 ; P3_U4441
g8239 nand P3_U3025 P3_U3074 ; P3_U4442
g8240 nand P3_U3907 P3_U4064 ; P3_U4443
g8241 nand P3_U3657 P3_U4440 ; P3_U4444
g8242 nand P3_U3020 P3_REG2_REG_22__SCAN_IN ; P3_U4445
g8243 nand P3_U3021 P3_REG1_REG_22__SCAN_IN ; P3_U4446
g8244 nand P3_U3022 P3_REG0_REG_22__SCAN_IN ; P3_U4447
g8245 nand P3_SUB_609_U17 P3_U3019 ; P3_U4448
g8246 not P3_U3060 ; P3_U4449
g8247 nand P3_U3033 P3_U3075 ; P3_U4450
g8248 nand P3_R1110_U14 P3_U3883 ; P3_U4451
g8249 nand P3_R1077_U14 P3_U3885 ; P3_U4452
g8250 nand P3_R1095_U113 P3_U3884 ; P3_U4453
g8251 nand P3_R1143_U14 P3_U3881 ; P3_U4454
g8252 nand P3_R1161_U14 P3_U3891 ; P3_U4455
g8253 nand P3_R1131_U113 P3_U3887 ; P3_U4456
g8254 nand P3_R1200_U113 P3_U3017 ; P3_U4457
g8255 not P3_U3337 ; P3_U4458
g8256 nand P3_R1179_U113 P3_U3026 ; P3_U4459
g8257 nand P3_U3025 P3_U3060 ; P3_U4460
g8258 nand P3_U3906 P3_U4064 ; P3_U4461
g8259 nand P3_U3660 P3_U4458 ; P3_U4462
g8260 nand P3_U3020 P3_REG2_REG_23__SCAN_IN ; P3_U4463
g8261 nand P3_U3021 P3_REG1_REG_23__SCAN_IN ; P3_U4464
g8262 nand P3_U3022 P3_REG0_REG_23__SCAN_IN ; P3_U4465
g8263 nand P3_SUB_609_U6 P3_U3019 ; P3_U4466
g8264 not P3_U3065 ; P3_U4467
g8265 nand P3_U3033 P3_U3074 ; P3_U4468
g8266 nand P3_R1110_U107 P3_U3883 ; P3_U4469
g8267 nand P3_R1077_U107 P3_U3885 ; P3_U4470
g8268 nand P3_R1095_U112 P3_U3884 ; P3_U4471
g8269 nand P3_R1143_U107 P3_U3881 ; P3_U4472
g8270 nand P3_R1161_U107 P3_U3891 ; P3_U4473
g8271 nand P3_R1131_U112 P3_U3887 ; P3_U4474
g8272 nand P3_R1200_U112 P3_U3017 ; P3_U4475
g8273 not P3_U3339 ; P3_U4476
g8274 nand P3_R1179_U112 P3_U3026 ; P3_U4477
g8275 nand P3_U3025 P3_U3065 ; P3_U4478
g8276 nand P3_U3905 P3_U4064 ; P3_U4479
g8277 nand P3_U3663 P3_U4476 ; P3_U4480
g8278 nand P3_U3020 P3_REG2_REG_24__SCAN_IN ; P3_U4481
g8279 nand P3_U3021 P3_REG1_REG_24__SCAN_IN ; P3_U4482
g8280 nand P3_U3022 P3_REG0_REG_24__SCAN_IN ; P3_U4483
g8281 nand P3_SUB_609_U10 P3_U3019 ; P3_U4484
g8282 not P3_U3064 ; P3_U4485
g8283 nand P3_U3033 P3_U3060 ; P3_U4486
g8284 nand P3_R1110_U106 P3_U3883 ; P3_U4487
g8285 nand P3_R1077_U106 P3_U3885 ; P3_U4488
g8286 nand P3_R1095_U18 P3_U3884 ; P3_U4489
g8287 nand P3_R1143_U106 P3_U3881 ; P3_U4490
g8288 nand P3_R1161_U106 P3_U3891 ; P3_U4491
g8289 nand P3_R1131_U18 P3_U3887 ; P3_U4492
g8290 nand P3_R1200_U18 P3_U3017 ; P3_U4493
g8291 not P3_U3341 ; P3_U4494
g8292 nand P3_R1179_U18 P3_U3026 ; P3_U4495
g8293 nand P3_U3025 P3_U3064 ; P3_U4496
g8294 nand P3_U3904 P3_U4064 ; P3_U4497
g8295 nand P3_U3666 P3_U4494 ; P3_U4498
g8296 nand P3_U3020 P3_REG2_REG_25__SCAN_IN ; P3_U4499
g8297 nand P3_U3021 P3_REG1_REG_25__SCAN_IN ; P3_U4500
g8298 nand P3_U3022 P3_REG0_REG_25__SCAN_IN ; P3_U4501
g8299 nand P3_SUB_609_U16 P3_U3019 ; P3_U4502
g8300 not P3_U3057 ; P3_U4503
g8301 nand P3_U3033 P3_U3065 ; P3_U4504
g8302 nand P3_R1110_U105 P3_U3883 ; P3_U4505
g8303 nand P3_R1077_U105 P3_U3885 ; P3_U4506
g8304 nand P3_R1095_U98 P3_U3884 ; P3_U4507
g8305 nand P3_R1143_U105 P3_U3881 ; P3_U4508
g8306 nand P3_R1161_U105 P3_U3891 ; P3_U4509
g8307 nand P3_R1131_U98 P3_U3887 ; P3_U4510
g8308 nand P3_R1200_U98 P3_U3017 ; P3_U4511
g8309 not P3_U3343 ; P3_U4512
g8310 nand P3_R1179_U98 P3_U3026 ; P3_U4513
g8311 nand P3_U3025 P3_U3057 ; P3_U4514
g8312 nand P3_U3903 P3_U4064 ; P3_U4515
g8313 nand P3_U3670 P3_U4512 ; P3_U4516
g8314 nand P3_U3020 P3_REG2_REG_26__SCAN_IN ; P3_U4517
g8315 nand P3_U3021 P3_REG1_REG_26__SCAN_IN ; P3_U4518
g8316 nand P3_U3022 P3_REG0_REG_26__SCAN_IN ; P3_U4519
g8317 nand P3_SUB_609_U26 P3_U3019 ; P3_U4520
g8318 not P3_U3056 ; P3_U4521
g8319 nand P3_U3033 P3_U3064 ; P3_U4522
g8320 nand P3_R1110_U104 P3_U3883 ; P3_U4523
g8321 nand P3_R1077_U104 P3_U3885 ; P3_U4524
g8322 nand P3_R1095_U97 P3_U3884 ; P3_U4525
g8323 nand P3_R1143_U104 P3_U3881 ; P3_U4526
g8324 nand P3_R1161_U104 P3_U3891 ; P3_U4527
g8325 nand P3_R1131_U97 P3_U3887 ; P3_U4528
g8326 nand P3_R1200_U97 P3_U3017 ; P3_U4529
g8327 not P3_U3345 ; P3_U4530
g8328 nand P3_R1179_U97 P3_U3026 ; P3_U4531
g8329 nand P3_U3025 P3_U3056 ; P3_U4532
g8330 nand P3_U3902 P3_U4064 ; P3_U4533
g8331 nand P3_U3674 P3_U4530 ; P3_U4534
g8332 nand P3_U3020 P3_REG2_REG_27__SCAN_IN ; P3_U4535
g8333 nand P3_U3021 P3_REG1_REG_27__SCAN_IN ; P3_U4536
g8334 nand P3_U3022 P3_REG0_REG_27__SCAN_IN ; P3_U4537
g8335 nand P3_SUB_609_U22 P3_U3019 ; P3_U4538
g8336 not P3_U3052 ; P3_U4539
g8337 nand P3_U3033 P3_U3057 ; P3_U4540
g8338 nand P3_R1110_U15 P3_U3883 ; P3_U4541
g8339 nand P3_R1077_U15 P3_U3885 ; P3_U4542
g8340 nand P3_R1095_U111 P3_U3884 ; P3_U4543
g8341 nand P3_R1143_U15 P3_U3881 ; P3_U4544
g8342 nand P3_R1161_U15 P3_U3891 ; P3_U4545
g8343 nand P3_R1131_U111 P3_U3887 ; P3_U4546
g8344 nand P3_R1200_U111 P3_U3017 ; P3_U4547
g8345 not P3_U3347 ; P3_U4548
g8346 nand P3_R1179_U111 P3_U3026 ; P3_U4549
g8347 nand P3_U3025 P3_U3052 ; P3_U4550
g8348 nand P3_U3901 P3_U4064 ; P3_U4551
g8349 nand P3_U3678 P3_U4548 ; P3_U4552
g8350 nand P3_U3020 P3_REG2_REG_28__SCAN_IN ; P3_U4553
g8351 nand P3_U3021 P3_REG1_REG_28__SCAN_IN ; P3_U4554
g8352 nand P3_U3022 P3_REG0_REG_28__SCAN_IN ; P3_U4555
g8353 nand P3_SUB_609_U28 P3_U3019 ; P3_U4556
g8354 not P3_U3053 ; P3_U4557
g8355 nand P3_U3033 P3_U3056 ; P3_U4558
g8356 nand P3_R1110_U103 P3_U3883 ; P3_U4559
g8357 nand P3_R1077_U103 P3_U3885 ; P3_U4560
g8358 nand P3_R1095_U19 P3_U3884 ; P3_U4561
g8359 nand P3_R1143_U103 P3_U3881 ; P3_U4562
g8360 nand P3_R1161_U103 P3_U3891 ; P3_U4563
g8361 nand P3_R1131_U19 P3_U3887 ; P3_U4564
g8362 nand P3_R1200_U19 P3_U3017 ; P3_U4565
g8363 not P3_U3349 ; P3_U4566
g8364 nand P3_R1179_U19 P3_U3026 ; P3_U4567
g8365 nand P3_U3025 P3_U3053 ; P3_U4568
g8366 nand P3_U3900 P3_U4064 ; P3_U4569
g8367 nand P3_U3682 P3_U4566 ; P3_U4570
g8368 nand P3_SUB_609_U92 P3_U3019 ; P3_U4571
g8369 nand P3_U3020 P3_REG2_REG_29__SCAN_IN ; P3_U4572
g8370 nand P3_U3021 P3_REG1_REG_29__SCAN_IN ; P3_U4573
g8371 nand P3_U3022 P3_REG0_REG_29__SCAN_IN ; P3_U4574
g8372 not P3_U3054 ; P3_U4575
g8373 nand P3_U3033 P3_U3052 ; P3_U4576
g8374 nand P3_R1110_U102 P3_U3883 ; P3_U4577
g8375 nand P3_R1077_U102 P3_U3885 ; P3_U4578
g8376 nand P3_R1095_U96 P3_U3884 ; P3_U4579
g8377 nand P3_R1143_U102 P3_U3881 ; P3_U4580
g8378 nand P3_R1161_U102 P3_U3891 ; P3_U4581
g8379 nand P3_R1131_U96 P3_U3887 ; P3_U4582
g8380 nand P3_R1200_U96 P3_U3017 ; P3_U4583
g8381 not P3_U3351 ; P3_U4584
g8382 nand P3_R1179_U96 P3_U3026 ; P3_U4585
g8383 nand P3_U3025 P3_U3054 ; P3_U4586
g8384 nand P3_U3899 P3_U4064 ; P3_U4587
g8385 nand P3_U3686 P3_U4584 ; P3_U4588
g8386 nand P3_U3020 P3_REG2_REG_30__SCAN_IN ; P3_U4589
g8387 nand P3_U3021 P3_REG1_REG_30__SCAN_IN ; P3_U4590
g8388 nand P3_U3022 P3_REG0_REG_30__SCAN_IN ; P3_U4591
g8389 nand P3_SUB_609_U92 P3_U3019 ; P3_U4592
g8390 not P3_U3058 ; P3_U4593
g8391 nand P3_U3892 P3_U3298 ; P3_U4594
g8392 nand P3_U3833 P3_U4594 ; P3_U4595
g8393 nand P3_U4595 P3_U3911 P3_U3058 ; P3_U4596
g8394 nand P3_U3033 P3_U3053 ; P3_U4597
g8395 nand P3_R1110_U101 P3_U3883 ; P3_U4598
g8396 nand P3_R1077_U101 P3_U3885 ; P3_U4599
g8397 nand P3_R1095_U20 P3_U3884 ; P3_U4600
g8398 nand P3_R1143_U101 P3_U3881 ; P3_U4601
g8399 nand P3_R1161_U101 P3_U3891 ; P3_U4602
g8400 nand P3_R1131_U20 P3_U3887 ; P3_U4603
g8401 nand P3_R1200_U20 P3_U3017 ; P3_U4604
g8402 not P3_U3354 ; P3_U4605
g8403 nand P3_R1179_U20 P3_U3026 ; P3_U4606
g8404 nand P3_U3908 P3_U4064 ; P3_U4607
g8405 nand P3_U3690 P3_U4605 ; P3_U4608
g8406 nand P3_SUB_609_U92 P3_U3019 ; P3_U4609
g8407 nand P3_U3020 P3_REG2_REG_31__SCAN_IN ; P3_U4610
g8408 nand P3_U3021 P3_REG1_REG_31__SCAN_IN ; P3_U4611
g8409 nand P3_U3022 P3_REG0_REG_31__SCAN_IN ; P3_U4612
g8410 not P3_U3055 ; P3_U4613
g8411 nand P3_U3873 P3_U4064 ; P3_U4614
g8412 nand P3_U3361 P3_U4614 ; P3_U4615
g8413 nand P3_U3872 P3_U4064 ; P3_U4616
g8414 nand P3_U3361 P3_U4616 ; P3_U4617
g8415 nand P3_U5641 P3_U5640 P3_U3302 ; P3_U4618
g8416 nand P3_U3888 P3_U3367 ; P3_U4619
g8417 nand P3_U3048 P3_U4619 ; P3_U4620
g8418 nand P3_U3047 P3_U4618 ; P3_U4621
g8419 nand P3_U4621 P3_U4620 ; P3_U4622
g8420 nand P3_U5456 P3_U3379 ; P3_U4623
g8421 nand P3_U4623 P3_U3380 P3_U3834 ; P3_U4624
g8422 nand P3_U3048 P3_U4624 ; P3_U4625
g8423 nand P3_U3047 P3_U4619 ; P3_U4626
g8424 nand P3_U4625 P3_U3360 P3_U4626 ; P3_U4627
g8425 not P3_U3365 ; P3_U4628
g8426 nand P3_U3034 P3_U3077 ; P3_U4629
g8427 nand P3_U3030 P3_R1179_U24 ; P3_U4630
g8428 nand P3_U3029 P3_U3387 ; P3_U4631
g8429 nand P3_U3028 P3_REG3_REG_0__SCAN_IN ; P3_U4632
g8430 nand P3_U3034 P3_U3067 ; P3_U4633
g8431 nand P3_U3030 P3_R1179_U100 ; P3_U4634
g8432 nand P3_U3029 P3_U3392 ; P3_U4635
g8433 nand P3_U3028 P3_REG3_REG_1__SCAN_IN ; P3_U4636
g8434 nand P3_U3034 P3_U3063 ; P3_U4637
g8435 nand P3_U3030 P3_R1179_U110 ; P3_U4638
g8436 nand P3_U3029 P3_U3395 ; P3_U4639
g8437 nand P3_U3028 P3_REG3_REG_2__SCAN_IN ; P3_U4640
g8438 nand P3_U3034 P3_U3059 ; P3_U4641
g8439 nand P3_U3030 P3_R1179_U21 ; P3_U4642
g8440 nand P3_U3029 P3_U3398 ; P3_U4643
g8441 nand P3_U3028 P3_SUB_609_U25 ; P3_U4644
g8442 nand P3_U3034 P3_U3066 ; P3_U4645
g8443 nand P3_U3030 P3_R1179_U109 ; P3_U4646
g8444 nand P3_U3029 P3_U3401 ; P3_U4647
g8445 nand P3_U3028 P3_SUB_609_U29 ; P3_U4648
g8446 nand P3_U3034 P3_U3070 ; P3_U4649
g8447 nand P3_U3030 P3_R1179_U108 ; P3_U4650
g8448 nand P3_U3029 P3_U3404 ; P3_U4651
g8449 nand P3_U3028 P3_SUB_609_U53 ; P3_U4652
g8450 nand P3_U3034 P3_U3069 ; P3_U4653
g8451 nand P3_U3030 P3_R1179_U22 ; P3_U4654
g8452 nand P3_U3029 P3_U3407 ; P3_U4655
g8453 nand P3_U3028 P3_SUB_609_U8 ; P3_U4656
g8454 nand P3_U3034 P3_U3083 ; P3_U4657
g8455 nand P3_U3030 P3_R1179_U107 ; P3_U4658
g8456 nand P3_U3029 P3_U3410 ; P3_U4659
g8457 nand P3_U3028 P3_SUB_609_U18 ; P3_U4660
g8458 nand P3_U3034 P3_U3082 ; P3_U4661
g8459 nand P3_U3030 P3_R1179_U23 ; P3_U4662
g8460 nand P3_U3029 P3_U3413 ; P3_U4663
g8461 nand P3_U3028 P3_SUB_609_U12 ; P3_U4664
g8462 nand P3_U3034 P3_U3061 ; P3_U4665
g8463 nand P3_U3030 P3_R1179_U106 ; P3_U4666
g8464 nand P3_U3029 P3_U3416 ; P3_U4667
g8465 nand P3_U3028 P3_SUB_609_U14 ; P3_U4668
g8466 nand P3_U3034 P3_U3062 ; P3_U4669
g8467 nand P3_U3030 P3_R1179_U116 ; P3_U4670
g8468 nand P3_U3029 P3_U3419 ; P3_U4671
g8469 nand P3_U3028 P3_SUB_609_U13 ; P3_U4672
g8470 nand P3_U3034 P3_U3071 ; P3_U4673
g8471 nand P3_U3030 P3_R1179_U16 ; P3_U4674
g8472 nand P3_U3029 P3_U3422 ; P3_U4675
g8473 nand P3_U3028 P3_SUB_609_U9 ; P3_U4676
g8474 nand P3_U3034 P3_U3079 ; P3_U4677
g8475 nand P3_U3030 P3_R1179_U105 ; P3_U4678
g8476 nand P3_U3029 P3_U3425 ; P3_U4679
g8477 nand P3_U3028 P3_SUB_609_U23 ; P3_U4680
g8478 nand P3_U3034 P3_U3078 ; P3_U4681
g8479 nand P3_U3030 P3_R1179_U104 ; P3_U4682
g8480 nand P3_U3029 P3_U3428 ; P3_U4683
g8481 nand P3_U3028 P3_SUB_609_U24 ; P3_U4684
g8482 nand P3_U3034 P3_U3073 ; P3_U4685
g8483 nand P3_U3030 P3_R1179_U115 ; P3_U4686
g8484 nand P3_U3029 P3_U3431 ; P3_U4687
g8485 nand P3_U3028 P3_SUB_609_U30 ; P3_U4688
g8486 nand P3_U3034 P3_U3072 ; P3_U4689
g8487 nand P3_U3030 P3_R1179_U114 ; P3_U4690
g8488 nand P3_U3029 P3_U3434 ; P3_U4691
g8489 nand P3_U3028 P3_SUB_609_U21 ; P3_U4692
g8490 nand P3_U3034 P3_U3068 ; P3_U4693
g8491 nand P3_U3030 P3_R1179_U17 ; P3_U4694
g8492 nand P3_U3029 P3_U3437 ; P3_U4695
g8493 nand P3_U3028 P3_SUB_609_U7 ; P3_U4696
g8494 nand P3_U3034 P3_U3081 ; P3_U4697
g8495 nand P3_U3030 P3_R1179_U103 ; P3_U4698
g8496 nand P3_U3029 P3_U3440 ; P3_U4699
g8497 nand P3_U3028 P3_SUB_609_U19 ; P3_U4700
g8498 nand P3_U3034 P3_U3080 ; P3_U4701
g8499 nand P3_U3030 P3_R1179_U102 ; P3_U4702
g8500 nand P3_U3029 P3_U3443 ; P3_U4703
g8501 nand P3_U3028 P3_SUB_609_U11 ; P3_U4704
g8502 nand P3_U3034 P3_U3075 ; P3_U4705
g8503 nand P3_U3030 P3_R1179_U101 ; P3_U4706
g8504 nand P3_U3029 P3_U3445 ; P3_U4707
g8505 nand P3_U3028 P3_SUB_609_U15 ; P3_U4708
g8506 nand P3_U3034 P3_U3074 ; P3_U4709
g8507 nand P3_U3030 P3_R1179_U99 ; P3_U4710
g8508 nand P3_U3029 P3_U3907 ; P3_U4711
g8509 nand P3_U3028 P3_SUB_609_U20 ; P3_U4712
g8510 nand P3_U3034 P3_U3060 ; P3_U4713
g8511 nand P3_U3030 P3_R1179_U113 ; P3_U4714
g8512 nand P3_U3029 P3_U3906 ; P3_U4715
g8513 nand P3_U3028 P3_SUB_609_U27 ; P3_U4716
g8514 nand P3_U3034 P3_U3065 ; P3_U4717
g8515 nand P3_U3030 P3_R1179_U112 ; P3_U4718
g8516 nand P3_U3029 P3_U3905 ; P3_U4719
g8517 nand P3_U3028 P3_SUB_609_U17 ; P3_U4720
g8518 nand P3_U3034 P3_U3064 ; P3_U4721
g8519 nand P3_U3030 P3_R1179_U18 ; P3_U4722
g8520 nand P3_U3029 P3_U3904 ; P3_U4723
g8521 nand P3_U3028 P3_SUB_609_U6 ; P3_U4724
g8522 nand P3_U3034 P3_U3057 ; P3_U4725
g8523 nand P3_U3030 P3_R1179_U98 ; P3_U4726
g8524 nand P3_U3029 P3_U3903 ; P3_U4727
g8525 nand P3_U3028 P3_SUB_609_U10 ; P3_U4728
g8526 nand P3_U3034 P3_U3056 ; P3_U4729
g8527 nand P3_U3030 P3_R1179_U97 ; P3_U4730
g8528 nand P3_U3029 P3_U3902 ; P3_U4731
g8529 nand P3_U3028 P3_SUB_609_U16 ; P3_U4732
g8530 nand P3_U3034 P3_U3052 ; P3_U4733
g8531 nand P3_U3030 P3_R1179_U111 ; P3_U4734
g8532 nand P3_U3029 P3_U3901 ; P3_U4735
g8533 nand P3_U3028 P3_SUB_609_U26 ; P3_U4736
g8534 nand P3_U3034 P3_U3053 ; P3_U4737
g8535 nand P3_U3030 P3_R1179_U19 ; P3_U4738
g8536 nand P3_U3029 P3_U3900 ; P3_U4739
g8537 nand P3_U3028 P3_SUB_609_U22 ; P3_U4740
g8538 nand P3_U3034 P3_U3054 ; P3_U4741
g8539 nand P3_U3030 P3_R1179_U96 ; P3_U4742
g8540 nand P3_U3029 P3_U3899 ; P3_U4743
g8541 nand P3_U3028 P3_SUB_609_U28 ; P3_U4744
g8542 nand P3_U3030 P3_R1179_U20 ; P3_U4745
g8543 nand P3_U3029 P3_U3908 ; P3_U4746
g8544 nand P3_U3028 P3_SUB_609_U92 ; P3_U4747
g8545 nand P3_U3028 P3_SUB_609_U92 ; P3_U4748
g8546 nand P3_U3916 P3_U3912 ; P3_U4749
g8547 nand P3_U3029 P3_U3873 ; P3_U4750
g8548 nand P3_U3358 P3_REG2_REG_30__SCAN_IN ; P3_U4751
g8549 nand P3_U3029 P3_U3872 ; P3_U4752
g8550 nand P3_U3358 P3_REG2_REG_31__SCAN_IN ; P3_U4753
g8551 nand P3_U4628 P3_U3359 P3_U3698 P3_U3697 ; P3_U4754
g8552 nand P3_R1212_U6 P3_U3040 ; P3_U4755
g8553 nand P3_U3039 P3_U3379 ; P3_U4756
g8554 nand P3_R1209_U6 P3_U3037 ; P3_U4757
g8555 nand P3_U4756 P3_U4755 P3_U4757 ; P3_U4758
g8556 nand P3_U3910 P3_U5440 ; P3_U4759
g8557 not P3_U3366 ; P3_U4760
g8558 nand P3_U3833 P3_U3896 ; P3_U4761
g8559 nand P3_R1054_U67 P3_U3051 ; P3_U4762
g8560 nand P3_U5768 P3_U3379 ; P3_U4763
g8561 nand P3_U3042 P3_U4758 ; P3_U4764
g8562 nand P3_U3041 P3_R1212_U6 ; P3_U4765
g8563 nand P3_U3151 P3_REG3_REG_19__SCAN_IN ; P3_U4766
g8564 nand P3_U3038 P3_R1209_U6 ; P3_U4767
g8565 nand P3_U4760 P3_ADDR_REG_19__SCAN_IN ; P3_U4768
g8566 nand P3_R1212_U58 P3_U3040 ; P3_U4769
g8567 nand P3_U3039 P3_U3442 ; P3_U4770
g8568 nand P3_R1209_U58 P3_U3037 ; P3_U4771
g8569 nand P3_U4770 P3_U4769 P3_U4771 ; P3_U4772
g8570 nand P3_R1054_U68 P3_U3051 ; P3_U4773
g8571 nand P3_U5768 P3_U3442 ; P3_U4774
g8572 nand P3_U3042 P3_U4772 ; P3_U4775
g8573 nand P3_R1212_U58 P3_U3041 ; P3_U4776
g8574 nand P3_U3151 P3_REG3_REG_18__SCAN_IN ; P3_U4777
g8575 nand P3_R1209_U58 P3_U3038 ; P3_U4778
g8576 nand P3_U4760 P3_ADDR_REG_18__SCAN_IN ; P3_U4779
g8577 nand P3_R1212_U59 P3_U3040 ; P3_U4780
g8578 nand P3_U3039 P3_U3439 ; P3_U4781
g8579 nand P3_R1209_U59 P3_U3037 ; P3_U4782
g8580 nand P3_U4781 P3_U4780 P3_U4782 ; P3_U4783
g8581 nand P3_R1054_U69 P3_U3051 ; P3_U4784
g8582 nand P3_U5768 P3_U3439 ; P3_U4785
g8583 nand P3_U3042 P3_U4783 ; P3_U4786
g8584 nand P3_R1212_U59 P3_U3041 ; P3_U4787
g8585 nand P3_U3151 P3_REG3_REG_17__SCAN_IN ; P3_U4788
g8586 nand P3_R1209_U59 P3_U3038 ; P3_U4789
g8587 nand P3_U4760 P3_ADDR_REG_17__SCAN_IN ; P3_U4790
g8588 nand P3_R1212_U60 P3_U3040 ; P3_U4791
g8589 nand P3_U3039 P3_U3436 ; P3_U4792
g8590 nand P3_R1209_U60 P3_U3037 ; P3_U4793
g8591 nand P3_U4792 P3_U4791 P3_U4793 ; P3_U4794
g8592 nand P3_R1054_U13 P3_U3051 ; P3_U4795
g8593 nand P3_U5768 P3_U3436 ; P3_U4796
g8594 nand P3_U3042 P3_U4794 ; P3_U4797
g8595 nand P3_R1212_U60 P3_U3041 ; P3_U4798
g8596 nand P3_U3151 P3_REG3_REG_16__SCAN_IN ; P3_U4799
g8597 nand P3_R1209_U60 P3_U3038 ; P3_U4800
g8598 nand P3_U4760 P3_ADDR_REG_16__SCAN_IN ; P3_U4801
g8599 nand P3_R1212_U61 P3_U3040 ; P3_U4802
g8600 nand P3_U3039 P3_U3433 ; P3_U4803
g8601 nand P3_R1209_U61 P3_U3037 ; P3_U4804
g8602 nand P3_U4803 P3_U4802 P3_U4804 ; P3_U4805
g8603 nand P3_R1054_U77 P3_U3051 ; P3_U4806
g8604 nand P3_U5768 P3_U3433 ; P3_U4807
g8605 nand P3_U3042 P3_U4805 ; P3_U4808
g8606 nand P3_R1212_U61 P3_U3041 ; P3_U4809
g8607 nand P3_U3151 P3_REG3_REG_15__SCAN_IN ; P3_U4810
g8608 nand P3_R1209_U61 P3_U3038 ; P3_U4811
g8609 nand P3_U4760 P3_ADDR_REG_15__SCAN_IN ; P3_U4812
g8610 nand P3_R1212_U62 P3_U3040 ; P3_U4813
g8611 nand P3_U3039 P3_U3430 ; P3_U4814
g8612 nand P3_R1209_U62 P3_U3037 ; P3_U4815
g8613 nand P3_U4814 P3_U4813 P3_U4815 ; P3_U4816
g8614 nand P3_R1054_U78 P3_U3051 ; P3_U4817
g8615 nand P3_U5768 P3_U3430 ; P3_U4818
g8616 nand P3_U3042 P3_U4816 ; P3_U4819
g8617 nand P3_R1212_U62 P3_U3041 ; P3_U4820
g8618 nand P3_U3151 P3_REG3_REG_14__SCAN_IN ; P3_U4821
g8619 nand P3_R1209_U62 P3_U3038 ; P3_U4822
g8620 nand P3_U4760 P3_ADDR_REG_14__SCAN_IN ; P3_U4823
g8621 nand P3_R1212_U63 P3_U3040 ; P3_U4824
g8622 nand P3_U3039 P3_U3427 ; P3_U4825
g8623 nand P3_R1209_U63 P3_U3037 ; P3_U4826
g8624 nand P3_U4825 P3_U4824 P3_U4826 ; P3_U4827
g8625 nand P3_R1054_U70 P3_U3051 ; P3_U4828
g8626 nand P3_U5768 P3_U3427 ; P3_U4829
g8627 nand P3_U3042 P3_U4827 ; P3_U4830
g8628 nand P3_R1212_U63 P3_U3041 ; P3_U4831
g8629 nand P3_U3151 P3_REG3_REG_13__SCAN_IN ; P3_U4832
g8630 nand P3_R1209_U63 P3_U3038 ; P3_U4833
g8631 nand P3_U4760 P3_ADDR_REG_13__SCAN_IN ; P3_U4834
g8632 nand P3_R1212_U64 P3_U3040 ; P3_U4835
g8633 nand P3_U3039 P3_U3424 ; P3_U4836
g8634 nand P3_R1209_U64 P3_U3037 ; P3_U4837
g8635 nand P3_U4836 P3_U4835 P3_U4837 ; P3_U4838
g8636 nand P3_R1054_U71 P3_U3051 ; P3_U4839
g8637 nand P3_U5768 P3_U3424 ; P3_U4840
g8638 nand P3_U3042 P3_U4838 ; P3_U4841
g8639 nand P3_R1212_U64 P3_U3041 ; P3_U4842
g8640 nand P3_U3151 P3_REG3_REG_12__SCAN_IN ; P3_U4843
g8641 nand P3_R1209_U64 P3_U3038 ; P3_U4844
g8642 nand P3_U4760 P3_ADDR_REG_12__SCAN_IN ; P3_U4845
g8643 nand P3_R1212_U65 P3_U3040 ; P3_U4846
g8644 nand P3_U3039 P3_U3421 ; P3_U4847
g8645 nand P3_R1209_U65 P3_U3037 ; P3_U4848
g8646 nand P3_U4847 P3_U4846 P3_U4848 ; P3_U4849
g8647 nand P3_R1054_U12 P3_U3051 ; P3_U4850
g8648 nand P3_U5768 P3_U3421 ; P3_U4851
g8649 nand P3_U3042 P3_U4849 ; P3_U4852
g8650 nand P3_R1212_U65 P3_U3041 ; P3_U4853
g8651 nand P3_U3151 P3_REG3_REG_11__SCAN_IN ; P3_U4854
g8652 nand P3_R1209_U65 P3_U3038 ; P3_U4855
g8653 nand P3_U4760 P3_ADDR_REG_11__SCAN_IN ; P3_U4856
g8654 nand P3_R1212_U66 P3_U3040 ; P3_U4857
g8655 nand P3_U3039 P3_U3418 ; P3_U4858
g8656 nand P3_R1209_U66 P3_U3037 ; P3_U4859
g8657 nand P3_U4858 P3_U4857 P3_U4859 ; P3_U4860
g8658 nand P3_R1054_U79 P3_U3051 ; P3_U4861
g8659 nand P3_U5768 P3_U3418 ; P3_U4862
g8660 nand P3_U3042 P3_U4860 ; P3_U4863
g8661 nand P3_R1212_U66 P3_U3041 ; P3_U4864
g8662 nand P3_U3151 P3_REG3_REG_10__SCAN_IN ; P3_U4865
g8663 nand P3_R1209_U66 P3_U3038 ; P3_U4866
g8664 nand P3_U4760 P3_ADDR_REG_10__SCAN_IN ; P3_U4867
g8665 nand P3_R1212_U49 P3_U3040 ; P3_U4868
g8666 nand P3_U3039 P3_U3415 ; P3_U4869
g8667 nand P3_R1209_U49 P3_U3037 ; P3_U4870
g8668 nand P3_U4869 P3_U4868 P3_U4870 ; P3_U4871
g8669 nand P3_R1054_U72 P3_U3051 ; P3_U4872
g8670 nand P3_U5768 P3_U3415 ; P3_U4873
g8671 nand P3_U3042 P3_U4871 ; P3_U4874
g8672 nand P3_R1212_U49 P3_U3041 ; P3_U4875
g8673 nand P3_U3151 P3_REG3_REG_9__SCAN_IN ; P3_U4876
g8674 nand P3_R1209_U49 P3_U3038 ; P3_U4877
g8675 nand P3_U4760 P3_ADDR_REG_9__SCAN_IN ; P3_U4878
g8676 nand P3_R1212_U50 P3_U3040 ; P3_U4879
g8677 nand P3_U3039 P3_U3412 ; P3_U4880
g8678 nand P3_R1209_U50 P3_U3037 ; P3_U4881
g8679 nand P3_U4880 P3_U4879 P3_U4881 ; P3_U4882
g8680 nand P3_R1054_U16 P3_U3051 ; P3_U4883
g8681 nand P3_U5768 P3_U3412 ; P3_U4884
g8682 nand P3_U3042 P3_U4882 ; P3_U4885
g8683 nand P3_R1212_U50 P3_U3041 ; P3_U4886
g8684 nand P3_U3151 P3_REG3_REG_8__SCAN_IN ; P3_U4887
g8685 nand P3_R1209_U50 P3_U3038 ; P3_U4888
g8686 nand P3_U4760 P3_ADDR_REG_8__SCAN_IN ; P3_U4889
g8687 nand P3_R1212_U51 P3_U3040 ; P3_U4890
g8688 nand P3_U3039 P3_U3409 ; P3_U4891
g8689 nand P3_R1209_U51 P3_U3037 ; P3_U4892
g8690 nand P3_U4891 P3_U4890 P3_U4892 ; P3_U4893
g8691 nand P3_R1054_U73 P3_U3051 ; P3_U4894
g8692 nand P3_U5768 P3_U3409 ; P3_U4895
g8693 nand P3_U3042 P3_U4893 ; P3_U4896
g8694 nand P3_R1212_U51 P3_U3041 ; P3_U4897
g8695 nand P3_U3151 P3_REG3_REG_7__SCAN_IN ; P3_U4898
g8696 nand P3_R1209_U51 P3_U3038 ; P3_U4899
g8697 nand P3_U4760 P3_ADDR_REG_7__SCAN_IN ; P3_U4900
g8698 nand P3_R1212_U52 P3_U3040 ; P3_U4901
g8699 nand P3_U3039 P3_U3406 ; P3_U4902
g8700 nand P3_R1209_U52 P3_U3037 ; P3_U4903
g8701 nand P3_U4902 P3_U4901 P3_U4903 ; P3_U4904
g8702 nand P3_R1054_U15 P3_U3051 ; P3_U4905
g8703 nand P3_U5768 P3_U3406 ; P3_U4906
g8704 nand P3_U3042 P3_U4904 ; P3_U4907
g8705 nand P3_R1212_U52 P3_U3041 ; P3_U4908
g8706 nand P3_U3151 P3_REG3_REG_6__SCAN_IN ; P3_U4909
g8707 nand P3_R1209_U52 P3_U3038 ; P3_U4910
g8708 nand P3_U4760 P3_ADDR_REG_6__SCAN_IN ; P3_U4911
g8709 nand P3_R1212_U53 P3_U3040 ; P3_U4912
g8710 nand P3_U3039 P3_U3403 ; P3_U4913
g8711 nand P3_R1209_U53 P3_U3037 ; P3_U4914
g8712 nand P3_U4913 P3_U4912 P3_U4914 ; P3_U4915
g8713 nand P3_R1054_U74 P3_U3051 ; P3_U4916
g8714 nand P3_U5768 P3_U3403 ; P3_U4917
g8715 nand P3_U3042 P3_U4915 ; P3_U4918
g8716 nand P3_R1212_U53 P3_U3041 ; P3_U4919
g8717 nand P3_U3151 P3_REG3_REG_5__SCAN_IN ; P3_U4920
g8718 nand P3_R1209_U53 P3_U3038 ; P3_U4921
g8719 nand P3_U4760 P3_ADDR_REG_5__SCAN_IN ; P3_U4922
g8720 nand P3_R1212_U54 P3_U3040 ; P3_U4923
g8721 nand P3_U3039 P3_U3400 ; P3_U4924
g8722 nand P3_R1209_U54 P3_U3037 ; P3_U4925
g8723 nand P3_U4924 P3_U4923 P3_U4925 ; P3_U4926
g8724 nand P3_R1054_U75 P3_U3051 ; P3_U4927
g8725 nand P3_U5768 P3_U3400 ; P3_U4928
g8726 nand P3_U3042 P3_U4926 ; P3_U4929
g8727 nand P3_R1212_U54 P3_U3041 ; P3_U4930
g8728 nand P3_U3151 P3_REG3_REG_4__SCAN_IN ; P3_U4931
g8729 nand P3_R1209_U54 P3_U3038 ; P3_U4932
g8730 nand P3_U4760 P3_ADDR_REG_4__SCAN_IN ; P3_U4933
g8731 nand P3_R1212_U55 P3_U3040 ; P3_U4934
g8732 nand P3_U3039 P3_U3397 ; P3_U4935
g8733 nand P3_R1209_U55 P3_U3037 ; P3_U4936
g8734 nand P3_U4935 P3_U4934 P3_U4936 ; P3_U4937
g8735 nand P3_R1054_U14 P3_U3051 ; P3_U4938
g8736 nand P3_U5768 P3_U3397 ; P3_U4939
g8737 nand P3_U3042 P3_U4937 ; P3_U4940
g8738 nand P3_R1212_U55 P3_U3041 ; P3_U4941
g8739 nand P3_U3151 P3_REG3_REG_3__SCAN_IN ; P3_U4942
g8740 nand P3_R1209_U55 P3_U3038 ; P3_U4943
g8741 nand P3_U4760 P3_ADDR_REG_3__SCAN_IN ; P3_U4944
g8742 nand P3_R1212_U56 P3_U3040 ; P3_U4945
g8743 nand P3_U3039 P3_U3394 ; P3_U4946
g8744 nand P3_R1209_U56 P3_U3037 ; P3_U4947
g8745 nand P3_U4946 P3_U4945 P3_U4947 ; P3_U4948
g8746 nand P3_R1054_U76 P3_U3051 ; P3_U4949
g8747 nand P3_U5768 P3_U3394 ; P3_U4950
g8748 nand P3_U3042 P3_U4948 ; P3_U4951
g8749 nand P3_R1212_U56 P3_U3041 ; P3_U4952
g8750 nand P3_U3151 P3_REG3_REG_2__SCAN_IN ; P3_U4953
g8751 nand P3_R1209_U56 P3_U3038 ; P3_U4954
g8752 nand P3_U4760 P3_ADDR_REG_2__SCAN_IN ; P3_U4955
g8753 nand P3_R1212_U57 P3_U3040 ; P3_U4956
g8754 nand P3_U3039 P3_U3391 ; P3_U4957
g8755 nand P3_R1209_U57 P3_U3037 ; P3_U4958
g8756 nand P3_U4957 P3_U4956 P3_U4958 ; P3_U4959
g8757 nand P3_R1054_U66 P3_U3051 ; P3_U4960
g8758 nand P3_U5768 P3_U3391 ; P3_U4961
g8759 nand P3_U3042 P3_U4959 ; P3_U4962
g8760 nand P3_R1212_U57 P3_U3041 ; P3_U4963
g8761 nand P3_U3151 P3_REG3_REG_1__SCAN_IN ; P3_U4964
g8762 nand P3_R1209_U57 P3_U3038 ; P3_U4965
g8763 nand P3_U4760 P3_ADDR_REG_1__SCAN_IN ; P3_U4966
g8764 nand P3_R1212_U7 P3_U3040 ; P3_U4967
g8765 nand P3_U3039 P3_U3386 ; P3_U4968
g8766 nand P3_R1209_U7 P3_U3037 ; P3_U4969
g8767 nand P3_U4968 P3_U4967 P3_U4969 ; P3_U4970
g8768 nand P3_R1054_U17 P3_U3051 ; P3_U4971
g8769 nand P3_U5768 P3_U3386 ; P3_U4972
g8770 nand P3_U3042 P3_U4970 ; P3_U4973
g8771 nand P3_R1212_U7 P3_U3041 ; P3_U4974
g8772 nand P3_U3151 P3_REG3_REG_0__SCAN_IN ; P3_U4975
g8773 nand P3_R1209_U7 P3_U3038 ; P3_U4976
g8774 nand P3_U4760 P3_ADDR_REG_0__SCAN_IN ; P3_U4977
g8775 not P3_U3868 ; P3_U4978
g8776 nand P3_U5942 P3_U5941 P3_U3050 ; P3_U4979
g8777 nand P3_U3023 P3_U3909 P3_U3867 ; P3_U4980
g8778 nand P3_U4979 P3_B_REG_SCAN_IN ; P3_U4981
g8779 nand P3_U3036 P3_U3078 ; P3_U4982
g8780 nand P3_U3032 P3_U3072 ; P3_U4983
g8781 nand P3_SUB_609_U21 P3_U3304 ; P3_U4984
g8782 nand P3_U4983 P3_U4982 P3_U4984 ; P3_U4985
g8783 nand P3_U3311 P3_U3875 P3_U3888 P3_U5425 P3_U3312 ; P3_U4986
g8784 nand P3_U3894 P3_U4986 ; P3_U4987
g8785 nand P3_U3889 P3_U3895 ; P3_U4988
g8786 nand P3_U4988 P3_U4987 ; P3_U4989
g8787 nand P3_U3911 P3_U3378 ; P3_U4990
g8788 nand P3_U3889 P3_U3304 ; P3_U4991
g8789 nand P3_U4986 P3_U3303 ; P3_U4992
g8790 not P3_U3370 ; P3_U4993
g8791 nand P3_U3434 P3_U5420 ; P3_U4994
g8792 nand P3_SUB_609_U21 P3_U3371 ; P3_U4995
g8793 nand P3_R1158_U114 P3_U3035 ; P3_U4996
g8794 nand P3_U3031 P3_U4985 ; P3_U4997
g8795 nand P3_U3151 P3_REG3_REG_15__SCAN_IN ; P3_U4998
g8796 nand P3_U3036 P3_U3057 ; P3_U4999
g8797 nand P3_U3032 P3_U3052 ; P3_U5000
g8798 nand P3_SUB_609_U26 P3_U3304 ; P3_U5001
g8799 nand P3_U5000 P3_U4999 P3_U5001 ; P3_U5002
g8800 nand P3_U3365 P3_U3303 ; P3_U5003
g8801 nand P3_U4993 P3_U5003 ; P3_U5004
g8802 nand P3_U3894 P3_U3365 ; P3_U5005
g8803 nand P3_U3360 P3_U5005 ; P3_U5006
g8804 nand P3_U3045 P3_U3901 ; P3_U5007
g8805 nand P3_U3044 P3_SUB_609_U26 ; P3_U5008
g8806 nand P3_R1158_U16 P3_U3035 ; P3_U5009
g8807 nand P3_U3031 P3_U5002 ; P3_U5010
g8808 nand P3_U3151 P3_REG3_REG_26__SCAN_IN ; P3_U5011
g8809 nand P3_U3036 P3_U3066 ; P3_U5012
g8810 nand P3_U3032 P3_U3069 ; P3_U5013
g8811 nand P3_SUB_609_U8 P3_U3304 ; P3_U5014
g8812 nand P3_U5013 P3_U5012 P3_U5014 ; P3_U5015
g8813 nand P3_U3407 P3_U5420 ; P3_U5016
g8814 nand P3_SUB_609_U8 P3_U3371 ; P3_U5017
g8815 nand P3_R1158_U97 P3_U3035 ; P3_U5018
g8816 nand P3_U3031 P3_U5015 ; P3_U5019
g8817 nand P3_U3151 P3_REG3_REG_6__SCAN_IN ; P3_U5020
g8818 nand P3_U3036 P3_U3068 ; P3_U5021
g8819 nand P3_U3032 P3_U3080 ; P3_U5022
g8820 nand P3_SUB_609_U11 P3_U3304 ; P3_U5023
g8821 nand P3_U5022 P3_U5021 P3_U5023 ; P3_U5024
g8822 nand P3_U3443 P3_U5420 ; P3_U5025
g8823 nand P3_SUB_609_U11 P3_U3371 ; P3_U5026
g8824 nand P3_R1158_U112 P3_U3035 ; P3_U5027
g8825 nand P3_U3031 P3_U5024 ; P3_U5028
g8826 nand P3_U3151 P3_REG3_REG_18__SCAN_IN ; P3_U5029
g8827 nand P3_U3036 P3_U3077 ; P3_U5030
g8828 nand P3_U3032 P3_U3063 ; P3_U5031
g8829 nand P3_U3304 P3_REG3_REG_2__SCAN_IN ; P3_U5032
g8830 nand P3_U5031 P3_U5030 P3_U5032 ; P3_U5033
g8831 nand P3_U3395 P3_U5420 ; P3_U5034
g8832 nand P3_U3371 P3_REG3_REG_2__SCAN_IN ; P3_U5035
g8833 nand P3_R1158_U100 P3_U3035 ; P3_U5036
g8834 nand P3_U3031 P3_U5033 ; P3_U5037
g8835 nand P3_U3151 P3_REG3_REG_2__SCAN_IN ; P3_U5038
g8836 nand P3_U3036 P3_U3061 ; P3_U5039
g8837 nand P3_U3032 P3_U3071 ; P3_U5040
g8838 nand P3_SUB_609_U9 P3_U3304 ; P3_U5041
g8839 nand P3_U5040 P3_U5039 P3_U5041 ; P3_U5042
g8840 nand P3_U3422 P3_U5420 ; P3_U5043
g8841 nand P3_SUB_609_U9 P3_U3371 ; P3_U5044
g8842 nand P3_R1158_U117 P3_U3035 ; P3_U5045
g8843 nand P3_U3031 P3_U5042 ; P3_U5046
g8844 nand P3_U3151 P3_REG3_REG_11__SCAN_IN ; P3_U5047
g8845 nand P3_U3036 P3_U3074 ; P3_U5048
g8846 nand P3_U3032 P3_U3065 ; P3_U5049
g8847 nand P3_SUB_609_U17 P3_U3304 ; P3_U5050
g8848 nand P3_U5049 P3_U5048 P3_U5050 ; P3_U5051
g8849 nand P3_U3045 P3_U3905 ; P3_U5052
g8850 nand P3_U3044 P3_SUB_609_U17 ; P3_U5053
g8851 nand P3_R1158_U108 P3_U3035 ; P3_U5054
g8852 nand P3_U3031 P3_U5051 ; P3_U5055
g8853 nand P3_U3151 P3_REG3_REG_22__SCAN_IN ; P3_U5056
g8854 nand P3_U3036 P3_U3071 ; P3_U5057
g8855 nand P3_U3032 P3_U3078 ; P3_U5058
g8856 nand P3_SUB_609_U24 P3_U3304 ; P3_U5059
g8857 nand P3_U5058 P3_U5057 P3_U5059 ; P3_U5060
g8858 nand P3_U3428 P3_U5420 ; P3_U5061
g8859 nand P3_SUB_609_U24 P3_U3371 ; P3_U5062
g8860 nand P3_R1158_U13 P3_U3035 ; P3_U5063
g8861 nand P3_U3031 P3_U5060 ; P3_U5064
g8862 nand P3_U3151 P3_REG3_REG_13__SCAN_IN ; P3_U5065
g8863 nand P3_U3036 P3_U3080 ; P3_U5066
g8864 nand P3_U3032 P3_U3074 ; P3_U5067
g8865 nand P3_SUB_609_U20 P3_U3304 ; P3_U5068
g8866 nand P3_U5067 P3_U5066 P3_U5068 ; P3_U5069
g8867 nand P3_U3045 P3_U3907 ; P3_U5070
g8868 nand P3_U3044 P3_SUB_609_U20 ; P3_U5071
g8869 nand P3_R1158_U109 P3_U3035 ; P3_U5072
g8870 nand P3_U3031 P3_U5069 ; P3_U5073
g8871 nand P3_U3151 P3_REG3_REG_20__SCAN_IN ; P3_U5074
g8872 nand P3_U3031 P3_U3304 ; P3_U5075
g8873 nand P3_U5419 P3_U5075 ; P3_U5076
g8874 nand P3_U3787 P3_U3032 ; P3_U5077
g8875 nand P3_U3387 P3_U5420 ; P3_U5078
g8876 nand P3_U5076 P3_REG3_REG_0__SCAN_IN ; P3_U5079
g8877 nand P3_R1158_U94 P3_U3035 ; P3_U5080
g8878 nand P3_U3151 P3_REG3_REG_0__SCAN_IN ; P3_U5081
g8879 nand P3_U3036 P3_U3083 ; P3_U5082
g8880 nand P3_U3032 P3_U3061 ; P3_U5083
g8881 nand P3_SUB_609_U14 P3_U3304 ; P3_U5084
g8882 nand P3_U5083 P3_U5082 P3_U5084 ; P3_U5085
g8883 nand P3_U3416 P3_U5420 ; P3_U5086
g8884 nand P3_SUB_609_U14 P3_U3371 ; P3_U5087
g8885 nand P3_R1158_U95 P3_U3035 ; P3_U5088
g8886 nand P3_U3031 P3_U5085 ; P3_U5089
g8887 nand P3_U3151 P3_REG3_REG_9__SCAN_IN ; P3_U5090
g8888 nand P3_U3036 P3_U3063 ; P3_U5091
g8889 nand P3_U3032 P3_U3066 ; P3_U5092
g8890 nand P3_SUB_609_U29 P3_U3304 ; P3_U5093
g8891 nand P3_U5092 P3_U5091 P3_U5093 ; P3_U5094
g8892 nand P3_U3401 P3_U5420 ; P3_U5095
g8893 nand P3_SUB_609_U29 P3_U3371 ; P3_U5096
g8894 nand P3_R1158_U99 P3_U3035 ; P3_U5097
g8895 nand P3_U3031 P3_U5094 ; P3_U5098
g8896 nand P3_U3151 P3_REG3_REG_4__SCAN_IN ; P3_U5099
g8897 nand P3_U3036 P3_U3065 ; P3_U5100
g8898 nand P3_U3032 P3_U3057 ; P3_U5101
g8899 nand P3_SUB_609_U10 P3_U3304 ; P3_U5102
g8900 nand P3_U5101 P3_U5100 P3_U5102 ; P3_U5103
g8901 nand P3_U3045 P3_U3903 ; P3_U5104
g8902 nand P3_U3044 P3_SUB_609_U10 ; P3_U5105
g8903 nand P3_R1158_U106 P3_U3035 ; P3_U5106
g8904 nand P3_U3031 P3_U5103 ; P3_U5107
g8905 nand P3_U3151 P3_REG3_REG_24__SCAN_IN ; P3_U5108
g8906 nand P3_U3036 P3_U3072 ; P3_U5109
g8907 nand P3_U3032 P3_U3081 ; P3_U5110
g8908 nand P3_SUB_609_U19 P3_U3304 ; P3_U5111
g8909 nand P3_U5110 P3_U5109 P3_U5111 ; P3_U5112
g8910 nand P3_U3440 P3_U5420 ; P3_U5113
g8911 nand P3_SUB_609_U19 P3_U3371 ; P3_U5114
g8912 nand P3_R1158_U14 P3_U3035 ; P3_U5115
g8913 nand P3_U3031 P3_U5112 ; P3_U5116
g8914 nand P3_U3151 P3_REG3_REG_17__SCAN_IN ; P3_U5117
g8915 nand P3_U3036 P3_U3059 ; P3_U5118
g8916 nand P3_U3032 P3_U3070 ; P3_U5119
g8917 nand P3_SUB_609_U53 P3_U3304 ; P3_U5120
g8918 nand P3_U5119 P3_U5118 P3_U5120 ; P3_U5121
g8919 nand P3_U3404 P3_U5420 ; P3_U5122
g8920 nand P3_SUB_609_U53 P3_U3371 ; P3_U5123
g8921 nand P3_R1158_U98 P3_U3035 ; P3_U5124
g8922 nand P3_U3031 P3_U5121 ; P3_U5125
g8923 nand P3_U3151 P3_REG3_REG_5__SCAN_IN ; P3_U5126
g8924 nand P3_U3036 P3_U3073 ; P3_U5127
g8925 nand P3_U3032 P3_U3068 ; P3_U5128
g8926 nand P3_SUB_609_U7 P3_U3304 ; P3_U5129
g8927 nand P3_U5128 P3_U5127 P3_U5129 ; P3_U5130
g8928 nand P3_U3437 P3_U5420 ; P3_U5131
g8929 nand P3_SUB_609_U7 P3_U3371 ; P3_U5132
g8930 nand P3_R1158_U113 P3_U3035 ; P3_U5133
g8931 nand P3_U3031 P3_U5130 ; P3_U5134
g8932 nand P3_U3151 P3_REG3_REG_16__SCAN_IN ; P3_U5135
g8933 nand P3_U3036 P3_U3064 ; P3_U5136
g8934 nand P3_U3032 P3_U3056 ; P3_U5137
g8935 nand P3_SUB_609_U16 P3_U3304 ; P3_U5138
g8936 nand P3_U5137 P3_U5136 P3_U5138 ; P3_U5139
g8937 nand P3_U3045 P3_U3902 ; P3_U5140
g8938 nand P3_U3044 P3_SUB_609_U16 ; P3_U5141
g8939 nand P3_R1158_U105 P3_U3035 ; P3_U5142
g8940 nand P3_U3031 P3_U5139 ; P3_U5143
g8941 nand P3_U3151 P3_REG3_REG_25__SCAN_IN ; P3_U5144
g8942 nand P3_U3036 P3_U3062 ; P3_U5145
g8943 nand P3_U3032 P3_U3079 ; P3_U5146
g8944 nand P3_SUB_609_U23 P3_U3304 ; P3_U5147
g8945 nand P3_U5146 P3_U5145 P3_U5147 ; P3_U5148
g8946 nand P3_U3425 P3_U5420 ; P3_U5149
g8947 nand P3_SUB_609_U23 P3_U3371 ; P3_U5150
g8948 nand P3_R1158_U116 P3_U3035 ; P3_U5151
g8949 nand P3_U3031 P3_U5148 ; P3_U5152
g8950 nand P3_U3151 P3_REG3_REG_12__SCAN_IN ; P3_U5153
g8951 nand P3_U3036 P3_U3075 ; P3_U5154
g8952 nand P3_U3032 P3_U3060 ; P3_U5155
g8953 nand P3_SUB_609_U27 P3_U3304 ; P3_U5156
g8954 nand P3_U5155 P3_U5154 P3_U5156 ; P3_U5157
g8955 nand P3_U3045 P3_U3906 ; P3_U5158
g8956 nand P3_U3044 P3_SUB_609_U27 ; P3_U5159
g8957 nand P3_R1158_U15 P3_U3035 ; P3_U5160
g8958 nand P3_U3031 P3_U5157 ; P3_U5161
g8959 nand P3_U3151 P3_REG3_REG_21__SCAN_IN ; P3_U5162
g8960 nand P3_U3036 P3_U3076 ; P3_U5163
g8961 nand P3_U3032 P3_U3067 ; P3_U5164
g8962 nand P3_U3304 P3_REG3_REG_1__SCAN_IN ; P3_U5165
g8963 nand P3_U5164 P3_U5163 P3_U5165 ; P3_U5166
g8964 nand P3_U3392 P3_U5420 ; P3_U5167
g8965 nand P3_U3371 P3_REG3_REG_1__SCAN_IN ; P3_U5168
g8966 nand P3_R1158_U110 P3_U3035 ; P3_U5169
g8967 nand P3_U3031 P3_U5166 ; P3_U5170
g8968 nand P3_U3151 P3_REG3_REG_1__SCAN_IN ; P3_U5171
g8969 nand P3_U3036 P3_U3069 ; P3_U5172
g8970 nand P3_U3032 P3_U3082 ; P3_U5173
g8971 nand P3_SUB_609_U12 P3_U3304 ; P3_U5174
g8972 nand P3_U5173 P3_U5172 P3_U5174 ; P3_U5175
g8973 nand P3_U3413 P3_U5420 ; P3_U5176
g8974 nand P3_SUB_609_U12 P3_U3371 ; P3_U5177
g8975 nand P3_R1158_U96 P3_U3035 ; P3_U5178
g8976 nand P3_U3031 P3_U5175 ; P3_U5179
g8977 nand P3_U3151 P3_REG3_REG_8__SCAN_IN ; P3_U5180
g8978 nand P3_U3036 P3_U3052 ; P3_U5181
g8979 nand P3_U3032 P3_U3054 ; P3_U5182
g8980 nand P3_SUB_609_U28 P3_U3304 ; P3_U5183
g8981 nand P3_U5182 P3_U5181 P3_U5183 ; P3_U5184
g8982 nand P3_U3045 P3_U3899 ; P3_U5185
g8983 nand P3_U3044 P3_SUB_609_U28 ; P3_U5186
g8984 nand P3_R1158_U101 P3_U3035 ; P3_U5187
g8985 nand P3_U3031 P3_U5184 ; P3_U5188
g8986 nand P3_U3151 P3_REG3_REG_28__SCAN_IN ; P3_U5189
g8987 nand P3_U3036 P3_U3081 ; P3_U5190
g8988 nand P3_U3032 P3_U3075 ; P3_U5191
g8989 nand P3_SUB_609_U15 P3_U3304 ; P3_U5192
g8990 nand P3_U5191 P3_U5190 P3_U5192 ; P3_U5193
g8991 nand P3_U3445 P3_U5420 ; P3_U5194
g8992 nand P3_SUB_609_U15 P3_U3371 ; P3_U5195
g8993 nand P3_R1158_U111 P3_U3035 ; P3_U5196
g8994 nand P3_U3031 P3_U5193 ; P3_U5197
g8995 nand P3_U3151 P3_REG3_REG_19__SCAN_IN ; P3_U5198
g8996 nand P3_U3036 P3_U3067 ; P3_U5199
g8997 nand P3_U3032 P3_U3059 ; P3_U5200
g8998 nand P3_SUB_609_U25 P3_U3304 ; P3_U5201
g8999 nand P3_U5200 P3_U5199 P3_U5201 ; P3_U5202
g9000 nand P3_U3398 P3_U5420 ; P3_U5203
g9001 nand P3_SUB_609_U25 P3_U3371 ; P3_U5204
g9002 nand P3_R1158_U17 P3_U3035 ; P3_U5205
g9003 nand P3_U3031 P3_U5202 ; P3_U5206
g9004 nand P3_U3151 P3_REG3_REG_3__SCAN_IN ; P3_U5207
g9005 nand P3_U3036 P3_U3082 ; P3_U5208
g9006 nand P3_U3032 P3_U3062 ; P3_U5209
g9007 nand P3_SUB_609_U13 P3_U3304 ; P3_U5210
g9008 nand P3_U5209 P3_U5208 P3_U5210 ; P3_U5211
g9009 nand P3_U3419 P3_U5420 ; P3_U5212
g9010 nand P3_SUB_609_U13 P3_U3371 ; P3_U5213
g9011 nand P3_R1158_U118 P3_U3035 ; P3_U5214
g9012 nand P3_U3031 P3_U5211 ; P3_U5215
g9013 nand P3_U3151 P3_REG3_REG_10__SCAN_IN ; P3_U5216
g9014 nand P3_U3036 P3_U3060 ; P3_U5217
g9015 nand P3_U3032 P3_U3064 ; P3_U5218
g9016 nand P3_SUB_609_U6 P3_U3304 ; P3_U5219
g9017 nand P3_U5218 P3_U5217 P3_U5219 ; P3_U5220
g9018 nand P3_U3045 P3_U3904 ; P3_U5221
g9019 nand P3_U3044 P3_SUB_609_U6 ; P3_U5222
g9020 nand P3_R1158_U107 P3_U3035 ; P3_U5223
g9021 nand P3_U3031 P3_U5220 ; P3_U5224
g9022 nand P3_U3151 P3_REG3_REG_23__SCAN_IN ; P3_U5225
g9023 nand P3_U3036 P3_U3079 ; P3_U5226
g9024 nand P3_U3032 P3_U3073 ; P3_U5227
g9025 nand P3_SUB_609_U30 P3_U3304 ; P3_U5228
g9026 nand P3_U5227 P3_U5226 P3_U5228 ; P3_U5229
g9027 nand P3_U3431 P3_U5420 ; P3_U5230
g9028 nand P3_SUB_609_U30 P3_U3371 ; P3_U5231
g9029 nand P3_R1158_U115 P3_U3035 ; P3_U5232
g9030 nand P3_U3031 P3_U5229 ; P3_U5233
g9031 nand P3_U3151 P3_REG3_REG_14__SCAN_IN ; P3_U5234
g9032 nand P3_U3036 P3_U3056 ; P3_U5235
g9033 nand P3_U3032 P3_U3053 ; P3_U5236
g9034 nand P3_SUB_609_U22 P3_U3304 ; P3_U5237
g9035 nand P3_U5236 P3_U5235 P3_U5237 ; P3_U5238
g9036 nand P3_U3045 P3_U3900 ; P3_U5239
g9037 nand P3_U3044 P3_SUB_609_U22 ; P3_U5240
g9038 nand P3_R1158_U102 P3_U3035 ; P3_U5241
g9039 nand P3_U3031 P3_U5238 ; P3_U5242
g9040 nand P3_U3151 P3_REG3_REG_27__SCAN_IN ; P3_U5243
g9041 nand P3_U3036 P3_U3070 ; P3_U5244
g9042 nand P3_U3032 P3_U3083 ; P3_U5245
g9043 nand P3_SUB_609_U18 P3_U3304 ; P3_U5246
g9044 nand P3_U5245 P3_U5244 P3_U5246 ; P3_U5247
g9045 nand P3_U3410 P3_U5420 ; P3_U5248
g9046 nand P3_SUB_609_U18 P3_U3371 ; P3_U5249
g9047 nand P3_R1158_U18 P3_U3035 ; P3_U5250
g9048 nand P3_U3031 P3_U5247 ; P3_U5251
g9049 nand P3_U3151 P3_REG3_REG_7__SCAN_IN ; P3_U5252
g9050 nand P3_U3898 P3_U3046 ; P3_U5253
g9051 nand P3_U3375 P3_U3833 ; P3_U5254
g9052 nand P3_U3816 P3_U3815 ; P3_U5255
g9053 nand P3_U3814 P3_U3013 ; P3_U5256
g9054 nand P3_U3880 P3_U5256 ; P3_U5257
g9055 nand P3_U3416 P3_U5257 ; P3_U5258
g9056 nand P3_U5255 P3_U3082 ; P3_U5259
g9057 nand P3_U3413 P3_U5257 ; P3_U5260
g9058 nand P3_U5255 P3_U3083 ; P3_U5261
g9059 nand P3_U3410 P3_U5257 ; P3_U5262
g9060 nand P3_U5255 P3_U3069 ; P3_U5263
g9061 nand P3_U3407 P3_U5257 ; P3_U5264
g9062 nand P3_U5255 P3_U3070 ; P3_U5265
g9063 nand P3_U3404 P3_U5257 ; P3_U5266
g9064 nand P3_U5255 P3_U3066 ; P3_U5267
g9065 nand P3_U3401 P3_U5257 ; P3_U5268
g9066 nand P3_U5255 P3_U3059 ; P3_U5269
g9067 nand P3_U3872 P3_U5257 ; P3_U5270
g9068 nand P3_U5255 P3_U3055 ; P3_U5271
g9069 nand P3_U3873 P3_U5257 ; P3_U5272
g9070 nand P3_U5255 P3_U3058 ; P3_U5273
g9071 nand P3_U3398 P3_U5257 ; P3_U5274
g9072 nand P3_U5255 P3_U3063 ; P3_U5275
g9073 nand P3_U3908 P3_U5257 ; P3_U5276
g9074 nand P3_U5255 P3_U3054 ; P3_U5277
g9075 nand P3_U3899 P3_U5257 ; P3_U5278
g9076 nand P3_U5255 P3_U3053 ; P3_U5279
g9077 nand P3_U3900 P3_U5257 ; P3_U5280
g9078 nand P3_U5255 P3_U3052 ; P3_U5281
g9079 nand P3_U3901 P3_U5257 ; P3_U5282
g9080 nand P3_U5255 P3_U3056 ; P3_U5283
g9081 nand P3_U3902 P3_U5257 ; P3_U5284
g9082 nand P3_U5255 P3_U3057 ; P3_U5285
g9083 nand P3_U3903 P3_U5257 ; P3_U5286
g9084 nand P3_U5255 P3_U3064 ; P3_U5287
g9085 nand P3_U3904 P3_U5257 ; P3_U5288
g9086 nand P3_U5255 P3_U3065 ; P3_U5289
g9087 nand P3_U3905 P3_U5257 ; P3_U5290
g9088 nand P3_U5255 P3_U3060 ; P3_U5291
g9089 nand P3_U3906 P3_U5257 ; P3_U5292
g9090 nand P3_U5255 P3_U3074 ; P3_U5293
g9091 nand P3_U3907 P3_U5257 ; P3_U5294
g9092 nand P3_U5255 P3_U3075 ; P3_U5295
g9093 nand P3_U3395 P3_U5257 ; P3_U5296
g9094 nand P3_U5255 P3_U3067 ; P3_U5297
g9095 nand P3_U3445 P3_U5257 ; P3_U5298
g9096 nand P3_U5255 P3_U3080 ; P3_U5299
g9097 nand P3_U3443 P3_U5257 ; P3_U5300
g9098 nand P3_U5255 P3_U3081 ; P3_U5301
g9099 nand P3_U3440 P3_U5257 ; P3_U5302
g9100 nand P3_U5255 P3_U3068 ; P3_U5303
g9101 nand P3_U3437 P3_U5257 ; P3_U5304
g9102 nand P3_U5255 P3_U3072 ; P3_U5305
g9103 nand P3_U3434 P3_U5257 ; P3_U5306
g9104 nand P3_U5255 P3_U3073 ; P3_U5307
g9105 nand P3_U3431 P3_U5257 ; P3_U5308
g9106 nand P3_U5255 P3_U3078 ; P3_U5309
g9107 nand P3_U3428 P3_U5257 ; P3_U5310
g9108 nand P3_U5255 P3_U3079 ; P3_U5311
g9109 nand P3_U3425 P3_U5257 ; P3_U5312
g9110 nand P3_U5255 P3_U3071 ; P3_U5313
g9111 nand P3_U3422 P3_U5257 ; P3_U5314
g9112 nand P3_U5255 P3_U3062 ; P3_U5315
g9113 nand P3_U3419 P3_U5257 ; P3_U5316
g9114 nand P3_U5255 P3_U3061 ; P3_U5317
g9115 nand P3_U3392 P3_U5257 ; P3_U5318
g9116 nand P3_U5255 P3_U3077 ; P3_U5319
g9117 nand P3_U3387 P3_U5257 ; P3_U5320
g9118 nand P3_U5255 P3_U3076 ; P3_U5321
g9119 nand P3_U3416 P3_U5255 ; P3_U5322
g9120 nand P3_U5257 P3_U3082 ; P3_U5323
g9121 nand P3_U5440 P3_U3083 ; P3_U5324
g9122 nand P3_U3413 P3_U5255 ; P3_U5325
g9123 nand P3_U5257 P3_U3083 ; P3_U5326
g9124 nand P3_U5440 P3_U3069 ; P3_U5327
g9125 nand P3_U3410 P3_U5255 ; P3_U5328
g9126 nand P3_U5257 P3_U3069 ; P3_U5329
g9127 nand P3_U5440 P3_U3070 ; P3_U5330
g9128 nand P3_U3407 P3_U5255 ; P3_U5331
g9129 nand P3_U5257 P3_U3070 ; P3_U5332
g9130 nand P3_U5440 P3_U3066 ; P3_U5333
g9131 nand P3_U3404 P3_U5255 ; P3_U5334
g9132 nand P3_U5257 P3_U3066 ; P3_U5335
g9133 nand P3_U5440 P3_U3059 ; P3_U5336
g9134 nand P3_U3401 P3_U5255 ; P3_U5337
g9135 nand P3_U5257 P3_U3059 ; P3_U5338
g9136 nand P3_U5440 P3_U3063 ; P3_U5339
g9137 nand P3_U5257 P3_U3055 ; P3_U5340
g9138 nand P3_U3872 P3_U5255 ; P3_U5341
g9139 nand P3_U5257 P3_U3058 ; P3_U5342
g9140 nand P3_U3873 P3_U5255 ; P3_U5343
g9141 nand P3_U3398 P3_U5255 ; P3_U5344
g9142 nand P3_U5257 P3_U3063 ; P3_U5345
g9143 nand P3_U5440 P3_U3067 ; P3_U5346
g9144 nand P3_U5257 P3_U3054 ; P3_U5347
g9145 nand P3_U3908 P3_U5255 ; P3_U5348
g9146 nand P3_U5440 P3_U3053 ; P3_U5349
g9147 nand P3_U5257 P3_U3053 ; P3_U5350
g9148 nand P3_U3899 P3_U5255 ; P3_U5351
g9149 nand P3_U5440 P3_U3052 ; P3_U5352
g9150 nand P3_U5257 P3_U3052 ; P3_U5353
g9151 nand P3_U3900 P3_U5255 ; P3_U5354
g9152 nand P3_U5440 P3_U3056 ; P3_U5355
g9153 nand P3_U5257 P3_U3056 ; P3_U5356
g9154 nand P3_U3901 P3_U5255 ; P3_U5357
g9155 nand P3_U5440 P3_U3057 ; P3_U5358
g9156 nand P3_U5257 P3_U3057 ; P3_U5359
g9157 nand P3_U3902 P3_U5255 ; P3_U5360
g9158 nand P3_U5440 P3_U3064 ; P3_U5361
g9159 nand P3_U5257 P3_U3064 ; P3_U5362
g9160 nand P3_U3903 P3_U5255 ; P3_U5363
g9161 nand P3_U5440 P3_U3065 ; P3_U5364
g9162 nand P3_U5257 P3_U3065 ; P3_U5365
g9163 nand P3_U3904 P3_U5255 ; P3_U5366
g9164 nand P3_U5440 P3_U3060 ; P3_U5367
g9165 nand P3_U5257 P3_U3060 ; P3_U5368
g9166 nand P3_U3905 P3_U5255 ; P3_U5369
g9167 nand P3_U5440 P3_U3074 ; P3_U5370
g9168 nand P3_U5257 P3_U3074 ; P3_U5371
g9169 nand P3_U3906 P3_U5255 ; P3_U5372
g9170 nand P3_U5440 P3_U3075 ; P3_U5373
g9171 nand P3_U5257 P3_U3075 ; P3_U5374
g9172 nand P3_U3907 P3_U5255 ; P3_U5375
g9173 nand P3_U5440 P3_U3080 ; P3_U5376
g9174 nand P3_U3395 P3_U5255 ; P3_U5377
g9175 nand P3_U5257 P3_U3067 ; P3_U5378
g9176 nand P3_U5440 P3_U3077 ; P3_U5379
g9177 nand P3_U3445 P3_U5255 ; P3_U5380
g9178 nand P3_U5257 P3_U3080 ; P3_U5381
g9179 nand P3_U5440 P3_U3081 ; P3_U5382
g9180 nand P3_U3443 P3_U5255 ; P3_U5383
g9181 nand P3_U5257 P3_U3081 ; P3_U5384
g9182 nand P3_U5440 P3_U3068 ; P3_U5385
g9183 nand P3_U3440 P3_U5255 ; P3_U5386
g9184 nand P3_U5257 P3_U3068 ; P3_U5387
g9185 nand P3_U5440 P3_U3072 ; P3_U5388
g9186 nand P3_U3437 P3_U5255 ; P3_U5389
g9187 nand P3_U5257 P3_U3072 ; P3_U5390
g9188 nand P3_U5440 P3_U3073 ; P3_U5391
g9189 nand P3_U3434 P3_U5255 ; P3_U5392
g9190 nand P3_U5257 P3_U3073 ; P3_U5393
g9191 nand P3_U5440 P3_U3078 ; P3_U5394
g9192 nand P3_U3431 P3_U5255 ; P3_U5395
g9193 nand P3_U5257 P3_U3078 ; P3_U5396
g9194 nand P3_U5440 P3_U3079 ; P3_U5397
g9195 nand P3_U3428 P3_U5255 ; P3_U5398
g9196 nand P3_U5257 P3_U3079 ; P3_U5399
g9197 nand P3_U5440 P3_U3071 ; P3_U5400
g9198 nand P3_U3425 P3_U5255 ; P3_U5401
g9199 nand P3_U5257 P3_U3071 ; P3_U5402
g9200 nand P3_U5440 P3_U3062 ; P3_U5403
g9201 nand P3_U3422 P3_U5255 ; P3_U5404
g9202 nand P3_U5257 P3_U3062 ; P3_U5405
g9203 nand P3_U5440 P3_U3061 ; P3_U5406
g9204 nand P3_U3419 P3_U5255 ; P3_U5407
g9205 nand P3_U5257 P3_U3061 ; P3_U5408
g9206 nand P3_U5440 P3_U3082 ; P3_U5409
g9207 nand P3_U3392 P3_U5255 ; P3_U5410
g9208 nand P3_U5257 P3_U3077 ; P3_U5411
g9209 nand P3_U5440 P3_U3076 ; P3_U5412
g9210 nand P3_U3387 P3_U5255 ; P3_U5413
g9211 nand P3_U5257 P3_U3076 ; P3_U5414
g9212 nand P3_U4981 P3_U3151 ; P3_U5415
g9213 nand P3_U4981 P3_U5440 P3_U4980 ; P3_U5416
g9214 nand P3_U3043 P3_U3303 ; P3_U5417
g9215 nand P3_U3043 P3_U3894 ; P3_U5418
g9216 not P3_U3371 ; P3_U5419
g9217 nand P3_U5418 P3_U3918 ; P3_U5420
g9218 nand P3_U5938 P3_U5937 P3_U3774 ; P3_U5421
g9219 nand P3_U5434 P3_U5428 ; P3_U5422
g9220 nand P3_U3879 P3_U3378 ; P3_U5423
g9221 nand P3_U3375 P3_U3833 ; P3_U5424
g9222 nand P3_U3876 P3_U5447 ; P3_U5425
g9223 nand P3_U3831 P3_IR_REG_24__SCAN_IN ; P3_U5426
g9224 nand P3_SUB_598_U18 P3_IR_REG_31__SCAN_IN ; P3_U5427
g9225 not P3_U3372 ; P3_U5428
g9226 nand P3_U3831 P3_IR_REG_25__SCAN_IN ; P3_U5429
g9227 nand P3_SUB_598_U81 P3_IR_REG_31__SCAN_IN ; P3_U5430
g9228 not P3_U3373 ; P3_U5431
g9229 nand P3_U3831 P3_IR_REG_26__SCAN_IN ; P3_U5432
g9230 nand P3_SUB_598_U19 P3_IR_REG_31__SCAN_IN ; P3_U5433
g9231 not P3_U3374 ; P3_U5434
g9232 nand P3_U5428 P3_B_REG_SCAN_IN ; P3_U5435
g9233 nand P3_U3372 P3_U3298 ; P3_U5436
g9234 nand P3_U5436 P3_U5435 ; P3_U5437
g9235 nand P3_U3831 P3_IR_REG_23__SCAN_IN ; P3_U5438
g9236 nand P3_SUB_598_U17 P3_IR_REG_31__SCAN_IN ; P3_U5439
g9237 not P3_U3375 ; P3_U5440
g9238 nand P3_U3832 P3_D_REG_0__SCAN_IN ; P3_U5441
g9239 nand P3_U3915 P3_U4020 ; P3_U5442
g9240 nand P3_U3832 P3_D_REG_1__SCAN_IN ; P3_U5443
g9241 nand P3_U3915 P3_U4021 ; P3_U5444
g9242 nand P3_U3831 P3_IR_REG_20__SCAN_IN ; P3_U5445
g9243 nand P3_SUB_598_U15 P3_IR_REG_31__SCAN_IN ; P3_U5446
g9244 not P3_U3378 ; P3_U5447
g9245 nand P3_U3831 P3_IR_REG_19__SCAN_IN ; P3_U5448
g9246 nand P3_SUB_598_U14 P3_IR_REG_31__SCAN_IN ; P3_U5449
g9247 not P3_U3379 ; P3_U5450
g9248 nand P3_U3831 P3_IR_REG_22__SCAN_IN ; P3_U5451
g9249 nand P3_SUB_598_U16 P3_IR_REG_31__SCAN_IN ; P3_U5452
g9250 not P3_U3380 ; P3_U5453
g9251 nand P3_U3831 P3_IR_REG_21__SCAN_IN ; P3_U5454
g9252 nand P3_SUB_598_U83 P3_IR_REG_31__SCAN_IN ; P3_U5455
g9253 not P3_U3385 ; P3_U5456
g9254 nand P3_U3831 P3_IR_REG_30__SCAN_IN ; P3_U5457
g9255 nand P3_SUB_598_U77 P3_IR_REG_31__SCAN_IN ; P3_U5458
g9256 not P3_U3381 ; P3_U5459
g9257 nand P3_U3831 P3_IR_REG_29__SCAN_IN ; P3_U5460
g9258 nand P3_SUB_598_U21 P3_IR_REG_31__SCAN_IN ; P3_U5461
g9259 not P3_U3382 ; P3_U5462
g9260 nand P3_U3831 P3_IR_REG_28__SCAN_IN ; P3_U5463
g9261 nand P3_SUB_598_U20 P3_IR_REG_31__SCAN_IN ; P3_U5464
g9262 not P3_U3383 ; P3_U5465
g9263 nand P3_U3831 P3_IR_REG_27__SCAN_IN ; P3_U5466
g9264 nand P3_SUB_598_U79 P3_IR_REG_31__SCAN_IN ; P3_U5467
g9265 not P3_U3384 ; P3_U5468
g9266 nand P3_U3831 P3_IR_REG_0__SCAN_IN ; P3_U5469
g9267 nand P3_IR_REG_0__SCAN_IN P3_IR_REG_31__SCAN_IN ; P3_U5470
g9268 nand U61 P3_U3833 ; P3_U5471
g9269 nand P3_U3893 P3_U3386 ; P3_U5472
g9270 not P3_U3387 ; P3_U5473
g9271 nand P3_U5422 P3_U3300 ; P3_U5474
g9272 nand P3_U4019 P3_D_REG_0__SCAN_IN ; P3_U5475
g9273 not P3_U3388 ; P3_U5476
g9274 nand P3_U4019 P3_D_REG_1__SCAN_IN ; P3_U5477
g9275 nand P3_U4021 P3_U3300 ; P3_U5478
g9276 not P3_U3389 ; P3_U5479
g9277 nand P3_U4052 P3_U5453 ; P3_U5480
g9278 nand P3_U3380 P3_U3834 ; P3_U5481
g9279 nand P3_U5481 P3_U5480 ; P3_U5482
g9280 nand P3_U3835 P3_REG0_REG_0__SCAN_IN ; P3_U5483
g9281 nand P3_U3914 P3_U4077 ; P3_U5484
g9282 nand P3_U3831 P3_IR_REG_1__SCAN_IN ; P3_U5485
g9283 nand P3_SUB_598_U51 P3_IR_REG_31__SCAN_IN ; P3_U5486
g9284 nand U50 P3_U3833 ; P3_U5487
g9285 nand P3_U3391 P3_U3893 ; P3_U5488
g9286 not P3_U3392 ; P3_U5489
g9287 nand P3_U3835 P3_REG0_REG_1__SCAN_IN ; P3_U5490
g9288 nand P3_U3914 P3_U4102 ; P3_U5491
g9289 nand P3_U3831 P3_IR_REG_2__SCAN_IN ; P3_U5492
g9290 nand P3_SUB_598_U22 P3_IR_REG_31__SCAN_IN ; P3_U5493
g9291 nand U39 P3_U3833 ; P3_U5494
g9292 nand P3_U3394 P3_U3893 ; P3_U5495
g9293 not P3_U3395 ; P3_U5496
g9294 nand P3_U3835 P3_REG0_REG_2__SCAN_IN ; P3_U5497
g9295 nand P3_U3914 P3_U4120 ; P3_U5498
g9296 nand P3_U3831 P3_IR_REG_3__SCAN_IN ; P3_U5499
g9297 nand P3_SUB_598_U23 P3_IR_REG_31__SCAN_IN ; P3_U5500
g9298 nand U36 P3_U3833 ; P3_U5501
g9299 nand P3_U3397 P3_U3893 ; P3_U5502
g9300 not P3_U3398 ; P3_U5503
g9301 nand P3_U3835 P3_REG0_REG_3__SCAN_IN ; P3_U5504
g9302 nand P3_U3914 P3_U4138 ; P3_U5505
g9303 nand P3_U3831 P3_IR_REG_4__SCAN_IN ; P3_U5506
g9304 nand P3_SUB_598_U24 P3_IR_REG_31__SCAN_IN ; P3_U5507
g9305 nand U35 P3_U3833 ; P3_U5508
g9306 nand P3_U3400 P3_U3893 ; P3_U5509
g9307 not P3_U3401 ; P3_U5510
g9308 nand P3_U3835 P3_REG0_REG_4__SCAN_IN ; P3_U5511
g9309 nand P3_U3914 P3_U4156 ; P3_U5512
g9310 nand P3_U3831 P3_IR_REG_5__SCAN_IN ; P3_U5513
g9311 nand P3_SUB_598_U74 P3_IR_REG_31__SCAN_IN ; P3_U5514
g9312 nand U34 P3_U3833 ; P3_U5515
g9313 nand P3_U3403 P3_U3893 ; P3_U5516
g9314 not P3_U3404 ; P3_U5517
g9315 nand P3_U3835 P3_REG0_REG_5__SCAN_IN ; P3_U5518
g9316 nand P3_U3914 P3_U4174 ; P3_U5519
g9317 nand P3_U3831 P3_IR_REG_6__SCAN_IN ; P3_U5520
g9318 nand P3_SUB_598_U25 P3_IR_REG_31__SCAN_IN ; P3_U5521
g9319 nand U33 P3_U3833 ; P3_U5522
g9320 nand P3_U3406 P3_U3893 ; P3_U5523
g9321 not P3_U3407 ; P3_U5524
g9322 nand P3_U3835 P3_REG0_REG_6__SCAN_IN ; P3_U5525
g9323 nand P3_U3914 P3_U4192 ; P3_U5526
g9324 nand P3_U3831 P3_IR_REG_7__SCAN_IN ; P3_U5527
g9325 nand P3_SUB_598_U26 P3_IR_REG_31__SCAN_IN ; P3_U5528
g9326 nand U32 P3_U3833 ; P3_U5529
g9327 nand P3_U3409 P3_U3893 ; P3_U5530
g9328 not P3_U3410 ; P3_U5531
g9329 nand P3_U3835 P3_REG0_REG_7__SCAN_IN ; P3_U5532
g9330 nand P3_U3914 P3_U4210 ; P3_U5533
g9331 nand P3_U3831 P3_IR_REG_8__SCAN_IN ; P3_U5534
g9332 nand P3_SUB_598_U27 P3_IR_REG_31__SCAN_IN ; P3_U5535
g9333 nand U31 P3_U3833 ; P3_U5536
g9334 nand P3_U3412 P3_U3893 ; P3_U5537
g9335 not P3_U3413 ; P3_U5538
g9336 nand P3_U3835 P3_REG0_REG_8__SCAN_IN ; P3_U5539
g9337 nand P3_U3914 P3_U4228 ; P3_U5540
g9338 nand P3_U3831 P3_IR_REG_9__SCAN_IN ; P3_U5541
g9339 nand P3_SUB_598_U72 P3_IR_REG_31__SCAN_IN ; P3_U5542
g9340 nand U30 P3_U3833 ; P3_U5543
g9341 nand P3_U3415 P3_U3893 ; P3_U5544
g9342 not P3_U3416 ; P3_U5545
g9343 nand P3_U3835 P3_REG0_REG_9__SCAN_IN ; P3_U5546
g9344 nand P3_U3914 P3_U4246 ; P3_U5547
g9345 nand P3_U3831 P3_IR_REG_10__SCAN_IN ; P3_U5548
g9346 nand P3_SUB_598_U7 P3_IR_REG_31__SCAN_IN ; P3_U5549
g9347 nand U60 P3_U3833 ; P3_U5550
g9348 nand P3_U3418 P3_U3893 ; P3_U5551
g9349 not P3_U3419 ; P3_U5552
g9350 nand P3_U3835 P3_REG0_REG_10__SCAN_IN ; P3_U5553
g9351 nand P3_U3914 P3_U4264 ; P3_U5554
g9352 nand P3_U3831 P3_IR_REG_11__SCAN_IN ; P3_U5555
g9353 nand P3_SUB_598_U8 P3_IR_REG_31__SCAN_IN ; P3_U5556
g9354 nand U59 P3_U3833 ; P3_U5557
g9355 nand P3_U3421 P3_U3893 ; P3_U5558
g9356 not P3_U3422 ; P3_U5559
g9357 nand P3_U3835 P3_REG0_REG_11__SCAN_IN ; P3_U5560
g9358 nand P3_U3914 P3_U4282 ; P3_U5561
g9359 nand P3_U3831 P3_IR_REG_12__SCAN_IN ; P3_U5562
g9360 nand P3_SUB_598_U9 P3_IR_REG_31__SCAN_IN ; P3_U5563
g9361 nand U58 P3_U3833 ; P3_U5564
g9362 nand P3_U3424 P3_U3893 ; P3_U5565
g9363 not P3_U3425 ; P3_U5566
g9364 nand P3_U3835 P3_REG0_REG_12__SCAN_IN ; P3_U5567
g9365 nand P3_U3914 P3_U4300 ; P3_U5568
g9366 nand P3_U3831 P3_IR_REG_13__SCAN_IN ; P3_U5569
g9367 nand P3_SUB_598_U89 P3_IR_REG_31__SCAN_IN ; P3_U5570
g9368 nand U57 P3_U3833 ; P3_U5571
g9369 nand P3_U3427 P3_U3893 ; P3_U5572
g9370 not P3_U3428 ; P3_U5573
g9371 nand P3_U3835 P3_REG0_REG_13__SCAN_IN ; P3_U5574
g9372 nand P3_U3914 P3_U4318 ; P3_U5575
g9373 nand P3_U3831 P3_IR_REG_14__SCAN_IN ; P3_U5576
g9374 nand P3_SUB_598_U10 P3_IR_REG_31__SCAN_IN ; P3_U5577
g9375 nand U56 P3_U3833 ; P3_U5578
g9376 nand P3_U3430 P3_U3893 ; P3_U5579
g9377 not P3_U3431 ; P3_U5580
g9378 nand P3_U3835 P3_REG0_REG_14__SCAN_IN ; P3_U5581
g9379 nand P3_U3914 P3_U4336 ; P3_U5582
g9380 nand P3_U3831 P3_IR_REG_15__SCAN_IN ; P3_U5583
g9381 nand P3_SUB_598_U11 P3_IR_REG_31__SCAN_IN ; P3_U5584
g9382 nand U55 P3_U3833 ; P3_U5585
g9383 nand P3_U3433 P3_U3893 ; P3_U5586
g9384 not P3_U3434 ; P3_U5587
g9385 nand P3_U3835 P3_REG0_REG_15__SCAN_IN ; P3_U5588
g9386 nand P3_U3914 P3_U4354 ; P3_U5589
g9387 nand P3_U3831 P3_IR_REG_16__SCAN_IN ; P3_U5590
g9388 nand P3_SUB_598_U12 P3_IR_REG_31__SCAN_IN ; P3_U5591
g9389 nand U54 P3_U3833 ; P3_U5592
g9390 nand P3_U3436 P3_U3893 ; P3_U5593
g9391 not P3_U3437 ; P3_U5594
g9392 nand P3_U3835 P3_REG0_REG_16__SCAN_IN ; P3_U5595
g9393 nand P3_U3914 P3_U4372 ; P3_U5596
g9394 nand P3_U3831 P3_IR_REG_17__SCAN_IN ; P3_U5597
g9395 nand P3_SUB_598_U87 P3_IR_REG_31__SCAN_IN ; P3_U5598
g9396 nand U53 P3_U3833 ; P3_U5599
g9397 nand P3_U3439 P3_U3893 ; P3_U5600
g9398 not P3_U3440 ; P3_U5601
g9399 nand P3_U3835 P3_REG0_REG_17__SCAN_IN ; P3_U5602
g9400 nand P3_U3914 P3_U4390 ; P3_U5603
g9401 nand P3_U3831 P3_IR_REG_18__SCAN_IN ; P3_U5604
g9402 nand P3_SUB_598_U13 P3_IR_REG_31__SCAN_IN ; P3_U5605
g9403 nand U52 P3_U3833 ; P3_U5606
g9404 nand P3_U3442 P3_U3893 ; P3_U5607
g9405 not P3_U3443 ; P3_U5608
g9406 nand P3_U3835 P3_REG0_REG_18__SCAN_IN ; P3_U5609
g9407 nand P3_U3914 P3_U4408 ; P3_U5610
g9408 nand U51 P3_U3833 ; P3_U5611
g9409 nand P3_U3893 P3_U3379 ; P3_U5612
g9410 not P3_U3445 ; P3_U5613
g9411 nand P3_U3835 P3_REG0_REG_19__SCAN_IN ; P3_U5614
g9412 nand P3_U3914 P3_U4426 ; P3_U5615
g9413 nand P3_U3835 P3_REG0_REG_20__SCAN_IN ; P3_U5616
g9414 nand P3_U3914 P3_U4444 ; P3_U5617
g9415 nand P3_U3835 P3_REG0_REG_21__SCAN_IN ; P3_U5618
g9416 nand P3_U3914 P3_U4462 ; P3_U5619
g9417 nand P3_U3835 P3_REG0_REG_22__SCAN_IN ; P3_U5620
g9418 nand P3_U3914 P3_U4480 ; P3_U5621
g9419 nand P3_U3835 P3_REG0_REG_23__SCAN_IN ; P3_U5622
g9420 nand P3_U3914 P3_U4498 ; P3_U5623
g9421 nand P3_U3835 P3_REG0_REG_24__SCAN_IN ; P3_U5624
g9422 nand P3_U3914 P3_U4516 ; P3_U5625
g9423 nand P3_U3835 P3_REG0_REG_25__SCAN_IN ; P3_U5626
g9424 nand P3_U3914 P3_U4534 ; P3_U5627
g9425 nand P3_U3835 P3_REG0_REG_26__SCAN_IN ; P3_U5628
g9426 nand P3_U3914 P3_U4552 ; P3_U5629
g9427 nand P3_U3835 P3_REG0_REG_27__SCAN_IN ; P3_U5630
g9428 nand P3_U3914 P3_U4570 ; P3_U5631
g9429 nand P3_U3835 P3_REG0_REG_28__SCAN_IN ; P3_U5632
g9430 nand P3_U3914 P3_U4588 ; P3_U5633
g9431 nand P3_U3835 P3_REG0_REG_29__SCAN_IN ; P3_U5634
g9432 nand P3_U3914 P3_U4608 ; P3_U5635
g9433 nand P3_U3835 P3_REG0_REG_30__SCAN_IN ; P3_U5636
g9434 nand P3_U3914 P3_U4615 ; P3_U5637
g9435 nand P3_U3835 P3_REG0_REG_31__SCAN_IN ; P3_U5638
g9436 nand P3_U3914 P3_U4617 ; P3_U5639
g9437 nand P3_U5453 P3_U3834 ; P3_U5640
g9438 nand P3_U4052 P3_U5450 ; P3_U5641
g9439 nand P3_U3836 P3_REG1_REG_0__SCAN_IN ; P3_U5642
g9440 nand P3_U3913 P3_U4077 ; P3_U5643
g9441 nand P3_U3836 P3_REG1_REG_1__SCAN_IN ; P3_U5644
g9442 nand P3_U3913 P3_U4102 ; P3_U5645
g9443 nand P3_U3836 P3_REG1_REG_2__SCAN_IN ; P3_U5646
g9444 nand P3_U3913 P3_U4120 ; P3_U5647
g9445 nand P3_U3836 P3_REG1_REG_3__SCAN_IN ; P3_U5648
g9446 nand P3_U3913 P3_U4138 ; P3_U5649
g9447 nand P3_U3836 P3_REG1_REG_4__SCAN_IN ; P3_U5650
g9448 nand P3_U3913 P3_U4156 ; P3_U5651
g9449 nand P3_U3836 P3_REG1_REG_5__SCAN_IN ; P3_U5652
g9450 nand P3_U3913 P3_U4174 ; P3_U5653
g9451 nand P3_U3836 P3_REG1_REG_6__SCAN_IN ; P3_U5654
g9452 nand P3_U3913 P3_U4192 ; P3_U5655
g9453 nand P3_U3836 P3_REG1_REG_7__SCAN_IN ; P3_U5656
g9454 nand P3_U3913 P3_U4210 ; P3_U5657
g9455 nand P3_U3836 P3_REG1_REG_8__SCAN_IN ; P3_U5658
g9456 nand P3_U3913 P3_U4228 ; P3_U5659
g9457 nand P3_U3836 P3_REG1_REG_9__SCAN_IN ; P3_U5660
g9458 nand P3_U3913 P3_U4246 ; P3_U5661
g9459 nand P3_U3836 P3_REG1_REG_10__SCAN_IN ; P3_U5662
g9460 nand P3_U3913 P3_U4264 ; P3_U5663
g9461 nand P3_U3836 P3_REG1_REG_11__SCAN_IN ; P3_U5664
g9462 nand P3_U3913 P3_U4282 ; P3_U5665
g9463 nand P3_U3836 P3_REG1_REG_12__SCAN_IN ; P3_U5666
g9464 nand P3_U3913 P3_U4300 ; P3_U5667
g9465 nand P3_U3836 P3_REG1_REG_13__SCAN_IN ; P3_U5668
g9466 nand P3_U3913 P3_U4318 ; P3_U5669
g9467 nand P3_U3836 P3_REG1_REG_14__SCAN_IN ; P3_U5670
g9468 nand P3_U3913 P3_U4336 ; P3_U5671
g9469 nand P3_U3836 P3_REG1_REG_15__SCAN_IN ; P3_U5672
g9470 nand P3_U3913 P3_U4354 ; P3_U5673
g9471 nand P3_U3836 P3_REG1_REG_16__SCAN_IN ; P3_U5674
g9472 nand P3_U3913 P3_U4372 ; P3_U5675
g9473 nand P3_U3836 P3_REG1_REG_17__SCAN_IN ; P3_U5676
g9474 nand P3_U3913 P3_U4390 ; P3_U5677
g9475 nand P3_U3836 P3_REG1_REG_18__SCAN_IN ; P3_U5678
g9476 nand P3_U3913 P3_U4408 ; P3_U5679
g9477 nand P3_U3836 P3_REG1_REG_19__SCAN_IN ; P3_U5680
g9478 nand P3_U3913 P3_U4426 ; P3_U5681
g9479 nand P3_U3836 P3_REG1_REG_20__SCAN_IN ; P3_U5682
g9480 nand P3_U3913 P3_U4444 ; P3_U5683
g9481 nand P3_U3836 P3_REG1_REG_21__SCAN_IN ; P3_U5684
g9482 nand P3_U3913 P3_U4462 ; P3_U5685
g9483 nand P3_U3836 P3_REG1_REG_22__SCAN_IN ; P3_U5686
g9484 nand P3_U3913 P3_U4480 ; P3_U5687
g9485 nand P3_U3836 P3_REG1_REG_23__SCAN_IN ; P3_U5688
g9486 nand P3_U3913 P3_U4498 ; P3_U5689
g9487 nand P3_U3836 P3_REG1_REG_24__SCAN_IN ; P3_U5690
g9488 nand P3_U3913 P3_U4516 ; P3_U5691
g9489 nand P3_U3836 P3_REG1_REG_25__SCAN_IN ; P3_U5692
g9490 nand P3_U3913 P3_U4534 ; P3_U5693
g9491 nand P3_U3836 P3_REG1_REG_26__SCAN_IN ; P3_U5694
g9492 nand P3_U3913 P3_U4552 ; P3_U5695
g9493 nand P3_U3836 P3_REG1_REG_27__SCAN_IN ; P3_U5696
g9494 nand P3_U3913 P3_U4570 ; P3_U5697
g9495 nand P3_U3836 P3_REG1_REG_28__SCAN_IN ; P3_U5698
g9496 nand P3_U3913 P3_U4588 ; P3_U5699
g9497 nand P3_U3836 P3_REG1_REG_29__SCAN_IN ; P3_U5700
g9498 nand P3_U3913 P3_U4608 ; P3_U5701
g9499 nand P3_U3836 P3_REG1_REG_30__SCAN_IN ; P3_U5702
g9500 nand P3_U3913 P3_U4615 ; P3_U5703
g9501 nand P3_U3836 P3_REG1_REG_31__SCAN_IN ; P3_U5704
g9502 nand P3_U3913 P3_U4617 ; P3_U5705
g9503 nand P3_U3358 P3_REG2_REG_0__SCAN_IN ; P3_U5706
g9504 nand P3_U3912 P3_U3314 ; P3_U5707
g9505 nand P3_U3358 P3_REG2_REG_1__SCAN_IN ; P3_U5708
g9506 nand P3_U3912 P3_U3315 ; P3_U5709
g9507 nand P3_U3358 P3_REG2_REG_2__SCAN_IN ; P3_U5710
g9508 nand P3_U3912 P3_U3316 ; P3_U5711
g9509 nand P3_U3358 P3_REG2_REG_3__SCAN_IN ; P3_U5712
g9510 nand P3_U3912 P3_U3317 ; P3_U5713
g9511 nand P3_U3358 P3_REG2_REG_4__SCAN_IN ; P3_U5714
g9512 nand P3_U3912 P3_U3318 ; P3_U5715
g9513 nand P3_U3358 P3_REG2_REG_5__SCAN_IN ; P3_U5716
g9514 nand P3_U3912 P3_U3319 ; P3_U5717
g9515 nand P3_U3358 P3_REG2_REG_6__SCAN_IN ; P3_U5718
g9516 nand P3_U3912 P3_U3320 ; P3_U5719
g9517 nand P3_U3358 P3_REG2_REG_7__SCAN_IN ; P3_U5720
g9518 nand P3_U3912 P3_U3321 ; P3_U5721
g9519 nand P3_U3358 P3_REG2_REG_8__SCAN_IN ; P3_U5722
g9520 nand P3_U3912 P3_U3322 ; P3_U5723
g9521 nand P3_U3358 P3_REG2_REG_9__SCAN_IN ; P3_U5724
g9522 nand P3_U3912 P3_U3323 ; P3_U5725
g9523 nand P3_U3358 P3_REG2_REG_10__SCAN_IN ; P3_U5726
g9524 nand P3_U3912 P3_U3324 ; P3_U5727
g9525 nand P3_U3358 P3_REG2_REG_11__SCAN_IN ; P3_U5728
g9526 nand P3_U3912 P3_U3325 ; P3_U5729
g9527 nand P3_U3358 P3_REG2_REG_12__SCAN_IN ; P3_U5730
g9528 nand P3_U3912 P3_U3326 ; P3_U5731
g9529 nand P3_U3358 P3_REG2_REG_13__SCAN_IN ; P3_U5732
g9530 nand P3_U3912 P3_U3327 ; P3_U5733
g9531 nand P3_U3358 P3_REG2_REG_14__SCAN_IN ; P3_U5734
g9532 nand P3_U3912 P3_U3328 ; P3_U5735
g9533 nand P3_U3358 P3_REG2_REG_15__SCAN_IN ; P3_U5736
g9534 nand P3_U3912 P3_U3329 ; P3_U5737
g9535 nand P3_U3358 P3_REG2_REG_16__SCAN_IN ; P3_U5738
g9536 nand P3_U3912 P3_U3330 ; P3_U5739
g9537 nand P3_U3358 P3_REG2_REG_17__SCAN_IN ; P3_U5740
g9538 nand P3_U3912 P3_U3331 ; P3_U5741
g9539 nand P3_U3358 P3_REG2_REG_18__SCAN_IN ; P3_U5742
g9540 nand P3_U3912 P3_U3332 ; P3_U5743
g9541 nand P3_U3358 P3_REG2_REG_19__SCAN_IN ; P3_U5744
g9542 nand P3_U3912 P3_U3333 ; P3_U5745
g9543 nand P3_U3358 P3_REG2_REG_20__SCAN_IN ; P3_U5746
g9544 nand P3_U3912 P3_U3335 ; P3_U5747
g9545 nand P3_U3358 P3_REG2_REG_21__SCAN_IN ; P3_U5748
g9546 nand P3_U3912 P3_U3337 ; P3_U5749
g9547 nand P3_U3358 P3_REG2_REG_22__SCAN_IN ; P3_U5750
g9548 nand P3_U3912 P3_U3339 ; P3_U5751
g9549 nand P3_U3358 P3_REG2_REG_23__SCAN_IN ; P3_U5752
g9550 nand P3_U3912 P3_U3341 ; P3_U5753
g9551 nand P3_U3358 P3_REG2_REG_24__SCAN_IN ; P3_U5754
g9552 nand P3_U3912 P3_U3343 ; P3_U5755
g9553 nand P3_U3358 P3_REG2_REG_25__SCAN_IN ; P3_U5756
g9554 nand P3_U3912 P3_U3345 ; P3_U5757
g9555 nand P3_U3358 P3_REG2_REG_26__SCAN_IN ; P3_U5758
g9556 nand P3_U3912 P3_U3347 ; P3_U5759
g9557 nand P3_U3358 P3_REG2_REG_27__SCAN_IN ; P3_U5760
g9558 nand P3_U3912 P3_U3349 ; P3_U5761
g9559 nand P3_U3358 P3_REG2_REG_28__SCAN_IN ; P3_U5762
g9560 nand P3_U3912 P3_U3351 ; P3_U5763
g9561 nand P3_U3358 P3_REG2_REG_29__SCAN_IN ; P3_U5764
g9562 nand P3_U3912 P3_U3354 ; P3_U5765
g9563 nand P3_U5465 P3_U3024 ; P3_U5766
g9564 nand P3_U3383 P3_U3897 ; P3_U5767
g9565 nand P3_U5767 P3_U5766 ; P3_U5768
g9566 nand P3_U3363 P3_DATAO_REG_0__SCAN_IN ; P3_U5769
g9567 nand P3_U3897 P3_U3076 ; P3_U5770
g9568 nand P3_U3363 P3_DATAO_REG_1__SCAN_IN ; P3_U5771
g9569 nand P3_U3897 P3_U3077 ; P3_U5772
g9570 nand P3_U3363 P3_DATAO_REG_2__SCAN_IN ; P3_U5773
g9571 nand P3_U3897 P3_U3067 ; P3_U5774
g9572 nand P3_U3363 P3_DATAO_REG_3__SCAN_IN ; P3_U5775
g9573 nand P3_U3897 P3_U3063 ; P3_U5776
g9574 nand P3_U3363 P3_DATAO_REG_4__SCAN_IN ; P3_U5777
g9575 nand P3_U3897 P3_U3059 ; P3_U5778
g9576 nand P3_U3363 P3_DATAO_REG_5__SCAN_IN ; P3_U5779
g9577 nand P3_U3897 P3_U3066 ; P3_U5780
g9578 nand P3_U3363 P3_DATAO_REG_6__SCAN_IN ; P3_U5781
g9579 nand P3_U3897 P3_U3070 ; P3_U5782
g9580 nand P3_U3363 P3_DATAO_REG_7__SCAN_IN ; P3_U5783
g9581 nand P3_U3897 P3_U3069 ; P3_U5784
g9582 nand P3_U3363 P3_DATAO_REG_8__SCAN_IN ; P3_U5785
g9583 nand P3_U3897 P3_U3083 ; P3_U5786
g9584 nand P3_U3363 P3_DATAO_REG_9__SCAN_IN ; P3_U5787
g9585 nand P3_U3897 P3_U3082 ; P3_U5788
g9586 nand P3_U3363 P3_DATAO_REG_10__SCAN_IN ; P3_U5789
g9587 nand P3_U3897 P3_U3061 ; P3_U5790
g9588 nand P3_U3363 P3_DATAO_REG_11__SCAN_IN ; P3_U5791
g9589 nand P3_U3897 P3_U3062 ; P3_U5792
g9590 nand P3_U3363 P3_DATAO_REG_12__SCAN_IN ; P3_U5793
g9591 nand P3_U3897 P3_U3071 ; P3_U5794
g9592 nand P3_U3363 P3_DATAO_REG_13__SCAN_IN ; P3_U5795
g9593 nand P3_U3897 P3_U3079 ; P3_U5796
g9594 nand P3_U3363 P3_DATAO_REG_14__SCAN_IN ; P3_U5797
g9595 nand P3_U3897 P3_U3078 ; P3_U5798
g9596 nand P3_U3363 P3_DATAO_REG_15__SCAN_IN ; P3_U5799
g9597 nand P3_U3897 P3_U3073 ; P3_U5800
g9598 nand P3_U3363 P3_DATAO_REG_16__SCAN_IN ; P3_U5801
g9599 nand P3_U3897 P3_U3072 ; P3_U5802
g9600 nand P3_U3363 P3_DATAO_REG_17__SCAN_IN ; P3_U5803
g9601 nand P3_U3897 P3_U3068 ; P3_U5804
g9602 nand P3_U3363 P3_DATAO_REG_18__SCAN_IN ; P3_U5805
g9603 nand P3_U3897 P3_U3081 ; P3_U5806
g9604 nand P3_U3363 P3_DATAO_REG_19__SCAN_IN ; P3_U5807
g9605 nand P3_U3897 P3_U3080 ; P3_U5808
g9606 nand P3_U3363 P3_DATAO_REG_20__SCAN_IN ; P3_U5809
g9607 nand P3_U3897 P3_U3075 ; P3_U5810
g9608 nand P3_U3363 P3_DATAO_REG_21__SCAN_IN ; P3_U5811
g9609 nand P3_U3897 P3_U3074 ; P3_U5812
g9610 nand P3_U3363 P3_DATAO_REG_22__SCAN_IN ; P3_U5813
g9611 nand P3_U3897 P3_U3060 ; P3_U5814
g9612 nand P3_U3363 P3_DATAO_REG_23__SCAN_IN ; P3_U5815
g9613 nand P3_U3897 P3_U3065 ; P3_U5816
g9614 nand P3_U3363 P3_DATAO_REG_24__SCAN_IN ; P3_U5817
g9615 nand P3_U3897 P3_U3064 ; P3_U5818
g9616 nand P3_U3363 P3_DATAO_REG_25__SCAN_IN ; P3_U5819
g9617 nand P3_U3897 P3_U3057 ; P3_U5820
g9618 nand P3_U3363 P3_DATAO_REG_26__SCAN_IN ; P3_U5821
g9619 nand P3_U3897 P3_U3056 ; P3_U5822
g9620 nand P3_U3363 P3_DATAO_REG_27__SCAN_IN ; P3_U5823
g9621 nand P3_U3897 P3_U3052 ; P3_U5824
g9622 nand P3_U3363 P3_DATAO_REG_28__SCAN_IN ; P3_U5825
g9623 nand P3_U3897 P3_U3053 ; P3_U5826
g9624 nand P3_U3363 P3_DATAO_REG_29__SCAN_IN ; P3_U5827
g9625 nand P3_U3897 P3_U3054 ; P3_U5828
g9626 nand P3_U3363 P3_DATAO_REG_30__SCAN_IN ; P3_U5829
g9627 nand P3_U3897 P3_U3058 ; P3_U5830
g9628 nand P3_U3363 P3_DATAO_REG_31__SCAN_IN ; P3_U5831
g9629 nand P3_U3897 P3_U3055 ; P3_U5832
g9630 nand P3_U3379 P3_U3313 ; P3_U5833
g9631 nand P3_U5450 P3_U3911 ; P3_U5834
g9632 not P3_U3760 ; P3_U5835
g9633 nand P3_R1269_U11 P3_U5835 ; P3_U5836
g9634 nand P3_U3760 P3_U3867 ; P3_U5837
g9635 nand P3_U3900 P3_U3052 ; P3_U5838
g9636 nand P3_U3348 P3_U4539 ; P3_U5839
g9637 nand P3_U5839 P3_U5838 ; P3_U5840
g9638 nand P3_U3899 P3_U3053 ; P3_U5841
g9639 nand P3_U3350 P3_U4557 ; P3_U5842
g9640 nand P3_U5842 P3_U5841 ; P3_U5843
g9641 nand P3_U3872 P3_U3055 ; P3_U5844
g9642 nand P3_U3356 P3_U4613 ; P3_U5845
g9643 nand P3_U5845 P3_U5844 ; P3_U5846
g9644 nand P3_U3908 P3_U3054 ; P3_U5847
g9645 nand P3_U3353 P3_U4575 ; P3_U5848
g9646 nand P3_U5848 P3_U5847 ; P3_U5849
g9647 nand P3_U3906 P3_U3074 ; P3_U5850
g9648 nand P3_U3336 P3_U4431 ; P3_U5851
g9649 nand P3_U5851 P3_U5850 ; P3_U5852
g9650 nand P3_U3907 P3_U3075 ; P3_U5853
g9651 nand P3_U3334 P3_U4413 ; P3_U5854
g9652 nand P3_U5854 P3_U5853 ; P3_U5855
g9653 nand P3_U5503 P3_U4107 ; P3_U5856
g9654 nand P3_U3398 P3_U3063 ; P3_U5857
g9655 nand P3_U5857 P3_U5856 ; P3_U5858
g9656 nand P3_U5559 P3_U4251 ; P3_U5859
g9657 nand P3_U3422 P3_U3062 ; P3_U5860
g9658 nand P3_U5860 P3_U5859 ; P3_U5861
g9659 nand P3_U5552 P3_U4233 ; P3_U5862
g9660 nand P3_U3419 P3_U3061 ; P3_U5863
g9661 nand P3_U5863 P3_U5862 ; P3_U5864
g9662 nand P3_U5510 P3_U4125 ; P3_U5865
g9663 nand P3_U3401 P3_U3059 ; P3_U5866
g9664 nand P3_U5866 P3_U5865 ; P3_U5867
g9665 nand P3_U3905 P3_U3060 ; P3_U5868
g9666 nand P3_U3338 P3_U4449 ; P3_U5869
g9667 nand P3_U5869 P3_U5868 ; P3_U5870
g9668 nand P3_U5601 P3_U4359 ; P3_U5871
g9669 nand P3_U3440 P3_U3068 ; P3_U5872
g9670 nand P3_U5872 P3_U5871 ; P3_U5873
g9671 nand P3_U5594 P3_U4341 ; P3_U5874
g9672 nand P3_U3437 P3_U3072 ; P3_U5875
g9673 nand P3_U5875 P3_U5874 ; P3_U5876
g9674 nand P3_U5587 P3_U4323 ; P3_U5877
g9675 nand P3_U3434 P3_U3073 ; P3_U5878
g9676 nand P3_U5878 P3_U5877 ; P3_U5879
g9677 nand P3_U5566 P3_U4269 ; P3_U5880
g9678 nand P3_U3425 P3_U3071 ; P3_U5881
g9679 nand P3_U5881 P3_U5880 ; P3_U5882
g9680 nand P3_U5524 P3_U4161 ; P3_U5883
g9681 nand P3_U3407 P3_U3070 ; P3_U5884
g9682 nand P3_U5884 P3_U5883 ; P3_U5885
g9683 nand P3_U5531 P3_U4179 ; P3_U5886
g9684 nand P3_U3410 P3_U3069 ; P3_U5887
g9685 nand P3_U5887 P3_U5886 ; P3_U5888
g9686 nand P3_U5496 P3_U4082 ; P3_U5889
g9687 nand P3_U3395 P3_U3067 ; P3_U5890
g9688 nand P3_U5890 P3_U5889 ; P3_U5891
g9689 nand P3_U5517 P3_U4143 ; P3_U5892
g9690 nand P3_U3404 P3_U3066 ; P3_U5893
g9691 nand P3_U5893 P3_U5892 ; P3_U5894
g9692 nand P3_U5608 P3_U4377 ; P3_U5895
g9693 nand P3_U3443 P3_U3081 ; P3_U5896
g9694 nand P3_U5896 P3_U5895 ; P3_U5897
g9695 nand P3_U5573 P3_U4287 ; P3_U5898
g9696 nand P3_U3428 P3_U3079 ; P3_U5899
g9697 nand P3_U5899 P3_U5898 ; P3_U5900
g9698 nand P3_U5580 P3_U4305 ; P3_U5901
g9699 nand P3_U3431 P3_U3078 ; P3_U5902
g9700 nand P3_U5902 P3_U5901 ; P3_U5903
g9701 nand P3_U5489 P3_U4063 ; P3_U5904
g9702 nand P3_U3392 P3_U3077 ; P3_U5905
g9703 nand P3_U5905 P3_U5904 ; P3_U5906
g9704 nand P3_U5473 P3_U4087 ; P3_U5907
g9705 nand P3_U3387 P3_U3076 ; P3_U5908
g9706 nand P3_U5908 P3_U5907 ; P3_U5909
g9707 nand P3_U5538 P3_U4197 ; P3_U5910
g9708 nand P3_U3413 P3_U3083 ; P3_U5911
g9709 nand P3_U5911 P3_U5910 ; P3_U5912
g9710 nand P3_U5545 P3_U4215 ; P3_U5913
g9711 nand P3_U3416 P3_U3082 ; P3_U5914
g9712 nand P3_U5914 P3_U5913 ; P3_U5915
g9713 nand P3_U5613 P3_U4395 ; P3_U5916
g9714 nand P3_U3445 P3_U3080 ; P3_U5917
g9715 nand P3_U5917 P3_U5916 ; P3_U5918
g9716 nand P3_U3901 P3_U3056 ; P3_U5919
g9717 nand P3_U3346 P3_U4521 ; P3_U5920
g9718 nand P3_U5920 P3_U5919 ; P3_U5921
g9719 nand P3_U3902 P3_U3057 ; P3_U5922
g9720 nand P3_U3344 P3_U4503 ; P3_U5923
g9721 nand P3_U5923 P3_U5922 ; P3_U5924
g9722 nand P3_U3904 P3_U3065 ; P3_U5925
g9723 nand P3_U3340 P3_U4467 ; P3_U5926
g9724 nand P3_U5926 P3_U5925 ; P3_U5927
g9725 nand P3_U3903 P3_U3064 ; P3_U5928
g9726 nand P3_U3342 P3_U4485 ; P3_U5929
g9727 nand P3_U5929 P3_U5928 ; P3_U5930
g9728 nand P3_U3873 P3_U3058 ; P3_U5931
g9729 nand P3_U3355 P3_U4593 ; P3_U5932
g9730 nand P3_U5932 P3_U5931 ; P3_U5933
g9731 nand P3_U4978 P3_U5450 ; P3_U5934
g9732 nand P3_U3379 P3_U3868 ; P3_U5935
g9733 nand P3_U5935 P3_U5934 ; P3_U5936
g9734 nand P3_U5837 P3_U5836 P3_U5447 ; P3_U5937
g9735 nand P3_U5456 P3_U5936 P3_U3378 ; P3_U5938
g9736 nand P3_U3881 P3_U3869 ; P3_U5939
g9737 nand P3_R693_U14 P3_U3891 ; P3_U5940
g9738 nand P3_U5440 P3_U3368 ; P3_U5941
g9739 nand P3_U3380 P3_U3375 ; P3_U5942
g9740 nand P3_U5450 P3_U5447 ; P3_U5943
g9741 nand P3_U3388 P3_U5456 P3_U3378 ; P3_U5944
g9742 nand P3_U3082 P3_R1297_U6 ; P3_U5945
g9743 nand P3_U3082 P3_U3871 ; P3_U5946
g9744 nand P3_U3083 P3_R1297_U6 ; P3_U5947
g9745 nand P3_U3083 P3_U3871 ; P3_U5948
g9746 nand P3_U3069 P3_R1297_U6 ; P3_U5949
g9747 nand P3_U3069 P3_U3871 ; P3_U5950
g9748 nand P3_U3070 P3_R1297_U6 ; P3_U5951
g9749 nand P3_U3070 P3_U3871 ; P3_U5952
g9750 nand P3_U3066 P3_R1297_U6 ; P3_U5953
g9751 nand P3_U3066 P3_U3871 ; P3_U5954
g9752 nand P3_U3059 P3_R1297_U6 ; P3_U5955
g9753 nand P3_U3059 P3_U3871 ; P3_U5956
g9754 nand P3_R1300_U8 P3_R1297_U6 ; P3_U5957
g9755 nand P3_U3055 P3_U3871 ; P3_U5958
g9756 nand P3_R1300_U6 P3_R1297_U6 ; P3_U5959
g9757 nand P3_U3058 P3_U3871 ; P3_U5960
g9758 nand P3_U3063 P3_R1297_U6 ; P3_U5961
g9759 nand P3_U3063 P3_U3871 ; P3_U5962
g9760 nand P3_U3054 P3_R1297_U6 ; P3_U5963
g9761 nand P3_U3054 P3_U3871 ; P3_U5964
g9762 nand P3_U3053 P3_R1297_U6 ; P3_U5965
g9763 nand P3_U3053 P3_U3871 ; P3_U5966
g9764 nand P3_U3052 P3_R1297_U6 ; P3_U5967
g9765 nand P3_U3052 P3_U3871 ; P3_U5968
g9766 nand P3_U3056 P3_R1297_U6 ; P3_U5969
g9767 nand P3_U3056 P3_U3871 ; P3_U5970
g9768 nand P3_U3057 P3_R1297_U6 ; P3_U5971
g9769 nand P3_U3057 P3_U3871 ; P3_U5972
g9770 nand P3_U3064 P3_R1297_U6 ; P3_U5973
g9771 nand P3_U3064 P3_U3871 ; P3_U5974
g9772 nand P3_U3065 P3_R1297_U6 ; P3_U5975
g9773 nand P3_U3065 P3_U3871 ; P3_U5976
g9774 nand P3_U3060 P3_R1297_U6 ; P3_U5977
g9775 nand P3_U3060 P3_U3871 ; P3_U5978
g9776 nand P3_U3074 P3_R1297_U6 ; P3_U5979
g9777 nand P3_U3074 P3_U3871 ; P3_U5980
g9778 nand P3_U3075 P3_R1297_U6 ; P3_U5981
g9779 nand P3_U3075 P3_U3871 ; P3_U5982
g9780 nand P3_U3067 P3_R1297_U6 ; P3_U5983
g9781 nand P3_U3067 P3_U3871 ; P3_U5984
g9782 nand P3_U3080 P3_R1297_U6 ; P3_U5985
g9783 nand P3_U3080 P3_U3871 ; P3_U5986
g9784 nand P3_U3081 P3_R1297_U6 ; P3_U5987
g9785 nand P3_U3081 P3_U3871 ; P3_U5988
g9786 nand P3_U3068 P3_R1297_U6 ; P3_U5989
g9787 nand P3_U3068 P3_U3871 ; P3_U5990
g9788 nand P3_U3072 P3_R1297_U6 ; P3_U5991
g9789 nand P3_U3072 P3_U3871 ; P3_U5992
g9790 nand P3_U3073 P3_R1297_U6 ; P3_U5993
g9791 nand P3_U3073 P3_U3871 ; P3_U5994
g9792 nand P3_U3078 P3_R1297_U6 ; P3_U5995
g9793 nand P3_U3078 P3_U3871 ; P3_U5996
g9794 nand P3_U3079 P3_R1297_U6 ; P3_U5997
g9795 nand P3_U3079 P3_U3871 ; P3_U5998
g9796 nand P3_U3071 P3_R1297_U6 ; P3_U5999
g9797 nand P3_U3071 P3_U3871 ; P3_U6000
g9798 nand P3_U3062 P3_R1297_U6 ; P3_U6001
g9799 nand P3_U3062 P3_U3871 ; P3_U6002
g9800 nand P3_U3061 P3_R1297_U6 ; P3_U6003
g9801 nand P3_U3061 P3_U3871 ; P3_U6004
g9802 nand P3_U3077 P3_R1297_U6 ; P3_U6005
g9803 nand P3_U3077 P3_U3871 ; P3_U6006
g9804 nand P3_U3076 P3_R1297_U6 ; P3_U6007
g9805 nand P3_U3076 P3_U3871 ; P3_U6008
g9806 nand P3_U5468 P3_REG1_REG_9__SCAN_IN ; P3_U6009
g9807 nand P3_U3384 P3_REG2_REG_9__SCAN_IN ; P3_U6010
g9808 nand P3_U5468 P3_REG1_REG_8__SCAN_IN ; P3_U6011
g9809 nand P3_U3384 P3_REG2_REG_8__SCAN_IN ; P3_U6012
g9810 nand P3_U5468 P3_REG1_REG_7__SCAN_IN ; P3_U6013
g9811 nand P3_U3384 P3_REG2_REG_7__SCAN_IN ; P3_U6014
g9812 nand P3_U5468 P3_REG1_REG_6__SCAN_IN ; P3_U6015
g9813 nand P3_U3384 P3_REG2_REG_6__SCAN_IN ; P3_U6016
g9814 nand P3_U5468 P3_REG1_REG_5__SCAN_IN ; P3_U6017
g9815 nand P3_U3384 P3_REG2_REG_5__SCAN_IN ; P3_U6018
g9816 nand P3_U5468 P3_REG1_REG_4__SCAN_IN ; P3_U6019
g9817 nand P3_U3384 P3_REG2_REG_4__SCAN_IN ; P3_U6020
g9818 nand P3_U5468 P3_REG1_REG_3__SCAN_IN ; P3_U6021
g9819 nand P3_U3384 P3_REG2_REG_3__SCAN_IN ; P3_U6022
g9820 nand P3_U5468 P3_REG1_REG_2__SCAN_IN ; P3_U6023
g9821 nand P3_U3384 P3_REG2_REG_2__SCAN_IN ; P3_U6024
g9822 nand P3_U5468 P3_REG1_REG_19__SCAN_IN ; P3_U6025
g9823 nand P3_U3384 P3_REG2_REG_19__SCAN_IN ; P3_U6026
g9824 nand P3_U5468 P3_REG1_REG_18__SCAN_IN ; P3_U6027
g9825 nand P3_U3384 P3_REG2_REG_18__SCAN_IN ; P3_U6028
g9826 nand P3_U5468 P3_REG1_REG_17__SCAN_IN ; P3_U6029
g9827 nand P3_U3384 P3_REG2_REG_17__SCAN_IN ; P3_U6030
g9828 nand P3_U5468 P3_REG1_REG_16__SCAN_IN ; P3_U6031
g9829 nand P3_U3384 P3_REG2_REG_16__SCAN_IN ; P3_U6032
g9830 nand P3_U5468 P3_REG1_REG_15__SCAN_IN ; P3_U6033
g9831 nand P3_U3384 P3_REG2_REG_15__SCAN_IN ; P3_U6034
g9832 nand P3_U5468 P3_REG1_REG_14__SCAN_IN ; P3_U6035
g9833 nand P3_U3384 P3_REG2_REG_14__SCAN_IN ; P3_U6036
g9834 nand P3_U5468 P3_REG1_REG_13__SCAN_IN ; P3_U6037
g9835 nand P3_U3384 P3_REG2_REG_13__SCAN_IN ; P3_U6038
g9836 nand P3_U5468 P3_REG1_REG_12__SCAN_IN ; P3_U6039
g9837 nand P3_U3384 P3_REG2_REG_12__SCAN_IN ; P3_U6040
g9838 nand P3_U5468 P3_REG1_REG_11__SCAN_IN ; P3_U6041
g9839 nand P3_U3384 P3_REG2_REG_11__SCAN_IN ; P3_U6042
g9840 nand P3_U5468 P3_REG1_REG_10__SCAN_IN ; P3_U6043
g9841 nand P3_U3384 P3_REG2_REG_10__SCAN_IN ; P3_U6044
g9842 nand P3_U5468 P3_REG1_REG_1__SCAN_IN ; P3_U6045
g9843 nand P3_U3384 P3_REG2_REG_1__SCAN_IN ; P3_U6046
g9844 nand P3_U5468 P3_REG1_REG_0__SCAN_IN ; P3_U6047
g9845 nand P3_U3384 P3_REG2_REG_0__SCAN_IN ; P3_U6048
g9846 and SUB_1605_U194 SUB_1605_U190 ; SUB_1605_U6
g9847 and SUB_1605_U202 SUB_1605_U200 ; SUB_1605_U7
g9848 and SUB_1605_U7 SUB_1605_U204 ; SUB_1605_U8
g9849 and SUB_1605_U212 SUB_1605_U208 ; SUB_1605_U9
g9850 and SUB_1605_U9 SUB_1605_U215 ; SUB_1605_U10
g9851 and SUB_1605_U363 SUB_1605_U362 ; SUB_1605_U11
g9852 nand SUB_1605_U128 SUB_1605_U323 ; SUB_1605_U12
g9853 nand SUB_1605_U175 SUB_1605_U291 ; SUB_1605_U13
g9854 not P1_DATAO_REG_8__SCAN_IN ; SUB_1605_U14
g9855 not P2_DATAO_REG_8__SCAN_IN ; SUB_1605_U15
g9856 not P2_DATAO_REG_7__SCAN_IN ; SUB_1605_U16
g9857 not P1_DATAO_REG_6__SCAN_IN ; SUB_1605_U17
g9858 not P1_DATAO_REG_7__SCAN_IN ; SUB_1605_U18
g9859 not P2_DATAO_REG_6__SCAN_IN ; SUB_1605_U19
g9860 not P1_DATAO_REG_5__SCAN_IN ; SUB_1605_U20
g9861 nand SUB_1605_U303 SUB_1605_U204 ; SUB_1605_U21
g9862 not P1_DATAO_REG_4__SCAN_IN ; SUB_1605_U22
g9863 not P2_DATAO_REG_0__SCAN_IN ; SUB_1605_U23
g9864 not P1_DATAO_REG_1__SCAN_IN ; SUB_1605_U24
g9865 not P2_DATAO_REG_4__SCAN_IN ; SUB_1605_U25
g9866 not P2_DATAO_REG_2__SCAN_IN ; SUB_1605_U26
g9867 not P2_DATAO_REG_3__SCAN_IN ; SUB_1605_U27
g9868 not P1_DATAO_REG_2__SCAN_IN ; SUB_1605_U28
g9869 not P1_DATAO_REG_3__SCAN_IN ; SUB_1605_U29
g9870 not P2_DATAO_REG_5__SCAN_IN ; SUB_1605_U30
g9871 not P2_DATAO_REG_9__SCAN_IN ; SUB_1605_U31
g9872 not P1_DATAO_REG_9__SCAN_IN ; SUB_1605_U32
g9873 not P1_DATAO_REG_12__SCAN_IN ; SUB_1605_U33
g9874 not P2_DATAO_REG_12__SCAN_IN ; SUB_1605_U34
g9875 not P2_DATAO_REG_11__SCAN_IN ; SUB_1605_U35
g9876 not P2_DATAO_REG_10__SCAN_IN ; SUB_1605_U36
g9877 not P1_DATAO_REG_11__SCAN_IN ; SUB_1605_U37
g9878 not P1_DATAO_REG_10__SCAN_IN ; SUB_1605_U38
g9879 nand SUB_1605_U31 P1_DATAO_REG_9__SCAN_IN ; SUB_1605_U39
g9880 not P2_DATAO_REG_13__SCAN_IN ; SUB_1605_U40
g9881 not P1_DATAO_REG_13__SCAN_IN ; SUB_1605_U41
g9882 not P2_DATAO_REG_14__SCAN_IN ; SUB_1605_U42
g9883 not P1_DATAO_REG_14__SCAN_IN ; SUB_1605_U43
g9884 not P2_DATAO_REG_15__SCAN_IN ; SUB_1605_U44
g9885 not P1_DATAO_REG_15__SCAN_IN ; SUB_1605_U45
g9886 not P2_DATAO_REG_16__SCAN_IN ; SUB_1605_U46
g9887 not P1_DATAO_REG_16__SCAN_IN ; SUB_1605_U47
g9888 not P2_DATAO_REG_17__SCAN_IN ; SUB_1605_U48
g9889 not P1_DATAO_REG_17__SCAN_IN ; SUB_1605_U49
g9890 not P2_DATAO_REG_18__SCAN_IN ; SUB_1605_U50
g9891 not P1_DATAO_REG_18__SCAN_IN ; SUB_1605_U51
g9892 not P2_DATAO_REG_19__SCAN_IN ; SUB_1605_U52
g9893 not P1_DATAO_REG_19__SCAN_IN ; SUB_1605_U53
g9894 not P2_DATAO_REG_20__SCAN_IN ; SUB_1605_U54
g9895 not P1_DATAO_REG_20__SCAN_IN ; SUB_1605_U55
g9896 not P2_DATAO_REG_21__SCAN_IN ; SUB_1605_U56
g9897 not P1_DATAO_REG_21__SCAN_IN ; SUB_1605_U57
g9898 not P2_DATAO_REG_22__SCAN_IN ; SUB_1605_U58
g9899 not P1_DATAO_REG_22__SCAN_IN ; SUB_1605_U59
g9900 not P2_DATAO_REG_23__SCAN_IN ; SUB_1605_U60
g9901 not P1_DATAO_REG_23__SCAN_IN ; SUB_1605_U61
g9902 not P2_DATAO_REG_24__SCAN_IN ; SUB_1605_U62
g9903 not P1_DATAO_REG_24__SCAN_IN ; SUB_1605_U63
g9904 not P2_DATAO_REG_25__SCAN_IN ; SUB_1605_U64
g9905 not P1_DATAO_REG_25__SCAN_IN ; SUB_1605_U65
g9906 not P2_DATAO_REG_26__SCAN_IN ; SUB_1605_U66
g9907 not P1_DATAO_REG_26__SCAN_IN ; SUB_1605_U67
g9908 not P2_DATAO_REG_27__SCAN_IN ; SUB_1605_U68
g9909 not P1_DATAO_REG_27__SCAN_IN ; SUB_1605_U69
g9910 not P2_DATAO_REG_28__SCAN_IN ; SUB_1605_U70
g9911 not P1_DATAO_REG_28__SCAN_IN ; SUB_1605_U71
g9912 not P2_DATAO_REG_29__SCAN_IN ; SUB_1605_U72
g9913 not P1_DATAO_REG_29__SCAN_IN ; SUB_1605_U73
g9914 not P1_DATAO_REG_30__SCAN_IN ; SUB_1605_U74
g9915 not P2_DATAO_REG_30__SCAN_IN ; SUB_1605_U75
g9916 nand SUB_1605_U308 SUB_1605_U216 ; SUB_1605_U76
g9917 nand SUB_1605_U305 SUB_1605_U213 ; SUB_1605_U77
g9918 not P1_DATAO_REG_0__SCAN_IN ; SUB_1605_U78
g9919 nand SUB_1605_U328 SUB_1605_U327 ; SUB_1605_U79
g9920 nand SUB_1605_U333 SUB_1605_U332 ; SUB_1605_U80
g9921 nand SUB_1605_U338 SUB_1605_U337 ; SUB_1605_U81
g9922 nand SUB_1605_U343 SUB_1605_U342 ; SUB_1605_U82
g9923 nand SUB_1605_U348 SUB_1605_U347 ; SUB_1605_U83
g9924 nand SUB_1605_U353 SUB_1605_U352 ; SUB_1605_U84
g9925 nand SUB_1605_U358 SUB_1605_U357 ; SUB_1605_U85
g9926 nand SUB_1605_U370 SUB_1605_U369 ; SUB_1605_U86
g9927 nand SUB_1605_U375 SUB_1605_U374 ; SUB_1605_U87
g9928 nand SUB_1605_U380 SUB_1605_U379 ; SUB_1605_U88
g9929 nand SUB_1605_U385 SUB_1605_U384 ; SUB_1605_U89
g9930 nand SUB_1605_U390 SUB_1605_U389 ; SUB_1605_U90
g9931 nand SUB_1605_U395 SUB_1605_U394 ; SUB_1605_U91
g9932 nand SUB_1605_U400 SUB_1605_U399 ; SUB_1605_U92
g9933 nand SUB_1605_U405 SUB_1605_U404 ; SUB_1605_U93
g9934 nand SUB_1605_U410 SUB_1605_U409 ; SUB_1605_U94
g9935 nand SUB_1605_U415 SUB_1605_U414 ; SUB_1605_U95
g9936 nand SUB_1605_U420 SUB_1605_U419 ; SUB_1605_U96
g9937 nand SUB_1605_U425 SUB_1605_U424 ; SUB_1605_U97
g9938 nand SUB_1605_U430 SUB_1605_U429 ; SUB_1605_U98
g9939 nand SUB_1605_U435 SUB_1605_U434 ; SUB_1605_U99
g9940 nand SUB_1605_U440 SUB_1605_U439 ; SUB_1605_U100
g9941 nand SUB_1605_U445 SUB_1605_U444 ; SUB_1605_U101
g9942 nand SUB_1605_U450 SUB_1605_U449 ; SUB_1605_U102
g9943 nand SUB_1605_U455 SUB_1605_U454 ; SUB_1605_U103
g9944 nand SUB_1605_U460 SUB_1605_U459 ; SUB_1605_U104
g9945 nand SUB_1605_U465 SUB_1605_U464 ; SUB_1605_U105
g9946 nand SUB_1605_U470 SUB_1605_U469 ; SUB_1605_U106
g9947 nand SUB_1605_U475 SUB_1605_U474 ; SUB_1605_U107
g9948 nand SUB_1605_U480 SUB_1605_U479 ; SUB_1605_U108
g9949 and SUB_1605_U30 P1_DATAO_REG_5__SCAN_IN ; SUB_1605_U109
g9950 and SUB_1605_U205 SUB_1605_U203 ; SUB_1605_U110
g9951 and SUB_1605_U197 SUB_1605_U6 ; SUB_1605_U111
g9952 and SUB_1605_U299 SUB_1605_U197 ; SUB_1605_U112
g9953 and SUB_1605_U298 SUB_1605_U198 ; SUB_1605_U113
g9954 and SUB_1605_U206 SUB_1605_U8 ; SUB_1605_U114
g9955 and SUB_1605_U302 SUB_1605_U207 ; SUB_1605_U115
g9956 nand SUB_1605_U325 SUB_1605_U324 ; SUB_1605_U116
g9957 nand SUB_1605_U330 SUB_1605_U329 ; SUB_1605_U117
g9958 and SUB_1605_U300 SUB_1605_U203 ; SUB_1605_U118
g9959 nand SUB_1605_U335 SUB_1605_U334 ; SUB_1605_U119
g9960 nand SUB_1605_U340 SUB_1605_U339 ; SUB_1605_U120
g9961 nand SUB_1605_U345 SUB_1605_U344 ; SUB_1605_U121
g9962 nand SUB_1605_U350 SUB_1605_U349 ; SUB_1605_U122
g9963 nand SUB_1605_U355 SUB_1605_U354 ; SUB_1605_U123
g9964 and SUB_1605_U10 SUB_1605_U218 ; SUB_1605_U124
g9965 and SUB_1605_U311 SUB_1605_U219 ; SUB_1605_U125
g9966 and SUB_1605_U11 SUB_1605_U290 SUB_1605_U287 ; SUB_1605_U126
g9967 and SUB_1605_U289 SUB_1605_U361 ; SUB_1605_U127
g9968 and SUB_1605_U161 SUB_1605_U293 ; SUB_1605_U128
g9969 nand SUB_1605_U367 SUB_1605_U366 ; SUB_1605_U129
g9970 nand SUB_1605_U372 SUB_1605_U371 ; SUB_1605_U130
g9971 nand SUB_1605_U377 SUB_1605_U376 ; SUB_1605_U131
g9972 nand SUB_1605_U382 SUB_1605_U381 ; SUB_1605_U132
g9973 nand SUB_1605_U387 SUB_1605_U386 ; SUB_1605_U133
g9974 nand SUB_1605_U392 SUB_1605_U391 ; SUB_1605_U134
g9975 nand SUB_1605_U397 SUB_1605_U396 ; SUB_1605_U135
g9976 nand SUB_1605_U402 SUB_1605_U401 ; SUB_1605_U136
g9977 nand SUB_1605_U407 SUB_1605_U406 ; SUB_1605_U137
g9978 nand SUB_1605_U412 SUB_1605_U411 ; SUB_1605_U138
g9979 nand SUB_1605_U417 SUB_1605_U416 ; SUB_1605_U139
g9980 nand SUB_1605_U422 SUB_1605_U421 ; SUB_1605_U140
g9981 nand SUB_1605_U427 SUB_1605_U426 ; SUB_1605_U141
g9982 nand SUB_1605_U432 SUB_1605_U431 ; SUB_1605_U142
g9983 nand SUB_1605_U437 SUB_1605_U436 ; SUB_1605_U143
g9984 nand SUB_1605_U442 SUB_1605_U441 ; SUB_1605_U144
g9985 nand SUB_1605_U447 SUB_1605_U446 ; SUB_1605_U145
g9986 nand SUB_1605_U452 SUB_1605_U451 ; SUB_1605_U146
g9987 nand SUB_1605_U457 SUB_1605_U456 ; SUB_1605_U147
g9988 nand SUB_1605_U462 SUB_1605_U461 ; SUB_1605_U148
g9989 nand SUB_1605_U467 SUB_1605_U466 ; SUB_1605_U149
g9990 nand SUB_1605_U472 SUB_1605_U471 ; SUB_1605_U150
g9991 nand SUB_1605_U477 SUB_1605_U476 ; SUB_1605_U151
g9992 nand SUB_1605_U115 SUB_1605_U321 ; SUB_1605_U152
g9993 nand SUB_1605_U319 SUB_1605_U21 ; SUB_1605_U153
g9994 nand SUB_1605_U118 SUB_1605_U317 ; SUB_1605_U154
g9995 nand SUB_1605_U315 SUB_1605_U201 ; SUB_1605_U155
g9996 nand SUB_1605_U113 SUB_1605_U297 ; SUB_1605_U156
g9997 nand SUB_1605_U296 SUB_1605_U294 ; SUB_1605_U157
g9998 nand SUB_1605_U192 SUB_1605_U191 ; SUB_1605_U158
g9999 not P2_DATAO_REG_31__SCAN_IN ; SUB_1605_U159
g10000 not P1_DATAO_REG_31__SCAN_IN ; SUB_1605_U160
g10001 and SUB_1605_U365 SUB_1605_U364 ; SUB_1605_U161
g10002 nand SUB_1605_U287 SUB_1605_U286 ; SUB_1605_U162
g10003 nand SUB_1605_U188 SUB_1605_U186 SUB_1605_U292 ; SUB_1605_U163
g10004 nand SUB_1605_U283 SUB_1605_U282 ; SUB_1605_U164
g10005 nand SUB_1605_U279 SUB_1605_U278 ; SUB_1605_U165
g10006 nand SUB_1605_U275 SUB_1605_U274 ; SUB_1605_U166
g10007 nand SUB_1605_U271 SUB_1605_U270 ; SUB_1605_U167
g10008 nand SUB_1605_U267 SUB_1605_U266 ; SUB_1605_U168
g10009 nand SUB_1605_U263 SUB_1605_U262 ; SUB_1605_U169
g10010 nand SUB_1605_U259 SUB_1605_U258 ; SUB_1605_U170
g10011 nand SUB_1605_U255 SUB_1605_U254 ; SUB_1605_U171
g10012 nand SUB_1605_U251 SUB_1605_U250 ; SUB_1605_U172
g10013 nand SUB_1605_U247 SUB_1605_U246 ; SUB_1605_U173
g10014 not P2_DATAO_REG_1__SCAN_IN ; SUB_1605_U174
g10015 nand SUB_1605_U78 P2_DATAO_REG_0__SCAN_IN ; SUB_1605_U175
g10016 nand SUB_1605_U243 SUB_1605_U242 ; SUB_1605_U176
g10017 nand SUB_1605_U239 SUB_1605_U238 ; SUB_1605_U177
g10018 nand SUB_1605_U235 SUB_1605_U234 ; SUB_1605_U178
g10019 nand SUB_1605_U231 SUB_1605_U230 ; SUB_1605_U179
g10020 nand SUB_1605_U227 SUB_1605_U226 ; SUB_1605_U180
g10021 nand SUB_1605_U223 SUB_1605_U222 ; SUB_1605_U181
g10022 nand SUB_1605_U125 SUB_1605_U310 ; SUB_1605_U182
g10023 nand SUB_1605_U309 SUB_1605_U307 ; SUB_1605_U183
g10024 nand SUB_1605_U306 SUB_1605_U304 ; SUB_1605_U184
g10025 nand SUB_1605_U39 SUB_1605_U209 ; SUB_1605_U185
g10026 nand SUB_1605_U175 SUB_1605_U174 ; SUB_1605_U186
g10027 not SUB_1605_U175 ; SUB_1605_U187
g10028 nand SUB_1605_U175 P1_DATAO_REG_1__SCAN_IN ; SUB_1605_U188
g10029 not SUB_1605_U163 ; SUB_1605_U189
g10030 nand SUB_1605_U28 P2_DATAO_REG_2__SCAN_IN ; SUB_1605_U190
g10031 nand SUB_1605_U190 SUB_1605_U312 ; SUB_1605_U191
g10032 nand SUB_1605_U26 P1_DATAO_REG_2__SCAN_IN ; SUB_1605_U192
g10033 not SUB_1605_U158 ; SUB_1605_U193
g10034 nand SUB_1605_U29 P2_DATAO_REG_3__SCAN_IN ; SUB_1605_U194
g10035 nand SUB_1605_U27 P1_DATAO_REG_3__SCAN_IN ; SUB_1605_U195
g10036 not SUB_1605_U157 ; SUB_1605_U196
g10037 nand SUB_1605_U22 P2_DATAO_REG_4__SCAN_IN ; SUB_1605_U197
g10038 nand SUB_1605_U25 P1_DATAO_REG_4__SCAN_IN ; SUB_1605_U198
g10039 not SUB_1605_U156 ; SUB_1605_U199
g10040 nand SUB_1605_U20 P2_DATAO_REG_5__SCAN_IN ; SUB_1605_U200
g10041 nand SUB_1605_U30 P1_DATAO_REG_5__SCAN_IN ; SUB_1605_U201
g10042 nand SUB_1605_U17 P2_DATAO_REG_6__SCAN_IN ; SUB_1605_U202
g10043 nand SUB_1605_U19 P1_DATAO_REG_6__SCAN_IN ; SUB_1605_U203
g10044 nand SUB_1605_U18 P2_DATAO_REG_7__SCAN_IN ; SUB_1605_U204
g10045 nand SUB_1605_U16 P1_DATAO_REG_7__SCAN_IN ; SUB_1605_U205
g10046 nand SUB_1605_U14 P2_DATAO_REG_8__SCAN_IN ; SUB_1605_U206
g10047 nand SUB_1605_U15 P1_DATAO_REG_8__SCAN_IN ; SUB_1605_U207
g10048 nand SUB_1605_U32 P2_DATAO_REG_9__SCAN_IN ; SUB_1605_U208
g10049 nand SUB_1605_U208 SUB_1605_U152 ; SUB_1605_U209
g10050 not SUB_1605_U39 ; SUB_1605_U210
g10051 not SUB_1605_U185 ; SUB_1605_U211
g10052 nand SUB_1605_U38 P2_DATAO_REG_10__SCAN_IN ; SUB_1605_U212
g10053 nand SUB_1605_U36 P1_DATAO_REG_10__SCAN_IN ; SUB_1605_U213
g10054 not SUB_1605_U184 ; SUB_1605_U214
g10055 nand SUB_1605_U37 P2_DATAO_REG_11__SCAN_IN ; SUB_1605_U215
g10056 nand SUB_1605_U35 P1_DATAO_REG_11__SCAN_IN ; SUB_1605_U216
g10057 not SUB_1605_U183 ; SUB_1605_U217
g10058 nand SUB_1605_U33 P2_DATAO_REG_12__SCAN_IN ; SUB_1605_U218
g10059 nand SUB_1605_U34 P1_DATAO_REG_12__SCAN_IN ; SUB_1605_U219
g10060 not SUB_1605_U182 ; SUB_1605_U220
g10061 nand SUB_1605_U41 P2_DATAO_REG_13__SCAN_IN ; SUB_1605_U221
g10062 nand SUB_1605_U221 SUB_1605_U182 ; SUB_1605_U222
g10063 nand SUB_1605_U40 P1_DATAO_REG_13__SCAN_IN ; SUB_1605_U223
g10064 not SUB_1605_U181 ; SUB_1605_U224
g10065 nand SUB_1605_U43 P2_DATAO_REG_14__SCAN_IN ; SUB_1605_U225
g10066 nand SUB_1605_U225 SUB_1605_U181 ; SUB_1605_U226
g10067 nand SUB_1605_U42 P1_DATAO_REG_14__SCAN_IN ; SUB_1605_U227
g10068 not SUB_1605_U180 ; SUB_1605_U228
g10069 nand SUB_1605_U45 P2_DATAO_REG_15__SCAN_IN ; SUB_1605_U229
g10070 nand SUB_1605_U229 SUB_1605_U180 ; SUB_1605_U230
g10071 nand SUB_1605_U44 P1_DATAO_REG_15__SCAN_IN ; SUB_1605_U231
g10072 not SUB_1605_U179 ; SUB_1605_U232
g10073 nand SUB_1605_U47 P2_DATAO_REG_16__SCAN_IN ; SUB_1605_U233
g10074 nand SUB_1605_U233 SUB_1605_U179 ; SUB_1605_U234
g10075 nand SUB_1605_U46 P1_DATAO_REG_16__SCAN_IN ; SUB_1605_U235
g10076 not SUB_1605_U178 ; SUB_1605_U236
g10077 nand SUB_1605_U49 P2_DATAO_REG_17__SCAN_IN ; SUB_1605_U237
g10078 nand SUB_1605_U237 SUB_1605_U178 ; SUB_1605_U238
g10079 nand SUB_1605_U48 P1_DATAO_REG_17__SCAN_IN ; SUB_1605_U239
g10080 not SUB_1605_U177 ; SUB_1605_U240
g10081 nand SUB_1605_U51 P2_DATAO_REG_18__SCAN_IN ; SUB_1605_U241
g10082 nand SUB_1605_U241 SUB_1605_U177 ; SUB_1605_U242
g10083 nand SUB_1605_U50 P1_DATAO_REG_18__SCAN_IN ; SUB_1605_U243
g10084 not SUB_1605_U176 ; SUB_1605_U244
g10085 nand SUB_1605_U53 P2_DATAO_REG_19__SCAN_IN ; SUB_1605_U245
g10086 nand SUB_1605_U245 SUB_1605_U176 ; SUB_1605_U246
g10087 nand SUB_1605_U52 P1_DATAO_REG_19__SCAN_IN ; SUB_1605_U247
g10088 not SUB_1605_U173 ; SUB_1605_U248
g10089 nand SUB_1605_U55 P2_DATAO_REG_20__SCAN_IN ; SUB_1605_U249
g10090 nand SUB_1605_U249 SUB_1605_U173 ; SUB_1605_U250
g10091 nand SUB_1605_U54 P1_DATAO_REG_20__SCAN_IN ; SUB_1605_U251
g10092 not SUB_1605_U172 ; SUB_1605_U252
g10093 nand SUB_1605_U57 P2_DATAO_REG_21__SCAN_IN ; SUB_1605_U253
g10094 nand SUB_1605_U253 SUB_1605_U172 ; SUB_1605_U254
g10095 nand SUB_1605_U56 P1_DATAO_REG_21__SCAN_IN ; SUB_1605_U255
g10096 not SUB_1605_U171 ; SUB_1605_U256
g10097 nand SUB_1605_U59 P2_DATAO_REG_22__SCAN_IN ; SUB_1605_U257
g10098 nand SUB_1605_U257 SUB_1605_U171 ; SUB_1605_U258
g10099 nand SUB_1605_U58 P1_DATAO_REG_22__SCAN_IN ; SUB_1605_U259
g10100 not SUB_1605_U170 ; SUB_1605_U260
g10101 nand SUB_1605_U61 P2_DATAO_REG_23__SCAN_IN ; SUB_1605_U261
g10102 nand SUB_1605_U261 SUB_1605_U170 ; SUB_1605_U262
g10103 nand SUB_1605_U60 P1_DATAO_REG_23__SCAN_IN ; SUB_1605_U263
g10104 not SUB_1605_U169 ; SUB_1605_U264
g10105 nand SUB_1605_U63 P2_DATAO_REG_24__SCAN_IN ; SUB_1605_U265
g10106 nand SUB_1605_U265 SUB_1605_U169 ; SUB_1605_U266
g10107 nand SUB_1605_U62 P1_DATAO_REG_24__SCAN_IN ; SUB_1605_U267
g10108 not SUB_1605_U168 ; SUB_1605_U268
g10109 nand SUB_1605_U65 P2_DATAO_REG_25__SCAN_IN ; SUB_1605_U269
g10110 nand SUB_1605_U269 SUB_1605_U168 ; SUB_1605_U270
g10111 nand SUB_1605_U64 P1_DATAO_REG_25__SCAN_IN ; SUB_1605_U271
g10112 not SUB_1605_U167 ; SUB_1605_U272
g10113 nand SUB_1605_U67 P2_DATAO_REG_26__SCAN_IN ; SUB_1605_U273
g10114 nand SUB_1605_U273 SUB_1605_U167 ; SUB_1605_U274
g10115 nand SUB_1605_U66 P1_DATAO_REG_26__SCAN_IN ; SUB_1605_U275
g10116 not SUB_1605_U166 ; SUB_1605_U276
g10117 nand SUB_1605_U69 P2_DATAO_REG_27__SCAN_IN ; SUB_1605_U277
g10118 nand SUB_1605_U277 SUB_1605_U166 ; SUB_1605_U278
g10119 nand SUB_1605_U68 P1_DATAO_REG_27__SCAN_IN ; SUB_1605_U279
g10120 not SUB_1605_U165 ; SUB_1605_U280
g10121 nand SUB_1605_U71 P2_DATAO_REG_28__SCAN_IN ; SUB_1605_U281
g10122 nand SUB_1605_U281 SUB_1605_U165 ; SUB_1605_U282
g10123 nand SUB_1605_U70 P1_DATAO_REG_28__SCAN_IN ; SUB_1605_U283
g10124 not SUB_1605_U164 ; SUB_1605_U284
g10125 nand SUB_1605_U73 P2_DATAO_REG_29__SCAN_IN ; SUB_1605_U285
g10126 nand SUB_1605_U285 SUB_1605_U164 ; SUB_1605_U286
g10127 nand SUB_1605_U72 P1_DATAO_REG_29__SCAN_IN ; SUB_1605_U287
g10128 not SUB_1605_U162 ; SUB_1605_U288
g10129 nand SUB_1605_U74 P2_DATAO_REG_30__SCAN_IN ; SUB_1605_U289
g10130 nand SUB_1605_U75 P1_DATAO_REG_30__SCAN_IN ; SUB_1605_U290
g10131 nand SUB_1605_U23 P1_DATAO_REG_0__SCAN_IN ; SUB_1605_U291
g10132 nand SUB_1605_U174 P1_DATAO_REG_1__SCAN_IN ; SUB_1605_U292
g10133 nand SUB_1605_U286 SUB_1605_U126 ; SUB_1605_U293
g10134 nand SUB_1605_U6 SUB_1605_U163 ; SUB_1605_U294
g10135 nand SUB_1605_U195 SUB_1605_U192 ; SUB_1605_U295
g10136 nand SUB_1605_U295 SUB_1605_U299 ; SUB_1605_U296
g10137 nand SUB_1605_U111 SUB_1605_U163 ; SUB_1605_U297
g10138 nand SUB_1605_U112 SUB_1605_U295 ; SUB_1605_U298
g10139 nand SUB_1605_U29 P2_DATAO_REG_3__SCAN_IN ; SUB_1605_U299
g10140 nand SUB_1605_U109 SUB_1605_U202 ; SUB_1605_U300
g10141 not SUB_1605_U21 ; SUB_1605_U301
g10142 nand SUB_1605_U301 SUB_1605_U206 ; SUB_1605_U302
g10143 nand SUB_1605_U110 SUB_1605_U300 ; SUB_1605_U303
g10144 nand SUB_1605_U9 SUB_1605_U152 ; SUB_1605_U304
g10145 nand SUB_1605_U210 SUB_1605_U212 ; SUB_1605_U305
g10146 not SUB_1605_U77 ; SUB_1605_U306
g10147 nand SUB_1605_U10 SUB_1605_U152 ; SUB_1605_U307
g10148 nand SUB_1605_U77 SUB_1605_U215 ; SUB_1605_U308
g10149 not SUB_1605_U76 ; SUB_1605_U309
g10150 nand SUB_1605_U124 SUB_1605_U152 ; SUB_1605_U310
g10151 nand SUB_1605_U76 SUB_1605_U218 ; SUB_1605_U311
g10152 nand SUB_1605_U313 SUB_1605_U292 SUB_1605_U314 ; SUB_1605_U312
g10153 nand SUB_1605_U175 P1_DATAO_REG_1__SCAN_IN ; SUB_1605_U313
g10154 nand SUB_1605_U175 SUB_1605_U174 ; SUB_1605_U314
g10155 nand SUB_1605_U200 SUB_1605_U156 ; SUB_1605_U315
g10156 not SUB_1605_U155 ; SUB_1605_U316
g10157 nand SUB_1605_U7 SUB_1605_U156 ; SUB_1605_U317
g10158 not SUB_1605_U154 ; SUB_1605_U318
g10159 nand SUB_1605_U8 SUB_1605_U156 ; SUB_1605_U319
g10160 not SUB_1605_U153 ; SUB_1605_U320
g10161 nand SUB_1605_U114 SUB_1605_U156 ; SUB_1605_U321
g10162 not SUB_1605_U152 ; SUB_1605_U322
g10163 nand SUB_1605_U127 SUB_1605_U162 ; SUB_1605_U323
g10164 nand SUB_1605_U32 P2_DATAO_REG_9__SCAN_IN ; SUB_1605_U324
g10165 nand SUB_1605_U31 P1_DATAO_REG_9__SCAN_IN ; SUB_1605_U325
g10166 not SUB_1605_U116 ; SUB_1605_U326
g10167 nand SUB_1605_U322 SUB_1605_U326 ; SUB_1605_U327
g10168 nand SUB_1605_U116 SUB_1605_U152 ; SUB_1605_U328
g10169 nand SUB_1605_U14 P2_DATAO_REG_8__SCAN_IN ; SUB_1605_U329
g10170 nand SUB_1605_U15 P1_DATAO_REG_8__SCAN_IN ; SUB_1605_U330
g10171 not SUB_1605_U117 ; SUB_1605_U331
g10172 nand SUB_1605_U320 SUB_1605_U331 ; SUB_1605_U332
g10173 nand SUB_1605_U117 SUB_1605_U153 ; SUB_1605_U333
g10174 nand SUB_1605_U18 P2_DATAO_REG_7__SCAN_IN ; SUB_1605_U334
g10175 nand SUB_1605_U16 P1_DATAO_REG_7__SCAN_IN ; SUB_1605_U335
g10176 not SUB_1605_U119 ; SUB_1605_U336
g10177 nand SUB_1605_U318 SUB_1605_U336 ; SUB_1605_U337
g10178 nand SUB_1605_U119 SUB_1605_U154 ; SUB_1605_U338
g10179 nand SUB_1605_U17 P2_DATAO_REG_6__SCAN_IN ; SUB_1605_U339
g10180 nand SUB_1605_U19 P1_DATAO_REG_6__SCAN_IN ; SUB_1605_U340
g10181 not SUB_1605_U120 ; SUB_1605_U341
g10182 nand SUB_1605_U316 SUB_1605_U341 ; SUB_1605_U342
g10183 nand SUB_1605_U120 SUB_1605_U155 ; SUB_1605_U343
g10184 nand SUB_1605_U20 P2_DATAO_REG_5__SCAN_IN ; SUB_1605_U344
g10185 nand SUB_1605_U30 P1_DATAO_REG_5__SCAN_IN ; SUB_1605_U345
g10186 not SUB_1605_U121 ; SUB_1605_U346
g10187 nand SUB_1605_U199 SUB_1605_U346 ; SUB_1605_U347
g10188 nand SUB_1605_U121 SUB_1605_U156 ; SUB_1605_U348
g10189 nand SUB_1605_U22 P2_DATAO_REG_4__SCAN_IN ; SUB_1605_U349
g10190 nand SUB_1605_U25 P1_DATAO_REG_4__SCAN_IN ; SUB_1605_U350
g10191 not SUB_1605_U122 ; SUB_1605_U351
g10192 nand SUB_1605_U196 SUB_1605_U351 ; SUB_1605_U352
g10193 nand SUB_1605_U122 SUB_1605_U157 ; SUB_1605_U353
g10194 nand SUB_1605_U29 P2_DATAO_REG_3__SCAN_IN ; SUB_1605_U354
g10195 nand SUB_1605_U27 P1_DATAO_REG_3__SCAN_IN ; SUB_1605_U355
g10196 not SUB_1605_U123 ; SUB_1605_U356
g10197 nand SUB_1605_U193 SUB_1605_U356 ; SUB_1605_U357
g10198 nand SUB_1605_U123 SUB_1605_U158 ; SUB_1605_U358
g10199 nand SUB_1605_U160 P2_DATAO_REG_31__SCAN_IN ; SUB_1605_U359
g10200 nand SUB_1605_U159 P1_DATAO_REG_31__SCAN_IN ; SUB_1605_U360
g10201 nand SUB_1605_U360 SUB_1605_U359 ; SUB_1605_U361
g10202 nand SUB_1605_U160 P2_DATAO_REG_31__SCAN_IN ; SUB_1605_U362
g10203 nand SUB_1605_U159 P1_DATAO_REG_31__SCAN_IN ; SUB_1605_U363
g10204 nand SUB_1605_U361 SUB_1605_U75 P1_DATAO_REG_30__SCAN_IN ; SUB_1605_U364
g10205 nand SUB_1605_U11 SUB_1605_U74 P2_DATAO_REG_30__SCAN_IN ; SUB_1605_U365
g10206 nand SUB_1605_U74 P2_DATAO_REG_30__SCAN_IN ; SUB_1605_U366
g10207 nand SUB_1605_U75 P1_DATAO_REG_30__SCAN_IN ; SUB_1605_U367
g10208 not SUB_1605_U129 ; SUB_1605_U368
g10209 nand SUB_1605_U288 SUB_1605_U368 ; SUB_1605_U369
g10210 nand SUB_1605_U129 SUB_1605_U162 ; SUB_1605_U370
g10211 nand SUB_1605_U28 P2_DATAO_REG_2__SCAN_IN ; SUB_1605_U371
g10212 nand SUB_1605_U26 P1_DATAO_REG_2__SCAN_IN ; SUB_1605_U372
g10213 not SUB_1605_U130 ; SUB_1605_U373
g10214 nand SUB_1605_U189 SUB_1605_U373 ; SUB_1605_U374
g10215 nand SUB_1605_U130 SUB_1605_U163 ; SUB_1605_U375
g10216 nand SUB_1605_U73 P2_DATAO_REG_29__SCAN_IN ; SUB_1605_U376
g10217 nand SUB_1605_U72 P1_DATAO_REG_29__SCAN_IN ; SUB_1605_U377
g10218 not SUB_1605_U131 ; SUB_1605_U378
g10219 nand SUB_1605_U284 SUB_1605_U378 ; SUB_1605_U379
g10220 nand SUB_1605_U131 SUB_1605_U164 ; SUB_1605_U380
g10221 nand SUB_1605_U71 P2_DATAO_REG_28__SCAN_IN ; SUB_1605_U381
g10222 nand SUB_1605_U70 P1_DATAO_REG_28__SCAN_IN ; SUB_1605_U382
g10223 not SUB_1605_U132 ; SUB_1605_U383
g10224 nand SUB_1605_U280 SUB_1605_U383 ; SUB_1605_U384
g10225 nand SUB_1605_U132 SUB_1605_U165 ; SUB_1605_U385
g10226 nand SUB_1605_U69 P2_DATAO_REG_27__SCAN_IN ; SUB_1605_U386
g10227 nand SUB_1605_U68 P1_DATAO_REG_27__SCAN_IN ; SUB_1605_U387
g10228 not SUB_1605_U133 ; SUB_1605_U388
g10229 nand SUB_1605_U276 SUB_1605_U388 ; SUB_1605_U389
g10230 nand SUB_1605_U133 SUB_1605_U166 ; SUB_1605_U390
g10231 nand SUB_1605_U67 P2_DATAO_REG_26__SCAN_IN ; SUB_1605_U391
g10232 nand SUB_1605_U66 P1_DATAO_REG_26__SCAN_IN ; SUB_1605_U392
g10233 not SUB_1605_U134 ; SUB_1605_U393
g10234 nand SUB_1605_U272 SUB_1605_U393 ; SUB_1605_U394
g10235 nand SUB_1605_U134 SUB_1605_U167 ; SUB_1605_U395
g10236 nand SUB_1605_U65 P2_DATAO_REG_25__SCAN_IN ; SUB_1605_U396
g10237 nand SUB_1605_U64 P1_DATAO_REG_25__SCAN_IN ; SUB_1605_U397
g10238 not SUB_1605_U135 ; SUB_1605_U398
g10239 nand SUB_1605_U268 SUB_1605_U398 ; SUB_1605_U399
g10240 nand SUB_1605_U135 SUB_1605_U168 ; SUB_1605_U400
g10241 nand SUB_1605_U63 P2_DATAO_REG_24__SCAN_IN ; SUB_1605_U401
g10242 nand SUB_1605_U62 P1_DATAO_REG_24__SCAN_IN ; SUB_1605_U402
g10243 not SUB_1605_U136 ; SUB_1605_U403
g10244 nand SUB_1605_U264 SUB_1605_U403 ; SUB_1605_U404
g10245 nand SUB_1605_U136 SUB_1605_U169 ; SUB_1605_U405
g10246 nand SUB_1605_U61 P2_DATAO_REG_23__SCAN_IN ; SUB_1605_U406
g10247 nand SUB_1605_U60 P1_DATAO_REG_23__SCAN_IN ; SUB_1605_U407
g10248 not SUB_1605_U137 ; SUB_1605_U408
g10249 nand SUB_1605_U260 SUB_1605_U408 ; SUB_1605_U409
g10250 nand SUB_1605_U137 SUB_1605_U170 ; SUB_1605_U410
g10251 nand SUB_1605_U59 P2_DATAO_REG_22__SCAN_IN ; SUB_1605_U411
g10252 nand SUB_1605_U58 P1_DATAO_REG_22__SCAN_IN ; SUB_1605_U412
g10253 not SUB_1605_U138 ; SUB_1605_U413
g10254 nand SUB_1605_U256 SUB_1605_U413 ; SUB_1605_U414
g10255 nand SUB_1605_U138 SUB_1605_U171 ; SUB_1605_U415
g10256 nand SUB_1605_U57 P2_DATAO_REG_21__SCAN_IN ; SUB_1605_U416
g10257 nand SUB_1605_U56 P1_DATAO_REG_21__SCAN_IN ; SUB_1605_U417
g10258 not SUB_1605_U139 ; SUB_1605_U418
g10259 nand SUB_1605_U252 SUB_1605_U418 ; SUB_1605_U419
g10260 nand SUB_1605_U139 SUB_1605_U172 ; SUB_1605_U420
g10261 nand SUB_1605_U55 P2_DATAO_REG_20__SCAN_IN ; SUB_1605_U421
g10262 nand SUB_1605_U54 P1_DATAO_REG_20__SCAN_IN ; SUB_1605_U422
g10263 not SUB_1605_U140 ; SUB_1605_U423
g10264 nand SUB_1605_U248 SUB_1605_U423 ; SUB_1605_U424
g10265 nand SUB_1605_U140 SUB_1605_U173 ; SUB_1605_U425
g10266 nand SUB_1605_U24 P2_DATAO_REG_1__SCAN_IN ; SUB_1605_U426
g10267 nand SUB_1605_U174 P1_DATAO_REG_1__SCAN_IN ; SUB_1605_U427
g10268 not SUB_1605_U141 ; SUB_1605_U428
g10269 nand SUB_1605_U187 SUB_1605_U428 ; SUB_1605_U429
g10270 nand SUB_1605_U141 SUB_1605_U175 ; SUB_1605_U430
g10271 nand SUB_1605_U53 P2_DATAO_REG_19__SCAN_IN ; SUB_1605_U431
g10272 nand SUB_1605_U52 P1_DATAO_REG_19__SCAN_IN ; SUB_1605_U432
g10273 not SUB_1605_U142 ; SUB_1605_U433
g10274 nand SUB_1605_U244 SUB_1605_U433 ; SUB_1605_U434
g10275 nand SUB_1605_U142 SUB_1605_U176 ; SUB_1605_U435
g10276 nand SUB_1605_U51 P2_DATAO_REG_18__SCAN_IN ; SUB_1605_U436
g10277 nand SUB_1605_U50 P1_DATAO_REG_18__SCAN_IN ; SUB_1605_U437
g10278 not SUB_1605_U143 ; SUB_1605_U438
g10279 nand SUB_1605_U240 SUB_1605_U438 ; SUB_1605_U439
g10280 nand SUB_1605_U143 SUB_1605_U177 ; SUB_1605_U440
g10281 nand SUB_1605_U49 P2_DATAO_REG_17__SCAN_IN ; SUB_1605_U441
g10282 nand SUB_1605_U48 P1_DATAO_REG_17__SCAN_IN ; SUB_1605_U442
g10283 not SUB_1605_U144 ; SUB_1605_U443
g10284 nand SUB_1605_U236 SUB_1605_U443 ; SUB_1605_U444
g10285 nand SUB_1605_U144 SUB_1605_U178 ; SUB_1605_U445
g10286 nand SUB_1605_U47 P2_DATAO_REG_16__SCAN_IN ; SUB_1605_U446
g10287 nand SUB_1605_U46 P1_DATAO_REG_16__SCAN_IN ; SUB_1605_U447
g10288 not SUB_1605_U145 ; SUB_1605_U448
g10289 nand SUB_1605_U232 SUB_1605_U448 ; SUB_1605_U449
g10290 nand SUB_1605_U145 SUB_1605_U179 ; SUB_1605_U450
g10291 nand SUB_1605_U45 P2_DATAO_REG_15__SCAN_IN ; SUB_1605_U451
g10292 nand SUB_1605_U44 P1_DATAO_REG_15__SCAN_IN ; SUB_1605_U452
g10293 not SUB_1605_U146 ; SUB_1605_U453
g10294 nand SUB_1605_U228 SUB_1605_U453 ; SUB_1605_U454
g10295 nand SUB_1605_U146 SUB_1605_U180 ; SUB_1605_U455
g10296 nand SUB_1605_U43 P2_DATAO_REG_14__SCAN_IN ; SUB_1605_U456
g10297 nand SUB_1605_U42 P1_DATAO_REG_14__SCAN_IN ; SUB_1605_U457
g10298 not SUB_1605_U147 ; SUB_1605_U458
g10299 nand SUB_1605_U224 SUB_1605_U458 ; SUB_1605_U459
g10300 nand SUB_1605_U147 SUB_1605_U181 ; SUB_1605_U460
g10301 nand SUB_1605_U41 P2_DATAO_REG_13__SCAN_IN ; SUB_1605_U461
g10302 nand SUB_1605_U40 P1_DATAO_REG_13__SCAN_IN ; SUB_1605_U462
g10303 not SUB_1605_U148 ; SUB_1605_U463
g10304 nand SUB_1605_U220 SUB_1605_U463 ; SUB_1605_U464
g10305 nand SUB_1605_U148 SUB_1605_U182 ; SUB_1605_U465
g10306 nand SUB_1605_U33 P2_DATAO_REG_12__SCAN_IN ; SUB_1605_U466
g10307 nand SUB_1605_U34 P1_DATAO_REG_12__SCAN_IN ; SUB_1605_U467
g10308 not SUB_1605_U149 ; SUB_1605_U468
g10309 nand SUB_1605_U217 SUB_1605_U468 ; SUB_1605_U469
g10310 nand SUB_1605_U149 SUB_1605_U183 ; SUB_1605_U470
g10311 nand SUB_1605_U37 P2_DATAO_REG_11__SCAN_IN ; SUB_1605_U471
g10312 nand SUB_1605_U35 P1_DATAO_REG_11__SCAN_IN ; SUB_1605_U472
g10313 not SUB_1605_U150 ; SUB_1605_U473
g10314 nand SUB_1605_U214 SUB_1605_U473 ; SUB_1605_U474
g10315 nand SUB_1605_U150 SUB_1605_U184 ; SUB_1605_U475
g10316 nand SUB_1605_U38 P2_DATAO_REG_10__SCAN_IN ; SUB_1605_U476
g10317 nand SUB_1605_U36 P1_DATAO_REG_10__SCAN_IN ; SUB_1605_U477
g10318 not SUB_1605_U151 ; SUB_1605_U478
g10319 nand SUB_1605_U211 SUB_1605_U478 ; SUB_1605_U479
g10320 nand SUB_1605_U151 SUB_1605_U185 ; SUB_1605_U480
g10321 and R152_U206 R152_U202 ; R152_U4
g10322 and R152_U214 R152_U212 ; R152_U5
g10323 and R152_U5 R152_U216 ; R152_U6
g10324 and R152_U222 R152_U220 ; R152_U7
g10325 and R152_U7 R152_U224 ; R152_U8
g10326 and R152_U8 R152_U226 ; R152_U9
g10327 and R152_U199 R152_U196 ; R152_U10
g10328 and R152_U391 R152_U390 ; R152_U11
g10329 and R152_U128 R152_U193 ; R152_U12
g10330 nand R152_U172 R152_U337 ; R152_U13
g10331 not SI_8_ ; R152_U14
g10332 not U127 ; R152_U15
g10333 not SI_7_ ; R152_U16
g10334 not U128 ; R152_U17
g10335 nand U128 SI_7_ ; R152_U18
g10336 not SI_6_ ; R152_U19
g10337 not U129 ; R152_U20
g10338 not SI_3_ ; R152_U21
g10339 not U134 ; R152_U22
g10340 not SI_1_ ; R152_U23
g10341 not SI_0_ ; R152_U24
g10342 not U157 ; R152_U25
g10343 not U156 ; R152_U26
g10344 not SI_2_ ; R152_U27
g10345 not U145 ; R152_U28
g10346 nand U145 SI_2_ ; R152_U29
g10347 not SI_5_ ; R152_U30
g10348 not U130 ; R152_U31
g10349 not SI_4_ ; R152_U32
g10350 not U131 ; R152_U33
g10351 nand U131 SI_4_ ; R152_U34
g10352 not U126 ; R152_U35
g10353 not SI_9_ ; R152_U36
g10354 nand R152_U294 R152_U207 ; R152_U37
g10355 not SI_15_ ; R152_U38
g10356 not U150 ; R152_U39
g10357 not SI_14_ ; R152_U40
g10358 not U151 ; R152_U41
g10359 not SI_13_ ; R152_U42
g10360 not U152 ; R152_U43
g10361 not SI_12_ ; R152_U44
g10362 not U153 ; R152_U45
g10363 not SI_11_ ; R152_U46
g10364 not U154 ; R152_U47
g10365 nand U154 SI_11_ ; R152_U48
g10366 not SI_10_ ; R152_U49
g10367 not U155 ; R152_U50
g10368 not SI_16_ ; R152_U51
g10369 not U149 ; R152_U52
g10370 not SI_17_ ; R152_U53
g10371 not U148 ; R152_U54
g10372 not SI_18_ ; R152_U55
g10373 not U147 ; R152_U56
g10374 not SI_19_ ; R152_U57
g10375 not U146 ; R152_U58
g10376 not SI_20_ ; R152_U59
g10377 not U144 ; R152_U60
g10378 not SI_21_ ; R152_U61
g10379 not U143 ; R152_U62
g10380 not SI_22_ ; R152_U63
g10381 not U142 ; R152_U64
g10382 not SI_23_ ; R152_U65
g10383 not U141 ; R152_U66
g10384 not SI_24_ ; R152_U67
g10385 not U140 ; R152_U68
g10386 not SI_25_ ; R152_U69
g10387 not U139 ; R152_U70
g10388 not SI_26_ ; R152_U71
g10389 not U138 ; R152_U72
g10390 not SI_27_ ; R152_U73
g10391 not U137 ; R152_U74
g10392 not SI_28_ ; R152_U75
g10393 not U136 ; R152_U76
g10394 not SI_29_ ; R152_U77
g10395 not U135 ; R152_U78
g10396 not SI_30_ ; R152_U79
g10397 not U133 ; R152_U80
g10398 nand R152_U307 R152_U227 ; R152_U81
g10399 nand R152_U305 R152_U225 ; R152_U82
g10400 nand R152_U300 R152_U217 ; R152_U83
g10401 nand R152_U554 R152_U553 ; R152_U84
g10402 nand R152_U344 R152_U343 ; R152_U85
g10403 nand R152_U351 R152_U350 ; R152_U86
g10404 nand R152_U358 R152_U357 ; R152_U87
g10405 nand R152_U365 R152_U364 ; R152_U88
g10406 nand R152_U372 R152_U371 ; R152_U89
g10407 nand R152_U379 R152_U378 ; R152_U90
g10408 nand R152_U386 R152_U385 ; R152_U91
g10409 nand R152_U400 R152_U399 ; R152_U92
g10410 nand R152_U407 R152_U406 ; R152_U93
g10411 nand R152_U414 R152_U413 ; R152_U94
g10412 nand R152_U421 R152_U420 ; R152_U95
g10413 nand R152_U428 R152_U427 ; R152_U96
g10414 nand R152_U435 R152_U434 ; R152_U97
g10415 nand R152_U442 R152_U441 ; R152_U98
g10416 nand R152_U449 R152_U448 ; R152_U99
g10417 nand R152_U456 R152_U455 ; R152_U100
g10418 nand R152_U463 R152_U462 ; R152_U101
g10419 nand R152_U470 R152_U469 ; R152_U102
g10420 nand R152_U477 R152_U476 ; R152_U103
g10421 nand R152_U489 R152_U488 ; R152_U104
g10422 nand R152_U496 R152_U495 ; R152_U105
g10423 nand R152_U503 R152_U502 ; R152_U106
g10424 nand R152_U510 R152_U509 ; R152_U107
g10425 nand R152_U517 R152_U516 ; R152_U108
g10426 nand R152_U524 R152_U523 ; R152_U109
g10427 nand R152_U531 R152_U530 ; R152_U110
g10428 nand R152_U538 R152_U537 ; R152_U111
g10429 nand R152_U545 R152_U544 ; R152_U112
g10430 nand R152_U552 R152_U551 ; R152_U113
g10431 and R152_U292 R152_U200 ; R152_U114
g10432 and R152_U209 R152_U4 ; R152_U115
g10433 and R152_U297 R152_U210 ; R152_U116
g10434 and R152_U298 R152_U215 ; R152_U117
g10435 and R152_U292 R152_U200 ; R152_U118
g10436 and U156 U157 ; R152_U119
g10437 and U157 SI_0_ ; R152_U120
g10438 and SI_1_ U156 ; R152_U121
g10439 and R152_U218 R152_U6 ; R152_U122
g10440 and R152_U302 R152_U219 ; R152_U123
g10441 and R152_U9 R152_U228 ; R152_U124
g10442 and R152_U309 R152_U229 ; R152_U125
g10443 and R152_U287 R152_U389 ; R152_U126
g10444 and R152_U11 R152_U286 R152_U284 ; R152_U127
g10445 and R152_U288 R152_U146 ; R152_U128
g10446 and R152_U303 R152_U223 ; R152_U129
g10447 and R152_U339 R152_U338 ; R152_U130
g10448 nand R152_U117 R152_U331 ; R152_U131
g10449 and R152_U346 R152_U345 ; R152_U132
g10450 nand R152_U329 R152_U18 ; R152_U133
g10451 and R152_U353 R152_U352 ; R152_U134
g10452 nand R152_U116 R152_U296 ; R152_U135
g10453 and R152_U360 R152_U359 ; R152_U136
g10454 nand R152_U295 R152_U293 ; R152_U137
g10455 and R152_U367 R152_U366 ; R152_U138
g10456 nand R152_U34 R152_U203 ; R152_U139
g10457 and R152_U374 R152_U373 ; R152_U140
g10458 nand R152_U118 R152_U315 ; R152_U141
g10459 and R152_U381 R152_U380 ; R152_U142
g10460 nand R152_U312 R152_U311 R152_U310 R152_U29 ; R152_U143
g10461 not U132 ; R152_U144
g10462 not SI_31_ ; R152_U145
g10463 and R152_U393 R152_U392 ; R152_U146
g10464 and R152_U395 R152_U394 ; R152_U147
g10465 nand R152_U284 R152_U283 ; R152_U148
g10466 nand R152_U290 R152_U171 R152_U289 ; R152_U149
g10467 and R152_U409 R152_U408 ; R152_U150
g10468 nand R152_U280 R152_U279 ; R152_U151
g10469 and R152_U416 R152_U415 ; R152_U152
g10470 nand R152_U276 R152_U275 ; R152_U153
g10471 and R152_U423 R152_U422 ; R152_U154
g10472 nand R152_U272 R152_U271 ; R152_U155
g10473 and R152_U430 R152_U429 ; R152_U156
g10474 nand R152_U268 R152_U267 ; R152_U157
g10475 and R152_U437 R152_U436 ; R152_U158
g10476 nand R152_U264 R152_U263 ; R152_U159
g10477 and R152_U444 R152_U443 ; R152_U160
g10478 nand R152_U260 R152_U259 ; R152_U161
g10479 and R152_U451 R152_U450 ; R152_U162
g10480 nand R152_U256 R152_U255 ; R152_U163
g10481 and R152_U458 R152_U457 ; R152_U164
g10482 nand R152_U252 R152_U251 ; R152_U165
g10483 and R152_U465 R152_U464 ; R152_U166
g10484 nand R152_U248 R152_U247 ; R152_U167
g10485 and R152_U472 R152_U471 ; R152_U168
g10486 nand R152_U244 R152_U243 ; R152_U169
g10487 nand U157 SI_0_ ; R152_U170
g10488 nand SI_0_ SI_1_ U157 ; R152_U171
g10489 and R152_U482 R152_U481 ; R152_U172
g10490 and R152_U484 R152_U483 ; R152_U173
g10491 nand R152_U240 R152_U239 ; R152_U174
g10492 and R152_U491 R152_U490 ; R152_U175
g10493 nand R152_U236 R152_U235 ; R152_U176
g10494 and R152_U498 R152_U497 ; R152_U177
g10495 nand R152_U232 R152_U231 ; R152_U178
g10496 and R152_U505 R152_U504 ; R152_U179
g10497 nand R152_U125 R152_U327 ; R152_U180
g10498 and R152_U512 R152_U511 ; R152_U181
g10499 nand R152_U308 R152_U325 ; R152_U182
g10500 and R152_U519 R152_U518 ; R152_U183
g10501 nand R152_U306 R152_U323 ; R152_U184
g10502 and R152_U526 R152_U525 ; R152_U185
g10503 nand R152_U129 R152_U321 ; R152_U186
g10504 and R152_U533 R152_U532 ; R152_U187
g10505 nand R152_U319 R152_U48 ; R152_U188
g10506 and R152_U540 R152_U539 ; R152_U189
g10507 nand R152_U123 R152_U335 ; R152_U190
g10508 and R152_U547 R152_U546 ; R152_U191
g10509 nand R152_U301 R152_U333 ; R152_U192
g10510 nand R152_U126 R152_U148 ; R152_U193
g10511 not R152_U171 ; R152_U194
g10512 not R152_U149 ; R152_U195
g10513 or SI_2_ U145 ; R152_U196
g10514 not R152_U29 ; R152_U197
g10515 not R152_U143 ; R152_U198
g10516 or SI_3_ U134 ; R152_U199
g10517 nand U134 SI_3_ ; R152_U200
g10518 nand R152_U114 R152_U291 ; R152_U201
g10519 or SI_4_ U131 ; R152_U202
g10520 nand R152_U202 R152_U201 ; R152_U203
g10521 not R152_U34 ; R152_U204
g10522 not R152_U139 ; R152_U205
g10523 or SI_5_ U130 ; R152_U206
g10524 nand U130 SI_5_ ; R152_U207
g10525 not R152_U137 ; R152_U208
g10526 or SI_6_ U129 ; R152_U209
g10527 nand U129 SI_6_ ; R152_U210
g10528 not R152_U135 ; R152_U211
g10529 or SI_7_ U128 ; R152_U212
g10530 not R152_U18 ; R152_U213
g10531 or SI_8_ U127 ; R152_U214
g10532 nand U127 SI_8_ ; R152_U215
g10533 or SI_9_ U126 ; R152_U216
g10534 nand SI_9_ U126 ; R152_U217
g10535 or SI_10_ U155 ; R152_U218
g10536 nand U155 SI_10_ ; R152_U219
g10537 or SI_11_ U154 ; R152_U220
g10538 not R152_U48 ; R152_U221
g10539 or SI_12_ U153 ; R152_U222
g10540 nand U153 SI_12_ ; R152_U223
g10541 or SI_13_ U152 ; R152_U224
g10542 nand U152 SI_13_ ; R152_U225
g10543 or SI_14_ U151 ; R152_U226
g10544 nand U151 SI_14_ ; R152_U227
g10545 or SI_15_ U150 ; R152_U228
g10546 nand U150 SI_15_ ; R152_U229
g10547 or SI_16_ U149 ; R152_U230
g10548 nand R152_U230 R152_U180 ; R152_U231
g10549 nand U149 SI_16_ ; R152_U232
g10550 not R152_U178 ; R152_U233
g10551 or SI_17_ U148 ; R152_U234
g10552 nand R152_U234 R152_U178 ; R152_U235
g10553 nand U148 SI_17_ ; R152_U236
g10554 not R152_U176 ; R152_U237
g10555 or SI_18_ U147 ; R152_U238
g10556 nand R152_U238 R152_U176 ; R152_U239
g10557 nand U147 SI_18_ ; R152_U240
g10558 not R152_U174 ; R152_U241
g10559 or SI_19_ U146 ; R152_U242
g10560 nand R152_U242 R152_U174 ; R152_U243
g10561 nand U146 SI_19_ ; R152_U244
g10562 not R152_U169 ; R152_U245
g10563 or SI_20_ U144 ; R152_U246
g10564 nand R152_U246 R152_U169 ; R152_U247
g10565 nand U144 SI_20_ ; R152_U248
g10566 not R152_U167 ; R152_U249
g10567 or SI_21_ U143 ; R152_U250
g10568 nand R152_U250 R152_U167 ; R152_U251
g10569 nand U143 SI_21_ ; R152_U252
g10570 not R152_U165 ; R152_U253
g10571 or SI_22_ U142 ; R152_U254
g10572 nand R152_U254 R152_U165 ; R152_U255
g10573 nand U142 SI_22_ ; R152_U256
g10574 not R152_U163 ; R152_U257
g10575 or SI_23_ U141 ; R152_U258
g10576 nand R152_U258 R152_U163 ; R152_U259
g10577 nand U141 SI_23_ ; R152_U260
g10578 not R152_U161 ; R152_U261
g10579 or SI_24_ U140 ; R152_U262
g10580 nand R152_U262 R152_U161 ; R152_U263
g10581 nand U140 SI_24_ ; R152_U264
g10582 not R152_U159 ; R152_U265
g10583 or SI_25_ U139 ; R152_U266
g10584 nand R152_U266 R152_U159 ; R152_U267
g10585 nand U139 SI_25_ ; R152_U268
g10586 not R152_U157 ; R152_U269
g10587 or SI_26_ U138 ; R152_U270
g10588 nand R152_U270 R152_U157 ; R152_U271
g10589 nand U138 SI_26_ ; R152_U272
g10590 not R152_U155 ; R152_U273
g10591 or SI_27_ U137 ; R152_U274
g10592 nand R152_U274 R152_U155 ; R152_U275
g10593 nand U137 SI_27_ ; R152_U276
g10594 not R152_U153 ; R152_U277
g10595 or SI_28_ U136 ; R152_U278
g10596 nand R152_U278 R152_U153 ; R152_U279
g10597 nand U136 SI_28_ ; R152_U280
g10598 not R152_U151 ; R152_U281
g10599 or SI_29_ U135 ; R152_U282
g10600 nand R152_U282 R152_U151 ; R152_U283
g10601 nand U135 SI_29_ ; R152_U284
g10602 not R152_U148 ; R152_U285
g10603 nand U133 SI_30_ ; R152_U286
g10604 or U133 SI_30_ ; R152_U287
g10605 nand R152_U283 R152_U127 ; R152_U288
g10606 nand U157 SI_0_ U156 ; R152_U289
g10607 nand U156 SI_1_ ; R152_U290
g10608 nand R152_U10 R152_U313 ; R152_U291
g10609 nand R152_U197 R152_U199 ; R152_U292
g10610 nand R152_U4 R152_U201 ; R152_U293
g10611 nand R152_U204 R152_U206 ; R152_U294
g10612 not R152_U37 ; R152_U295
g10613 nand R152_U115 R152_U201 ; R152_U296
g10614 nand R152_U37 R152_U209 ; R152_U297
g10615 nand R152_U213 R152_U214 ; R152_U298
g10616 nand R152_U298 R152_U215 ; R152_U299
g10617 nand R152_U299 R152_U216 ; R152_U300
g10618 not R152_U83 ; R152_U301
g10619 nand R152_U83 R152_U218 ; R152_U302
g10620 nand R152_U221 R152_U222 ; R152_U303
g10621 nand R152_U303 R152_U223 ; R152_U304
g10622 nand R152_U304 R152_U224 ; R152_U305
g10623 not R152_U82 ; R152_U306
g10624 nand R152_U82 R152_U226 ; R152_U307
g10625 not R152_U81 ; R152_U308
g10626 nand R152_U81 R152_U228 ; R152_U309
g10627 nand SI_0_ R152_U196 R152_U119 ; R152_U310
g10628 nand SI_1_ R152_U196 R152_U120 ; R152_U311
g10629 nand R152_U121 R152_U196 ; R152_U312
g10630 nand R152_U290 R152_U171 R152_U289 ; R152_U313
g10631 not R152_U141 ; R152_U314
g10632 nand R152_U10 R152_U316 ; R152_U315
g10633 nand R152_U318 R152_U290 R152_U317 ; R152_U316
g10634 nand U157 SI_0_ U156 ; R152_U317
g10635 nand SI_0_ SI_1_ U157 ; R152_U318
g10636 nand R152_U220 R152_U190 ; R152_U319
g10637 not R152_U188 ; R152_U320
g10638 nand R152_U7 R152_U190 ; R152_U321
g10639 not R152_U186 ; R152_U322
g10640 nand R152_U8 R152_U190 ; R152_U323
g10641 not R152_U184 ; R152_U324
g10642 nand R152_U9 R152_U190 ; R152_U325
g10643 not R152_U182 ; R152_U326
g10644 nand R152_U124 R152_U190 ; R152_U327
g10645 not R152_U180 ; R152_U328
g10646 nand R152_U212 R152_U135 ; R152_U329
g10647 not R152_U133 ; R152_U330
g10648 nand R152_U5 R152_U135 ; R152_U331
g10649 not R152_U131 ; R152_U332
g10650 nand R152_U6 R152_U135 ; R152_U333
g10651 not R152_U192 ; R152_U334
g10652 nand R152_U122 R152_U135 ; R152_U335
g10653 not R152_U190 ; R152_U336
g10654 nand R152_U480 R152_U23 ; R152_U337
g10655 nand U126 R152_U36 ; R152_U338
g10656 nand SI_9_ R152_U35 ; R152_U339
g10657 nand U126 R152_U36 ; R152_U340
g10658 nand SI_9_ R152_U35 ; R152_U341
g10659 nand R152_U341 R152_U340 ; R152_U342
g10660 nand R152_U130 R152_U131 ; R152_U343
g10661 nand R152_U332 R152_U342 ; R152_U344
g10662 nand U127 R152_U14 ; R152_U345
g10663 nand SI_8_ R152_U15 ; R152_U346
g10664 nand U127 R152_U14 ; R152_U347
g10665 nand SI_8_ R152_U15 ; R152_U348
g10666 nand R152_U348 R152_U347 ; R152_U349
g10667 nand R152_U132 R152_U133 ; R152_U350
g10668 nand R152_U330 R152_U349 ; R152_U351
g10669 nand U128 R152_U16 ; R152_U352
g10670 nand SI_7_ R152_U17 ; R152_U353
g10671 nand U128 R152_U16 ; R152_U354
g10672 nand SI_7_ R152_U17 ; R152_U355
g10673 nand R152_U355 R152_U354 ; R152_U356
g10674 nand R152_U134 R152_U135 ; R152_U357
g10675 nand R152_U211 R152_U356 ; R152_U358
g10676 nand U129 R152_U19 ; R152_U359
g10677 nand SI_6_ R152_U20 ; R152_U360
g10678 nand U129 R152_U19 ; R152_U361
g10679 nand SI_6_ R152_U20 ; R152_U362
g10680 nand R152_U362 R152_U361 ; R152_U363
g10681 nand R152_U136 R152_U137 ; R152_U364
g10682 nand R152_U208 R152_U363 ; R152_U365
g10683 nand U130 R152_U30 ; R152_U366
g10684 nand SI_5_ R152_U31 ; R152_U367
g10685 nand U130 R152_U30 ; R152_U368
g10686 nand SI_5_ R152_U31 ; R152_U369
g10687 nand R152_U369 R152_U368 ; R152_U370
g10688 nand R152_U138 R152_U139 ; R152_U371
g10689 nand R152_U205 R152_U370 ; R152_U372
g10690 nand U131 R152_U32 ; R152_U373
g10691 nand SI_4_ R152_U33 ; R152_U374
g10692 nand U131 R152_U32 ; R152_U375
g10693 nand SI_4_ R152_U33 ; R152_U376
g10694 nand R152_U376 R152_U375 ; R152_U377
g10695 nand R152_U140 R152_U141 ; R152_U378
g10696 nand R152_U314 R152_U377 ; R152_U379
g10697 nand U134 R152_U21 ; R152_U380
g10698 nand SI_3_ R152_U22 ; R152_U381
g10699 nand U134 R152_U21 ; R152_U382
g10700 nand SI_3_ R152_U22 ; R152_U383
g10701 nand R152_U383 R152_U382 ; R152_U384
g10702 nand R152_U142 R152_U143 ; R152_U385
g10703 nand R152_U198 R152_U384 ; R152_U386
g10704 nand U132 R152_U145 ; R152_U387
g10705 nand SI_31_ R152_U144 ; R152_U388
g10706 nand R152_U388 R152_U387 ; R152_U389
g10707 nand U132 R152_U145 ; R152_U390
g10708 nand SI_31_ R152_U144 ; R152_U391
g10709 nand R152_U11 R152_U79 R152_U80 ; R152_U392
g10710 nand SI_30_ R152_U389 U133 ; R152_U393
g10711 nand U133 R152_U79 ; R152_U394
g10712 nand SI_30_ R152_U80 ; R152_U395
g10713 nand U133 R152_U79 ; R152_U396
g10714 nand SI_30_ R152_U80 ; R152_U397
g10715 nand R152_U397 R152_U396 ; R152_U398
g10716 nand R152_U147 R152_U148 ; R152_U399
g10717 nand R152_U285 R152_U398 ; R152_U400
g10718 nand U145 R152_U27 ; R152_U401
g10719 nand SI_2_ R152_U28 ; R152_U402
g10720 nand U145 R152_U27 ; R152_U403
g10721 nand SI_2_ R152_U28 ; R152_U404
g10722 nand R152_U404 R152_U403 ; R152_U405
g10723 nand R152_U402 R152_U401 R152_U149 ; R152_U406
g10724 nand R152_U195 R152_U405 ; R152_U407
g10725 nand U135 R152_U77 ; R152_U408
g10726 nand SI_29_ R152_U78 ; R152_U409
g10727 nand U135 R152_U77 ; R152_U410
g10728 nand SI_29_ R152_U78 ; R152_U411
g10729 nand R152_U411 R152_U410 ; R152_U412
g10730 nand R152_U150 R152_U151 ; R152_U413
g10731 nand R152_U281 R152_U412 ; R152_U414
g10732 nand U136 R152_U75 ; R152_U415
g10733 nand SI_28_ R152_U76 ; R152_U416
g10734 nand U136 R152_U75 ; R152_U417
g10735 nand SI_28_ R152_U76 ; R152_U418
g10736 nand R152_U418 R152_U417 ; R152_U419
g10737 nand R152_U152 R152_U153 ; R152_U420
g10738 nand R152_U277 R152_U419 ; R152_U421
g10739 nand U137 R152_U73 ; R152_U422
g10740 nand SI_27_ R152_U74 ; R152_U423
g10741 nand U137 R152_U73 ; R152_U424
g10742 nand SI_27_ R152_U74 ; R152_U425
g10743 nand R152_U425 R152_U424 ; R152_U426
g10744 nand R152_U154 R152_U155 ; R152_U427
g10745 nand R152_U273 R152_U426 ; R152_U428
g10746 nand U138 R152_U71 ; R152_U429
g10747 nand SI_26_ R152_U72 ; R152_U430
g10748 nand U138 R152_U71 ; R152_U431
g10749 nand SI_26_ R152_U72 ; R152_U432
g10750 nand R152_U432 R152_U431 ; R152_U433
g10751 nand R152_U156 R152_U157 ; R152_U434
g10752 nand R152_U269 R152_U433 ; R152_U435
g10753 nand U139 R152_U69 ; R152_U436
g10754 nand SI_25_ R152_U70 ; R152_U437
g10755 nand U139 R152_U69 ; R152_U438
g10756 nand SI_25_ R152_U70 ; R152_U439
g10757 nand R152_U439 R152_U438 ; R152_U440
g10758 nand R152_U158 R152_U159 ; R152_U441
g10759 nand R152_U265 R152_U440 ; R152_U442
g10760 nand U140 R152_U67 ; R152_U443
g10761 nand SI_24_ R152_U68 ; R152_U444
g10762 nand U140 R152_U67 ; R152_U445
g10763 nand SI_24_ R152_U68 ; R152_U446
g10764 nand R152_U446 R152_U445 ; R152_U447
g10765 nand R152_U160 R152_U161 ; R152_U448
g10766 nand R152_U261 R152_U447 ; R152_U449
g10767 nand U141 R152_U65 ; R152_U450
g10768 nand SI_23_ R152_U66 ; R152_U451
g10769 nand U141 R152_U65 ; R152_U452
g10770 nand SI_23_ R152_U66 ; R152_U453
g10771 nand R152_U453 R152_U452 ; R152_U454
g10772 nand R152_U162 R152_U163 ; R152_U455
g10773 nand R152_U257 R152_U454 ; R152_U456
g10774 nand U142 R152_U63 ; R152_U457
g10775 nand SI_22_ R152_U64 ; R152_U458
g10776 nand U142 R152_U63 ; R152_U459
g10777 nand SI_22_ R152_U64 ; R152_U460
g10778 nand R152_U460 R152_U459 ; R152_U461
g10779 nand R152_U164 R152_U165 ; R152_U462
g10780 nand R152_U253 R152_U461 ; R152_U463
g10781 nand U143 R152_U61 ; R152_U464
g10782 nand SI_21_ R152_U62 ; R152_U465
g10783 nand U143 R152_U61 ; R152_U466
g10784 nand SI_21_ R152_U62 ; R152_U467
g10785 nand R152_U467 R152_U466 ; R152_U468
g10786 nand R152_U166 R152_U167 ; R152_U469
g10787 nand R152_U249 R152_U468 ; R152_U470
g10788 nand U144 R152_U59 ; R152_U471
g10789 nand SI_20_ R152_U60 ; R152_U472
g10790 nand U144 R152_U59 ; R152_U473
g10791 nand SI_20_ R152_U60 ; R152_U474
g10792 nand R152_U474 R152_U473 ; R152_U475
g10793 nand R152_U168 R152_U169 ; R152_U476
g10794 nand R152_U245 R152_U475 ; R152_U477
g10795 nand U156 R152_U170 ; R152_U478
g10796 nand R152_U120 R152_U26 ; R152_U479
g10797 nand R152_U479 R152_U478 ; R152_U480
g10798 nand SI_1_ R152_U170 R152_U26 ; R152_U481
g10799 nand R152_U194 U156 ; R152_U482
g10800 nand U146 R152_U57 ; R152_U483
g10801 nand SI_19_ R152_U58 ; R152_U484
g10802 nand U146 R152_U57 ; R152_U485
g10803 nand SI_19_ R152_U58 ; R152_U486
g10804 nand R152_U486 R152_U485 ; R152_U487
g10805 nand R152_U173 R152_U174 ; R152_U488
g10806 nand R152_U241 R152_U487 ; R152_U489
g10807 nand U147 R152_U55 ; R152_U490
g10808 nand SI_18_ R152_U56 ; R152_U491
g10809 nand U147 R152_U55 ; R152_U492
g10810 nand SI_18_ R152_U56 ; R152_U493
g10811 nand R152_U493 R152_U492 ; R152_U494
g10812 nand R152_U175 R152_U176 ; R152_U495
g10813 nand R152_U237 R152_U494 ; R152_U496
g10814 nand U148 R152_U53 ; R152_U497
g10815 nand SI_17_ R152_U54 ; R152_U498
g10816 nand U148 R152_U53 ; R152_U499
g10817 nand SI_17_ R152_U54 ; R152_U500
g10818 nand R152_U500 R152_U499 ; R152_U501
g10819 nand R152_U177 R152_U178 ; R152_U502
g10820 nand R152_U233 R152_U501 ; R152_U503
g10821 nand U149 R152_U51 ; R152_U504
g10822 nand SI_16_ R152_U52 ; R152_U505
g10823 nand U149 R152_U51 ; R152_U506
g10824 nand SI_16_ R152_U52 ; R152_U507
g10825 nand R152_U507 R152_U506 ; R152_U508
g10826 nand R152_U179 R152_U180 ; R152_U509
g10827 nand R152_U328 R152_U508 ; R152_U510
g10828 nand U150 R152_U38 ; R152_U511
g10829 nand SI_15_ R152_U39 ; R152_U512
g10830 nand U150 R152_U38 ; R152_U513
g10831 nand SI_15_ R152_U39 ; R152_U514
g10832 nand R152_U514 R152_U513 ; R152_U515
g10833 nand R152_U181 R152_U182 ; R152_U516
g10834 nand R152_U326 R152_U515 ; R152_U517
g10835 nand U151 R152_U40 ; R152_U518
g10836 nand SI_14_ R152_U41 ; R152_U519
g10837 nand U151 R152_U40 ; R152_U520
g10838 nand SI_14_ R152_U41 ; R152_U521
g10839 nand R152_U521 R152_U520 ; R152_U522
g10840 nand R152_U183 R152_U184 ; R152_U523
g10841 nand R152_U324 R152_U522 ; R152_U524
g10842 nand U152 R152_U42 ; R152_U525
g10843 nand SI_13_ R152_U43 ; R152_U526
g10844 nand U152 R152_U42 ; R152_U527
g10845 nand SI_13_ R152_U43 ; R152_U528
g10846 nand R152_U528 R152_U527 ; R152_U529
g10847 nand R152_U185 R152_U186 ; R152_U530
g10848 nand R152_U322 R152_U529 ; R152_U531
g10849 nand U153 R152_U44 ; R152_U532
g10850 nand SI_12_ R152_U45 ; R152_U533
g10851 nand U153 R152_U44 ; R152_U534
g10852 nand SI_12_ R152_U45 ; R152_U535
g10853 nand R152_U535 R152_U534 ; R152_U536
g10854 nand R152_U187 R152_U188 ; R152_U537
g10855 nand R152_U320 R152_U536 ; R152_U538
g10856 nand U154 R152_U46 ; R152_U539
g10857 nand SI_11_ R152_U47 ; R152_U540
g10858 nand U154 R152_U46 ; R152_U541
g10859 nand SI_11_ R152_U47 ; R152_U542
g10860 nand R152_U542 R152_U541 ; R152_U543
g10861 nand R152_U189 R152_U190 ; R152_U544
g10862 nand R152_U336 R152_U543 ; R152_U545
g10863 nand U155 R152_U49 ; R152_U546
g10864 nand SI_10_ R152_U50 ; R152_U547
g10865 nand U155 R152_U49 ; R152_U548
g10866 nand SI_10_ R152_U50 ; R152_U549
g10867 nand R152_U549 R152_U548 ; R152_U550
g10868 nand R152_U191 R152_U192 ; R152_U551
g10869 nand R152_U334 R152_U550 ; R152_U552
g10870 nand U157 R152_U24 ; R152_U553
g10871 nand SI_0_ R152_U25 ; R152_U554
g10872 not P3_ADDR_REG_19__SCAN_IN ; LT_1602_U6
g10873 not P1_ADDR_REG_19__SCAN_IN ; LT_1601_U6
g10874 and SUB_1596_U159 SUB_1596_U155 ; SUB_1596_U4
g10875 nand SUB_1596_U221 SUB_1596_U220 SUB_1596_U160 ; SUB_1596_U5
g10876 not ADD_1596_U7 ; SUB_1596_U6
g10877 not P2_ADDR_REG_0__SCAN_IN ; SUB_1596_U7
g10878 not P2_ADDR_REG_1__SCAN_IN ; SUB_1596_U8
g10879 nand ADD_1596_U7 P2_ADDR_REG_0__SCAN_IN ; SUB_1596_U9
g10880 not ADD_1596_U55 ; SUB_1596_U10
g10881 not ADD_1596_U54 ; SUB_1596_U11
g10882 not P2_ADDR_REG_2__SCAN_IN ; SUB_1596_U12
g10883 nand SUB_1596_U90 SUB_1596_U89 ; SUB_1596_U13
g10884 not ADD_1596_U53 ; SUB_1596_U14
g10885 not P2_ADDR_REG_3__SCAN_IN ; SUB_1596_U15
g10886 not ADD_1596_U52 ; SUB_1596_U16
g10887 not P2_ADDR_REG_4__SCAN_IN ; SUB_1596_U17
g10888 nand SUB_1596_U98 SUB_1596_U97 ; SUB_1596_U18
g10889 not ADD_1596_U51 ; SUB_1596_U19
g10890 not P2_ADDR_REG_5__SCAN_IN ; SUB_1596_U20
g10891 not ADD_1596_U50 ; SUB_1596_U21
g10892 not P2_ADDR_REG_6__SCAN_IN ; SUB_1596_U22
g10893 not ADD_1596_U49 ; SUB_1596_U23
g10894 not P2_ADDR_REG_7__SCAN_IN ; SUB_1596_U24
g10895 nand SUB_1596_U110 SUB_1596_U109 ; SUB_1596_U25
g10896 not ADD_1596_U48 ; SUB_1596_U26
g10897 not P2_ADDR_REG_8__SCAN_IN ; SUB_1596_U27
g10898 not P2_ADDR_REG_9__SCAN_IN ; SUB_1596_U28
g10899 not ADD_1596_U47 ; SUB_1596_U29
g10900 nand SUB_1596_U118 SUB_1596_U117 ; SUB_1596_U30
g10901 not ADD_1596_U64 ; SUB_1596_U31
g10902 not P2_ADDR_REG_10__SCAN_IN ; SUB_1596_U32
g10903 not ADD_1596_U63 ; SUB_1596_U33
g10904 not P2_ADDR_REG_11__SCAN_IN ; SUB_1596_U34
g10905 not ADD_1596_U62 ; SUB_1596_U35
g10906 not P2_ADDR_REG_12__SCAN_IN ; SUB_1596_U36
g10907 nand SUB_1596_U130 SUB_1596_U129 ; SUB_1596_U37
g10908 not ADD_1596_U61 ; SUB_1596_U38
g10909 not P2_ADDR_REG_13__SCAN_IN ; SUB_1596_U39
g10910 nand SUB_1596_U134 SUB_1596_U133 ; SUB_1596_U40
g10911 not ADD_1596_U60 ; SUB_1596_U41
g10912 not P2_ADDR_REG_14__SCAN_IN ; SUB_1596_U42
g10913 nand SUB_1596_U138 SUB_1596_U137 ; SUB_1596_U43
g10914 not ADD_1596_U59 ; SUB_1596_U44
g10915 not P2_ADDR_REG_15__SCAN_IN ; SUB_1596_U45
g10916 not ADD_1596_U58 ; SUB_1596_U46
g10917 not P2_ADDR_REG_16__SCAN_IN ; SUB_1596_U47
g10918 not ADD_1596_U57 ; SUB_1596_U48
g10919 not P2_ADDR_REG_17__SCAN_IN ; SUB_1596_U49
g10920 nand SUB_1596_U150 SUB_1596_U149 ; SUB_1596_U50
g10921 not ADD_1596_U56 ; SUB_1596_U51
g10922 not P2_ADDR_REG_18__SCAN_IN ; SUB_1596_U52
g10923 nand SUB_1596_U291 SUB_1596_U290 ; SUB_1596_U53
g10924 nand SUB_1596_U167 SUB_1596_U166 ; SUB_1596_U54
g10925 nand SUB_1596_U174 SUB_1596_U173 ; SUB_1596_U55
g10926 nand SUB_1596_U181 SUB_1596_U180 ; SUB_1596_U56
g10927 nand SUB_1596_U188 SUB_1596_U187 ; SUB_1596_U57
g10928 nand SUB_1596_U195 SUB_1596_U194 ; SUB_1596_U58
g10929 nand SUB_1596_U202 SUB_1596_U201 ; SUB_1596_U59
g10930 nand SUB_1596_U209 SUB_1596_U208 ; SUB_1596_U60
g10931 nand SUB_1596_U216 SUB_1596_U215 ; SUB_1596_U61
g10932 nand SUB_1596_U233 SUB_1596_U232 ; SUB_1596_U62
g10933 nand SUB_1596_U240 SUB_1596_U239 ; SUB_1596_U63
g10934 nand SUB_1596_U247 SUB_1596_U246 ; SUB_1596_U64
g10935 nand SUB_1596_U254 SUB_1596_U253 ; SUB_1596_U65
g10936 nand SUB_1596_U261 SUB_1596_U260 ; SUB_1596_U66
g10937 nand SUB_1596_U268 SUB_1596_U267 ; SUB_1596_U67
g10938 nand SUB_1596_U275 SUB_1596_U274 ; SUB_1596_U68
g10939 nand SUB_1596_U282 SUB_1596_U281 ; SUB_1596_U69
g10940 nand SUB_1596_U289 SUB_1596_U288 ; SUB_1596_U70
g10941 nand SUB_1596_U114 SUB_1596_U113 ; SUB_1596_U71
g10942 nand SUB_1596_U106 SUB_1596_U105 ; SUB_1596_U72
g10943 nand SUB_1596_U102 SUB_1596_U101 ; SUB_1596_U73
g10944 nand SUB_1596_U94 SUB_1596_U93 ; SUB_1596_U74
g10945 nand SUB_1596_U76 SUB_1596_U86 ; SUB_1596_U75
g10946 nand ADD_1596_U55 SUB_1596_U84 ; SUB_1596_U76
g10947 not P2_ADDR_REG_19__SCAN_IN ; SUB_1596_U77
g10948 not ADD_1596_U6 ; SUB_1596_U78
g10949 nand SUB_1596_U146 SUB_1596_U145 ; SUB_1596_U79
g10950 nand SUB_1596_U142 SUB_1596_U141 ; SUB_1596_U80
g10951 nand SUB_1596_U126 SUB_1596_U125 ; SUB_1596_U81
g10952 nand SUB_1596_U122 SUB_1596_U121 ; SUB_1596_U82
g10953 not SUB_1596_U76 ; SUB_1596_U83
g10954 not SUB_1596_U9 ; SUB_1596_U84
g10955 nand SUB_1596_U10 SUB_1596_U9 ; SUB_1596_U85
g10956 nand SUB_1596_U85 P2_ADDR_REG_1__SCAN_IN ; SUB_1596_U86
g10957 not SUB_1596_U75 ; SUB_1596_U87
g10958 or ADD_1596_U54 P2_ADDR_REG_2__SCAN_IN ; SUB_1596_U88
g10959 nand SUB_1596_U88 SUB_1596_U75 ; SUB_1596_U89
g10960 nand ADD_1596_U54 P2_ADDR_REG_2__SCAN_IN ; SUB_1596_U90
g10961 not SUB_1596_U13 ; SUB_1596_U91
g10962 nand SUB_1596_U91 SUB_1596_U15 ; SUB_1596_U92
g10963 nand ADD_1596_U53 SUB_1596_U92 ; SUB_1596_U93
g10964 nand SUB_1596_U13 P2_ADDR_REG_3__SCAN_IN ; SUB_1596_U94
g10965 not SUB_1596_U74 ; SUB_1596_U95
g10966 or ADD_1596_U52 P2_ADDR_REG_4__SCAN_IN ; SUB_1596_U96
g10967 nand SUB_1596_U96 SUB_1596_U74 ; SUB_1596_U97
g10968 nand ADD_1596_U52 P2_ADDR_REG_4__SCAN_IN ; SUB_1596_U98
g10969 not SUB_1596_U18 ; SUB_1596_U99
g10970 nand SUB_1596_U99 SUB_1596_U20 ; SUB_1596_U100
g10971 nand ADD_1596_U51 SUB_1596_U100 ; SUB_1596_U101
g10972 nand SUB_1596_U18 P2_ADDR_REG_5__SCAN_IN ; SUB_1596_U102
g10973 not SUB_1596_U73 ; SUB_1596_U103
g10974 or ADD_1596_U50 P2_ADDR_REG_6__SCAN_IN ; SUB_1596_U104
g10975 nand SUB_1596_U104 SUB_1596_U73 ; SUB_1596_U105
g10976 nand ADD_1596_U50 P2_ADDR_REG_6__SCAN_IN ; SUB_1596_U106
g10977 not SUB_1596_U72 ; SUB_1596_U107
g10978 or ADD_1596_U49 P2_ADDR_REG_7__SCAN_IN ; SUB_1596_U108
g10979 nand SUB_1596_U108 SUB_1596_U72 ; SUB_1596_U109
g10980 nand ADD_1596_U49 P2_ADDR_REG_7__SCAN_IN ; SUB_1596_U110
g10981 not SUB_1596_U25 ; SUB_1596_U111
g10982 nand SUB_1596_U111 SUB_1596_U27 ; SUB_1596_U112
g10983 nand ADD_1596_U48 SUB_1596_U112 ; SUB_1596_U113
g10984 nand SUB_1596_U25 P2_ADDR_REG_8__SCAN_IN ; SUB_1596_U114
g10985 not SUB_1596_U71 ; SUB_1596_U115
g10986 or ADD_1596_U47 P2_ADDR_REG_9__SCAN_IN ; SUB_1596_U116
g10987 nand SUB_1596_U116 SUB_1596_U71 ; SUB_1596_U117
g10988 nand ADD_1596_U47 P2_ADDR_REG_9__SCAN_IN ; SUB_1596_U118
g10989 not SUB_1596_U30 ; SUB_1596_U119
g10990 nand SUB_1596_U119 SUB_1596_U32 ; SUB_1596_U120
g10991 nand ADD_1596_U64 SUB_1596_U120 ; SUB_1596_U121
g10992 nand SUB_1596_U30 P2_ADDR_REG_10__SCAN_IN ; SUB_1596_U122
g10993 not SUB_1596_U82 ; SUB_1596_U123
g10994 or ADD_1596_U63 P2_ADDR_REG_11__SCAN_IN ; SUB_1596_U124
g10995 nand SUB_1596_U124 SUB_1596_U82 ; SUB_1596_U125
g10996 nand ADD_1596_U63 P2_ADDR_REG_11__SCAN_IN ; SUB_1596_U126
g10997 not SUB_1596_U81 ; SUB_1596_U127
g10998 or ADD_1596_U62 P2_ADDR_REG_12__SCAN_IN ; SUB_1596_U128
g10999 nand SUB_1596_U128 SUB_1596_U81 ; SUB_1596_U129
g11000 nand ADD_1596_U62 P2_ADDR_REG_12__SCAN_IN ; SUB_1596_U130
g11001 not SUB_1596_U37 ; SUB_1596_U131
g11002 nand SUB_1596_U131 SUB_1596_U39 ; SUB_1596_U132
g11003 nand ADD_1596_U61 SUB_1596_U132 ; SUB_1596_U133
g11004 nand SUB_1596_U37 P2_ADDR_REG_13__SCAN_IN ; SUB_1596_U134
g11005 not SUB_1596_U40 ; SUB_1596_U135
g11006 nand SUB_1596_U135 SUB_1596_U42 ; SUB_1596_U136
g11007 nand ADD_1596_U60 SUB_1596_U136 ; SUB_1596_U137
g11008 nand SUB_1596_U40 P2_ADDR_REG_14__SCAN_IN ; SUB_1596_U138
g11009 not SUB_1596_U43 ; SUB_1596_U139
g11010 nand SUB_1596_U139 SUB_1596_U45 ; SUB_1596_U140
g11011 nand ADD_1596_U59 SUB_1596_U140 ; SUB_1596_U141
g11012 nand SUB_1596_U43 P2_ADDR_REG_15__SCAN_IN ; SUB_1596_U142
g11013 not SUB_1596_U80 ; SUB_1596_U143
g11014 or ADD_1596_U58 P2_ADDR_REG_16__SCAN_IN ; SUB_1596_U144
g11015 nand SUB_1596_U144 SUB_1596_U80 ; SUB_1596_U145
g11016 nand ADD_1596_U58 P2_ADDR_REG_16__SCAN_IN ; SUB_1596_U146
g11017 not SUB_1596_U79 ; SUB_1596_U147
g11018 or ADD_1596_U57 P2_ADDR_REG_17__SCAN_IN ; SUB_1596_U148
g11019 nand SUB_1596_U148 SUB_1596_U79 ; SUB_1596_U149
g11020 nand ADD_1596_U57 P2_ADDR_REG_17__SCAN_IN ; SUB_1596_U150
g11021 not SUB_1596_U50 ; SUB_1596_U151
g11022 nand SUB_1596_U151 SUB_1596_U52 ; SUB_1596_U152
g11023 nand ADD_1596_U56 SUB_1596_U152 ; SUB_1596_U153
g11024 nand SUB_1596_U50 P2_ADDR_REG_18__SCAN_IN ; SUB_1596_U154
g11025 nand SUB_1596_U154 SUB_1596_U153 SUB_1596_U223 SUB_1596_U222 ; SUB_1596_U155
g11026 nand SUB_1596_U50 P2_ADDR_REG_18__SCAN_IN ; SUB_1596_U156
g11027 nand SUB_1596_U156 SUB_1596_U51 ; SUB_1596_U157
g11028 nand SUB_1596_U151 SUB_1596_U52 ; SUB_1596_U158
g11029 nand SUB_1596_U158 SUB_1596_U157 SUB_1596_U226 ; SUB_1596_U159
g11030 nand SUB_1596_U219 SUB_1596_U10 ; SUB_1596_U160
g11031 nand SUB_1596_U29 P2_ADDR_REG_9__SCAN_IN ; SUB_1596_U161
g11032 nand ADD_1596_U47 SUB_1596_U28 ; SUB_1596_U162
g11033 nand SUB_1596_U29 P2_ADDR_REG_9__SCAN_IN ; SUB_1596_U163
g11034 nand ADD_1596_U47 SUB_1596_U28 ; SUB_1596_U164
g11035 nand SUB_1596_U164 SUB_1596_U163 ; SUB_1596_U165
g11036 nand SUB_1596_U162 SUB_1596_U161 SUB_1596_U71 ; SUB_1596_U166
g11037 nand SUB_1596_U115 SUB_1596_U165 ; SUB_1596_U167
g11038 nand SUB_1596_U25 P2_ADDR_REG_8__SCAN_IN ; SUB_1596_U168
g11039 nand SUB_1596_U111 SUB_1596_U27 ; SUB_1596_U169
g11040 nand SUB_1596_U25 P2_ADDR_REG_8__SCAN_IN ; SUB_1596_U170
g11041 nand SUB_1596_U111 SUB_1596_U27 ; SUB_1596_U171
g11042 nand SUB_1596_U171 SUB_1596_U170 ; SUB_1596_U172
g11043 nand SUB_1596_U169 SUB_1596_U168 SUB_1596_U26 ; SUB_1596_U173
g11044 nand SUB_1596_U172 ADD_1596_U48 ; SUB_1596_U174
g11045 nand SUB_1596_U23 P2_ADDR_REG_7__SCAN_IN ; SUB_1596_U175
g11046 nand ADD_1596_U49 SUB_1596_U24 ; SUB_1596_U176
g11047 nand SUB_1596_U23 P2_ADDR_REG_7__SCAN_IN ; SUB_1596_U177
g11048 nand ADD_1596_U49 SUB_1596_U24 ; SUB_1596_U178
g11049 nand SUB_1596_U178 SUB_1596_U177 ; SUB_1596_U179
g11050 nand SUB_1596_U176 SUB_1596_U175 SUB_1596_U72 ; SUB_1596_U180
g11051 nand SUB_1596_U107 SUB_1596_U179 ; SUB_1596_U181
g11052 nand SUB_1596_U21 P2_ADDR_REG_6__SCAN_IN ; SUB_1596_U182
g11053 nand ADD_1596_U50 SUB_1596_U22 ; SUB_1596_U183
g11054 nand SUB_1596_U21 P2_ADDR_REG_6__SCAN_IN ; SUB_1596_U184
g11055 nand ADD_1596_U50 SUB_1596_U22 ; SUB_1596_U185
g11056 nand SUB_1596_U185 SUB_1596_U184 ; SUB_1596_U186
g11057 nand SUB_1596_U183 SUB_1596_U182 SUB_1596_U73 ; SUB_1596_U187
g11058 nand SUB_1596_U103 SUB_1596_U186 ; SUB_1596_U188
g11059 nand SUB_1596_U18 P2_ADDR_REG_5__SCAN_IN ; SUB_1596_U189
g11060 nand SUB_1596_U99 SUB_1596_U20 ; SUB_1596_U190
g11061 nand SUB_1596_U18 P2_ADDR_REG_5__SCAN_IN ; SUB_1596_U191
g11062 nand SUB_1596_U99 SUB_1596_U20 ; SUB_1596_U192
g11063 nand SUB_1596_U192 SUB_1596_U191 ; SUB_1596_U193
g11064 nand SUB_1596_U190 SUB_1596_U189 SUB_1596_U19 ; SUB_1596_U194
g11065 nand SUB_1596_U193 ADD_1596_U51 ; SUB_1596_U195
g11066 nand SUB_1596_U16 P2_ADDR_REG_4__SCAN_IN ; SUB_1596_U196
g11067 nand ADD_1596_U52 SUB_1596_U17 ; SUB_1596_U197
g11068 nand SUB_1596_U16 P2_ADDR_REG_4__SCAN_IN ; SUB_1596_U198
g11069 nand ADD_1596_U52 SUB_1596_U17 ; SUB_1596_U199
g11070 nand SUB_1596_U199 SUB_1596_U198 ; SUB_1596_U200
g11071 nand SUB_1596_U197 SUB_1596_U196 SUB_1596_U74 ; SUB_1596_U201
g11072 nand SUB_1596_U95 SUB_1596_U200 ; SUB_1596_U202
g11073 nand SUB_1596_U13 P2_ADDR_REG_3__SCAN_IN ; SUB_1596_U203
g11074 nand SUB_1596_U91 SUB_1596_U15 ; SUB_1596_U204
g11075 nand SUB_1596_U13 P2_ADDR_REG_3__SCAN_IN ; SUB_1596_U205
g11076 nand SUB_1596_U91 SUB_1596_U15 ; SUB_1596_U206
g11077 nand SUB_1596_U206 SUB_1596_U205 ; SUB_1596_U207
g11078 nand SUB_1596_U204 SUB_1596_U203 SUB_1596_U14 ; SUB_1596_U208
g11079 nand SUB_1596_U207 ADD_1596_U53 ; SUB_1596_U209
g11080 nand SUB_1596_U11 P2_ADDR_REG_2__SCAN_IN ; SUB_1596_U210
g11081 nand ADD_1596_U54 SUB_1596_U12 ; SUB_1596_U211
g11082 nand SUB_1596_U11 P2_ADDR_REG_2__SCAN_IN ; SUB_1596_U212
g11083 nand ADD_1596_U54 SUB_1596_U12 ; SUB_1596_U213
g11084 nand SUB_1596_U213 SUB_1596_U212 ; SUB_1596_U214
g11085 nand SUB_1596_U211 SUB_1596_U210 SUB_1596_U75 ; SUB_1596_U215
g11086 nand SUB_1596_U87 SUB_1596_U214 ; SUB_1596_U216
g11087 nand SUB_1596_U9 P2_ADDR_REG_1__SCAN_IN ; SUB_1596_U217
g11088 nand SUB_1596_U84 SUB_1596_U8 ; SUB_1596_U218
g11089 nand SUB_1596_U218 SUB_1596_U217 ; SUB_1596_U219
g11090 nand ADD_1596_U55 SUB_1596_U9 SUB_1596_U8 ; SUB_1596_U220
g11091 nand SUB_1596_U83 P2_ADDR_REG_1__SCAN_IN ; SUB_1596_U221
g11092 nand SUB_1596_U78 P2_ADDR_REG_19__SCAN_IN ; SUB_1596_U222
g11093 nand ADD_1596_U6 SUB_1596_U77 ; SUB_1596_U223
g11094 nand SUB_1596_U78 P2_ADDR_REG_19__SCAN_IN ; SUB_1596_U224
g11095 nand ADD_1596_U6 SUB_1596_U77 ; SUB_1596_U225
g11096 nand SUB_1596_U225 SUB_1596_U224 ; SUB_1596_U226
g11097 nand SUB_1596_U50 P2_ADDR_REG_18__SCAN_IN ; SUB_1596_U227
g11098 nand SUB_1596_U151 SUB_1596_U52 ; SUB_1596_U228
g11099 nand SUB_1596_U50 P2_ADDR_REG_18__SCAN_IN ; SUB_1596_U229
g11100 nand SUB_1596_U151 SUB_1596_U52 ; SUB_1596_U230
g11101 nand SUB_1596_U230 SUB_1596_U229 ; SUB_1596_U231
g11102 nand SUB_1596_U228 SUB_1596_U227 SUB_1596_U51 ; SUB_1596_U232
g11103 nand SUB_1596_U231 ADD_1596_U56 ; SUB_1596_U233
g11104 nand SUB_1596_U48 P2_ADDR_REG_17__SCAN_IN ; SUB_1596_U234
g11105 nand ADD_1596_U57 SUB_1596_U49 ; SUB_1596_U235
g11106 nand SUB_1596_U48 P2_ADDR_REG_17__SCAN_IN ; SUB_1596_U236
g11107 nand ADD_1596_U57 SUB_1596_U49 ; SUB_1596_U237
g11108 nand SUB_1596_U237 SUB_1596_U236 ; SUB_1596_U238
g11109 nand SUB_1596_U235 SUB_1596_U234 SUB_1596_U79 ; SUB_1596_U239
g11110 nand SUB_1596_U147 SUB_1596_U238 ; SUB_1596_U240
g11111 nand SUB_1596_U46 P2_ADDR_REG_16__SCAN_IN ; SUB_1596_U241
g11112 nand ADD_1596_U58 SUB_1596_U47 ; SUB_1596_U242
g11113 nand SUB_1596_U46 P2_ADDR_REG_16__SCAN_IN ; SUB_1596_U243
g11114 nand ADD_1596_U58 SUB_1596_U47 ; SUB_1596_U244
g11115 nand SUB_1596_U244 SUB_1596_U243 ; SUB_1596_U245
g11116 nand SUB_1596_U242 SUB_1596_U241 SUB_1596_U80 ; SUB_1596_U246
g11117 nand SUB_1596_U143 SUB_1596_U245 ; SUB_1596_U247
g11118 nand SUB_1596_U43 P2_ADDR_REG_15__SCAN_IN ; SUB_1596_U248
g11119 nand SUB_1596_U139 SUB_1596_U45 ; SUB_1596_U249
g11120 nand SUB_1596_U43 P2_ADDR_REG_15__SCAN_IN ; SUB_1596_U250
g11121 nand SUB_1596_U139 SUB_1596_U45 ; SUB_1596_U251
g11122 nand SUB_1596_U251 SUB_1596_U250 ; SUB_1596_U252
g11123 nand SUB_1596_U249 SUB_1596_U248 SUB_1596_U44 ; SUB_1596_U253
g11124 nand SUB_1596_U252 ADD_1596_U59 ; SUB_1596_U254
g11125 nand SUB_1596_U40 P2_ADDR_REG_14__SCAN_IN ; SUB_1596_U255
g11126 nand SUB_1596_U135 SUB_1596_U42 ; SUB_1596_U256
g11127 nand SUB_1596_U40 P2_ADDR_REG_14__SCAN_IN ; SUB_1596_U257
g11128 nand SUB_1596_U135 SUB_1596_U42 ; SUB_1596_U258
g11129 nand SUB_1596_U258 SUB_1596_U257 ; SUB_1596_U259
g11130 nand SUB_1596_U256 SUB_1596_U255 SUB_1596_U41 ; SUB_1596_U260
g11131 nand SUB_1596_U259 ADD_1596_U60 ; SUB_1596_U261
g11132 nand SUB_1596_U37 P2_ADDR_REG_13__SCAN_IN ; SUB_1596_U262
g11133 nand SUB_1596_U131 SUB_1596_U39 ; SUB_1596_U263
g11134 nand SUB_1596_U37 P2_ADDR_REG_13__SCAN_IN ; SUB_1596_U264
g11135 nand SUB_1596_U131 SUB_1596_U39 ; SUB_1596_U265
g11136 nand SUB_1596_U265 SUB_1596_U264 ; SUB_1596_U266
g11137 nand SUB_1596_U263 SUB_1596_U262 SUB_1596_U38 ; SUB_1596_U267
g11138 nand SUB_1596_U266 ADD_1596_U61 ; SUB_1596_U268
g11139 nand SUB_1596_U35 P2_ADDR_REG_12__SCAN_IN ; SUB_1596_U269
g11140 nand ADD_1596_U62 SUB_1596_U36 ; SUB_1596_U270
g11141 nand SUB_1596_U35 P2_ADDR_REG_12__SCAN_IN ; SUB_1596_U271
g11142 nand ADD_1596_U62 SUB_1596_U36 ; SUB_1596_U272
g11143 nand SUB_1596_U272 SUB_1596_U271 ; SUB_1596_U273
g11144 nand SUB_1596_U270 SUB_1596_U269 SUB_1596_U81 ; SUB_1596_U274
g11145 nand SUB_1596_U127 SUB_1596_U273 ; SUB_1596_U275
g11146 nand SUB_1596_U33 P2_ADDR_REG_11__SCAN_IN ; SUB_1596_U276
g11147 nand ADD_1596_U63 SUB_1596_U34 ; SUB_1596_U277
g11148 nand SUB_1596_U33 P2_ADDR_REG_11__SCAN_IN ; SUB_1596_U278
g11149 nand ADD_1596_U63 SUB_1596_U34 ; SUB_1596_U279
g11150 nand SUB_1596_U279 SUB_1596_U278 ; SUB_1596_U280
g11151 nand SUB_1596_U277 SUB_1596_U276 SUB_1596_U82 ; SUB_1596_U281
g11152 nand SUB_1596_U123 SUB_1596_U280 ; SUB_1596_U282
g11153 nand SUB_1596_U30 P2_ADDR_REG_10__SCAN_IN ; SUB_1596_U283
g11154 nand SUB_1596_U119 SUB_1596_U32 ; SUB_1596_U284
g11155 nand SUB_1596_U30 P2_ADDR_REG_10__SCAN_IN ; SUB_1596_U285
g11156 nand SUB_1596_U119 SUB_1596_U32 ; SUB_1596_U286
g11157 nand SUB_1596_U286 SUB_1596_U285 ; SUB_1596_U287
g11158 nand SUB_1596_U284 SUB_1596_U283 SUB_1596_U31 ; SUB_1596_U288
g11159 nand SUB_1596_U287 ADD_1596_U64 ; SUB_1596_U289
g11160 nand SUB_1596_U6 P2_ADDR_REG_0__SCAN_IN ; SUB_1596_U290
g11161 nand ADD_1596_U7 SUB_1596_U7 ; SUB_1596_U291
g11162 nand ADD_1596_U174 ADD_1596_U178 ; ADD_1596_U6
g11163 nand ADD_1596_U9 ADD_1596_U179 ; ADD_1596_U7
g11164 not P3_ADDR_REG_0__SCAN_IN ; ADD_1596_U8
g11165 nand ADD_1596_U46 P3_ADDR_REG_0__SCAN_IN ; ADD_1596_U9
g11166 not P1_ADDR_REG_1__SCAN_IN ; ADD_1596_U10
g11167 not P3_ADDR_REG_2__SCAN_IN ; ADD_1596_U11
g11168 not P1_ADDR_REG_2__SCAN_IN ; ADD_1596_U12
g11169 not P3_ADDR_REG_3__SCAN_IN ; ADD_1596_U13
g11170 not P1_ADDR_REG_3__SCAN_IN ; ADD_1596_U14
g11171 not P3_ADDR_REG_4__SCAN_IN ; ADD_1596_U15
g11172 not P1_ADDR_REG_4__SCAN_IN ; ADD_1596_U16
g11173 not P3_ADDR_REG_5__SCAN_IN ; ADD_1596_U17
g11174 not P1_ADDR_REG_5__SCAN_IN ; ADD_1596_U18
g11175 not P3_ADDR_REG_6__SCAN_IN ; ADD_1596_U19
g11176 not P1_ADDR_REG_6__SCAN_IN ; ADD_1596_U20
g11177 not P3_ADDR_REG_7__SCAN_IN ; ADD_1596_U21
g11178 not P1_ADDR_REG_7__SCAN_IN ; ADD_1596_U22
g11179 not P3_ADDR_REG_8__SCAN_IN ; ADD_1596_U23
g11180 not P1_ADDR_REG_8__SCAN_IN ; ADD_1596_U24
g11181 not P3_ADDR_REG_9__SCAN_IN ; ADD_1596_U25
g11182 not P1_ADDR_REG_9__SCAN_IN ; ADD_1596_U26
g11183 not P3_ADDR_REG_10__SCAN_IN ; ADD_1596_U27
g11184 not P1_ADDR_REG_10__SCAN_IN ; ADD_1596_U28
g11185 not P3_ADDR_REG_11__SCAN_IN ; ADD_1596_U29
g11186 not P1_ADDR_REG_11__SCAN_IN ; ADD_1596_U30
g11187 not P3_ADDR_REG_12__SCAN_IN ; ADD_1596_U31
g11188 not P1_ADDR_REG_12__SCAN_IN ; ADD_1596_U32
g11189 not P3_ADDR_REG_13__SCAN_IN ; ADD_1596_U33
g11190 not P1_ADDR_REG_13__SCAN_IN ; ADD_1596_U34
g11191 not P3_ADDR_REG_14__SCAN_IN ; ADD_1596_U35
g11192 not P1_ADDR_REG_14__SCAN_IN ; ADD_1596_U36
g11193 not P3_ADDR_REG_15__SCAN_IN ; ADD_1596_U37
g11194 not P1_ADDR_REG_15__SCAN_IN ; ADD_1596_U38
g11195 not P3_ADDR_REG_16__SCAN_IN ; ADD_1596_U39
g11196 not P1_ADDR_REG_16__SCAN_IN ; ADD_1596_U40
g11197 not P3_ADDR_REG_17__SCAN_IN ; ADD_1596_U41
g11198 not P1_ADDR_REG_17__SCAN_IN ; ADD_1596_U42
g11199 not P3_ADDR_REG_18__SCAN_IN ; ADD_1596_U43
g11200 not P1_ADDR_REG_18__SCAN_IN ; ADD_1596_U44
g11201 nand ADD_1596_U169 ADD_1596_U168 ; ADD_1596_U45
g11202 not P1_ADDR_REG_0__SCAN_IN ; ADD_1596_U46
g11203 nand ADD_1596_U184 ADD_1596_U183 ; ADD_1596_U47
g11204 nand ADD_1596_U189 ADD_1596_U188 ; ADD_1596_U48
g11205 nand ADD_1596_U194 ADD_1596_U193 ; ADD_1596_U49
g11206 nand ADD_1596_U199 ADD_1596_U198 ; ADD_1596_U50
g11207 nand ADD_1596_U204 ADD_1596_U203 ; ADD_1596_U51
g11208 nand ADD_1596_U209 ADD_1596_U208 ; ADD_1596_U52
g11209 nand ADD_1596_U214 ADD_1596_U213 ; ADD_1596_U53
g11210 nand ADD_1596_U219 ADD_1596_U218 ; ADD_1596_U54
g11211 nand ADD_1596_U224 ADD_1596_U223 ; ADD_1596_U55
g11212 nand ADD_1596_U234 ADD_1596_U233 ; ADD_1596_U56
g11213 nand ADD_1596_U239 ADD_1596_U238 ; ADD_1596_U57
g11214 nand ADD_1596_U244 ADD_1596_U243 ; ADD_1596_U58
g11215 nand ADD_1596_U249 ADD_1596_U248 ; ADD_1596_U59
g11216 nand ADD_1596_U254 ADD_1596_U253 ; ADD_1596_U60
g11217 nand ADD_1596_U259 ADD_1596_U258 ; ADD_1596_U61
g11218 nand ADD_1596_U264 ADD_1596_U263 ; ADD_1596_U62
g11219 nand ADD_1596_U269 ADD_1596_U268 ; ADD_1596_U63
g11220 nand ADD_1596_U274 ADD_1596_U273 ; ADD_1596_U64
g11221 nand ADD_1596_U181 ADD_1596_U180 ; ADD_1596_U65
g11222 nand ADD_1596_U186 ADD_1596_U185 ; ADD_1596_U66
g11223 nand ADD_1596_U191 ADD_1596_U190 ; ADD_1596_U67
g11224 nand ADD_1596_U196 ADD_1596_U195 ; ADD_1596_U68
g11225 nand ADD_1596_U201 ADD_1596_U200 ; ADD_1596_U69
g11226 nand ADD_1596_U206 ADD_1596_U205 ; ADD_1596_U70
g11227 nand ADD_1596_U211 ADD_1596_U210 ; ADD_1596_U71
g11228 nand ADD_1596_U216 ADD_1596_U215 ; ADD_1596_U72
g11229 nand ADD_1596_U221 ADD_1596_U220 ; ADD_1596_U73
g11230 nand ADD_1596_U231 ADD_1596_U230 ; ADD_1596_U74
g11231 nand ADD_1596_U236 ADD_1596_U235 ; ADD_1596_U75
g11232 nand ADD_1596_U241 ADD_1596_U240 ; ADD_1596_U76
g11233 nand ADD_1596_U246 ADD_1596_U245 ; ADD_1596_U77
g11234 nand ADD_1596_U251 ADD_1596_U250 ; ADD_1596_U78
g11235 nand ADD_1596_U256 ADD_1596_U255 ; ADD_1596_U79
g11236 nand ADD_1596_U261 ADD_1596_U260 ; ADD_1596_U80
g11237 nand ADD_1596_U266 ADD_1596_U265 ; ADD_1596_U81
g11238 nand ADD_1596_U271 ADD_1596_U270 ; ADD_1596_U82
g11239 nand ADD_1596_U133 ADD_1596_U132 ; ADD_1596_U83
g11240 nand ADD_1596_U129 ADD_1596_U128 ; ADD_1596_U84
g11241 nand ADD_1596_U125 ADD_1596_U124 ; ADD_1596_U85
g11242 nand ADD_1596_U121 ADD_1596_U120 ; ADD_1596_U86
g11243 nand ADD_1596_U117 ADD_1596_U116 ; ADD_1596_U87
g11244 nand ADD_1596_U113 ADD_1596_U112 ; ADD_1596_U88
g11245 nand ADD_1596_U109 ADD_1596_U108 ; ADD_1596_U89
g11246 nand ADD_1596_U105 ADD_1596_U104 ; ADD_1596_U90
g11247 not P3_ADDR_REG_1__SCAN_IN ; ADD_1596_U91
g11248 not P3_ADDR_REG_19__SCAN_IN ; ADD_1596_U92
g11249 not P1_ADDR_REG_19__SCAN_IN ; ADD_1596_U93
g11250 nand ADD_1596_U165 ADD_1596_U164 ; ADD_1596_U94
g11251 nand ADD_1596_U161 ADD_1596_U160 ; ADD_1596_U95
g11252 nand ADD_1596_U157 ADD_1596_U156 ; ADD_1596_U96
g11253 nand ADD_1596_U153 ADD_1596_U152 ; ADD_1596_U97
g11254 nand ADD_1596_U149 ADD_1596_U148 ; ADD_1596_U98
g11255 nand ADD_1596_U145 ADD_1596_U144 ; ADD_1596_U99
g11256 nand ADD_1596_U141 ADD_1596_U140 ; ADD_1596_U100
g11257 nand ADD_1596_U137 ADD_1596_U136 ; ADD_1596_U101
g11258 not ADD_1596_U9 ; ADD_1596_U102
g11259 nand ADD_1596_U102 ADD_1596_U10 ; ADD_1596_U103
g11260 nand ADD_1596_U103 ADD_1596_U91 ; ADD_1596_U104
g11261 nand ADD_1596_U9 P1_ADDR_REG_1__SCAN_IN ; ADD_1596_U105
g11262 not ADD_1596_U90 ; ADD_1596_U106
g11263 nand ADD_1596_U12 P3_ADDR_REG_2__SCAN_IN ; ADD_1596_U107
g11264 nand ADD_1596_U107 ADD_1596_U90 ; ADD_1596_U108
g11265 nand ADD_1596_U11 P1_ADDR_REG_2__SCAN_IN ; ADD_1596_U109
g11266 not ADD_1596_U89 ; ADD_1596_U110
g11267 nand ADD_1596_U14 P3_ADDR_REG_3__SCAN_IN ; ADD_1596_U111
g11268 nand ADD_1596_U111 ADD_1596_U89 ; ADD_1596_U112
g11269 nand ADD_1596_U13 P1_ADDR_REG_3__SCAN_IN ; ADD_1596_U113
g11270 not ADD_1596_U88 ; ADD_1596_U114
g11271 nand ADD_1596_U16 P3_ADDR_REG_4__SCAN_IN ; ADD_1596_U115
g11272 nand ADD_1596_U115 ADD_1596_U88 ; ADD_1596_U116
g11273 nand ADD_1596_U15 P1_ADDR_REG_4__SCAN_IN ; ADD_1596_U117
g11274 not ADD_1596_U87 ; ADD_1596_U118
g11275 nand ADD_1596_U18 P3_ADDR_REG_5__SCAN_IN ; ADD_1596_U119
g11276 nand ADD_1596_U119 ADD_1596_U87 ; ADD_1596_U120
g11277 nand ADD_1596_U17 P1_ADDR_REG_5__SCAN_IN ; ADD_1596_U121
g11278 not ADD_1596_U86 ; ADD_1596_U122
g11279 nand ADD_1596_U20 P3_ADDR_REG_6__SCAN_IN ; ADD_1596_U123
g11280 nand ADD_1596_U123 ADD_1596_U86 ; ADD_1596_U124
g11281 nand ADD_1596_U19 P1_ADDR_REG_6__SCAN_IN ; ADD_1596_U125
g11282 not ADD_1596_U85 ; ADD_1596_U126
g11283 nand ADD_1596_U22 P3_ADDR_REG_7__SCAN_IN ; ADD_1596_U127
g11284 nand ADD_1596_U127 ADD_1596_U85 ; ADD_1596_U128
g11285 nand ADD_1596_U21 P1_ADDR_REG_7__SCAN_IN ; ADD_1596_U129
g11286 not ADD_1596_U84 ; ADD_1596_U130
g11287 nand ADD_1596_U24 P3_ADDR_REG_8__SCAN_IN ; ADD_1596_U131
g11288 nand ADD_1596_U131 ADD_1596_U84 ; ADD_1596_U132
g11289 nand ADD_1596_U23 P1_ADDR_REG_8__SCAN_IN ; ADD_1596_U133
g11290 not ADD_1596_U83 ; ADD_1596_U134
g11291 nand ADD_1596_U26 P3_ADDR_REG_9__SCAN_IN ; ADD_1596_U135
g11292 nand ADD_1596_U135 ADD_1596_U83 ; ADD_1596_U136
g11293 nand ADD_1596_U25 P1_ADDR_REG_9__SCAN_IN ; ADD_1596_U137
g11294 not ADD_1596_U101 ; ADD_1596_U138
g11295 nand ADD_1596_U28 P3_ADDR_REG_10__SCAN_IN ; ADD_1596_U139
g11296 nand ADD_1596_U139 ADD_1596_U101 ; ADD_1596_U140
g11297 nand ADD_1596_U27 P1_ADDR_REG_10__SCAN_IN ; ADD_1596_U141
g11298 not ADD_1596_U100 ; ADD_1596_U142
g11299 nand ADD_1596_U30 P3_ADDR_REG_11__SCAN_IN ; ADD_1596_U143
g11300 nand ADD_1596_U143 ADD_1596_U100 ; ADD_1596_U144
g11301 nand ADD_1596_U29 P1_ADDR_REG_11__SCAN_IN ; ADD_1596_U145
g11302 not ADD_1596_U99 ; ADD_1596_U146
g11303 nand ADD_1596_U32 P3_ADDR_REG_12__SCAN_IN ; ADD_1596_U147
g11304 nand ADD_1596_U147 ADD_1596_U99 ; ADD_1596_U148
g11305 nand ADD_1596_U31 P1_ADDR_REG_12__SCAN_IN ; ADD_1596_U149
g11306 not ADD_1596_U98 ; ADD_1596_U150
g11307 nand ADD_1596_U34 P3_ADDR_REG_13__SCAN_IN ; ADD_1596_U151
g11308 nand ADD_1596_U151 ADD_1596_U98 ; ADD_1596_U152
g11309 nand ADD_1596_U33 P1_ADDR_REG_13__SCAN_IN ; ADD_1596_U153
g11310 not ADD_1596_U97 ; ADD_1596_U154
g11311 nand ADD_1596_U36 P3_ADDR_REG_14__SCAN_IN ; ADD_1596_U155
g11312 nand ADD_1596_U155 ADD_1596_U97 ; ADD_1596_U156
g11313 nand ADD_1596_U35 P1_ADDR_REG_14__SCAN_IN ; ADD_1596_U157
g11314 not ADD_1596_U96 ; ADD_1596_U158
g11315 nand ADD_1596_U38 P3_ADDR_REG_15__SCAN_IN ; ADD_1596_U159
g11316 nand ADD_1596_U159 ADD_1596_U96 ; ADD_1596_U160
g11317 nand ADD_1596_U37 P1_ADDR_REG_15__SCAN_IN ; ADD_1596_U161
g11318 not ADD_1596_U95 ; ADD_1596_U162
g11319 nand ADD_1596_U40 P3_ADDR_REG_16__SCAN_IN ; ADD_1596_U163
g11320 nand ADD_1596_U163 ADD_1596_U95 ; ADD_1596_U164
g11321 nand ADD_1596_U39 P1_ADDR_REG_16__SCAN_IN ; ADD_1596_U165
g11322 not ADD_1596_U94 ; ADD_1596_U166
g11323 nand ADD_1596_U42 P3_ADDR_REG_17__SCAN_IN ; ADD_1596_U167
g11324 nand ADD_1596_U167 ADD_1596_U94 ; ADD_1596_U168
g11325 nand ADD_1596_U41 P1_ADDR_REG_17__SCAN_IN ; ADD_1596_U169
g11326 not ADD_1596_U45 ; ADD_1596_U170
g11327 nand ADD_1596_U43 P1_ADDR_REG_18__SCAN_IN ; ADD_1596_U171
g11328 nand ADD_1596_U170 ADD_1596_U171 ; ADD_1596_U172
g11329 nand ADD_1596_U44 P3_ADDR_REG_18__SCAN_IN ; ADD_1596_U173
g11330 nand ADD_1596_U173 ADD_1596_U229 ADD_1596_U172 ; ADD_1596_U174
g11331 nand ADD_1596_U44 P3_ADDR_REG_18__SCAN_IN ; ADD_1596_U175
g11332 nand ADD_1596_U175 ADD_1596_U45 ; ADD_1596_U176
g11333 nand ADD_1596_U43 P1_ADDR_REG_18__SCAN_IN ; ADD_1596_U177
g11334 nand ADD_1596_U226 ADD_1596_U225 ADD_1596_U177 ADD_1596_U176 ; ADD_1596_U178
g11335 nand ADD_1596_U8 P1_ADDR_REG_0__SCAN_IN ; ADD_1596_U179
g11336 nand ADD_1596_U26 P3_ADDR_REG_9__SCAN_IN ; ADD_1596_U180
g11337 nand ADD_1596_U25 P1_ADDR_REG_9__SCAN_IN ; ADD_1596_U181
g11338 not ADD_1596_U65 ; ADD_1596_U182
g11339 nand ADD_1596_U134 ADD_1596_U182 ; ADD_1596_U183
g11340 nand ADD_1596_U65 ADD_1596_U83 ; ADD_1596_U184
g11341 nand ADD_1596_U24 P3_ADDR_REG_8__SCAN_IN ; ADD_1596_U185
g11342 nand ADD_1596_U23 P1_ADDR_REG_8__SCAN_IN ; ADD_1596_U186
g11343 not ADD_1596_U66 ; ADD_1596_U187
g11344 nand ADD_1596_U130 ADD_1596_U187 ; ADD_1596_U188
g11345 nand ADD_1596_U66 ADD_1596_U84 ; ADD_1596_U189
g11346 nand ADD_1596_U22 P3_ADDR_REG_7__SCAN_IN ; ADD_1596_U190
g11347 nand ADD_1596_U21 P1_ADDR_REG_7__SCAN_IN ; ADD_1596_U191
g11348 not ADD_1596_U67 ; ADD_1596_U192
g11349 nand ADD_1596_U126 ADD_1596_U192 ; ADD_1596_U193
g11350 nand ADD_1596_U67 ADD_1596_U85 ; ADD_1596_U194
g11351 nand ADD_1596_U20 P3_ADDR_REG_6__SCAN_IN ; ADD_1596_U195
g11352 nand ADD_1596_U19 P1_ADDR_REG_6__SCAN_IN ; ADD_1596_U196
g11353 not ADD_1596_U68 ; ADD_1596_U197
g11354 nand ADD_1596_U122 ADD_1596_U197 ; ADD_1596_U198
g11355 nand ADD_1596_U68 ADD_1596_U86 ; ADD_1596_U199
g11356 nand ADD_1596_U18 P3_ADDR_REG_5__SCAN_IN ; ADD_1596_U200
g11357 nand ADD_1596_U17 P1_ADDR_REG_5__SCAN_IN ; ADD_1596_U201
g11358 not ADD_1596_U69 ; ADD_1596_U202
g11359 nand ADD_1596_U118 ADD_1596_U202 ; ADD_1596_U203
g11360 nand ADD_1596_U69 ADD_1596_U87 ; ADD_1596_U204
g11361 nand ADD_1596_U16 P3_ADDR_REG_4__SCAN_IN ; ADD_1596_U205
g11362 nand ADD_1596_U15 P1_ADDR_REG_4__SCAN_IN ; ADD_1596_U206
g11363 not ADD_1596_U70 ; ADD_1596_U207
g11364 nand ADD_1596_U114 ADD_1596_U207 ; ADD_1596_U208
g11365 nand ADD_1596_U70 ADD_1596_U88 ; ADD_1596_U209
g11366 nand ADD_1596_U14 P3_ADDR_REG_3__SCAN_IN ; ADD_1596_U210
g11367 nand ADD_1596_U13 P1_ADDR_REG_3__SCAN_IN ; ADD_1596_U211
g11368 not ADD_1596_U71 ; ADD_1596_U212
g11369 nand ADD_1596_U110 ADD_1596_U212 ; ADD_1596_U213
g11370 nand ADD_1596_U71 ADD_1596_U89 ; ADD_1596_U214
g11371 nand ADD_1596_U12 P3_ADDR_REG_2__SCAN_IN ; ADD_1596_U215
g11372 nand ADD_1596_U11 P1_ADDR_REG_2__SCAN_IN ; ADD_1596_U216
g11373 not ADD_1596_U72 ; ADD_1596_U217
g11374 nand ADD_1596_U106 ADD_1596_U217 ; ADD_1596_U218
g11375 nand ADD_1596_U72 ADD_1596_U90 ; ADD_1596_U219
g11376 nand ADD_1596_U10 P3_ADDR_REG_1__SCAN_IN ; ADD_1596_U220
g11377 nand ADD_1596_U91 P1_ADDR_REG_1__SCAN_IN ; ADD_1596_U221
g11378 not ADD_1596_U73 ; ADD_1596_U222
g11379 nand ADD_1596_U222 ADD_1596_U102 ; ADD_1596_U223
g11380 nand ADD_1596_U73 ADD_1596_U9 ; ADD_1596_U224
g11381 nand ADD_1596_U93 P3_ADDR_REG_19__SCAN_IN ; ADD_1596_U225
g11382 nand ADD_1596_U92 P1_ADDR_REG_19__SCAN_IN ; ADD_1596_U226
g11383 nand ADD_1596_U93 P3_ADDR_REG_19__SCAN_IN ; ADD_1596_U227
g11384 nand ADD_1596_U92 P1_ADDR_REG_19__SCAN_IN ; ADD_1596_U228
g11385 nand ADD_1596_U228 ADD_1596_U227 ; ADD_1596_U229
g11386 nand ADD_1596_U44 P3_ADDR_REG_18__SCAN_IN ; ADD_1596_U230
g11387 nand ADD_1596_U43 P1_ADDR_REG_18__SCAN_IN ; ADD_1596_U231
g11388 not ADD_1596_U74 ; ADD_1596_U232
g11389 nand ADD_1596_U232 ADD_1596_U170 ; ADD_1596_U233
g11390 nand ADD_1596_U74 ADD_1596_U45 ; ADD_1596_U234
g11391 nand ADD_1596_U42 P3_ADDR_REG_17__SCAN_IN ; ADD_1596_U235
g11392 nand ADD_1596_U41 P1_ADDR_REG_17__SCAN_IN ; ADD_1596_U236
g11393 not ADD_1596_U75 ; ADD_1596_U237
g11394 nand ADD_1596_U166 ADD_1596_U237 ; ADD_1596_U238
g11395 nand ADD_1596_U75 ADD_1596_U94 ; ADD_1596_U239
g11396 nand ADD_1596_U40 P3_ADDR_REG_16__SCAN_IN ; ADD_1596_U240
g11397 nand ADD_1596_U39 P1_ADDR_REG_16__SCAN_IN ; ADD_1596_U241
g11398 not ADD_1596_U76 ; ADD_1596_U242
g11399 nand ADD_1596_U162 ADD_1596_U242 ; ADD_1596_U243
g11400 nand ADD_1596_U76 ADD_1596_U95 ; ADD_1596_U244
g11401 nand ADD_1596_U38 P3_ADDR_REG_15__SCAN_IN ; ADD_1596_U245
g11402 nand ADD_1596_U37 P1_ADDR_REG_15__SCAN_IN ; ADD_1596_U246
g11403 not ADD_1596_U77 ; ADD_1596_U247
g11404 nand ADD_1596_U158 ADD_1596_U247 ; ADD_1596_U248
g11405 nand ADD_1596_U77 ADD_1596_U96 ; ADD_1596_U249
g11406 nand ADD_1596_U36 P3_ADDR_REG_14__SCAN_IN ; ADD_1596_U250
g11407 nand ADD_1596_U35 P1_ADDR_REG_14__SCAN_IN ; ADD_1596_U251
g11408 not ADD_1596_U78 ; ADD_1596_U252
g11409 nand ADD_1596_U154 ADD_1596_U252 ; ADD_1596_U253
g11410 nand ADD_1596_U78 ADD_1596_U97 ; ADD_1596_U254
g11411 nand ADD_1596_U34 P3_ADDR_REG_13__SCAN_IN ; ADD_1596_U255
g11412 nand ADD_1596_U33 P1_ADDR_REG_13__SCAN_IN ; ADD_1596_U256
g11413 not ADD_1596_U79 ; ADD_1596_U257
g11414 nand ADD_1596_U150 ADD_1596_U257 ; ADD_1596_U258
g11415 nand ADD_1596_U79 ADD_1596_U98 ; ADD_1596_U259
g11416 nand ADD_1596_U32 P3_ADDR_REG_12__SCAN_IN ; ADD_1596_U260
g11417 nand ADD_1596_U31 P1_ADDR_REG_12__SCAN_IN ; ADD_1596_U261
g11418 not ADD_1596_U80 ; ADD_1596_U262
g11419 nand ADD_1596_U146 ADD_1596_U262 ; ADD_1596_U263
g11420 nand ADD_1596_U80 ADD_1596_U99 ; ADD_1596_U264
g11421 nand ADD_1596_U30 P3_ADDR_REG_11__SCAN_IN ; ADD_1596_U265
g11422 nand ADD_1596_U29 P1_ADDR_REG_11__SCAN_IN ; ADD_1596_U266
g11423 not ADD_1596_U81 ; ADD_1596_U267
g11424 nand ADD_1596_U142 ADD_1596_U267 ; ADD_1596_U268
g11425 nand ADD_1596_U81 ADD_1596_U100 ; ADD_1596_U269
g11426 nand ADD_1596_U28 P3_ADDR_REG_10__SCAN_IN ; ADD_1596_U270
g11427 nand ADD_1596_U27 P1_ADDR_REG_10__SCAN_IN ; ADD_1596_U271
g11428 not ADD_1596_U82 ; ADD_1596_U272
g11429 nand ADD_1596_U138 ADD_1596_U272 ; ADD_1596_U273
g11430 nand ADD_1596_U82 ADD_1596_U101 ; ADD_1596_U274
g11431 not P2_ADDR_REG_19__SCAN_IN ; LT_1601_21_U6
g11432 not P1_REG3_REG_3__SCAN_IN ; P1_ADD_99_U4
g11433 and P1_ADD_99_U102 P1_REG3_REG_28__SCAN_IN P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U5
g11434 not P1_REG3_REG_4__SCAN_IN ; P1_ADD_99_U6
g11435 nand P1_REG3_REG_4__SCAN_IN P1_REG3_REG_3__SCAN_IN ; P1_ADD_99_U7
g11436 not P1_REG3_REG_5__SCAN_IN ; P1_ADD_99_U8
g11437 nand P1_ADD_99_U80 P1_REG3_REG_5__SCAN_IN ; P1_ADD_99_U9
g11438 not P1_REG3_REG_6__SCAN_IN ; P1_ADD_99_U10
g11439 nand P1_ADD_99_U81 P1_REG3_REG_6__SCAN_IN ; P1_ADD_99_U11
g11440 not P1_REG3_REG_7__SCAN_IN ; P1_ADD_99_U12
g11441 nand P1_ADD_99_U82 P1_REG3_REG_7__SCAN_IN ; P1_ADD_99_U13
g11442 not P1_REG3_REG_8__SCAN_IN ; P1_ADD_99_U14
g11443 not P1_REG3_REG_9__SCAN_IN ; P1_ADD_99_U15
g11444 nand P1_ADD_99_U83 P1_REG3_REG_8__SCAN_IN ; P1_ADD_99_U16
g11445 nand P1_ADD_99_U84 P1_REG3_REG_9__SCAN_IN ; P1_ADD_99_U17
g11446 not P1_REG3_REG_10__SCAN_IN ; P1_ADD_99_U18
g11447 nand P1_ADD_99_U85 P1_REG3_REG_10__SCAN_IN ; P1_ADD_99_U19
g11448 not P1_REG3_REG_11__SCAN_IN ; P1_ADD_99_U20
g11449 nand P1_ADD_99_U86 P1_REG3_REG_11__SCAN_IN ; P1_ADD_99_U21
g11450 not P1_REG3_REG_12__SCAN_IN ; P1_ADD_99_U22
g11451 nand P1_ADD_99_U87 P1_REG3_REG_12__SCAN_IN ; P1_ADD_99_U23
g11452 not P1_REG3_REG_13__SCAN_IN ; P1_ADD_99_U24
g11453 nand P1_ADD_99_U88 P1_REG3_REG_13__SCAN_IN ; P1_ADD_99_U25
g11454 not P1_REG3_REG_14__SCAN_IN ; P1_ADD_99_U26
g11455 nand P1_ADD_99_U89 P1_REG3_REG_14__SCAN_IN ; P1_ADD_99_U27
g11456 not P1_REG3_REG_15__SCAN_IN ; P1_ADD_99_U28
g11457 nand P1_ADD_99_U90 P1_REG3_REG_15__SCAN_IN ; P1_ADD_99_U29
g11458 not P1_REG3_REG_16__SCAN_IN ; P1_ADD_99_U30
g11459 nand P1_ADD_99_U91 P1_REG3_REG_16__SCAN_IN ; P1_ADD_99_U31
g11460 not P1_REG3_REG_17__SCAN_IN ; P1_ADD_99_U32
g11461 nand P1_ADD_99_U92 P1_REG3_REG_17__SCAN_IN ; P1_ADD_99_U33
g11462 not P1_REG3_REG_18__SCAN_IN ; P1_ADD_99_U34
g11463 nand P1_ADD_99_U93 P1_REG3_REG_18__SCAN_IN ; P1_ADD_99_U35
g11464 not P1_REG3_REG_19__SCAN_IN ; P1_ADD_99_U36
g11465 nand P1_ADD_99_U94 P1_REG3_REG_19__SCAN_IN ; P1_ADD_99_U37
g11466 not P1_REG3_REG_20__SCAN_IN ; P1_ADD_99_U38
g11467 nand P1_ADD_99_U95 P1_REG3_REG_20__SCAN_IN ; P1_ADD_99_U39
g11468 not P1_REG3_REG_21__SCAN_IN ; P1_ADD_99_U40
g11469 nand P1_ADD_99_U96 P1_REG3_REG_21__SCAN_IN ; P1_ADD_99_U41
g11470 not P1_REG3_REG_22__SCAN_IN ; P1_ADD_99_U42
g11471 nand P1_ADD_99_U97 P1_REG3_REG_22__SCAN_IN ; P1_ADD_99_U43
g11472 not P1_REG3_REG_23__SCAN_IN ; P1_ADD_99_U44
g11473 nand P1_ADD_99_U98 P1_REG3_REG_23__SCAN_IN ; P1_ADD_99_U45
g11474 not P1_REG3_REG_24__SCAN_IN ; P1_ADD_99_U46
g11475 nand P1_ADD_99_U99 P1_REG3_REG_24__SCAN_IN ; P1_ADD_99_U47
g11476 not P1_REG3_REG_25__SCAN_IN ; P1_ADD_99_U48
g11477 nand P1_ADD_99_U100 P1_REG3_REG_25__SCAN_IN ; P1_ADD_99_U49
g11478 not P1_REG3_REG_26__SCAN_IN ; P1_ADD_99_U50
g11479 nand P1_ADD_99_U101 P1_REG3_REG_26__SCAN_IN ; P1_ADD_99_U51
g11480 not P1_REG3_REG_28__SCAN_IN ; P1_ADD_99_U52
g11481 not P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U53
g11482 nand P1_ADD_99_U105 P1_ADD_99_U104 ; P1_ADD_99_U54
g11483 nand P1_ADD_99_U107 P1_ADD_99_U106 ; P1_ADD_99_U55
g11484 nand P1_ADD_99_U109 P1_ADD_99_U108 ; P1_ADD_99_U56
g11485 nand P1_ADD_99_U111 P1_ADD_99_U110 ; P1_ADD_99_U57
g11486 nand P1_ADD_99_U113 P1_ADD_99_U112 ; P1_ADD_99_U58
g11487 nand P1_ADD_99_U115 P1_ADD_99_U114 ; P1_ADD_99_U59
g11488 nand P1_ADD_99_U117 P1_ADD_99_U116 ; P1_ADD_99_U60
g11489 nand P1_ADD_99_U119 P1_ADD_99_U118 ; P1_ADD_99_U61
g11490 nand P1_ADD_99_U121 P1_ADD_99_U120 ; P1_ADD_99_U62
g11491 nand P1_ADD_99_U123 P1_ADD_99_U122 ; P1_ADD_99_U63
g11492 nand P1_ADD_99_U125 P1_ADD_99_U124 ; P1_ADD_99_U64
g11493 nand P1_ADD_99_U127 P1_ADD_99_U126 ; P1_ADD_99_U65
g11494 nand P1_ADD_99_U129 P1_ADD_99_U128 ; P1_ADD_99_U66
g11495 nand P1_ADD_99_U131 P1_ADD_99_U130 ; P1_ADD_99_U67
g11496 nand P1_ADD_99_U133 P1_ADD_99_U132 ; P1_ADD_99_U68
g11497 nand P1_ADD_99_U135 P1_ADD_99_U134 ; P1_ADD_99_U69
g11498 nand P1_ADD_99_U137 P1_ADD_99_U136 ; P1_ADD_99_U70
g11499 nand P1_ADD_99_U139 P1_ADD_99_U138 ; P1_ADD_99_U71
g11500 nand P1_ADD_99_U141 P1_ADD_99_U140 ; P1_ADD_99_U72
g11501 nand P1_ADD_99_U143 P1_ADD_99_U142 ; P1_ADD_99_U73
g11502 nand P1_ADD_99_U145 P1_ADD_99_U144 ; P1_ADD_99_U74
g11503 nand P1_ADD_99_U147 P1_ADD_99_U146 ; P1_ADD_99_U75
g11504 nand P1_ADD_99_U149 P1_ADD_99_U148 ; P1_ADD_99_U76
g11505 nand P1_ADD_99_U151 P1_ADD_99_U150 ; P1_ADD_99_U77
g11506 nand P1_ADD_99_U153 P1_ADD_99_U152 ; P1_ADD_99_U78
g11507 nand P1_ADD_99_U102 P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U79
g11508 not P1_ADD_99_U7 ; P1_ADD_99_U80
g11509 not P1_ADD_99_U9 ; P1_ADD_99_U81
g11510 not P1_ADD_99_U11 ; P1_ADD_99_U82
g11511 not P1_ADD_99_U13 ; P1_ADD_99_U83
g11512 not P1_ADD_99_U16 ; P1_ADD_99_U84
g11513 not P1_ADD_99_U17 ; P1_ADD_99_U85
g11514 not P1_ADD_99_U19 ; P1_ADD_99_U86
g11515 not P1_ADD_99_U21 ; P1_ADD_99_U87
g11516 not P1_ADD_99_U23 ; P1_ADD_99_U88
g11517 not P1_ADD_99_U25 ; P1_ADD_99_U89
g11518 not P1_ADD_99_U27 ; P1_ADD_99_U90
g11519 not P1_ADD_99_U29 ; P1_ADD_99_U91
g11520 not P1_ADD_99_U31 ; P1_ADD_99_U92
g11521 not P1_ADD_99_U33 ; P1_ADD_99_U93
g11522 not P1_ADD_99_U35 ; P1_ADD_99_U94
g11523 not P1_ADD_99_U37 ; P1_ADD_99_U95
g11524 not P1_ADD_99_U39 ; P1_ADD_99_U96
g11525 not P1_ADD_99_U41 ; P1_ADD_99_U97
g11526 not P1_ADD_99_U43 ; P1_ADD_99_U98
g11527 not P1_ADD_99_U45 ; P1_ADD_99_U99
g11528 not P1_ADD_99_U47 ; P1_ADD_99_U100
g11529 not P1_ADD_99_U49 ; P1_ADD_99_U101
g11530 not P1_ADD_99_U51 ; P1_ADD_99_U102
g11531 not P1_ADD_99_U79 ; P1_ADD_99_U103
g11532 nand P1_ADD_99_U16 P1_REG3_REG_9__SCAN_IN ; P1_ADD_99_U104
g11533 nand P1_ADD_99_U84 P1_ADD_99_U15 ; P1_ADD_99_U105
g11534 nand P1_ADD_99_U13 P1_REG3_REG_8__SCAN_IN ; P1_ADD_99_U106
g11535 nand P1_ADD_99_U83 P1_ADD_99_U14 ; P1_ADD_99_U107
g11536 nand P1_ADD_99_U11 P1_REG3_REG_7__SCAN_IN ; P1_ADD_99_U108
g11537 nand P1_ADD_99_U82 P1_ADD_99_U12 ; P1_ADD_99_U109
g11538 nand P1_ADD_99_U9 P1_REG3_REG_6__SCAN_IN ; P1_ADD_99_U110
g11539 nand P1_ADD_99_U81 P1_ADD_99_U10 ; P1_ADD_99_U111
g11540 nand P1_ADD_99_U7 P1_REG3_REG_5__SCAN_IN ; P1_ADD_99_U112
g11541 nand P1_ADD_99_U80 P1_ADD_99_U8 ; P1_ADD_99_U113
g11542 nand P1_ADD_99_U4 P1_REG3_REG_4__SCAN_IN ; P1_ADD_99_U114
g11543 nand P1_ADD_99_U6 P1_REG3_REG_3__SCAN_IN ; P1_ADD_99_U115
g11544 nand P1_ADD_99_U79 P1_REG3_REG_28__SCAN_IN ; P1_ADD_99_U116
g11545 nand P1_ADD_99_U103 P1_ADD_99_U52 ; P1_ADD_99_U117
g11546 nand P1_ADD_99_U51 P1_REG3_REG_27__SCAN_IN ; P1_ADD_99_U118
g11547 nand P1_ADD_99_U102 P1_ADD_99_U53 ; P1_ADD_99_U119
g11548 nand P1_ADD_99_U49 P1_REG3_REG_26__SCAN_IN ; P1_ADD_99_U120
g11549 nand P1_ADD_99_U101 P1_ADD_99_U50 ; P1_ADD_99_U121
g11550 nand P1_ADD_99_U47 P1_REG3_REG_25__SCAN_IN ; P1_ADD_99_U122
g11551 nand P1_ADD_99_U100 P1_ADD_99_U48 ; P1_ADD_99_U123
g11552 nand P1_ADD_99_U45 P1_REG3_REG_24__SCAN_IN ; P1_ADD_99_U124
g11553 nand P1_ADD_99_U99 P1_ADD_99_U46 ; P1_ADD_99_U125
g11554 nand P1_ADD_99_U43 P1_REG3_REG_23__SCAN_IN ; P1_ADD_99_U126
g11555 nand P1_ADD_99_U98 P1_ADD_99_U44 ; P1_ADD_99_U127
g11556 nand P1_ADD_99_U41 P1_REG3_REG_22__SCAN_IN ; P1_ADD_99_U128
g11557 nand P1_ADD_99_U97 P1_ADD_99_U42 ; P1_ADD_99_U129
g11558 nand P1_ADD_99_U39 P1_REG3_REG_21__SCAN_IN ; P1_ADD_99_U130
g11559 nand P1_ADD_99_U96 P1_ADD_99_U40 ; P1_ADD_99_U131
g11560 nand P1_ADD_99_U37 P1_REG3_REG_20__SCAN_IN ; P1_ADD_99_U132
g11561 nand P1_ADD_99_U95 P1_ADD_99_U38 ; P1_ADD_99_U133
g11562 nand P1_ADD_99_U35 P1_REG3_REG_19__SCAN_IN ; P1_ADD_99_U134
g11563 nand P1_ADD_99_U94 P1_ADD_99_U36 ; P1_ADD_99_U135
g11564 nand P1_ADD_99_U33 P1_REG3_REG_18__SCAN_IN ; P1_ADD_99_U136
g11565 nand P1_ADD_99_U93 P1_ADD_99_U34 ; P1_ADD_99_U137
g11566 nand P1_ADD_99_U31 P1_REG3_REG_17__SCAN_IN ; P1_ADD_99_U138
g11567 nand P1_ADD_99_U92 P1_ADD_99_U32 ; P1_ADD_99_U139
g11568 nand P1_ADD_99_U29 P1_REG3_REG_16__SCAN_IN ; P1_ADD_99_U140
g11569 nand P1_ADD_99_U91 P1_ADD_99_U30 ; P1_ADD_99_U141
g11570 nand P1_ADD_99_U27 P1_REG3_REG_15__SCAN_IN ; P1_ADD_99_U142
g11571 nand P1_ADD_99_U90 P1_ADD_99_U28 ; P1_ADD_99_U143
g11572 nand P1_ADD_99_U25 P1_REG3_REG_14__SCAN_IN ; P1_ADD_99_U144
g11573 nand P1_ADD_99_U89 P1_ADD_99_U26 ; P1_ADD_99_U145
g11574 nand P1_ADD_99_U23 P1_REG3_REG_13__SCAN_IN ; P1_ADD_99_U146
g11575 nand P1_ADD_99_U88 P1_ADD_99_U24 ; P1_ADD_99_U147
g11576 nand P1_ADD_99_U21 P1_REG3_REG_12__SCAN_IN ; P1_ADD_99_U148
g11577 nand P1_ADD_99_U87 P1_ADD_99_U22 ; P1_ADD_99_U149
g11578 nand P1_ADD_99_U19 P1_REG3_REG_11__SCAN_IN ; P1_ADD_99_U150
g11579 nand P1_ADD_99_U86 P1_ADD_99_U20 ; P1_ADD_99_U151
g11580 nand P1_ADD_99_U17 P1_REG3_REG_10__SCAN_IN ; P1_ADD_99_U152
g11581 nand P1_ADD_99_U85 P1_ADD_99_U18 ; P1_ADD_99_U153
g11582 and P1_R1105_U95 P1_R1105_U94 ; P1_R1105_U4
g11583 and P1_R1105_U96 P1_R1105_U97 ; P1_R1105_U5
g11584 and P1_R1105_U113 P1_R1105_U112 ; P1_R1105_U6
g11585 and P1_R1105_U155 P1_R1105_U154 ; P1_R1105_U7
g11586 and P1_R1105_U164 P1_R1105_U163 ; P1_R1105_U8
g11587 and P1_R1105_U182 P1_R1105_U181 ; P1_R1105_U9
g11588 and P1_R1105_U218 P1_R1105_U215 ; P1_R1105_U10
g11589 and P1_R1105_U211 P1_R1105_U208 ; P1_R1105_U11
g11590 and P1_R1105_U202 P1_R1105_U199 ; P1_R1105_U12
g11591 and P1_R1105_U196 P1_R1105_U192 ; P1_R1105_U13
g11592 and P1_R1105_U151 P1_R1105_U148 ; P1_R1105_U14
g11593 and P1_R1105_U143 P1_R1105_U140 ; P1_R1105_U15
g11594 and P1_R1105_U129 P1_R1105_U126 ; P1_R1105_U16
g11595 not P1_REG2_REG_6__SCAN_IN ; P1_R1105_U17
g11596 not P1_U3475 ; P1_R1105_U18
g11597 not P1_U3478 ; P1_R1105_U19
g11598 nand P1_U3475 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U20
g11599 not P1_REG2_REG_7__SCAN_IN ; P1_R1105_U21
g11600 not P1_REG2_REG_4__SCAN_IN ; P1_R1105_U22
g11601 not P1_U3469 ; P1_R1105_U23
g11602 not P1_U3472 ; P1_R1105_U24
g11603 not P1_REG2_REG_2__SCAN_IN ; P1_R1105_U25
g11604 not P1_U3463 ; P1_R1105_U26
g11605 not P1_REG2_REG_0__SCAN_IN ; P1_R1105_U27
g11606 not P1_U3454 ; P1_R1105_U28
g11607 nand P1_U3454 P1_REG2_REG_0__SCAN_IN ; P1_R1105_U29
g11608 not P1_REG2_REG_3__SCAN_IN ; P1_R1105_U30
g11609 not P1_U3466 ; P1_R1105_U31
g11610 nand P1_U3469 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U32
g11611 not P1_REG2_REG_5__SCAN_IN ; P1_R1105_U33
g11612 not P1_REG2_REG_8__SCAN_IN ; P1_R1105_U34
g11613 not P1_U3481 ; P1_R1105_U35
g11614 not P1_U3484 ; P1_R1105_U36
g11615 not P1_REG2_REG_9__SCAN_IN ; P1_R1105_U37
g11616 nand P1_R1105_U49 P1_R1105_U121 ; P1_R1105_U38
g11617 nand P1_R1105_U110 P1_R1105_U108 P1_R1105_U109 ; P1_R1105_U39
g11618 nand P1_R1105_U98 P1_R1105_U99 ; P1_R1105_U40
g11619 nand P1_U3460 P1_REG2_REG_1__SCAN_IN ; P1_R1105_U41
g11620 nand P1_R1105_U136 P1_R1105_U134 P1_R1105_U135 ; P1_R1105_U42
g11621 nand P1_R1105_U132 P1_R1105_U131 ; P1_R1105_U43
g11622 not P1_REG2_REG_16__SCAN_IN ; P1_R1105_U44
g11623 not P1_U3505 ; P1_R1105_U45
g11624 not P1_U3508 ; P1_R1105_U46
g11625 nand P1_U3505 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U47
g11626 not P1_REG2_REG_17__SCAN_IN ; P1_R1105_U48
g11627 nand P1_U3481 P1_REG2_REG_8__SCAN_IN ; P1_R1105_U49
g11628 not P1_REG2_REG_10__SCAN_IN ; P1_R1105_U50
g11629 not P1_U3487 ; P1_R1105_U51
g11630 not P1_REG2_REG_12__SCAN_IN ; P1_R1105_U52
g11631 not P1_U3493 ; P1_R1105_U53
g11632 not P1_REG2_REG_11__SCAN_IN ; P1_R1105_U54
g11633 not P1_U3490 ; P1_R1105_U55
g11634 nand P1_U3490 P1_REG2_REG_11__SCAN_IN ; P1_R1105_U56
g11635 not P1_REG2_REG_13__SCAN_IN ; P1_R1105_U57
g11636 not P1_U3496 ; P1_R1105_U58
g11637 not P1_REG2_REG_14__SCAN_IN ; P1_R1105_U59
g11638 not P1_U3499 ; P1_R1105_U60
g11639 not P1_REG2_REG_15__SCAN_IN ; P1_R1105_U61
g11640 not P1_U3502 ; P1_R1105_U62
g11641 not P1_REG2_REG_18__SCAN_IN ; P1_R1105_U63
g11642 not P1_U3511 ; P1_R1105_U64
g11643 nand P1_R1105_U186 P1_R1105_U185 P1_R1105_U187 ; P1_R1105_U65
g11644 nand P1_R1105_U179 P1_R1105_U178 ; P1_R1105_U66
g11645 nand P1_R1105_U56 P1_R1105_U204 ; P1_R1105_U67
g11646 nand P1_R1105_U259 P1_R1105_U258 ; P1_R1105_U68
g11647 nand P1_R1105_U308 P1_R1105_U307 ; P1_R1105_U69
g11648 nand P1_R1105_U231 P1_R1105_U230 ; P1_R1105_U70
g11649 nand P1_R1105_U236 P1_R1105_U235 ; P1_R1105_U71
g11650 nand P1_R1105_U243 P1_R1105_U242 ; P1_R1105_U72
g11651 nand P1_R1105_U250 P1_R1105_U249 ; P1_R1105_U73
g11652 nand P1_R1105_U255 P1_R1105_U254 ; P1_R1105_U74
g11653 nand P1_R1105_U271 P1_R1105_U270 ; P1_R1105_U75
g11654 nand P1_R1105_U278 P1_R1105_U277 ; P1_R1105_U76
g11655 nand P1_R1105_U285 P1_R1105_U284 ; P1_R1105_U77
g11656 nand P1_R1105_U292 P1_R1105_U291 ; P1_R1105_U78
g11657 nand P1_R1105_U299 P1_R1105_U298 ; P1_R1105_U79
g11658 nand P1_R1105_U304 P1_R1105_U303 ; P1_R1105_U80
g11659 nand P1_R1105_U117 P1_R1105_U116 P1_R1105_U118 ; P1_R1105_U81
g11660 nand P1_R1105_U133 P1_R1105_U145 ; P1_R1105_U82
g11661 nand P1_R1105_U41 P1_R1105_U152 ; P1_R1105_U83
g11662 not P1_U3452 ; P1_R1105_U84
g11663 not P1_REG2_REG_19__SCAN_IN ; P1_R1105_U85
g11664 nand P1_R1105_U175 P1_R1105_U174 ; P1_R1105_U86
g11665 nand P1_R1105_U171 P1_R1105_U170 ; P1_R1105_U87
g11666 nand P1_R1105_U161 P1_R1105_U160 ; P1_R1105_U88
g11667 not P1_R1105_U32 ; P1_R1105_U89
g11668 nand P1_U3484 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U90
g11669 nand P1_U3493 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U91
g11670 not P1_R1105_U56 ; P1_R1105_U92
g11671 not P1_R1105_U49 ; P1_R1105_U93
g11672 or P1_U3472 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U94
g11673 or P1_U3469 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U95
g11674 or P1_U3466 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U96
g11675 or P1_U3463 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U97
g11676 not P1_R1105_U29 ; P1_R1105_U98
g11677 or P1_U3460 P1_REG2_REG_1__SCAN_IN ; P1_R1105_U99
g11678 not P1_R1105_U40 ; P1_R1105_U100
g11679 not P1_R1105_U41 ; P1_R1105_U101
g11680 nand P1_R1105_U40 P1_R1105_U41 ; P1_R1105_U102
g11681 nand P1_U3463 P1_R1105_U96 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U103
g11682 nand P1_R1105_U5 P1_R1105_U102 ; P1_R1105_U104
g11683 nand P1_U3466 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U105
g11684 nand P1_R1105_U105 P1_R1105_U103 P1_R1105_U104 ; P1_R1105_U106
g11685 nand P1_R1105_U33 P1_R1105_U32 ; P1_R1105_U107
g11686 nand P1_U3472 P1_R1105_U107 ; P1_R1105_U108
g11687 nand P1_R1105_U4 P1_R1105_U106 ; P1_R1105_U109
g11688 nand P1_R1105_U89 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U110
g11689 not P1_R1105_U39 ; P1_R1105_U111
g11690 or P1_U3478 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U112
g11691 or P1_U3475 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U113
g11692 not P1_R1105_U20 ; P1_R1105_U114
g11693 nand P1_R1105_U21 P1_R1105_U20 ; P1_R1105_U115
g11694 nand P1_U3478 P1_R1105_U115 ; P1_R1105_U116
g11695 nand P1_R1105_U114 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U117
g11696 nand P1_R1105_U6 P1_R1105_U39 ; P1_R1105_U118
g11697 not P1_R1105_U81 ; P1_R1105_U119
g11698 or P1_U3481 P1_REG2_REG_8__SCAN_IN ; P1_R1105_U120
g11699 nand P1_R1105_U120 P1_R1105_U81 ; P1_R1105_U121
g11700 not P1_R1105_U38 ; P1_R1105_U122
g11701 or P1_U3484 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U123
g11702 or P1_U3475 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U124
g11703 nand P1_R1105_U124 P1_R1105_U39 ; P1_R1105_U125
g11704 nand P1_R1105_U238 P1_R1105_U237 P1_R1105_U20 P1_R1105_U125 ; P1_R1105_U126
g11705 nand P1_R1105_U111 P1_R1105_U20 ; P1_R1105_U127
g11706 nand P1_U3478 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U128
g11707 nand P1_R1105_U128 P1_R1105_U6 P1_R1105_U127 ; P1_R1105_U129
g11708 or P1_U3475 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U130
g11709 nand P1_R1105_U101 P1_R1105_U97 ; P1_R1105_U131
g11710 nand P1_U3463 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U132
g11711 not P1_R1105_U43 ; P1_R1105_U133
g11712 nand P1_R1105_U100 P1_R1105_U5 ; P1_R1105_U134
g11713 nand P1_R1105_U43 P1_R1105_U96 ; P1_R1105_U135
g11714 nand P1_U3466 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U136
g11715 not P1_R1105_U42 ; P1_R1105_U137
g11716 or P1_U3469 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U138
g11717 nand P1_R1105_U138 P1_R1105_U42 ; P1_R1105_U139
g11718 nand P1_R1105_U245 P1_R1105_U244 P1_R1105_U32 P1_R1105_U139 ; P1_R1105_U140
g11719 nand P1_R1105_U137 P1_R1105_U32 ; P1_R1105_U141
g11720 nand P1_U3472 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U142
g11721 nand P1_R1105_U142 P1_R1105_U4 P1_R1105_U141 ; P1_R1105_U143
g11722 or P1_U3469 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U144
g11723 nand P1_R1105_U100 P1_R1105_U97 ; P1_R1105_U145
g11724 not P1_R1105_U82 ; P1_R1105_U146
g11725 nand P1_U3466 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U147
g11726 nand P1_R1105_U41 P1_R1105_U40 P1_R1105_U257 P1_R1105_U256 ; P1_R1105_U148
g11727 nand P1_R1105_U41 P1_R1105_U40 ; P1_R1105_U149
g11728 nand P1_U3463 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U150
g11729 nand P1_R1105_U150 P1_R1105_U97 P1_R1105_U149 ; P1_R1105_U151
g11730 or P1_U3460 P1_REG2_REG_1__SCAN_IN ; P1_R1105_U152
g11731 not P1_R1105_U83 ; P1_R1105_U153
g11732 or P1_U3484 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U154
g11733 or P1_U3487 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U155
g11734 nand P1_R1105_U93 P1_R1105_U7 ; P1_R1105_U156
g11735 nand P1_U3487 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U157
g11736 nand P1_R1105_U157 P1_R1105_U90 P1_R1105_U156 ; P1_R1105_U158
g11737 or P1_U3487 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U159
g11738 nand P1_R1105_U120 P1_R1105_U7 P1_R1105_U81 ; P1_R1105_U160
g11739 nand P1_R1105_U159 P1_R1105_U158 ; P1_R1105_U161
g11740 not P1_R1105_U88 ; P1_R1105_U162
g11741 or P1_U3496 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U163
g11742 or P1_U3493 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U164
g11743 nand P1_R1105_U92 P1_R1105_U8 ; P1_R1105_U165
g11744 nand P1_U3496 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U166
g11745 nand P1_R1105_U166 P1_R1105_U91 P1_R1105_U165 ; P1_R1105_U167
g11746 or P1_U3490 P1_REG2_REG_11__SCAN_IN ; P1_R1105_U168
g11747 or P1_U3496 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U169
g11748 nand P1_R1105_U168 P1_R1105_U8 P1_R1105_U88 ; P1_R1105_U170
g11749 nand P1_R1105_U169 P1_R1105_U167 ; P1_R1105_U171
g11750 not P1_R1105_U87 ; P1_R1105_U172
g11751 or P1_U3499 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U173
g11752 nand P1_R1105_U173 P1_R1105_U87 ; P1_R1105_U174
g11753 nand P1_U3499 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U175
g11754 not P1_R1105_U86 ; P1_R1105_U176
g11755 or P1_U3502 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U177
g11756 nand P1_R1105_U177 P1_R1105_U86 ; P1_R1105_U178
g11757 nand P1_U3502 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U179
g11758 not P1_R1105_U66 ; P1_R1105_U180
g11759 or P1_U3508 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U181
g11760 or P1_U3505 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U182
g11761 not P1_R1105_U47 ; P1_R1105_U183
g11762 nand P1_R1105_U48 P1_R1105_U47 ; P1_R1105_U184
g11763 nand P1_U3508 P1_R1105_U184 ; P1_R1105_U185
g11764 nand P1_R1105_U183 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U186
g11765 nand P1_R1105_U9 P1_R1105_U66 ; P1_R1105_U187
g11766 not P1_R1105_U65 ; P1_R1105_U188
g11767 or P1_U3511 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U189
g11768 nand P1_R1105_U189 P1_R1105_U65 ; P1_R1105_U190
g11769 nand P1_U3511 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U191
g11770 nand P1_R1105_U261 P1_R1105_U260 P1_R1105_U191 P1_R1105_U190 ; P1_R1105_U192
g11771 nand P1_U3511 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U193
g11772 nand P1_R1105_U188 P1_R1105_U193 ; P1_R1105_U194
g11773 or P1_U3511 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U195
g11774 nand P1_R1105_U195 P1_R1105_U264 P1_R1105_U194 ; P1_R1105_U196
g11775 or P1_U3505 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U197
g11776 nand P1_R1105_U197 P1_R1105_U66 ; P1_R1105_U198
g11777 nand P1_R1105_U273 P1_R1105_U272 P1_R1105_U47 P1_R1105_U198 ; P1_R1105_U199
g11778 nand P1_R1105_U180 P1_R1105_U47 ; P1_R1105_U200
g11779 nand P1_U3508 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U201
g11780 nand P1_R1105_U201 P1_R1105_U9 P1_R1105_U200 ; P1_R1105_U202
g11781 or P1_U3505 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U203
g11782 nand P1_R1105_U168 P1_R1105_U88 ; P1_R1105_U204
g11783 not P1_R1105_U67 ; P1_R1105_U205
g11784 or P1_U3493 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U206
g11785 nand P1_R1105_U206 P1_R1105_U67 ; P1_R1105_U207
g11786 nand P1_R1105_U294 P1_R1105_U293 P1_R1105_U91 P1_R1105_U207 ; P1_R1105_U208
g11787 nand P1_R1105_U205 P1_R1105_U91 ; P1_R1105_U209
g11788 nand P1_U3496 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U210
g11789 nand P1_R1105_U210 P1_R1105_U8 P1_R1105_U209 ; P1_R1105_U211
g11790 or P1_U3493 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U212
g11791 or P1_U3484 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U213
g11792 nand P1_R1105_U213 P1_R1105_U38 ; P1_R1105_U214
g11793 nand P1_R1105_U306 P1_R1105_U305 P1_R1105_U90 P1_R1105_U214 ; P1_R1105_U215
g11794 nand P1_R1105_U122 P1_R1105_U90 ; P1_R1105_U216
g11795 nand P1_U3487 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U217
g11796 nand P1_R1105_U217 P1_R1105_U7 P1_R1105_U216 ; P1_R1105_U218
g11797 nand P1_R1105_U123 P1_R1105_U90 ; P1_R1105_U219
g11798 nand P1_R1105_U120 P1_R1105_U49 ; P1_R1105_U220
g11799 nand P1_R1105_U130 P1_R1105_U20 ; P1_R1105_U221
g11800 nand P1_R1105_U144 P1_R1105_U32 ; P1_R1105_U222
g11801 nand P1_R1105_U147 P1_R1105_U96 ; P1_R1105_U223
g11802 nand P1_R1105_U203 P1_R1105_U47 ; P1_R1105_U224
g11803 nand P1_R1105_U212 P1_R1105_U91 ; P1_R1105_U225
g11804 nand P1_R1105_U168 P1_R1105_U56 ; P1_R1105_U226
g11805 nand P1_U3484 P1_R1105_U37 ; P1_R1105_U227
g11806 nand P1_R1105_U36 P1_REG2_REG_9__SCAN_IN ; P1_R1105_U228
g11807 nand P1_R1105_U228 P1_R1105_U227 ; P1_R1105_U229
g11808 nand P1_R1105_U219 P1_R1105_U38 ; P1_R1105_U230
g11809 nand P1_R1105_U229 P1_R1105_U122 ; P1_R1105_U231
g11810 nand P1_U3481 P1_R1105_U34 ; P1_R1105_U232
g11811 nand P1_R1105_U35 P1_REG2_REG_8__SCAN_IN ; P1_R1105_U233
g11812 nand P1_R1105_U233 P1_R1105_U232 ; P1_R1105_U234
g11813 nand P1_R1105_U220 P1_R1105_U81 ; P1_R1105_U235
g11814 nand P1_R1105_U119 P1_R1105_U234 ; P1_R1105_U236
g11815 nand P1_U3478 P1_R1105_U21 ; P1_R1105_U237
g11816 nand P1_R1105_U19 P1_REG2_REG_7__SCAN_IN ; P1_R1105_U238
g11817 nand P1_U3475 P1_R1105_U17 ; P1_R1105_U239
g11818 nand P1_R1105_U18 P1_REG2_REG_6__SCAN_IN ; P1_R1105_U240
g11819 nand P1_R1105_U240 P1_R1105_U239 ; P1_R1105_U241
g11820 nand P1_R1105_U221 P1_R1105_U39 ; P1_R1105_U242
g11821 nand P1_R1105_U241 P1_R1105_U111 ; P1_R1105_U243
g11822 nand P1_U3472 P1_R1105_U33 ; P1_R1105_U244
g11823 nand P1_R1105_U24 P1_REG2_REG_5__SCAN_IN ; P1_R1105_U245
g11824 nand P1_U3469 P1_R1105_U22 ; P1_R1105_U246
g11825 nand P1_R1105_U23 P1_REG2_REG_4__SCAN_IN ; P1_R1105_U247
g11826 nand P1_R1105_U247 P1_R1105_U246 ; P1_R1105_U248
g11827 nand P1_R1105_U222 P1_R1105_U42 ; P1_R1105_U249
g11828 nand P1_R1105_U248 P1_R1105_U137 ; P1_R1105_U250
g11829 nand P1_U3466 P1_R1105_U30 ; P1_R1105_U251
g11830 nand P1_R1105_U31 P1_REG2_REG_3__SCAN_IN ; P1_R1105_U252
g11831 nand P1_R1105_U252 P1_R1105_U251 ; P1_R1105_U253
g11832 nand P1_R1105_U223 P1_R1105_U82 ; P1_R1105_U254
g11833 nand P1_R1105_U146 P1_R1105_U253 ; P1_R1105_U255
g11834 nand P1_U3463 P1_R1105_U25 ; P1_R1105_U256
g11835 nand P1_R1105_U26 P1_REG2_REG_2__SCAN_IN ; P1_R1105_U257
g11836 nand P1_R1105_U98 P1_R1105_U83 ; P1_R1105_U258
g11837 nand P1_R1105_U153 P1_R1105_U29 ; P1_R1105_U259
g11838 nand P1_U3452 P1_R1105_U85 ; P1_R1105_U260
g11839 nand P1_R1105_U84 P1_REG2_REG_19__SCAN_IN ; P1_R1105_U261
g11840 nand P1_U3452 P1_R1105_U85 ; P1_R1105_U262
g11841 nand P1_R1105_U84 P1_REG2_REG_19__SCAN_IN ; P1_R1105_U263
g11842 nand P1_R1105_U263 P1_R1105_U262 ; P1_R1105_U264
g11843 nand P1_U3511 P1_R1105_U63 ; P1_R1105_U265
g11844 nand P1_R1105_U64 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U266
g11845 nand P1_U3511 P1_R1105_U63 ; P1_R1105_U267
g11846 nand P1_R1105_U64 P1_REG2_REG_18__SCAN_IN ; P1_R1105_U268
g11847 nand P1_R1105_U268 P1_R1105_U267 ; P1_R1105_U269
g11848 nand P1_R1105_U266 P1_R1105_U265 P1_R1105_U65 ; P1_R1105_U270
g11849 nand P1_R1105_U269 P1_R1105_U188 ; P1_R1105_U271
g11850 nand P1_U3508 P1_R1105_U48 ; P1_R1105_U272
g11851 nand P1_R1105_U46 P1_REG2_REG_17__SCAN_IN ; P1_R1105_U273
g11852 nand P1_U3505 P1_R1105_U44 ; P1_R1105_U274
g11853 nand P1_R1105_U45 P1_REG2_REG_16__SCAN_IN ; P1_R1105_U275
g11854 nand P1_R1105_U275 P1_R1105_U274 ; P1_R1105_U276
g11855 nand P1_R1105_U224 P1_R1105_U66 ; P1_R1105_U277
g11856 nand P1_R1105_U276 P1_R1105_U180 ; P1_R1105_U278
g11857 nand P1_U3502 P1_R1105_U61 ; P1_R1105_U279
g11858 nand P1_R1105_U62 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U280
g11859 nand P1_U3502 P1_R1105_U61 ; P1_R1105_U281
g11860 nand P1_R1105_U62 P1_REG2_REG_15__SCAN_IN ; P1_R1105_U282
g11861 nand P1_R1105_U282 P1_R1105_U281 ; P1_R1105_U283
g11862 nand P1_R1105_U280 P1_R1105_U279 P1_R1105_U86 ; P1_R1105_U284
g11863 nand P1_R1105_U176 P1_R1105_U283 ; P1_R1105_U285
g11864 nand P1_U3499 P1_R1105_U59 ; P1_R1105_U286
g11865 nand P1_R1105_U60 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U287
g11866 nand P1_U3499 P1_R1105_U59 ; P1_R1105_U288
g11867 nand P1_R1105_U60 P1_REG2_REG_14__SCAN_IN ; P1_R1105_U289
g11868 nand P1_R1105_U289 P1_R1105_U288 ; P1_R1105_U290
g11869 nand P1_R1105_U287 P1_R1105_U286 P1_R1105_U87 ; P1_R1105_U291
g11870 nand P1_R1105_U172 P1_R1105_U290 ; P1_R1105_U292
g11871 nand P1_U3496 P1_R1105_U57 ; P1_R1105_U293
g11872 nand P1_R1105_U58 P1_REG2_REG_13__SCAN_IN ; P1_R1105_U294
g11873 nand P1_U3493 P1_R1105_U52 ; P1_R1105_U295
g11874 nand P1_R1105_U53 P1_REG2_REG_12__SCAN_IN ; P1_R1105_U296
g11875 nand P1_R1105_U296 P1_R1105_U295 ; P1_R1105_U297
g11876 nand P1_R1105_U225 P1_R1105_U67 ; P1_R1105_U298
g11877 nand P1_R1105_U297 P1_R1105_U205 ; P1_R1105_U299
g11878 nand P1_U3490 P1_R1105_U54 ; P1_R1105_U300
g11879 nand P1_R1105_U55 P1_REG2_REG_11__SCAN_IN ; P1_R1105_U301
g11880 nand P1_R1105_U301 P1_R1105_U300 ; P1_R1105_U302
g11881 nand P1_R1105_U226 P1_R1105_U88 ; P1_R1105_U303
g11882 nand P1_R1105_U162 P1_R1105_U302 ; P1_R1105_U304
g11883 nand P1_U3487 P1_R1105_U50 ; P1_R1105_U305
g11884 nand P1_R1105_U51 P1_REG2_REG_10__SCAN_IN ; P1_R1105_U306
g11885 nand P1_U3454 P1_R1105_U27 ; P1_R1105_U307
g11886 nand P1_R1105_U28 P1_REG2_REG_0__SCAN_IN ; P1_R1105_U308
g11887 and P1_SUB_88_U227 P1_SUB_88_U38 ; P1_SUB_88_U6
g11888 and P1_SUB_88_U225 P1_SUB_88_U192 ; P1_SUB_88_U7
g11889 and P1_SUB_88_U224 P1_SUB_88_U35 ; P1_SUB_88_U8
g11890 and P1_SUB_88_U223 P1_SUB_88_U36 ; P1_SUB_88_U9
g11891 and P1_SUB_88_U221 P1_SUB_88_U195 ; P1_SUB_88_U10
g11892 and P1_SUB_88_U220 P1_SUB_88_U34 ; P1_SUB_88_U11
g11893 and P1_SUB_88_U219 P1_SUB_88_U197 ; P1_SUB_88_U12
g11894 and P1_SUB_88_U217 P1_SUB_88_U198 ; P1_SUB_88_U13
g11895 and P1_SUB_88_U216 P1_SUB_88_U172 ; P1_SUB_88_U14
g11896 and P1_SUB_88_U215 P1_SUB_88_U200 ; P1_SUB_88_U15
g11897 and P1_SUB_88_U213 P1_SUB_88_U201 ; P1_SUB_88_U16
g11898 and P1_SUB_88_U212 P1_SUB_88_U169 ; P1_SUB_88_U17
g11899 and P1_SUB_88_U211 P1_SUB_88_U167 ; P1_SUB_88_U18
g11900 and P1_SUB_88_U209 P1_SUB_88_U204 ; P1_SUB_88_U19
g11901 and P1_SUB_88_U208 P1_SUB_88_U33 ; P1_SUB_88_U20
g11902 and P1_SUB_88_U207 P1_SUB_88_U27 ; P1_SUB_88_U21
g11903 and P1_SUB_88_U190 P1_SUB_88_U180 ; P1_SUB_88_U22
g11904 and P1_SUB_88_U189 P1_SUB_88_U29 ; P1_SUB_88_U23
g11905 and P1_SUB_88_U188 P1_SUB_88_U30 ; P1_SUB_88_U24
g11906 and P1_SUB_88_U186 P1_SUB_88_U183 ; P1_SUB_88_U25
g11907 and P1_SUB_88_U185 P1_SUB_88_U28 ; P1_SUB_88_U26
g11908 or P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_2__SCAN_IN ; P1_SUB_88_U27
g11909 nand P1_SUB_88_U44 P1_SUB_88_U230 P1_SUB_88_U43 ; P1_SUB_88_U28
g11910 nand P1_SUB_88_U45 P1_SUB_88_U230 ; P1_SUB_88_U29
g11911 nand P1_SUB_88_U46 P1_SUB_88_U181 ; P1_SUB_88_U30
g11912 not P1_IR_REG_7__SCAN_IN ; P1_SUB_88_U31
g11913 not P1_IR_REG_3__SCAN_IN ; P1_SUB_88_U32
g11914 nand P1_SUB_88_U56 P1_SUB_88_U51 ; P1_SUB_88_U33
g11915 nand P1_SUB_88_U130 P1_SUB_88_U129 P1_SUB_88_U128 P1_SUB_88_U127 ; P1_SUB_88_U34
g11916 nand P1_SUB_88_U156 P1_SUB_88_U184 ; P1_SUB_88_U35
g11917 nand P1_SUB_88_U157 P1_SUB_88_U193 ; P1_SUB_88_U36
g11918 not P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U37
g11919 nand P1_SUB_88_U158 P1_SUB_88_U184 ; P1_SUB_88_U38
g11920 not P1_IR_REG_11__SCAN_IN ; P1_SUB_88_U39
g11921 nand P1_SUB_88_U247 P1_SUB_88_U246 ; P1_SUB_88_U40
g11922 nand P1_SUB_88_U237 P1_SUB_88_U236 ; P1_SUB_88_U41
g11923 nand P1_SUB_88_U241 P1_SUB_88_U240 ; P1_SUB_88_U42
g11924 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U43
g11925 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN ; P1_SUB_88_U44
g11926 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U45
g11927 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U46
g11928 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U47
g11929 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U48
g11930 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U49
g11931 nor P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U50
g11932 and P1_SUB_88_U50 P1_SUB_88_U49 P1_SUB_88_U48 P1_SUB_88_U47 ; P1_SUB_88_U51
g11933 nor P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U52
g11934 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_27__SCAN_IN P1_IR_REG_28__SCAN_IN P1_IR_REG_29__SCAN_IN ; P1_SUB_88_U53
g11935 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U54
g11936 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U55
g11937 and P1_SUB_88_U55 P1_SUB_88_U54 P1_SUB_88_U53 P1_SUB_88_U52 ; P1_SUB_88_U56
g11938 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U57
g11939 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U58
g11940 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U59
g11941 nor P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U60
g11942 and P1_SUB_88_U60 P1_SUB_88_U59 P1_SUB_88_U58 P1_SUB_88_U57 ; P1_SUB_88_U61
g11943 nor P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U62
g11944 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_27__SCAN_IN P1_IR_REG_28__SCAN_IN ; P1_SUB_88_U63
g11945 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U64
g11946 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U65
g11947 and P1_SUB_88_U65 P1_SUB_88_U64 P1_SUB_88_U63 P1_SUB_88_U62 ; P1_SUB_88_U66
g11948 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U67
g11949 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U68
g11950 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U69
g11951 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U70
g11952 and P1_SUB_88_U70 P1_SUB_88_U69 P1_SUB_88_U68 P1_SUB_88_U67 ; P1_SUB_88_U71
g11953 nor P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U72
g11954 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_26__SCAN_IN P1_IR_REG_27__SCAN_IN ; P1_SUB_88_U73
g11955 nor P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U74
g11956 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U75
g11957 and P1_SUB_88_U75 P1_SUB_88_U74 P1_SUB_88_U73 P1_SUB_88_U72 ; P1_SUB_88_U76
g11958 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U77
g11959 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U78
g11960 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U79
g11961 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U80
g11962 and P1_SUB_88_U80 P1_SUB_88_U79 P1_SUB_88_U78 P1_SUB_88_U77 ; P1_SUB_88_U81
g11963 nor P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U82
g11964 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U83
g11965 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U84
g11966 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U85
g11967 and P1_SUB_88_U85 P1_SUB_88_U84 P1_SUB_88_U83 P1_SUB_88_U82 ; P1_SUB_88_U86
g11968 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U87
g11969 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U88
g11970 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U89
g11971 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U90
g11972 and P1_SUB_88_U90 P1_SUB_88_U89 P1_SUB_88_U88 P1_SUB_88_U87 ; P1_SUB_88_U91
g11973 nor P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U92
g11974 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U93
g11975 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U94
g11976 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U95
g11977 and P1_SUB_88_U95 P1_SUB_88_U94 P1_SUB_88_U93 P1_SUB_88_U92 ; P1_SUB_88_U96
g11978 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U97
g11979 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U98
g11980 nor P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U99
g11981 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U100
g11982 and P1_SUB_88_U100 P1_SUB_88_U99 P1_SUB_88_U98 P1_SUB_88_U97 ; P1_SUB_88_U101
g11983 nor P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN P1_IR_REG_24__SCAN_IN ; P1_SUB_88_U102
g11984 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U103
g11985 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U104
g11986 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U105
g11987 and P1_SUB_88_U105 P1_SUB_88_U104 P1_SUB_88_U103 P1_SUB_88_U102 ; P1_SUB_88_U106
g11988 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U107
g11989 nor P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U108
g11990 nor P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U109
g11991 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U110
g11992 and P1_SUB_88_U110 P1_SUB_88_U109 P1_SUB_88_U108 P1_SUB_88_U107 ; P1_SUB_88_U111
g11993 nor P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN P1_IR_REG_23__SCAN_IN ; P1_SUB_88_U112
g11994 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_24__SCAN_IN ; P1_SUB_88_U113
g11995 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U114
g11996 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U115
g11997 and P1_SUB_88_U115 P1_SUB_88_U114 P1_SUB_88_U113 P1_SUB_88_U112 ; P1_SUB_88_U116
g11998 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U117
g11999 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U118
g12000 nor P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U119
g12001 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U120
g12002 and P1_SUB_88_U120 P1_SUB_88_U119 P1_SUB_88_U118 P1_SUB_88_U117 ; P1_SUB_88_U121
g12003 nor P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U122
g12004 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_23__SCAN_IN ; P1_SUB_88_U123
g12005 nor P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U124
g12006 nor P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U125
g12007 and P1_SUB_88_U125 P1_SUB_88_U124 P1_SUB_88_U123 P1_SUB_88_U122 ; P1_SUB_88_U126
g12008 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U127
g12009 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U128
g12010 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U129
g12011 nor P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U130
g12012 nor P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U131
g12013 nor P1_IR_REG_19__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U132
g12014 nor P1_IR_REG_21__SCAN_IN P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U133
g12015 and P1_SUB_88_U132 P1_SUB_88_U131 P1_SUB_88_U133 ; P1_SUB_88_U134
g12016 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U135
g12017 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U136
g12018 and P1_SUB_88_U136 P1_SUB_88_U135 ; P1_SUB_88_U137
g12019 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U138
g12020 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_20__SCAN_IN P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U139
g12021 nor P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U140
g12022 and P1_SUB_88_U140 P1_SUB_88_U139 ; P1_SUB_88_U141
g12023 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U142
g12024 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U143
g12025 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U144
g12026 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U145
g12027 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U146
g12028 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U147
g12029 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U148
g12030 nor P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U149
g12031 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U150
g12032 nor P1_IR_REG_5__SCAN_IN P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U151
g12033 nor P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U152
g12034 nor P1_IR_REG_1__SCAN_IN P1_IR_REG_15__SCAN_IN P1_IR_REG_16__SCAN_IN P1_IR_REG_17__SCAN_IN P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U153
g12035 nor P1_IR_REG_0__SCAN_IN P1_IR_REG_2__SCAN_IN P1_IR_REG_3__SCAN_IN P1_IR_REG_4__SCAN_IN P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U154
g12036 nor P1_IR_REG_6__SCAN_IN P1_IR_REG_7__SCAN_IN P1_IR_REG_8__SCAN_IN P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U155
g12037 nor P1_IR_REG_9__SCAN_IN P1_IR_REG_10__SCAN_IN P1_IR_REG_11__SCAN_IN P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U156
g12038 nor P1_IR_REG_13__SCAN_IN P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U157
g12039 nor P1_IR_REG_9__SCAN_IN P1_IR_REG_10__SCAN_IN ; P1_SUB_88_U158
g12040 not P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U159
g12041 and P1_SUB_88_U233 P1_SUB_88_U232 ; P1_SUB_88_U160
g12042 not P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U161
g12043 and P1_SUB_88_U235 P1_SUB_88_U234 ; P1_SUB_88_U162
g12044 not P1_IR_REG_31__SCAN_IN ; P1_SUB_88_U163
g12045 not P1_IR_REG_30__SCAN_IN ; P1_SUB_88_U164
g12046 and P1_SUB_88_U239 P1_SUB_88_U238 ; P1_SUB_88_U165
g12047 not P1_IR_REG_27__SCAN_IN ; P1_SUB_88_U166
g12048 nand P1_SUB_88_U96 P1_SUB_88_U91 ; P1_SUB_88_U167
g12049 not P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U168
g12050 nand P1_SUB_88_U116 P1_SUB_88_U111 ; P1_SUB_88_U169
g12051 and P1_SUB_88_U243 P1_SUB_88_U242 ; P1_SUB_88_U170
g12052 not P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U171
g12053 nand P1_SUB_88_U144 P1_SUB_88_U143 P1_SUB_88_U145 P1_SUB_88_U147 P1_SUB_88_U146 ; P1_SUB_88_U172
g12054 and P1_SUB_88_U245 P1_SUB_88_U244 ; P1_SUB_88_U173
g12055 not P1_IR_REG_1__SCAN_IN ; P1_SUB_88_U174
g12056 not P1_IR_REG_0__SCAN_IN ; P1_SUB_88_U175
g12057 not P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U176
g12058 and P1_SUB_88_U249 P1_SUB_88_U248 ; P1_SUB_88_U177
g12059 not P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U178
g12060 and P1_SUB_88_U251 P1_SUB_88_U250 ; P1_SUB_88_U179
g12061 nand P1_SUB_88_U230 P1_SUB_88_U32 ; P1_SUB_88_U180
g12062 not P1_SUB_88_U29 ; P1_SUB_88_U181
g12063 not P1_SUB_88_U30 ; P1_SUB_88_U182
g12064 nand P1_SUB_88_U182 P1_SUB_88_U31 ; P1_SUB_88_U183
g12065 not P1_SUB_88_U28 ; P1_SUB_88_U184
g12066 nand P1_SUB_88_U183 P1_IR_REG_8__SCAN_IN ; P1_SUB_88_U185
g12067 nand P1_SUB_88_U30 P1_IR_REG_7__SCAN_IN ; P1_SUB_88_U186
g12068 nand P1_SUB_88_U181 P1_SUB_88_U161 ; P1_SUB_88_U187
g12069 nand P1_SUB_88_U187 P1_IR_REG_6__SCAN_IN ; P1_SUB_88_U188
g12070 nand P1_SUB_88_U180 P1_IR_REG_4__SCAN_IN ; P1_SUB_88_U189
g12071 nand P1_SUB_88_U27 P1_IR_REG_3__SCAN_IN ; P1_SUB_88_U190
g12072 not P1_SUB_88_U38 ; P1_SUB_88_U191
g12073 nand P1_SUB_88_U191 P1_SUB_88_U39 ; P1_SUB_88_U192
g12074 not P1_SUB_88_U35 ; P1_SUB_88_U193
g12075 not P1_SUB_88_U36 ; P1_SUB_88_U194
g12076 nand P1_SUB_88_U194 P1_SUB_88_U37 ; P1_SUB_88_U195
g12077 not P1_SUB_88_U34 ; P1_SUB_88_U196
g12078 nand P1_SUB_88_U155 P1_SUB_88_U154 P1_SUB_88_U153 P1_SUB_88_U152 ; P1_SUB_88_U197
g12079 nand P1_SUB_88_U151 P1_SUB_88_U150 P1_SUB_88_U149 P1_SUB_88_U148 ; P1_SUB_88_U198
g12080 not P1_SUB_88_U172 ; P1_SUB_88_U199
g12081 nand P1_SUB_88_U134 P1_SUB_88_U196 ; P1_SUB_88_U200
g12082 nand P1_SUB_88_U126 P1_SUB_88_U121 ; P1_SUB_88_U201
g12083 not P1_SUB_88_U169 ; P1_SUB_88_U202
g12084 not P1_SUB_88_U167 ; P1_SUB_88_U203
g12085 nand P1_SUB_88_U66 P1_SUB_88_U61 ; P1_SUB_88_U204
g12086 not P1_SUB_88_U33 ; P1_SUB_88_U205
g12087 or P1_IR_REG_0__SCAN_IN P1_IR_REG_1__SCAN_IN ; P1_SUB_88_U206
g12088 nand P1_SUB_88_U206 P1_IR_REG_2__SCAN_IN ; P1_SUB_88_U207
g12089 nand P1_SUB_88_U204 P1_IR_REG_29__SCAN_IN ; P1_SUB_88_U208
g12090 nand P1_SUB_88_U229 P1_IR_REG_28__SCAN_IN ; P1_SUB_88_U209
g12091 nand P1_SUB_88_U106 P1_SUB_88_U101 ; P1_SUB_88_U210
g12092 nand P1_SUB_88_U210 P1_IR_REG_26__SCAN_IN ; P1_SUB_88_U211
g12093 nand P1_SUB_88_U201 P1_IR_REG_24__SCAN_IN ; P1_SUB_88_U212
g12094 nand P1_SUB_88_U200 P1_IR_REG_23__SCAN_IN ; P1_SUB_88_U213
g12095 nand P1_SUB_88_U142 P1_SUB_88_U141 P1_SUB_88_U138 P1_SUB_88_U137 ; P1_SUB_88_U214
g12096 nand P1_SUB_88_U214 P1_IR_REG_22__SCAN_IN ; P1_SUB_88_U215
g12097 nand P1_SUB_88_U198 P1_IR_REG_20__SCAN_IN ; P1_SUB_88_U216
g12098 nand P1_SUB_88_U197 P1_IR_REG_19__SCAN_IN ; P1_SUB_88_U217
g12099 nand P1_SUB_88_U196 P1_SUB_88_U176 ; P1_SUB_88_U218
g12100 nand P1_SUB_88_U218 P1_IR_REG_18__SCAN_IN ; P1_SUB_88_U219
g12101 nand P1_SUB_88_U195 P1_IR_REG_16__SCAN_IN ; P1_SUB_88_U220
g12102 nand P1_SUB_88_U36 P1_IR_REG_15__SCAN_IN ; P1_SUB_88_U221
g12103 nand P1_SUB_88_U193 P1_SUB_88_U178 ; P1_SUB_88_U222
g12104 nand P1_SUB_88_U222 P1_IR_REG_14__SCAN_IN ; P1_SUB_88_U223
g12105 nand P1_SUB_88_U192 P1_IR_REG_12__SCAN_IN ; P1_SUB_88_U224
g12106 nand P1_SUB_88_U38 P1_IR_REG_11__SCAN_IN ; P1_SUB_88_U225
g12107 nand P1_SUB_88_U184 P1_SUB_88_U159 ; P1_SUB_88_U226
g12108 nand P1_SUB_88_U226 P1_IR_REG_10__SCAN_IN ; P1_SUB_88_U227
g12109 nand P1_SUB_88_U205 P1_SUB_88_U164 ; P1_SUB_88_U228
g12110 nand P1_SUB_88_U76 P1_SUB_88_U71 ; P1_SUB_88_U229
g12111 not P1_SUB_88_U27 ; P1_SUB_88_U230
g12112 nand P1_SUB_88_U86 P1_SUB_88_U81 ; P1_SUB_88_U231
g12113 nand P1_SUB_88_U28 P1_IR_REG_9__SCAN_IN ; P1_SUB_88_U232
g12114 nand P1_SUB_88_U184 P1_SUB_88_U159 ; P1_SUB_88_U233
g12115 nand P1_SUB_88_U29 P1_IR_REG_5__SCAN_IN ; P1_SUB_88_U234
g12116 nand P1_SUB_88_U181 P1_SUB_88_U161 ; P1_SUB_88_U235
g12117 nand P1_SUB_88_U228 P1_SUB_88_U163 ; P1_SUB_88_U236
g12118 nand P1_SUB_88_U205 P1_SUB_88_U164 P1_IR_REG_31__SCAN_IN ; P1_SUB_88_U237
g12119 nand P1_SUB_88_U33 P1_IR_REG_30__SCAN_IN ; P1_SUB_88_U238
g12120 nand P1_SUB_88_U205 P1_SUB_88_U164 ; P1_SUB_88_U239
g12121 nand P1_SUB_88_U203 P1_IR_REG_27__SCAN_IN ; P1_SUB_88_U240
g12122 nand P1_SUB_88_U231 P1_SUB_88_U166 ; P1_SUB_88_U241
g12123 nand P1_SUB_88_U169 P1_IR_REG_25__SCAN_IN ; P1_SUB_88_U242
g12124 nand P1_SUB_88_U202 P1_SUB_88_U168 ; P1_SUB_88_U243
g12125 nand P1_SUB_88_U172 P1_IR_REG_21__SCAN_IN ; P1_SUB_88_U244
g12126 nand P1_SUB_88_U199 P1_SUB_88_U171 ; P1_SUB_88_U245
g12127 nand P1_SUB_88_U175 P1_IR_REG_1__SCAN_IN ; P1_SUB_88_U246
g12128 nand P1_SUB_88_U174 P1_IR_REG_0__SCAN_IN ; P1_SUB_88_U247
g12129 nand P1_SUB_88_U34 P1_IR_REG_17__SCAN_IN ; P1_SUB_88_U248
g12130 nand P1_SUB_88_U196 P1_SUB_88_U176 ; P1_SUB_88_U249
g12131 nand P1_SUB_88_U35 P1_IR_REG_13__SCAN_IN ; P1_SUB_88_U250
g12132 nand P1_SUB_88_U193 P1_SUB_88_U178 ; P1_SUB_88_U251
g12133 not P1_U3059 ; P1_R1309_U6
g12134 not P1_U3056 ; P1_R1309_U7
g12135 and P1_R1309_U10 P1_R1309_U9 ; P1_R1309_U8
g12136 nand P1_U3056 P1_R1309_U6 ; P1_R1309_U9
g12137 nand P1_U3059 P1_R1309_U7 ; P1_R1309_U10
g12138 and P1_R1282_U135 P1_R1282_U35 ; P1_R1282_U6
g12139 and P1_R1282_U133 P1_R1282_U36 ; P1_R1282_U7
g12140 and P1_R1282_U132 P1_R1282_U37 ; P1_R1282_U8
g12141 and P1_R1282_U131 P1_R1282_U38 ; P1_R1282_U9
g12142 and P1_R1282_U129 P1_R1282_U39 ; P1_R1282_U10
g12143 and P1_R1282_U128 P1_R1282_U40 ; P1_R1282_U11
g12144 and P1_R1282_U127 P1_R1282_U41 ; P1_R1282_U12
g12145 and P1_R1282_U125 P1_R1282_U42 ; P1_R1282_U13
g12146 and P1_R1282_U123 P1_R1282_U43 ; P1_R1282_U14
g12147 and P1_R1282_U121 P1_R1282_U44 ; P1_R1282_U15
g12148 and P1_R1282_U119 P1_R1282_U45 ; P1_R1282_U16
g12149 and P1_R1282_U117 P1_R1282_U46 ; P1_R1282_U17
g12150 and P1_R1282_U115 P1_R1282_U25 ; P1_R1282_U18
g12151 and P1_R1282_U113 P1_R1282_U67 ; P1_R1282_U19
g12152 and P1_R1282_U98 P1_R1282_U26 ; P1_R1282_U20
g12153 and P1_R1282_U97 P1_R1282_U27 ; P1_R1282_U21
g12154 and P1_R1282_U96 P1_R1282_U28 ; P1_R1282_U22
g12155 and P1_R1282_U94 P1_R1282_U29 ; P1_R1282_U23
g12156 and P1_R1282_U93 P1_R1282_U30 ; P1_R1282_U24
g12157 or P1_U3461 P1_U3456 P1_U3464 ; P1_R1282_U25
g12158 nand P1_R1282_U87 P1_R1282_U34 ; P1_R1282_U26
g12159 nand P1_R1282_U88 P1_R1282_U33 ; P1_R1282_U27
g12160 nand P1_R1282_U57 P1_R1282_U89 ; P1_R1282_U28
g12161 nand P1_R1282_U90 P1_R1282_U32 ; P1_R1282_U29
g12162 nand P1_R1282_U91 P1_R1282_U31 ; P1_R1282_U30
g12163 not P1_U3482 ; P1_R1282_U31
g12164 not P1_U3479 ; P1_R1282_U32
g12165 not P1_U3470 ; P1_R1282_U33
g12166 not P1_U3467 ; P1_R1282_U34
g12167 nand P1_R1282_U58 P1_R1282_U92 ; P1_R1282_U35
g12168 nand P1_R1282_U99 P1_R1282_U55 ; P1_R1282_U36
g12169 nand P1_R1282_U100 P1_R1282_U54 ; P1_R1282_U37
g12170 nand P1_R1282_U59 P1_R1282_U101 ; P1_R1282_U38
g12171 nand P1_R1282_U102 P1_R1282_U53 ; P1_R1282_U39
g12172 nand P1_R1282_U103 P1_R1282_U52 ; P1_R1282_U40
g12173 nand P1_R1282_U60 P1_R1282_U104 ; P1_R1282_U41
g12174 nand P1_R1282_U61 P1_R1282_U105 ; P1_R1282_U42
g12175 nand P1_R1282_U106 P1_R1282_U77 P1_R1282_U51 ; P1_R1282_U43
g12176 nand P1_R1282_U107 P1_R1282_U75 P1_R1282_U50 ; P1_R1282_U44
g12177 nand P1_R1282_U108 P1_R1282_U73 P1_R1282_U49 ; P1_R1282_U45
g12178 nand P1_R1282_U109 P1_R1282_U71 P1_R1282_U48 ; P1_R1282_U46
g12179 not P1_U4027 ; P1_R1282_U47
g12180 not P1_U4017 ; P1_R1282_U48
g12181 not P1_U4019 ; P1_R1282_U49
g12182 not P1_U4021 ; P1_R1282_U50
g12183 not P1_U4023 ; P1_R1282_U51
g12184 not P1_U3506 ; P1_R1282_U52
g12185 not P1_U3503 ; P1_R1282_U53
g12186 not P1_U3494 ; P1_R1282_U54
g12187 not P1_U3491 ; P1_R1282_U55
g12188 nand P1_R1282_U153 P1_R1282_U152 ; P1_R1282_U56
g12189 nor P1_U3473 P1_U3476 ; P1_R1282_U57
g12190 nor P1_U3488 P1_U3485 ; P1_R1282_U58
g12191 nor P1_U3497 P1_U3500 ; P1_R1282_U59
g12192 nor P1_U3509 P1_U3512 ; P1_R1282_U60
g12193 nor P1_U3514 P1_U4025 ; P1_R1282_U61
g12194 not P1_U3485 ; P1_R1282_U62
g12195 and P1_R1282_U137 P1_R1282_U136 ; P1_R1282_U63
g12196 not P1_U3473 ; P1_R1282_U64
g12197 and P1_R1282_U139 P1_R1282_U138 ; P1_R1282_U65
g12198 not P1_U4026 ; P1_R1282_U66
g12199 nand P1_R1282_U110 P1_R1282_U69 P1_R1282_U47 ; P1_R1282_U67
g12200 and P1_R1282_U141 P1_R1282_U140 ; P1_R1282_U68
g12201 not P1_U4028 ; P1_R1282_U69
g12202 and P1_R1282_U143 P1_R1282_U142 ; P1_R1282_U70
g12203 not P1_U4018 ; P1_R1282_U71
g12204 and P1_R1282_U145 P1_R1282_U144 ; P1_R1282_U72
g12205 not P1_U4020 ; P1_R1282_U73
g12206 and P1_R1282_U147 P1_R1282_U146 ; P1_R1282_U74
g12207 not P1_U4022 ; P1_R1282_U75
g12208 and P1_R1282_U149 P1_R1282_U148 ; P1_R1282_U76
g12209 not P1_U4024 ; P1_R1282_U77
g12210 and P1_R1282_U151 P1_R1282_U150 ; P1_R1282_U78
g12211 not P1_U3461 ; P1_R1282_U79
g12212 not P1_U3456 ; P1_R1282_U80
g12213 not P1_U3514 ; P1_R1282_U81
g12214 and P1_R1282_U155 P1_R1282_U154 ; P1_R1282_U82
g12215 not P1_U3509 ; P1_R1282_U83
g12216 and P1_R1282_U157 P1_R1282_U156 ; P1_R1282_U84
g12217 not P1_U3497 ; P1_R1282_U85
g12218 and P1_R1282_U159 P1_R1282_U158 ; P1_R1282_U86
g12219 not P1_R1282_U25 ; P1_R1282_U87
g12220 not P1_R1282_U26 ; P1_R1282_U88
g12221 not P1_R1282_U27 ; P1_R1282_U89
g12222 not P1_R1282_U28 ; P1_R1282_U90
g12223 not P1_R1282_U29 ; P1_R1282_U91
g12224 not P1_R1282_U30 ; P1_R1282_U92
g12225 nand P1_U3482 P1_R1282_U29 ; P1_R1282_U93
g12226 nand P1_U3479 P1_R1282_U28 ; P1_R1282_U94
g12227 nand P1_R1282_U89 P1_R1282_U64 ; P1_R1282_U95
g12228 nand P1_U3476 P1_R1282_U95 ; P1_R1282_U96
g12229 nand P1_U3470 P1_R1282_U26 ; P1_R1282_U97
g12230 nand P1_U3467 P1_R1282_U25 ; P1_R1282_U98
g12231 not P1_R1282_U35 ; P1_R1282_U99
g12232 not P1_R1282_U36 ; P1_R1282_U100
g12233 not P1_R1282_U37 ; P1_R1282_U101
g12234 not P1_R1282_U38 ; P1_R1282_U102
g12235 not P1_R1282_U39 ; P1_R1282_U103
g12236 not P1_R1282_U40 ; P1_R1282_U104
g12237 not P1_R1282_U41 ; P1_R1282_U105
g12238 not P1_R1282_U42 ; P1_R1282_U106
g12239 not P1_R1282_U43 ; P1_R1282_U107
g12240 not P1_R1282_U44 ; P1_R1282_U108
g12241 not P1_R1282_U45 ; P1_R1282_U109
g12242 not P1_R1282_U46 ; P1_R1282_U110
g12243 not P1_R1282_U67 ; P1_R1282_U111
g12244 nand P1_R1282_U110 P1_R1282_U69 ; P1_R1282_U112
g12245 nand P1_U4027 P1_R1282_U112 ; P1_R1282_U113
g12246 or P1_U3461 P1_U3456 ; P1_R1282_U114
g12247 nand P1_U3464 P1_R1282_U114 ; P1_R1282_U115
g12248 nand P1_R1282_U109 P1_R1282_U71 ; P1_R1282_U116
g12249 nand P1_U4017 P1_R1282_U116 ; P1_R1282_U117
g12250 nand P1_R1282_U108 P1_R1282_U73 ; P1_R1282_U118
g12251 nand P1_U4019 P1_R1282_U118 ; P1_R1282_U119
g12252 nand P1_R1282_U107 P1_R1282_U75 ; P1_R1282_U120
g12253 nand P1_U4021 P1_R1282_U120 ; P1_R1282_U121
g12254 nand P1_R1282_U106 P1_R1282_U77 ; P1_R1282_U122
g12255 nand P1_U4023 P1_R1282_U122 ; P1_R1282_U123
g12256 nand P1_R1282_U105 P1_R1282_U81 ; P1_R1282_U124
g12257 nand P1_U4025 P1_R1282_U124 ; P1_R1282_U125
g12258 nand P1_R1282_U104 P1_R1282_U83 ; P1_R1282_U126
g12259 nand P1_U3512 P1_R1282_U126 ; P1_R1282_U127
g12260 nand P1_U3506 P1_R1282_U39 ; P1_R1282_U128
g12261 nand P1_U3503 P1_R1282_U38 ; P1_R1282_U129
g12262 nand P1_R1282_U101 P1_R1282_U85 ; P1_R1282_U130
g12263 nand P1_U3500 P1_R1282_U130 ; P1_R1282_U131
g12264 nand P1_U3494 P1_R1282_U36 ; P1_R1282_U132
g12265 nand P1_U3491 P1_R1282_U35 ; P1_R1282_U133
g12266 nand P1_R1282_U92 P1_R1282_U62 ; P1_R1282_U134
g12267 nand P1_U3488 P1_R1282_U134 ; P1_R1282_U135
g12268 nand P1_U3485 P1_R1282_U30 ; P1_R1282_U136
g12269 nand P1_R1282_U92 P1_R1282_U62 ; P1_R1282_U137
g12270 nand P1_U3473 P1_R1282_U27 ; P1_R1282_U138
g12271 nand P1_R1282_U89 P1_R1282_U64 ; P1_R1282_U139
g12272 nand P1_U4026 P1_R1282_U67 ; P1_R1282_U140
g12273 nand P1_R1282_U111 P1_R1282_U66 ; P1_R1282_U141
g12274 nand P1_U4028 P1_R1282_U46 ; P1_R1282_U142
g12275 nand P1_R1282_U110 P1_R1282_U69 ; P1_R1282_U143
g12276 nand P1_U4018 P1_R1282_U45 ; P1_R1282_U144
g12277 nand P1_R1282_U109 P1_R1282_U71 ; P1_R1282_U145
g12278 nand P1_U4020 P1_R1282_U44 ; P1_R1282_U146
g12279 nand P1_R1282_U108 P1_R1282_U73 ; P1_R1282_U147
g12280 nand P1_U4022 P1_R1282_U43 ; P1_R1282_U148
g12281 nand P1_R1282_U107 P1_R1282_U75 ; P1_R1282_U149
g12282 nand P1_U4024 P1_R1282_U42 ; P1_R1282_U150
g12283 nand P1_R1282_U106 P1_R1282_U77 ; P1_R1282_U151
g12284 nand P1_U3461 P1_R1282_U80 ; P1_R1282_U152
g12285 nand P1_U3456 P1_R1282_U79 ; P1_R1282_U153
g12286 nand P1_U3514 P1_R1282_U41 ; P1_R1282_U154
g12287 nand P1_R1282_U105 P1_R1282_U81 ; P1_R1282_U155
g12288 nand P1_U3509 P1_R1282_U40 ; P1_R1282_U156
g12289 nand P1_R1282_U104 P1_R1282_U83 ; P1_R1282_U157
g12290 nand P1_U3497 P1_R1282_U37 ; P1_R1282_U158
g12291 nand P1_R1282_U101 P1_R1282_U85 ; P1_R1282_U159
g12292 and P1_R1240_U176 P1_R1240_U175 ; P1_R1240_U4
g12293 and P1_R1240_U177 P1_R1240_U178 ; P1_R1240_U5
g12294 and P1_R1240_U194 P1_R1240_U193 ; P1_R1240_U6
g12295 and P1_R1240_U234 P1_R1240_U233 ; P1_R1240_U7
g12296 and P1_R1240_U243 P1_R1240_U242 ; P1_R1240_U8
g12297 and P1_R1240_U261 P1_R1240_U260 ; P1_R1240_U9
g12298 and P1_R1240_U269 P1_R1240_U268 ; P1_R1240_U10
g12299 and P1_R1240_U348 P1_R1240_U345 ; P1_R1240_U11
g12300 and P1_R1240_U341 P1_R1240_U338 ; P1_R1240_U12
g12301 and P1_R1240_U332 P1_R1240_U329 ; P1_R1240_U13
g12302 and P1_R1240_U323 P1_R1240_U320 ; P1_R1240_U14
g12303 and P1_R1240_U317 P1_R1240_U315 ; P1_R1240_U15
g12304 and P1_R1240_U310 P1_R1240_U307 ; P1_R1240_U16
g12305 and P1_R1240_U232 P1_R1240_U229 ; P1_R1240_U17
g12306 and P1_R1240_U224 P1_R1240_U221 ; P1_R1240_U18
g12307 and P1_R1240_U210 P1_R1240_U207 ; P1_R1240_U19
g12308 not P1_U3476 ; P1_R1240_U20
g12309 not P1_U3071 ; P1_R1240_U21
g12310 not P1_U3070 ; P1_R1240_U22
g12311 nand P1_U3071 P1_U3476 ; P1_R1240_U23
g12312 not P1_U3479 ; P1_R1240_U24
g12313 not P1_U3470 ; P1_R1240_U25
g12314 not P1_U3060 ; P1_R1240_U26
g12315 not P1_U3067 ; P1_R1240_U27
g12316 not P1_U3464 ; P1_R1240_U28
g12317 not P1_U3068 ; P1_R1240_U29
g12318 not P1_U3456 ; P1_R1240_U30
g12319 not P1_U3077 ; P1_R1240_U31
g12320 nand P1_U3077 P1_U3456 ; P1_R1240_U32
g12321 not P1_U3467 ; P1_R1240_U33
g12322 not P1_U3064 ; P1_R1240_U34
g12323 nand P1_U3060 P1_U3470 ; P1_R1240_U35
g12324 not P1_U3473 ; P1_R1240_U36
g12325 not P1_U3482 ; P1_R1240_U37
g12326 not P1_U3084 ; P1_R1240_U38
g12327 not P1_U3083 ; P1_R1240_U39
g12328 not P1_U3485 ; P1_R1240_U40
g12329 nand P1_R1240_U62 P1_R1240_U202 ; P1_R1240_U41
g12330 nand P1_R1240_U118 P1_R1240_U190 ; P1_R1240_U42
g12331 nand P1_R1240_U179 P1_R1240_U180 ; P1_R1240_U43
g12332 nand P1_U3461 P1_U3078 ; P1_R1240_U44
g12333 nand P1_R1240_U122 P1_R1240_U216 ; P1_R1240_U45
g12334 nand P1_R1240_U213 P1_R1240_U212 ; P1_R1240_U46
g12335 not P1_U4018 ; P1_R1240_U47
g12336 not P1_U3053 ; P1_R1240_U48
g12337 not P1_U3057 ; P1_R1240_U49
g12338 not P1_U4019 ; P1_R1240_U50
g12339 not P1_U4020 ; P1_R1240_U51
g12340 not P1_U3058 ; P1_R1240_U52
g12341 not P1_U4021 ; P1_R1240_U53
g12342 not P1_U3065 ; P1_R1240_U54
g12343 not P1_U4024 ; P1_R1240_U55
g12344 not P1_U3075 ; P1_R1240_U56
g12345 not P1_U3506 ; P1_R1240_U57
g12346 not P1_U3073 ; P1_R1240_U58
g12347 not P1_U3069 ; P1_R1240_U59
g12348 nand P1_U3073 P1_U3506 ; P1_R1240_U60
g12349 not P1_U3509 ; P1_R1240_U61
g12350 nand P1_U3084 P1_U3482 ; P1_R1240_U62
g12351 not P1_U3488 ; P1_R1240_U63
g12352 not P1_U3062 ; P1_R1240_U64
g12353 not P1_U3494 ; P1_R1240_U65
g12354 not P1_U3072 ; P1_R1240_U66
g12355 not P1_U3491 ; P1_R1240_U67
g12356 not P1_U3063 ; P1_R1240_U68
g12357 nand P1_U3063 P1_U3491 ; P1_R1240_U69
g12358 not P1_U3497 ; P1_R1240_U70
g12359 not P1_U3080 ; P1_R1240_U71
g12360 not P1_U3500 ; P1_R1240_U72
g12361 not P1_U3079 ; P1_R1240_U73
g12362 not P1_U3503 ; P1_R1240_U74
g12363 not P1_U3074 ; P1_R1240_U75
g12364 not P1_U3512 ; P1_R1240_U76
g12365 not P1_U3082 ; P1_R1240_U77
g12366 nand P1_U3082 P1_U3512 ; P1_R1240_U78
g12367 not P1_U3514 ; P1_R1240_U79
g12368 not P1_U3081 ; P1_R1240_U80
g12369 nand P1_U3081 P1_U3514 ; P1_R1240_U81
g12370 not P1_U4025 ; P1_R1240_U82
g12371 not P1_U4023 ; P1_R1240_U83
g12372 not P1_U3061 ; P1_R1240_U84
g12373 not P1_U4022 ; P1_R1240_U85
g12374 not P1_U3066 ; P1_R1240_U86
g12375 nand P1_U4019 P1_U3057 ; P1_R1240_U87
g12376 not P1_U3054 ; P1_R1240_U88
g12377 not P1_U4017 ; P1_R1240_U89
g12378 nand P1_R1240_U303 P1_R1240_U173 ; P1_R1240_U90
g12379 not P1_U3076 ; P1_R1240_U91
g12380 nand P1_R1240_U78 P1_R1240_U312 ; P1_R1240_U92
g12381 nand P1_R1240_U258 P1_R1240_U257 ; P1_R1240_U93
g12382 nand P1_R1240_U69 P1_R1240_U334 ; P1_R1240_U94
g12383 nand P1_R1240_U454 P1_R1240_U453 ; P1_R1240_U95
g12384 nand P1_R1240_U501 P1_R1240_U500 ; P1_R1240_U96
g12385 nand P1_R1240_U372 P1_R1240_U371 ; P1_R1240_U97
g12386 nand P1_R1240_U377 P1_R1240_U376 ; P1_R1240_U98
g12387 nand P1_R1240_U384 P1_R1240_U383 ; P1_R1240_U99
g12388 nand P1_R1240_U391 P1_R1240_U390 ; P1_R1240_U100
g12389 nand P1_R1240_U396 P1_R1240_U395 ; P1_R1240_U101
g12390 nand P1_R1240_U405 P1_R1240_U404 ; P1_R1240_U102
g12391 nand P1_R1240_U412 P1_R1240_U411 ; P1_R1240_U103
g12392 nand P1_R1240_U419 P1_R1240_U418 ; P1_R1240_U104
g12393 nand P1_R1240_U426 P1_R1240_U425 ; P1_R1240_U105
g12394 nand P1_R1240_U431 P1_R1240_U430 ; P1_R1240_U106
g12395 nand P1_R1240_U438 P1_R1240_U437 ; P1_R1240_U107
g12396 nand P1_R1240_U445 P1_R1240_U444 ; P1_R1240_U108
g12397 nand P1_R1240_U459 P1_R1240_U458 ; P1_R1240_U109
g12398 nand P1_R1240_U464 P1_R1240_U463 ; P1_R1240_U110
g12399 nand P1_R1240_U471 P1_R1240_U470 ; P1_R1240_U111
g12400 nand P1_R1240_U478 P1_R1240_U477 ; P1_R1240_U112
g12401 nand P1_R1240_U485 P1_R1240_U484 ; P1_R1240_U113
g12402 nand P1_R1240_U492 P1_R1240_U491 ; P1_R1240_U114
g12403 nand P1_R1240_U497 P1_R1240_U496 ; P1_R1240_U115
g12404 and P1_U3464 P1_U3068 ; P1_R1240_U116
g12405 and P1_R1240_U186 P1_R1240_U184 ; P1_R1240_U117
g12406 and P1_R1240_U191 P1_R1240_U189 ; P1_R1240_U118
g12407 and P1_R1240_U198 P1_R1240_U197 ; P1_R1240_U119
g12408 and P1_R1240_U379 P1_R1240_U378 P1_R1240_U23 ; P1_R1240_U120
g12409 and P1_R1240_U209 P1_R1240_U6 ; P1_R1240_U121
g12410 and P1_R1240_U217 P1_R1240_U215 ; P1_R1240_U122
g12411 and P1_R1240_U386 P1_R1240_U385 P1_R1240_U35 ; P1_R1240_U123
g12412 and P1_R1240_U223 P1_R1240_U4 ; P1_R1240_U124
g12413 and P1_R1240_U231 P1_R1240_U178 ; P1_R1240_U125
g12414 and P1_R1240_U201 P1_R1240_U7 ; P1_R1240_U126
g12415 and P1_R1240_U236 P1_R1240_U168 ; P1_R1240_U127
g12416 and P1_R1240_U245 P1_R1240_U169 ; P1_R1240_U128
g12417 and P1_R1240_U265 P1_R1240_U264 ; P1_R1240_U129
g12418 and P1_R1240_U10 P1_R1240_U279 ; P1_R1240_U130
g12419 and P1_R1240_U282 P1_R1240_U277 ; P1_R1240_U131
g12420 and P1_R1240_U298 P1_R1240_U295 ; P1_R1240_U132
g12421 and P1_R1240_U365 P1_R1240_U299 ; P1_R1240_U133
g12422 and P1_R1240_U156 P1_R1240_U275 ; P1_R1240_U134
g12423 and P1_R1240_U466 P1_R1240_U465 P1_R1240_U60 ; P1_R1240_U135
g12424 and P1_R1240_U487 P1_R1240_U486 P1_R1240_U169 ; P1_R1240_U136
g12425 and P1_R1240_U340 P1_R1240_U8 ; P1_R1240_U137
g12426 and P1_R1240_U499 P1_R1240_U498 P1_R1240_U168 ; P1_R1240_U138
g12427 and P1_R1240_U347 P1_R1240_U7 ; P1_R1240_U139
g12428 nand P1_R1240_U119 P1_R1240_U199 ; P1_R1240_U140
g12429 nand P1_R1240_U214 P1_R1240_U226 ; P1_R1240_U141
g12430 not P1_U3055 ; P1_R1240_U142
g12431 not P1_U4028 ; P1_R1240_U143
g12432 and P1_R1240_U400 P1_R1240_U399 ; P1_R1240_U144
g12433 nand P1_R1240_U301 P1_R1240_U166 P1_R1240_U361 ; P1_R1240_U145
g12434 and P1_R1240_U407 P1_R1240_U406 ; P1_R1240_U146
g12435 nand P1_R1240_U367 P1_R1240_U366 P1_R1240_U133 ; P1_R1240_U147
g12436 and P1_R1240_U414 P1_R1240_U413 ; P1_R1240_U148
g12437 nand P1_R1240_U362 P1_R1240_U296 P1_R1240_U87 ; P1_R1240_U149
g12438 and P1_R1240_U421 P1_R1240_U420 ; P1_R1240_U150
g12439 nand P1_R1240_U290 P1_R1240_U289 ; P1_R1240_U151
g12440 and P1_R1240_U433 P1_R1240_U432 ; P1_R1240_U152
g12441 nand P1_R1240_U286 P1_R1240_U285 ; P1_R1240_U153
g12442 and P1_R1240_U440 P1_R1240_U439 ; P1_R1240_U154
g12443 nand P1_R1240_U131 P1_R1240_U281 ; P1_R1240_U155
g12444 and P1_R1240_U447 P1_R1240_U446 ; P1_R1240_U156
g12445 and P1_R1240_U452 P1_R1240_U451 ; P1_R1240_U157
g12446 nand P1_R1240_U44 P1_R1240_U324 ; P1_R1240_U158
g12447 nand P1_R1240_U129 P1_R1240_U266 ; P1_R1240_U159
g12448 and P1_R1240_U473 P1_R1240_U472 ; P1_R1240_U160
g12449 nand P1_R1240_U254 P1_R1240_U253 ; P1_R1240_U161
g12450 and P1_R1240_U480 P1_R1240_U479 ; P1_R1240_U162
g12451 nand P1_R1240_U250 P1_R1240_U249 ; P1_R1240_U163
g12452 nand P1_R1240_U240 P1_R1240_U239 ; P1_R1240_U164
g12453 nand P1_R1240_U364 P1_R1240_U363 ; P1_R1240_U165
g12454 nand P1_U3054 P1_R1240_U147 ; P1_R1240_U166
g12455 not P1_R1240_U35 ; P1_R1240_U167
g12456 nand P1_U3485 P1_U3083 ; P1_R1240_U168
g12457 nand P1_U3072 P1_U3494 ; P1_R1240_U169
g12458 nand P1_U3058 P1_U4020 ; P1_R1240_U170
g12459 not P1_R1240_U69 ; P1_R1240_U171
g12460 not P1_R1240_U78 ; P1_R1240_U172
g12461 nand P1_U3065 P1_U4021 ; P1_R1240_U173
g12462 not P1_R1240_U62 ; P1_R1240_U174
g12463 or P1_U3067 P1_U3473 ; P1_R1240_U175
g12464 or P1_U3060 P1_U3470 ; P1_R1240_U176
g12465 or P1_U3467 P1_U3064 ; P1_R1240_U177
g12466 or P1_U3464 P1_U3068 ; P1_R1240_U178
g12467 not P1_R1240_U32 ; P1_R1240_U179
g12468 or P1_U3461 P1_U3078 ; P1_R1240_U180
g12469 not P1_R1240_U43 ; P1_R1240_U181
g12470 not P1_R1240_U44 ; P1_R1240_U182
g12471 nand P1_R1240_U43 P1_R1240_U44 ; P1_R1240_U183
g12472 nand P1_R1240_U116 P1_R1240_U177 ; P1_R1240_U184
g12473 nand P1_R1240_U5 P1_R1240_U183 ; P1_R1240_U185
g12474 nand P1_U3064 P1_U3467 ; P1_R1240_U186
g12475 nand P1_R1240_U117 P1_R1240_U185 ; P1_R1240_U187
g12476 nand P1_R1240_U36 P1_R1240_U35 ; P1_R1240_U188
g12477 nand P1_U3067 P1_R1240_U188 ; P1_R1240_U189
g12478 nand P1_R1240_U4 P1_R1240_U187 ; P1_R1240_U190
g12479 nand P1_U3473 P1_R1240_U167 ; P1_R1240_U191
g12480 not P1_R1240_U42 ; P1_R1240_U192
g12481 or P1_U3070 P1_U3479 ; P1_R1240_U193
g12482 or P1_U3071 P1_U3476 ; P1_R1240_U194
g12483 not P1_R1240_U23 ; P1_R1240_U195
g12484 nand P1_R1240_U24 P1_R1240_U23 ; P1_R1240_U196
g12485 nand P1_U3070 P1_R1240_U196 ; P1_R1240_U197
g12486 nand P1_U3479 P1_R1240_U195 ; P1_R1240_U198
g12487 nand P1_R1240_U6 P1_R1240_U42 ; P1_R1240_U199
g12488 not P1_R1240_U140 ; P1_R1240_U200
g12489 or P1_U3482 P1_U3084 ; P1_R1240_U201
g12490 nand P1_R1240_U201 P1_R1240_U140 ; P1_R1240_U202
g12491 not P1_R1240_U41 ; P1_R1240_U203
g12492 or P1_U3083 P1_U3485 ; P1_R1240_U204
g12493 or P1_U3476 P1_U3071 ; P1_R1240_U205
g12494 nand P1_R1240_U205 P1_R1240_U42 ; P1_R1240_U206
g12495 nand P1_R1240_U120 P1_R1240_U206 ; P1_R1240_U207
g12496 nand P1_R1240_U192 P1_R1240_U23 ; P1_R1240_U208
g12497 nand P1_U3479 P1_U3070 ; P1_R1240_U209
g12498 nand P1_R1240_U121 P1_R1240_U208 ; P1_R1240_U210
g12499 or P1_U3071 P1_U3476 ; P1_R1240_U211
g12500 nand P1_R1240_U182 P1_R1240_U178 ; P1_R1240_U212
g12501 nand P1_U3068 P1_U3464 ; P1_R1240_U213
g12502 not P1_R1240_U46 ; P1_R1240_U214
g12503 nand P1_R1240_U181 P1_R1240_U5 ; P1_R1240_U215
g12504 nand P1_R1240_U46 P1_R1240_U177 ; P1_R1240_U216
g12505 nand P1_U3064 P1_U3467 ; P1_R1240_U217
g12506 not P1_R1240_U45 ; P1_R1240_U218
g12507 or P1_U3470 P1_U3060 ; P1_R1240_U219
g12508 nand P1_R1240_U219 P1_R1240_U45 ; P1_R1240_U220
g12509 nand P1_R1240_U123 P1_R1240_U220 ; P1_R1240_U221
g12510 nand P1_R1240_U218 P1_R1240_U35 ; P1_R1240_U222
g12511 nand P1_U3473 P1_U3067 ; P1_R1240_U223
g12512 nand P1_R1240_U124 P1_R1240_U222 ; P1_R1240_U224
g12513 or P1_U3060 P1_U3470 ; P1_R1240_U225
g12514 nand P1_R1240_U181 P1_R1240_U178 ; P1_R1240_U226
g12515 not P1_R1240_U141 ; P1_R1240_U227
g12516 nand P1_U3064 P1_U3467 ; P1_R1240_U228
g12517 nand P1_R1240_U398 P1_R1240_U397 P1_R1240_U44 P1_R1240_U43 ; P1_R1240_U229
g12518 nand P1_R1240_U44 P1_R1240_U43 ; P1_R1240_U230
g12519 nand P1_U3068 P1_U3464 ; P1_R1240_U231
g12520 nand P1_R1240_U125 P1_R1240_U230 ; P1_R1240_U232
g12521 or P1_U3083 P1_U3485 ; P1_R1240_U233
g12522 or P1_U3062 P1_U3488 ; P1_R1240_U234
g12523 nand P1_R1240_U174 P1_R1240_U7 ; P1_R1240_U235
g12524 nand P1_U3062 P1_U3488 ; P1_R1240_U236
g12525 nand P1_R1240_U127 P1_R1240_U235 ; P1_R1240_U237
g12526 or P1_U3488 P1_U3062 ; P1_R1240_U238
g12527 nand P1_R1240_U126 P1_R1240_U140 ; P1_R1240_U239
g12528 nand P1_R1240_U238 P1_R1240_U237 ; P1_R1240_U240
g12529 not P1_R1240_U164 ; P1_R1240_U241
g12530 or P1_U3080 P1_U3497 ; P1_R1240_U242
g12531 or P1_U3072 P1_U3494 ; P1_R1240_U243
g12532 nand P1_R1240_U171 P1_R1240_U8 ; P1_R1240_U244
g12533 nand P1_U3080 P1_U3497 ; P1_R1240_U245
g12534 nand P1_R1240_U128 P1_R1240_U244 ; P1_R1240_U246
g12535 or P1_U3491 P1_U3063 ; P1_R1240_U247
g12536 or P1_U3497 P1_U3080 ; P1_R1240_U248
g12537 nand P1_R1240_U247 P1_R1240_U164 P1_R1240_U8 ; P1_R1240_U249
g12538 nand P1_R1240_U248 P1_R1240_U246 ; P1_R1240_U250
g12539 not P1_R1240_U163 ; P1_R1240_U251
g12540 or P1_U3500 P1_U3079 ; P1_R1240_U252
g12541 nand P1_R1240_U252 P1_R1240_U163 ; P1_R1240_U253
g12542 nand P1_U3079 P1_U3500 ; P1_R1240_U254
g12543 not P1_R1240_U161 ; P1_R1240_U255
g12544 or P1_U3503 P1_U3074 ; P1_R1240_U256
g12545 nand P1_R1240_U256 P1_R1240_U161 ; P1_R1240_U257
g12546 nand P1_U3074 P1_U3503 ; P1_R1240_U258
g12547 not P1_R1240_U93 ; P1_R1240_U259
g12548 or P1_U3069 P1_U3509 ; P1_R1240_U260
g12549 or P1_U3073 P1_U3506 ; P1_R1240_U261
g12550 not P1_R1240_U60 ; P1_R1240_U262
g12551 nand P1_R1240_U61 P1_R1240_U60 ; P1_R1240_U263
g12552 nand P1_U3069 P1_R1240_U263 ; P1_R1240_U264
g12553 nand P1_U3509 P1_R1240_U262 ; P1_R1240_U265
g12554 nand P1_R1240_U9 P1_R1240_U93 ; P1_R1240_U266
g12555 not P1_R1240_U159 ; P1_R1240_U267
g12556 or P1_U3076 P1_U4025 ; P1_R1240_U268
g12557 or P1_U3081 P1_U3514 ; P1_R1240_U269
g12558 or P1_U3075 P1_U4024 ; P1_R1240_U270
g12559 not P1_R1240_U81 ; P1_R1240_U271
g12560 nand P1_U4025 P1_R1240_U271 ; P1_R1240_U272
g12561 nand P1_R1240_U272 P1_R1240_U91 ; P1_R1240_U273
g12562 nand P1_R1240_U81 P1_R1240_U82 ; P1_R1240_U274
g12563 nand P1_R1240_U274 P1_R1240_U273 ; P1_R1240_U275
g12564 nand P1_R1240_U172 P1_R1240_U10 ; P1_R1240_U276
g12565 nand P1_U3075 P1_U4024 ; P1_R1240_U277
g12566 nand P1_R1240_U275 P1_R1240_U276 ; P1_R1240_U278
g12567 or P1_U3512 P1_U3082 ; P1_R1240_U279
g12568 or P1_U4024 P1_U3075 ; P1_R1240_U280
g12569 nand P1_R1240_U270 P1_R1240_U159 P1_R1240_U130 ; P1_R1240_U281
g12570 nand P1_R1240_U280 P1_R1240_U278 ; P1_R1240_U282
g12571 not P1_R1240_U155 ; P1_R1240_U283
g12572 or P1_U4023 P1_U3061 ; P1_R1240_U284
g12573 nand P1_R1240_U284 P1_R1240_U155 ; P1_R1240_U285
g12574 nand P1_U3061 P1_U4023 ; P1_R1240_U286
g12575 not P1_R1240_U153 ; P1_R1240_U287
g12576 or P1_U4022 P1_U3066 ; P1_R1240_U288
g12577 nand P1_R1240_U288 P1_R1240_U153 ; P1_R1240_U289
g12578 nand P1_U3066 P1_U4022 ; P1_R1240_U290
g12579 not P1_R1240_U151 ; P1_R1240_U291
g12580 or P1_U3058 P1_U4020 ; P1_R1240_U292
g12581 nand P1_R1240_U173 P1_R1240_U170 ; P1_R1240_U293
g12582 not P1_R1240_U87 ; P1_R1240_U294
g12583 or P1_U4021 P1_U3065 ; P1_R1240_U295
g12584 nand P1_R1240_U151 P1_R1240_U295 P1_R1240_U165 ; P1_R1240_U296
g12585 not P1_R1240_U149 ; P1_R1240_U297
g12586 or P1_U4018 P1_U3053 ; P1_R1240_U298
g12587 nand P1_U3053 P1_U4018 ; P1_R1240_U299
g12588 not P1_R1240_U147 ; P1_R1240_U300
g12589 nand P1_U4017 P1_R1240_U147 ; P1_R1240_U301
g12590 not P1_R1240_U145 ; P1_R1240_U302
g12591 nand P1_R1240_U295 P1_R1240_U151 ; P1_R1240_U303
g12592 not P1_R1240_U90 ; P1_R1240_U304
g12593 or P1_U4020 P1_U3058 ; P1_R1240_U305
g12594 nand P1_R1240_U305 P1_R1240_U90 ; P1_R1240_U306
g12595 nand P1_R1240_U306 P1_R1240_U170 P1_R1240_U150 ; P1_R1240_U307
g12596 nand P1_R1240_U304 P1_R1240_U170 ; P1_R1240_U308
g12597 nand P1_U4019 P1_U3057 ; P1_R1240_U309
g12598 nand P1_R1240_U308 P1_R1240_U309 P1_R1240_U165 ; P1_R1240_U310
g12599 or P1_U3058 P1_U4020 ; P1_R1240_U311
g12600 nand P1_R1240_U279 P1_R1240_U159 ; P1_R1240_U312
g12601 not P1_R1240_U92 ; P1_R1240_U313
g12602 nand P1_R1240_U10 P1_R1240_U92 ; P1_R1240_U314
g12603 nand P1_R1240_U134 P1_R1240_U314 ; P1_R1240_U315
g12604 nand P1_R1240_U314 P1_R1240_U275 ; P1_R1240_U316
g12605 nand P1_R1240_U450 P1_R1240_U316 ; P1_R1240_U317
g12606 or P1_U3514 P1_U3081 ; P1_R1240_U318
g12607 nand P1_R1240_U318 P1_R1240_U92 ; P1_R1240_U319
g12608 nand P1_R1240_U319 P1_R1240_U81 P1_R1240_U157 ; P1_R1240_U320
g12609 nand P1_R1240_U313 P1_R1240_U81 ; P1_R1240_U321
g12610 nand P1_U3076 P1_U4025 ; P1_R1240_U322
g12611 nand P1_R1240_U322 P1_R1240_U321 P1_R1240_U10 ; P1_R1240_U323
g12612 or P1_U3461 P1_U3078 ; P1_R1240_U324
g12613 not P1_R1240_U158 ; P1_R1240_U325
g12614 or P1_U3081 P1_U3514 ; P1_R1240_U326
g12615 or P1_U3506 P1_U3073 ; P1_R1240_U327
g12616 nand P1_R1240_U327 P1_R1240_U93 ; P1_R1240_U328
g12617 nand P1_R1240_U135 P1_R1240_U328 ; P1_R1240_U329
g12618 nand P1_R1240_U259 P1_R1240_U60 ; P1_R1240_U330
g12619 nand P1_U3509 P1_U3069 ; P1_R1240_U331
g12620 nand P1_R1240_U331 P1_R1240_U330 P1_R1240_U9 ; P1_R1240_U332
g12621 or P1_U3073 P1_U3506 ; P1_R1240_U333
g12622 nand P1_R1240_U247 P1_R1240_U164 ; P1_R1240_U334
g12623 not P1_R1240_U94 ; P1_R1240_U335
g12624 or P1_U3494 P1_U3072 ; P1_R1240_U336
g12625 nand P1_R1240_U336 P1_R1240_U94 ; P1_R1240_U337
g12626 nand P1_R1240_U136 P1_R1240_U337 ; P1_R1240_U338
g12627 nand P1_R1240_U335 P1_R1240_U169 ; P1_R1240_U339
g12628 nand P1_U3080 P1_U3497 ; P1_R1240_U340
g12629 nand P1_R1240_U137 P1_R1240_U339 ; P1_R1240_U341
g12630 or P1_U3072 P1_U3494 ; P1_R1240_U342
g12631 or P1_U3485 P1_U3083 ; P1_R1240_U343
g12632 nand P1_R1240_U343 P1_R1240_U41 ; P1_R1240_U344
g12633 nand P1_R1240_U138 P1_R1240_U344 ; P1_R1240_U345
g12634 nand P1_R1240_U203 P1_R1240_U168 ; P1_R1240_U346
g12635 nand P1_U3062 P1_U3488 ; P1_R1240_U347
g12636 nand P1_R1240_U139 P1_R1240_U346 ; P1_R1240_U348
g12637 nand P1_R1240_U204 P1_R1240_U168 ; P1_R1240_U349
g12638 nand P1_R1240_U201 P1_R1240_U62 ; P1_R1240_U350
g12639 nand P1_R1240_U211 P1_R1240_U23 ; P1_R1240_U351
g12640 nand P1_R1240_U225 P1_R1240_U35 ; P1_R1240_U352
g12641 nand P1_R1240_U228 P1_R1240_U177 ; P1_R1240_U353
g12642 nand P1_R1240_U311 P1_R1240_U170 ; P1_R1240_U354
g12643 nand P1_R1240_U295 P1_R1240_U173 ; P1_R1240_U355
g12644 nand P1_R1240_U326 P1_R1240_U81 ; P1_R1240_U356
g12645 nand P1_R1240_U279 P1_R1240_U78 ; P1_R1240_U357
g12646 nand P1_R1240_U333 P1_R1240_U60 ; P1_R1240_U358
g12647 nand P1_R1240_U342 P1_R1240_U169 ; P1_R1240_U359
g12648 nand P1_R1240_U247 P1_R1240_U69 ; P1_R1240_U360
g12649 nand P1_U4017 P1_U3054 ; P1_R1240_U361
g12650 nand P1_R1240_U293 P1_R1240_U165 ; P1_R1240_U362
g12651 nand P1_U3057 P1_R1240_U292 ; P1_R1240_U363
g12652 nand P1_U4019 P1_R1240_U292 ; P1_R1240_U364
g12653 nand P1_R1240_U293 P1_R1240_U165 P1_R1240_U298 ; P1_R1240_U365
g12654 nand P1_R1240_U151 P1_R1240_U165 P1_R1240_U132 ; P1_R1240_U366
g12655 nand P1_R1240_U294 P1_R1240_U298 ; P1_R1240_U367
g12656 nand P1_U3083 P1_R1240_U40 ; P1_R1240_U368
g12657 nand P1_U3485 P1_R1240_U39 ; P1_R1240_U369
g12658 nand P1_R1240_U369 P1_R1240_U368 ; P1_R1240_U370
g12659 nand P1_R1240_U349 P1_R1240_U41 ; P1_R1240_U371
g12660 nand P1_R1240_U370 P1_R1240_U203 ; P1_R1240_U372
g12661 nand P1_U3084 P1_R1240_U37 ; P1_R1240_U373
g12662 nand P1_U3482 P1_R1240_U38 ; P1_R1240_U374
g12663 nand P1_R1240_U374 P1_R1240_U373 ; P1_R1240_U375
g12664 nand P1_R1240_U350 P1_R1240_U140 ; P1_R1240_U376
g12665 nand P1_R1240_U200 P1_R1240_U375 ; P1_R1240_U377
g12666 nand P1_U3070 P1_R1240_U24 ; P1_R1240_U378
g12667 nand P1_U3479 P1_R1240_U22 ; P1_R1240_U379
g12668 nand P1_U3071 P1_R1240_U20 ; P1_R1240_U380
g12669 nand P1_U3476 P1_R1240_U21 ; P1_R1240_U381
g12670 nand P1_R1240_U381 P1_R1240_U380 ; P1_R1240_U382
g12671 nand P1_R1240_U351 P1_R1240_U42 ; P1_R1240_U383
g12672 nand P1_R1240_U382 P1_R1240_U192 ; P1_R1240_U384
g12673 nand P1_U3067 P1_R1240_U36 ; P1_R1240_U385
g12674 nand P1_U3473 P1_R1240_U27 ; P1_R1240_U386
g12675 nand P1_U3060 P1_R1240_U25 ; P1_R1240_U387
g12676 nand P1_U3470 P1_R1240_U26 ; P1_R1240_U388
g12677 nand P1_R1240_U388 P1_R1240_U387 ; P1_R1240_U389
g12678 nand P1_R1240_U352 P1_R1240_U45 ; P1_R1240_U390
g12679 nand P1_R1240_U389 P1_R1240_U218 ; P1_R1240_U391
g12680 nand P1_U3064 P1_R1240_U33 ; P1_R1240_U392
g12681 nand P1_U3467 P1_R1240_U34 ; P1_R1240_U393
g12682 nand P1_R1240_U393 P1_R1240_U392 ; P1_R1240_U394
g12683 nand P1_R1240_U353 P1_R1240_U141 ; P1_R1240_U395
g12684 nand P1_R1240_U227 P1_R1240_U394 ; P1_R1240_U396
g12685 nand P1_U3068 P1_R1240_U28 ; P1_R1240_U397
g12686 nand P1_U3464 P1_R1240_U29 ; P1_R1240_U398
g12687 nand P1_U3055 P1_R1240_U143 ; P1_R1240_U399
g12688 nand P1_U4028 P1_R1240_U142 ; P1_R1240_U400
g12689 nand P1_U3055 P1_R1240_U143 ; P1_R1240_U401
g12690 nand P1_U4028 P1_R1240_U142 ; P1_R1240_U402
g12691 nand P1_R1240_U402 P1_R1240_U401 ; P1_R1240_U403
g12692 nand P1_R1240_U144 P1_R1240_U145 ; P1_R1240_U404
g12693 nand P1_R1240_U302 P1_R1240_U403 ; P1_R1240_U405
g12694 nand P1_U3054 P1_R1240_U89 ; P1_R1240_U406
g12695 nand P1_U4017 P1_R1240_U88 ; P1_R1240_U407
g12696 nand P1_U3054 P1_R1240_U89 ; P1_R1240_U408
g12697 nand P1_U4017 P1_R1240_U88 ; P1_R1240_U409
g12698 nand P1_R1240_U409 P1_R1240_U408 ; P1_R1240_U410
g12699 nand P1_R1240_U146 P1_R1240_U147 ; P1_R1240_U411
g12700 nand P1_R1240_U300 P1_R1240_U410 ; P1_R1240_U412
g12701 nand P1_U3053 P1_R1240_U47 ; P1_R1240_U413
g12702 nand P1_U4018 P1_R1240_U48 ; P1_R1240_U414
g12703 nand P1_U3053 P1_R1240_U47 ; P1_R1240_U415
g12704 nand P1_U4018 P1_R1240_U48 ; P1_R1240_U416
g12705 nand P1_R1240_U416 P1_R1240_U415 ; P1_R1240_U417
g12706 nand P1_R1240_U148 P1_R1240_U149 ; P1_R1240_U418
g12707 nand P1_R1240_U297 P1_R1240_U417 ; P1_R1240_U419
g12708 nand P1_U3057 P1_R1240_U50 ; P1_R1240_U420
g12709 nand P1_U4019 P1_R1240_U49 ; P1_R1240_U421
g12710 nand P1_U3058 P1_R1240_U51 ; P1_R1240_U422
g12711 nand P1_U4020 P1_R1240_U52 ; P1_R1240_U423
g12712 nand P1_R1240_U423 P1_R1240_U422 ; P1_R1240_U424
g12713 nand P1_R1240_U354 P1_R1240_U90 ; P1_R1240_U425
g12714 nand P1_R1240_U424 P1_R1240_U304 ; P1_R1240_U426
g12715 nand P1_U3065 P1_R1240_U53 ; P1_R1240_U427
g12716 nand P1_U4021 P1_R1240_U54 ; P1_R1240_U428
g12717 nand P1_R1240_U428 P1_R1240_U427 ; P1_R1240_U429
g12718 nand P1_R1240_U355 P1_R1240_U151 ; P1_R1240_U430
g12719 nand P1_R1240_U291 P1_R1240_U429 ; P1_R1240_U431
g12720 nand P1_U3066 P1_R1240_U85 ; P1_R1240_U432
g12721 nand P1_U4022 P1_R1240_U86 ; P1_R1240_U433
g12722 nand P1_U3066 P1_R1240_U85 ; P1_R1240_U434
g12723 nand P1_U4022 P1_R1240_U86 ; P1_R1240_U435
g12724 nand P1_R1240_U435 P1_R1240_U434 ; P1_R1240_U436
g12725 nand P1_R1240_U152 P1_R1240_U153 ; P1_R1240_U437
g12726 nand P1_R1240_U287 P1_R1240_U436 ; P1_R1240_U438
g12727 nand P1_U3061 P1_R1240_U83 ; P1_R1240_U439
g12728 nand P1_U4023 P1_R1240_U84 ; P1_R1240_U440
g12729 nand P1_U3061 P1_R1240_U83 ; P1_R1240_U441
g12730 nand P1_U4023 P1_R1240_U84 ; P1_R1240_U442
g12731 nand P1_R1240_U442 P1_R1240_U441 ; P1_R1240_U443
g12732 nand P1_R1240_U154 P1_R1240_U155 ; P1_R1240_U444
g12733 nand P1_R1240_U283 P1_R1240_U443 ; P1_R1240_U445
g12734 nand P1_U3075 P1_R1240_U55 ; P1_R1240_U446
g12735 nand P1_U4024 P1_R1240_U56 ; P1_R1240_U447
g12736 nand P1_U3075 P1_R1240_U55 ; P1_R1240_U448
g12737 nand P1_U4024 P1_R1240_U56 ; P1_R1240_U449
g12738 nand P1_R1240_U449 P1_R1240_U448 ; P1_R1240_U450
g12739 nand P1_U3076 P1_R1240_U82 ; P1_R1240_U451
g12740 nand P1_U4025 P1_R1240_U91 ; P1_R1240_U452
g12741 nand P1_R1240_U179 P1_R1240_U158 ; P1_R1240_U453
g12742 nand P1_R1240_U325 P1_R1240_U32 ; P1_R1240_U454
g12743 nand P1_U3081 P1_R1240_U79 ; P1_R1240_U455
g12744 nand P1_U3514 P1_R1240_U80 ; P1_R1240_U456
g12745 nand P1_R1240_U456 P1_R1240_U455 ; P1_R1240_U457
g12746 nand P1_R1240_U356 P1_R1240_U92 ; P1_R1240_U458
g12747 nand P1_R1240_U457 P1_R1240_U313 ; P1_R1240_U459
g12748 nand P1_U3082 P1_R1240_U76 ; P1_R1240_U460
g12749 nand P1_U3512 P1_R1240_U77 ; P1_R1240_U461
g12750 nand P1_R1240_U461 P1_R1240_U460 ; P1_R1240_U462
g12751 nand P1_R1240_U357 P1_R1240_U159 ; P1_R1240_U463
g12752 nand P1_R1240_U267 P1_R1240_U462 ; P1_R1240_U464
g12753 nand P1_U3069 P1_R1240_U61 ; P1_R1240_U465
g12754 nand P1_U3509 P1_R1240_U59 ; P1_R1240_U466
g12755 nand P1_U3073 P1_R1240_U57 ; P1_R1240_U467
g12756 nand P1_U3506 P1_R1240_U58 ; P1_R1240_U468
g12757 nand P1_R1240_U468 P1_R1240_U467 ; P1_R1240_U469
g12758 nand P1_R1240_U358 P1_R1240_U93 ; P1_R1240_U470
g12759 nand P1_R1240_U469 P1_R1240_U259 ; P1_R1240_U471
g12760 nand P1_U3074 P1_R1240_U74 ; P1_R1240_U472
g12761 nand P1_U3503 P1_R1240_U75 ; P1_R1240_U473
g12762 nand P1_U3074 P1_R1240_U74 ; P1_R1240_U474
g12763 nand P1_U3503 P1_R1240_U75 ; P1_R1240_U475
g12764 nand P1_R1240_U475 P1_R1240_U474 ; P1_R1240_U476
g12765 nand P1_R1240_U160 P1_R1240_U161 ; P1_R1240_U477
g12766 nand P1_R1240_U255 P1_R1240_U476 ; P1_R1240_U478
g12767 nand P1_U3079 P1_R1240_U72 ; P1_R1240_U479
g12768 nand P1_U3500 P1_R1240_U73 ; P1_R1240_U480
g12769 nand P1_U3079 P1_R1240_U72 ; P1_R1240_U481
g12770 nand P1_U3500 P1_R1240_U73 ; P1_R1240_U482
g12771 nand P1_R1240_U482 P1_R1240_U481 ; P1_R1240_U483
g12772 nand P1_R1240_U162 P1_R1240_U163 ; P1_R1240_U484
g12773 nand P1_R1240_U251 P1_R1240_U483 ; P1_R1240_U485
g12774 nand P1_U3080 P1_R1240_U70 ; P1_R1240_U486
g12775 nand P1_U3497 P1_R1240_U71 ; P1_R1240_U487
g12776 nand P1_U3072 P1_R1240_U65 ; P1_R1240_U488
g12777 nand P1_U3494 P1_R1240_U66 ; P1_R1240_U489
g12778 nand P1_R1240_U489 P1_R1240_U488 ; P1_R1240_U490
g12779 nand P1_R1240_U359 P1_R1240_U94 ; P1_R1240_U491
g12780 nand P1_R1240_U490 P1_R1240_U335 ; P1_R1240_U492
g12781 nand P1_U3063 P1_R1240_U67 ; P1_R1240_U493
g12782 nand P1_U3491 P1_R1240_U68 ; P1_R1240_U494
g12783 nand P1_R1240_U494 P1_R1240_U493 ; P1_R1240_U495
g12784 nand P1_R1240_U360 P1_R1240_U164 ; P1_R1240_U496
g12785 nand P1_R1240_U241 P1_R1240_U495 ; P1_R1240_U497
g12786 nand P1_U3062 P1_R1240_U63 ; P1_R1240_U498
g12787 nand P1_U3488 P1_R1240_U64 ; P1_R1240_U499
g12788 nand P1_U3077 P1_R1240_U30 ; P1_R1240_U500
g12789 nand P1_U3456 P1_R1240_U31 ; P1_R1240_U501
g12790 and P1_R1162_U95 P1_R1162_U94 ; P1_R1162_U4
g12791 and P1_R1162_U96 P1_R1162_U97 ; P1_R1162_U5
g12792 and P1_R1162_U113 P1_R1162_U112 ; P1_R1162_U6
g12793 and P1_R1162_U155 P1_R1162_U154 ; P1_R1162_U7
g12794 and P1_R1162_U164 P1_R1162_U163 ; P1_R1162_U8
g12795 and P1_R1162_U182 P1_R1162_U181 ; P1_R1162_U9
g12796 and P1_R1162_U218 P1_R1162_U215 ; P1_R1162_U10
g12797 and P1_R1162_U211 P1_R1162_U208 ; P1_R1162_U11
g12798 and P1_R1162_U202 P1_R1162_U199 ; P1_R1162_U12
g12799 and P1_R1162_U196 P1_R1162_U192 ; P1_R1162_U13
g12800 and P1_R1162_U151 P1_R1162_U148 ; P1_R1162_U14
g12801 and P1_R1162_U143 P1_R1162_U140 ; P1_R1162_U15
g12802 and P1_R1162_U129 P1_R1162_U126 ; P1_R1162_U16
g12803 not P1_REG1_REG_6__SCAN_IN ; P1_R1162_U17
g12804 not P1_U3475 ; P1_R1162_U18
g12805 not P1_U3478 ; P1_R1162_U19
g12806 nand P1_U3475 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U20
g12807 not P1_REG1_REG_7__SCAN_IN ; P1_R1162_U21
g12808 not P1_REG1_REG_4__SCAN_IN ; P1_R1162_U22
g12809 not P1_U3469 ; P1_R1162_U23
g12810 not P1_U3472 ; P1_R1162_U24
g12811 not P1_REG1_REG_2__SCAN_IN ; P1_R1162_U25
g12812 not P1_U3463 ; P1_R1162_U26
g12813 not P1_REG1_REG_0__SCAN_IN ; P1_R1162_U27
g12814 not P1_U3454 ; P1_R1162_U28
g12815 nand P1_U3454 P1_REG1_REG_0__SCAN_IN ; P1_R1162_U29
g12816 not P1_REG1_REG_3__SCAN_IN ; P1_R1162_U30
g12817 not P1_U3466 ; P1_R1162_U31
g12818 nand P1_U3469 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U32
g12819 not P1_REG1_REG_5__SCAN_IN ; P1_R1162_U33
g12820 not P1_REG1_REG_8__SCAN_IN ; P1_R1162_U34
g12821 not P1_U3481 ; P1_R1162_U35
g12822 not P1_U3484 ; P1_R1162_U36
g12823 not P1_REG1_REG_9__SCAN_IN ; P1_R1162_U37
g12824 nand P1_R1162_U49 P1_R1162_U121 ; P1_R1162_U38
g12825 nand P1_R1162_U110 P1_R1162_U108 P1_R1162_U109 ; P1_R1162_U39
g12826 nand P1_R1162_U98 P1_R1162_U99 ; P1_R1162_U40
g12827 nand P1_U3460 P1_REG1_REG_1__SCAN_IN ; P1_R1162_U41
g12828 nand P1_R1162_U136 P1_R1162_U134 P1_R1162_U135 ; P1_R1162_U42
g12829 nand P1_R1162_U132 P1_R1162_U131 ; P1_R1162_U43
g12830 not P1_REG1_REG_16__SCAN_IN ; P1_R1162_U44
g12831 not P1_U3505 ; P1_R1162_U45
g12832 not P1_U3508 ; P1_R1162_U46
g12833 nand P1_U3505 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U47
g12834 not P1_REG1_REG_17__SCAN_IN ; P1_R1162_U48
g12835 nand P1_U3481 P1_REG1_REG_8__SCAN_IN ; P1_R1162_U49
g12836 not P1_REG1_REG_10__SCAN_IN ; P1_R1162_U50
g12837 not P1_U3487 ; P1_R1162_U51
g12838 not P1_REG1_REG_12__SCAN_IN ; P1_R1162_U52
g12839 not P1_U3493 ; P1_R1162_U53
g12840 not P1_REG1_REG_11__SCAN_IN ; P1_R1162_U54
g12841 not P1_U3490 ; P1_R1162_U55
g12842 nand P1_U3490 P1_REG1_REG_11__SCAN_IN ; P1_R1162_U56
g12843 not P1_REG1_REG_13__SCAN_IN ; P1_R1162_U57
g12844 not P1_U3496 ; P1_R1162_U58
g12845 not P1_REG1_REG_14__SCAN_IN ; P1_R1162_U59
g12846 not P1_U3499 ; P1_R1162_U60
g12847 not P1_REG1_REG_15__SCAN_IN ; P1_R1162_U61
g12848 not P1_U3502 ; P1_R1162_U62
g12849 not P1_REG1_REG_18__SCAN_IN ; P1_R1162_U63
g12850 not P1_U3511 ; P1_R1162_U64
g12851 nand P1_R1162_U186 P1_R1162_U185 P1_R1162_U187 ; P1_R1162_U65
g12852 nand P1_R1162_U179 P1_R1162_U178 ; P1_R1162_U66
g12853 nand P1_R1162_U56 P1_R1162_U204 ; P1_R1162_U67
g12854 nand P1_R1162_U259 P1_R1162_U258 ; P1_R1162_U68
g12855 nand P1_R1162_U308 P1_R1162_U307 ; P1_R1162_U69
g12856 nand P1_R1162_U231 P1_R1162_U230 ; P1_R1162_U70
g12857 nand P1_R1162_U236 P1_R1162_U235 ; P1_R1162_U71
g12858 nand P1_R1162_U243 P1_R1162_U242 ; P1_R1162_U72
g12859 nand P1_R1162_U250 P1_R1162_U249 ; P1_R1162_U73
g12860 nand P1_R1162_U255 P1_R1162_U254 ; P1_R1162_U74
g12861 nand P1_R1162_U271 P1_R1162_U270 ; P1_R1162_U75
g12862 nand P1_R1162_U278 P1_R1162_U277 ; P1_R1162_U76
g12863 nand P1_R1162_U285 P1_R1162_U284 ; P1_R1162_U77
g12864 nand P1_R1162_U292 P1_R1162_U291 ; P1_R1162_U78
g12865 nand P1_R1162_U299 P1_R1162_U298 ; P1_R1162_U79
g12866 nand P1_R1162_U304 P1_R1162_U303 ; P1_R1162_U80
g12867 nand P1_R1162_U117 P1_R1162_U116 P1_R1162_U118 ; P1_R1162_U81
g12868 nand P1_R1162_U133 P1_R1162_U145 ; P1_R1162_U82
g12869 nand P1_R1162_U41 P1_R1162_U152 ; P1_R1162_U83
g12870 not P1_U3452 ; P1_R1162_U84
g12871 not P1_REG1_REG_19__SCAN_IN ; P1_R1162_U85
g12872 nand P1_R1162_U175 P1_R1162_U174 ; P1_R1162_U86
g12873 nand P1_R1162_U171 P1_R1162_U170 ; P1_R1162_U87
g12874 nand P1_R1162_U161 P1_R1162_U160 ; P1_R1162_U88
g12875 not P1_R1162_U32 ; P1_R1162_U89
g12876 nand P1_U3484 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U90
g12877 nand P1_U3493 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U91
g12878 not P1_R1162_U56 ; P1_R1162_U92
g12879 not P1_R1162_U49 ; P1_R1162_U93
g12880 or P1_U3472 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U94
g12881 or P1_U3469 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U95
g12882 or P1_U3466 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U96
g12883 or P1_U3463 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U97
g12884 not P1_R1162_U29 ; P1_R1162_U98
g12885 or P1_U3460 P1_REG1_REG_1__SCAN_IN ; P1_R1162_U99
g12886 not P1_R1162_U40 ; P1_R1162_U100
g12887 not P1_R1162_U41 ; P1_R1162_U101
g12888 nand P1_R1162_U40 P1_R1162_U41 ; P1_R1162_U102
g12889 nand P1_U3463 P1_R1162_U96 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U103
g12890 nand P1_R1162_U5 P1_R1162_U102 ; P1_R1162_U104
g12891 nand P1_U3466 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U105
g12892 nand P1_R1162_U105 P1_R1162_U103 P1_R1162_U104 ; P1_R1162_U106
g12893 nand P1_R1162_U33 P1_R1162_U32 ; P1_R1162_U107
g12894 nand P1_U3472 P1_R1162_U107 ; P1_R1162_U108
g12895 nand P1_R1162_U4 P1_R1162_U106 ; P1_R1162_U109
g12896 nand P1_R1162_U89 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U110
g12897 not P1_R1162_U39 ; P1_R1162_U111
g12898 or P1_U3478 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U112
g12899 or P1_U3475 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U113
g12900 not P1_R1162_U20 ; P1_R1162_U114
g12901 nand P1_R1162_U21 P1_R1162_U20 ; P1_R1162_U115
g12902 nand P1_U3478 P1_R1162_U115 ; P1_R1162_U116
g12903 nand P1_R1162_U114 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U117
g12904 nand P1_R1162_U6 P1_R1162_U39 ; P1_R1162_U118
g12905 not P1_R1162_U81 ; P1_R1162_U119
g12906 or P1_U3481 P1_REG1_REG_8__SCAN_IN ; P1_R1162_U120
g12907 nand P1_R1162_U120 P1_R1162_U81 ; P1_R1162_U121
g12908 not P1_R1162_U38 ; P1_R1162_U122
g12909 or P1_U3484 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U123
g12910 or P1_U3475 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U124
g12911 nand P1_R1162_U124 P1_R1162_U39 ; P1_R1162_U125
g12912 nand P1_R1162_U238 P1_R1162_U237 P1_R1162_U20 P1_R1162_U125 ; P1_R1162_U126
g12913 nand P1_R1162_U111 P1_R1162_U20 ; P1_R1162_U127
g12914 nand P1_U3478 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U128
g12915 nand P1_R1162_U128 P1_R1162_U6 P1_R1162_U127 ; P1_R1162_U129
g12916 or P1_U3475 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U130
g12917 nand P1_R1162_U101 P1_R1162_U97 ; P1_R1162_U131
g12918 nand P1_U3463 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U132
g12919 not P1_R1162_U43 ; P1_R1162_U133
g12920 nand P1_R1162_U100 P1_R1162_U5 ; P1_R1162_U134
g12921 nand P1_R1162_U43 P1_R1162_U96 ; P1_R1162_U135
g12922 nand P1_U3466 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U136
g12923 not P1_R1162_U42 ; P1_R1162_U137
g12924 or P1_U3469 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U138
g12925 nand P1_R1162_U138 P1_R1162_U42 ; P1_R1162_U139
g12926 nand P1_R1162_U245 P1_R1162_U244 P1_R1162_U32 P1_R1162_U139 ; P1_R1162_U140
g12927 nand P1_R1162_U137 P1_R1162_U32 ; P1_R1162_U141
g12928 nand P1_U3472 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U142
g12929 nand P1_R1162_U142 P1_R1162_U4 P1_R1162_U141 ; P1_R1162_U143
g12930 or P1_U3469 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U144
g12931 nand P1_R1162_U100 P1_R1162_U97 ; P1_R1162_U145
g12932 not P1_R1162_U82 ; P1_R1162_U146
g12933 nand P1_U3466 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U147
g12934 nand P1_R1162_U257 P1_R1162_U256 P1_R1162_U41 P1_R1162_U40 ; P1_R1162_U148
g12935 nand P1_R1162_U41 P1_R1162_U40 ; P1_R1162_U149
g12936 nand P1_U3463 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U150
g12937 nand P1_R1162_U150 P1_R1162_U97 P1_R1162_U149 ; P1_R1162_U151
g12938 or P1_U3460 P1_REG1_REG_1__SCAN_IN ; P1_R1162_U152
g12939 not P1_R1162_U83 ; P1_R1162_U153
g12940 or P1_U3484 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U154
g12941 or P1_U3487 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U155
g12942 nand P1_R1162_U93 P1_R1162_U7 ; P1_R1162_U156
g12943 nand P1_U3487 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U157
g12944 nand P1_R1162_U157 P1_R1162_U90 P1_R1162_U156 ; P1_R1162_U158
g12945 or P1_U3487 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U159
g12946 nand P1_R1162_U120 P1_R1162_U7 P1_R1162_U81 ; P1_R1162_U160
g12947 nand P1_R1162_U159 P1_R1162_U158 ; P1_R1162_U161
g12948 not P1_R1162_U88 ; P1_R1162_U162
g12949 or P1_U3496 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U163
g12950 or P1_U3493 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U164
g12951 nand P1_R1162_U92 P1_R1162_U8 ; P1_R1162_U165
g12952 nand P1_U3496 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U166
g12953 nand P1_R1162_U166 P1_R1162_U91 P1_R1162_U165 ; P1_R1162_U167
g12954 or P1_U3490 P1_REG1_REG_11__SCAN_IN ; P1_R1162_U168
g12955 or P1_U3496 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U169
g12956 nand P1_R1162_U168 P1_R1162_U8 P1_R1162_U88 ; P1_R1162_U170
g12957 nand P1_R1162_U169 P1_R1162_U167 ; P1_R1162_U171
g12958 not P1_R1162_U87 ; P1_R1162_U172
g12959 or P1_U3499 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U173
g12960 nand P1_R1162_U173 P1_R1162_U87 ; P1_R1162_U174
g12961 nand P1_U3499 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U175
g12962 not P1_R1162_U86 ; P1_R1162_U176
g12963 or P1_U3502 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U177
g12964 nand P1_R1162_U177 P1_R1162_U86 ; P1_R1162_U178
g12965 nand P1_U3502 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U179
g12966 not P1_R1162_U66 ; P1_R1162_U180
g12967 or P1_U3508 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U181
g12968 or P1_U3505 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U182
g12969 not P1_R1162_U47 ; P1_R1162_U183
g12970 nand P1_R1162_U48 P1_R1162_U47 ; P1_R1162_U184
g12971 nand P1_U3508 P1_R1162_U184 ; P1_R1162_U185
g12972 nand P1_R1162_U183 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U186
g12973 nand P1_R1162_U9 P1_R1162_U66 ; P1_R1162_U187
g12974 not P1_R1162_U65 ; P1_R1162_U188
g12975 or P1_U3511 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U189
g12976 nand P1_R1162_U189 P1_R1162_U65 ; P1_R1162_U190
g12977 nand P1_U3511 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U191
g12978 nand P1_R1162_U261 P1_R1162_U260 P1_R1162_U191 P1_R1162_U190 ; P1_R1162_U192
g12979 nand P1_U3511 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U193
g12980 nand P1_R1162_U188 P1_R1162_U193 ; P1_R1162_U194
g12981 or P1_U3511 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U195
g12982 nand P1_R1162_U195 P1_R1162_U264 P1_R1162_U194 ; P1_R1162_U196
g12983 or P1_U3505 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U197
g12984 nand P1_R1162_U197 P1_R1162_U66 ; P1_R1162_U198
g12985 nand P1_R1162_U273 P1_R1162_U272 P1_R1162_U47 P1_R1162_U198 ; P1_R1162_U199
g12986 nand P1_R1162_U180 P1_R1162_U47 ; P1_R1162_U200
g12987 nand P1_U3508 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U201
g12988 nand P1_R1162_U201 P1_R1162_U9 P1_R1162_U200 ; P1_R1162_U202
g12989 or P1_U3505 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U203
g12990 nand P1_R1162_U168 P1_R1162_U88 ; P1_R1162_U204
g12991 not P1_R1162_U67 ; P1_R1162_U205
g12992 or P1_U3493 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U206
g12993 nand P1_R1162_U206 P1_R1162_U67 ; P1_R1162_U207
g12994 nand P1_R1162_U294 P1_R1162_U293 P1_R1162_U91 P1_R1162_U207 ; P1_R1162_U208
g12995 nand P1_R1162_U205 P1_R1162_U91 ; P1_R1162_U209
g12996 nand P1_U3496 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U210
g12997 nand P1_R1162_U210 P1_R1162_U8 P1_R1162_U209 ; P1_R1162_U211
g12998 or P1_U3493 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U212
g12999 or P1_U3484 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U213
g13000 nand P1_R1162_U213 P1_R1162_U38 ; P1_R1162_U214
g13001 nand P1_R1162_U306 P1_R1162_U305 P1_R1162_U90 P1_R1162_U214 ; P1_R1162_U215
g13002 nand P1_R1162_U122 P1_R1162_U90 ; P1_R1162_U216
g13003 nand P1_U3487 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U217
g13004 nand P1_R1162_U217 P1_R1162_U7 P1_R1162_U216 ; P1_R1162_U218
g13005 nand P1_R1162_U123 P1_R1162_U90 ; P1_R1162_U219
g13006 nand P1_R1162_U120 P1_R1162_U49 ; P1_R1162_U220
g13007 nand P1_R1162_U130 P1_R1162_U20 ; P1_R1162_U221
g13008 nand P1_R1162_U144 P1_R1162_U32 ; P1_R1162_U222
g13009 nand P1_R1162_U147 P1_R1162_U96 ; P1_R1162_U223
g13010 nand P1_R1162_U203 P1_R1162_U47 ; P1_R1162_U224
g13011 nand P1_R1162_U212 P1_R1162_U91 ; P1_R1162_U225
g13012 nand P1_R1162_U168 P1_R1162_U56 ; P1_R1162_U226
g13013 nand P1_U3484 P1_R1162_U37 ; P1_R1162_U227
g13014 nand P1_R1162_U36 P1_REG1_REG_9__SCAN_IN ; P1_R1162_U228
g13015 nand P1_R1162_U228 P1_R1162_U227 ; P1_R1162_U229
g13016 nand P1_R1162_U219 P1_R1162_U38 ; P1_R1162_U230
g13017 nand P1_R1162_U229 P1_R1162_U122 ; P1_R1162_U231
g13018 nand P1_U3481 P1_R1162_U34 ; P1_R1162_U232
g13019 nand P1_R1162_U35 P1_REG1_REG_8__SCAN_IN ; P1_R1162_U233
g13020 nand P1_R1162_U233 P1_R1162_U232 ; P1_R1162_U234
g13021 nand P1_R1162_U220 P1_R1162_U81 ; P1_R1162_U235
g13022 nand P1_R1162_U119 P1_R1162_U234 ; P1_R1162_U236
g13023 nand P1_U3478 P1_R1162_U21 ; P1_R1162_U237
g13024 nand P1_R1162_U19 P1_REG1_REG_7__SCAN_IN ; P1_R1162_U238
g13025 nand P1_U3475 P1_R1162_U17 ; P1_R1162_U239
g13026 nand P1_R1162_U18 P1_REG1_REG_6__SCAN_IN ; P1_R1162_U240
g13027 nand P1_R1162_U240 P1_R1162_U239 ; P1_R1162_U241
g13028 nand P1_R1162_U221 P1_R1162_U39 ; P1_R1162_U242
g13029 nand P1_R1162_U241 P1_R1162_U111 ; P1_R1162_U243
g13030 nand P1_U3472 P1_R1162_U33 ; P1_R1162_U244
g13031 nand P1_R1162_U24 P1_REG1_REG_5__SCAN_IN ; P1_R1162_U245
g13032 nand P1_U3469 P1_R1162_U22 ; P1_R1162_U246
g13033 nand P1_R1162_U23 P1_REG1_REG_4__SCAN_IN ; P1_R1162_U247
g13034 nand P1_R1162_U247 P1_R1162_U246 ; P1_R1162_U248
g13035 nand P1_R1162_U222 P1_R1162_U42 ; P1_R1162_U249
g13036 nand P1_R1162_U248 P1_R1162_U137 ; P1_R1162_U250
g13037 nand P1_U3466 P1_R1162_U30 ; P1_R1162_U251
g13038 nand P1_R1162_U31 P1_REG1_REG_3__SCAN_IN ; P1_R1162_U252
g13039 nand P1_R1162_U252 P1_R1162_U251 ; P1_R1162_U253
g13040 nand P1_R1162_U223 P1_R1162_U82 ; P1_R1162_U254
g13041 nand P1_R1162_U146 P1_R1162_U253 ; P1_R1162_U255
g13042 nand P1_U3463 P1_R1162_U25 ; P1_R1162_U256
g13043 nand P1_R1162_U26 P1_REG1_REG_2__SCAN_IN ; P1_R1162_U257
g13044 nand P1_R1162_U98 P1_R1162_U83 ; P1_R1162_U258
g13045 nand P1_R1162_U153 P1_R1162_U29 ; P1_R1162_U259
g13046 nand P1_U3452 P1_R1162_U85 ; P1_R1162_U260
g13047 nand P1_R1162_U84 P1_REG1_REG_19__SCAN_IN ; P1_R1162_U261
g13048 nand P1_U3452 P1_R1162_U85 ; P1_R1162_U262
g13049 nand P1_R1162_U84 P1_REG1_REG_19__SCAN_IN ; P1_R1162_U263
g13050 nand P1_R1162_U263 P1_R1162_U262 ; P1_R1162_U264
g13051 nand P1_U3511 P1_R1162_U63 ; P1_R1162_U265
g13052 nand P1_R1162_U64 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U266
g13053 nand P1_U3511 P1_R1162_U63 ; P1_R1162_U267
g13054 nand P1_R1162_U64 P1_REG1_REG_18__SCAN_IN ; P1_R1162_U268
g13055 nand P1_R1162_U268 P1_R1162_U267 ; P1_R1162_U269
g13056 nand P1_R1162_U266 P1_R1162_U265 P1_R1162_U65 ; P1_R1162_U270
g13057 nand P1_R1162_U269 P1_R1162_U188 ; P1_R1162_U271
g13058 nand P1_U3508 P1_R1162_U48 ; P1_R1162_U272
g13059 nand P1_R1162_U46 P1_REG1_REG_17__SCAN_IN ; P1_R1162_U273
g13060 nand P1_U3505 P1_R1162_U44 ; P1_R1162_U274
g13061 nand P1_R1162_U45 P1_REG1_REG_16__SCAN_IN ; P1_R1162_U275
g13062 nand P1_R1162_U275 P1_R1162_U274 ; P1_R1162_U276
g13063 nand P1_R1162_U224 P1_R1162_U66 ; P1_R1162_U277
g13064 nand P1_R1162_U276 P1_R1162_U180 ; P1_R1162_U278
g13065 nand P1_U3502 P1_R1162_U61 ; P1_R1162_U279
g13066 nand P1_R1162_U62 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U280
g13067 nand P1_U3502 P1_R1162_U61 ; P1_R1162_U281
g13068 nand P1_R1162_U62 P1_REG1_REG_15__SCAN_IN ; P1_R1162_U282
g13069 nand P1_R1162_U282 P1_R1162_U281 ; P1_R1162_U283
g13070 nand P1_R1162_U280 P1_R1162_U279 P1_R1162_U86 ; P1_R1162_U284
g13071 nand P1_R1162_U176 P1_R1162_U283 ; P1_R1162_U285
g13072 nand P1_U3499 P1_R1162_U59 ; P1_R1162_U286
g13073 nand P1_R1162_U60 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U287
g13074 nand P1_U3499 P1_R1162_U59 ; P1_R1162_U288
g13075 nand P1_R1162_U60 P1_REG1_REG_14__SCAN_IN ; P1_R1162_U289
g13076 nand P1_R1162_U289 P1_R1162_U288 ; P1_R1162_U290
g13077 nand P1_R1162_U287 P1_R1162_U286 P1_R1162_U87 ; P1_R1162_U291
g13078 nand P1_R1162_U172 P1_R1162_U290 ; P1_R1162_U292
g13079 nand P1_U3496 P1_R1162_U57 ; P1_R1162_U293
g13080 nand P1_R1162_U58 P1_REG1_REG_13__SCAN_IN ; P1_R1162_U294
g13081 nand P1_U3493 P1_R1162_U52 ; P1_R1162_U295
g13082 nand P1_R1162_U53 P1_REG1_REG_12__SCAN_IN ; P1_R1162_U296
g13083 nand P1_R1162_U296 P1_R1162_U295 ; P1_R1162_U297
g13084 nand P1_R1162_U225 P1_R1162_U67 ; P1_R1162_U298
g13085 nand P1_R1162_U297 P1_R1162_U205 ; P1_R1162_U299
g13086 nand P1_U3490 P1_R1162_U54 ; P1_R1162_U300
g13087 nand P1_R1162_U55 P1_REG1_REG_11__SCAN_IN ; P1_R1162_U301
g13088 nand P1_R1162_U301 P1_R1162_U300 ; P1_R1162_U302
g13089 nand P1_R1162_U226 P1_R1162_U88 ; P1_R1162_U303
g13090 nand P1_R1162_U162 P1_R1162_U302 ; P1_R1162_U304
g13091 nand P1_U3487 P1_R1162_U50 ; P1_R1162_U305
g13092 nand P1_R1162_U51 P1_REG1_REG_10__SCAN_IN ; P1_R1162_U306
g13093 nand P1_U3454 P1_R1162_U27 ; P1_R1162_U307
g13094 nand P1_R1162_U28 P1_REG1_REG_0__SCAN_IN ; P1_R1162_U308
g13095 and P1_R1117_U184 P1_R1117_U201 ; P1_R1117_U6
g13096 and P1_R1117_U203 P1_R1117_U202 ; P1_R1117_U7
g13097 and P1_R1117_U179 P1_R1117_U240 ; P1_R1117_U8
g13098 and P1_R1117_U242 P1_R1117_U241 ; P1_R1117_U9
g13099 and P1_R1117_U259 P1_R1117_U258 ; P1_R1117_U10
g13100 and P1_R1117_U285 P1_R1117_U284 ; P1_R1117_U11
g13101 and P1_R1117_U383 P1_R1117_U382 ; P1_R1117_U12
g13102 nand P1_R1117_U340 P1_R1117_U343 ; P1_R1117_U13
g13103 nand P1_R1117_U329 P1_R1117_U332 ; P1_R1117_U14
g13104 nand P1_R1117_U318 P1_R1117_U321 ; P1_R1117_U15
g13105 nand P1_R1117_U310 P1_R1117_U312 ; P1_R1117_U16
g13106 nand P1_R1117_U156 P1_R1117_U175 P1_R1117_U348 ; P1_R1117_U17
g13107 nand P1_R1117_U236 P1_R1117_U238 ; P1_R1117_U18
g13108 nand P1_R1117_U228 P1_R1117_U231 ; P1_R1117_U19
g13109 nand P1_R1117_U220 P1_R1117_U222 ; P1_R1117_U20
g13110 nand P1_R1117_U25 P1_R1117_U346 ; P1_R1117_U21
g13111 not P1_U3479 ; P1_R1117_U22
g13112 not P1_U3464 ; P1_R1117_U23
g13113 not P1_U3456 ; P1_R1117_U24
g13114 nand P1_U3456 P1_R1117_U93 ; P1_R1117_U25
g13115 not P1_U3078 ; P1_R1117_U26
g13116 not P1_U3467 ; P1_R1117_U27
g13117 not P1_U3068 ; P1_R1117_U28
g13118 nand P1_U3068 P1_R1117_U23 ; P1_R1117_U29
g13119 not P1_U3064 ; P1_R1117_U30
g13120 not P1_U3476 ; P1_R1117_U31
g13121 not P1_U3473 ; P1_R1117_U32
g13122 not P1_U3470 ; P1_R1117_U33
g13123 not P1_U3071 ; P1_R1117_U34
g13124 not P1_U3067 ; P1_R1117_U35
g13125 not P1_U3060 ; P1_R1117_U36
g13126 nand P1_U3060 P1_R1117_U33 ; P1_R1117_U37
g13127 not P1_U3482 ; P1_R1117_U38
g13128 not P1_U3070 ; P1_R1117_U39
g13129 nand P1_U3070 P1_R1117_U22 ; P1_R1117_U40
g13130 not P1_U3084 ; P1_R1117_U41
g13131 not P1_U3485 ; P1_R1117_U42
g13132 not P1_U3083 ; P1_R1117_U43
g13133 nand P1_R1117_U209 P1_R1117_U208 ; P1_R1117_U44
g13134 nand P1_R1117_U37 P1_R1117_U224 ; P1_R1117_U45
g13135 nand P1_R1117_U193 P1_R1117_U192 ; P1_R1117_U46
g13136 not P1_U4019 ; P1_R1117_U47
g13137 not P1_U4023 ; P1_R1117_U48
g13138 not P1_U3503 ; P1_R1117_U49
g13139 not P1_U3491 ; P1_R1117_U50
g13140 not P1_U3488 ; P1_R1117_U51
g13141 not P1_U3063 ; P1_R1117_U52
g13142 not P1_U3062 ; P1_R1117_U53
g13143 nand P1_U3083 P1_R1117_U42 ; P1_R1117_U54
g13144 not P1_U3494 ; P1_R1117_U55
g13145 not P1_U3072 ; P1_R1117_U56
g13146 not P1_U3497 ; P1_R1117_U57
g13147 not P1_U3080 ; P1_R1117_U58
g13148 not P1_U3506 ; P1_R1117_U59
g13149 not P1_U3500 ; P1_R1117_U60
g13150 not P1_U3073 ; P1_R1117_U61
g13151 not P1_U3074 ; P1_R1117_U62
g13152 not P1_U3079 ; P1_R1117_U63
g13153 nand P1_U3079 P1_R1117_U60 ; P1_R1117_U64
g13154 not P1_U3509 ; P1_R1117_U65
g13155 not P1_U3069 ; P1_R1117_U66
g13156 nand P1_R1117_U269 P1_R1117_U268 ; P1_R1117_U67
g13157 not P1_U3082 ; P1_R1117_U68
g13158 not P1_U3514 ; P1_R1117_U69
g13159 not P1_U3081 ; P1_R1117_U70
g13160 not P1_U4025 ; P1_R1117_U71
g13161 not P1_U3076 ; P1_R1117_U72
g13162 not P1_U4022 ; P1_R1117_U73
g13163 not P1_U4024 ; P1_R1117_U74
g13164 not P1_U3066 ; P1_R1117_U75
g13165 not P1_U3061 ; P1_R1117_U76
g13166 not P1_U3075 ; P1_R1117_U77
g13167 nand P1_U3075 P1_R1117_U74 ; P1_R1117_U78
g13168 not P1_U4021 ; P1_R1117_U79
g13169 not P1_U3065 ; P1_R1117_U80
g13170 not P1_U4020 ; P1_R1117_U81
g13171 not P1_U3058 ; P1_R1117_U82
g13172 not P1_U4018 ; P1_R1117_U83
g13173 not P1_U3057 ; P1_R1117_U84
g13174 nand P1_U3057 P1_R1117_U47 ; P1_R1117_U85
g13175 not P1_U3053 ; P1_R1117_U86
g13176 not P1_U4017 ; P1_R1117_U87
g13177 not P1_U3054 ; P1_R1117_U88
g13178 nand P1_R1117_U299 P1_R1117_U298 ; P1_R1117_U89
g13179 nand P1_R1117_U78 P1_R1117_U314 ; P1_R1117_U90
g13180 nand P1_R1117_U64 P1_R1117_U325 ; P1_R1117_U91
g13181 nand P1_R1117_U54 P1_R1117_U336 ; P1_R1117_U92
g13182 not P1_U3077 ; P1_R1117_U93
g13183 nand P1_R1117_U393 P1_R1117_U392 ; P1_R1117_U94
g13184 nand P1_R1117_U407 P1_R1117_U406 ; P1_R1117_U95
g13185 nand P1_R1117_U412 P1_R1117_U411 ; P1_R1117_U96
g13186 nand P1_R1117_U428 P1_R1117_U427 ; P1_R1117_U97
g13187 nand P1_R1117_U433 P1_R1117_U432 ; P1_R1117_U98
g13188 nand P1_R1117_U438 P1_R1117_U437 ; P1_R1117_U99
g13189 nand P1_R1117_U443 P1_R1117_U442 ; P1_R1117_U100
g13190 nand P1_R1117_U448 P1_R1117_U447 ; P1_R1117_U101
g13191 nand P1_R1117_U464 P1_R1117_U463 ; P1_R1117_U102
g13192 nand P1_R1117_U469 P1_R1117_U468 ; P1_R1117_U103
g13193 nand P1_R1117_U352 P1_R1117_U351 ; P1_R1117_U104
g13194 nand P1_R1117_U361 P1_R1117_U360 ; P1_R1117_U105
g13195 nand P1_R1117_U368 P1_R1117_U367 ; P1_R1117_U106
g13196 nand P1_R1117_U372 P1_R1117_U371 ; P1_R1117_U107
g13197 nand P1_R1117_U381 P1_R1117_U380 ; P1_R1117_U108
g13198 nand P1_R1117_U402 P1_R1117_U401 ; P1_R1117_U109
g13199 nand P1_R1117_U419 P1_R1117_U418 ; P1_R1117_U110
g13200 nand P1_R1117_U423 P1_R1117_U422 ; P1_R1117_U111
g13201 nand P1_R1117_U455 P1_R1117_U454 ; P1_R1117_U112
g13202 nand P1_R1117_U459 P1_R1117_U458 ; P1_R1117_U113
g13203 nand P1_R1117_U476 P1_R1117_U475 ; P1_R1117_U114
g13204 and P1_R1117_U195 P1_R1117_U183 ; P1_R1117_U115
g13205 and P1_R1117_U198 P1_R1117_U199 ; P1_R1117_U116
g13206 and P1_R1117_U211 P1_R1117_U185 ; P1_R1117_U117
g13207 and P1_R1117_U214 P1_R1117_U215 ; P1_R1117_U118
g13208 and P1_R1117_U354 P1_R1117_U353 P1_R1117_U40 ; P1_R1117_U119
g13209 and P1_R1117_U357 P1_R1117_U185 ; P1_R1117_U120
g13210 and P1_R1117_U230 P1_R1117_U7 ; P1_R1117_U121
g13211 and P1_R1117_U364 P1_R1117_U184 ; P1_R1117_U122
g13212 and P1_R1117_U374 P1_R1117_U373 P1_R1117_U29 ; P1_R1117_U123
g13213 and P1_R1117_U377 P1_R1117_U183 ; P1_R1117_U124
g13214 and P1_R1117_U217 P1_R1117_U8 ; P1_R1117_U125
g13215 and P1_R1117_U262 P1_R1117_U180 ; P1_R1117_U126
g13216 and P1_R1117_U288 P1_R1117_U181 ; P1_R1117_U127
g13217 and P1_R1117_U304 P1_R1117_U305 ; P1_R1117_U128
g13218 and P1_R1117_U307 P1_R1117_U386 ; P1_R1117_U129
g13219 and P1_R1117_U305 P1_R1117_U304 P1_R1117_U308 ; P1_R1117_U130
g13220 nand P1_R1117_U390 P1_R1117_U389 ; P1_R1117_U131
g13221 and P1_R1117_U395 P1_R1117_U394 P1_R1117_U85 ; P1_R1117_U132
g13222 and P1_R1117_U398 P1_R1117_U182 ; P1_R1117_U133
g13223 nand P1_R1117_U404 P1_R1117_U403 ; P1_R1117_U134
g13224 nand P1_R1117_U409 P1_R1117_U408 ; P1_R1117_U135
g13225 and P1_R1117_U415 P1_R1117_U181 ; P1_R1117_U136
g13226 nand P1_R1117_U425 P1_R1117_U424 ; P1_R1117_U137
g13227 nand P1_R1117_U430 P1_R1117_U429 ; P1_R1117_U138
g13228 nand P1_R1117_U435 P1_R1117_U434 ; P1_R1117_U139
g13229 nand P1_R1117_U440 P1_R1117_U439 ; P1_R1117_U140
g13230 nand P1_R1117_U445 P1_R1117_U444 ; P1_R1117_U141
g13231 and P1_R1117_U451 P1_R1117_U180 ; P1_R1117_U142
g13232 nand P1_R1117_U461 P1_R1117_U460 ; P1_R1117_U143
g13233 nand P1_R1117_U466 P1_R1117_U465 ; P1_R1117_U144
g13234 and P1_R1117_U342 P1_R1117_U9 ; P1_R1117_U145
g13235 and P1_R1117_U472 P1_R1117_U179 ; P1_R1117_U146
g13236 and P1_R1117_U350 P1_R1117_U349 ; P1_R1117_U147
g13237 nand P1_R1117_U118 P1_R1117_U212 ; P1_R1117_U148
g13238 and P1_R1117_U359 P1_R1117_U358 ; P1_R1117_U149
g13239 and P1_R1117_U366 P1_R1117_U365 ; P1_R1117_U150
g13240 and P1_R1117_U370 P1_R1117_U369 ; P1_R1117_U151
g13241 nand P1_R1117_U116 P1_R1117_U196 ; P1_R1117_U152
g13242 and P1_R1117_U379 P1_R1117_U378 ; P1_R1117_U153
g13243 not P1_U4028 ; P1_R1117_U154
g13244 not P1_U3055 ; P1_R1117_U155
g13245 and P1_R1117_U388 P1_R1117_U387 ; P1_R1117_U156
g13246 nand P1_R1117_U128 P1_R1117_U302 ; P1_R1117_U157
g13247 and P1_R1117_U400 P1_R1117_U399 ; P1_R1117_U158
g13248 nand P1_R1117_U295 P1_R1117_U294 ; P1_R1117_U159
g13249 nand P1_R1117_U291 P1_R1117_U290 ; P1_R1117_U160
g13250 and P1_R1117_U417 P1_R1117_U416 ; P1_R1117_U161
g13251 and P1_R1117_U421 P1_R1117_U420 ; P1_R1117_U162
g13252 nand P1_R1117_U281 P1_R1117_U280 ; P1_R1117_U163
g13253 nand P1_R1117_U277 P1_R1117_U276 ; P1_R1117_U164
g13254 not P1_U3461 ; P1_R1117_U165
g13255 nand P1_R1117_U273 P1_R1117_U272 ; P1_R1117_U166
g13256 not P1_U3512 ; P1_R1117_U167
g13257 nand P1_R1117_U265 P1_R1117_U264 ; P1_R1117_U168
g13258 and P1_R1117_U453 P1_R1117_U452 ; P1_R1117_U169
g13259 and P1_R1117_U457 P1_R1117_U456 ; P1_R1117_U170
g13260 nand P1_R1117_U255 P1_R1117_U254 ; P1_R1117_U171
g13261 nand P1_R1117_U251 P1_R1117_U250 ; P1_R1117_U172
g13262 nand P1_R1117_U247 P1_R1117_U246 ; P1_R1117_U173
g13263 and P1_R1117_U474 P1_R1117_U473 ; P1_R1117_U174
g13264 nand P1_R1117_U129 P1_R1117_U157 ; P1_R1117_U175
g13265 not P1_R1117_U85 ; P1_R1117_U176
g13266 not P1_R1117_U29 ; P1_R1117_U177
g13267 not P1_R1117_U40 ; P1_R1117_U178
g13268 nand P1_U3488 P1_R1117_U53 ; P1_R1117_U179
g13269 nand P1_U3503 P1_R1117_U62 ; P1_R1117_U180
g13270 nand P1_U4023 P1_R1117_U76 ; P1_R1117_U181
g13271 nand P1_U4019 P1_R1117_U84 ; P1_R1117_U182
g13272 nand P1_U3464 P1_R1117_U28 ; P1_R1117_U183
g13273 nand P1_U3473 P1_R1117_U35 ; P1_R1117_U184
g13274 nand P1_U3479 P1_R1117_U39 ; P1_R1117_U185
g13275 not P1_R1117_U64 ; P1_R1117_U186
g13276 not P1_R1117_U78 ; P1_R1117_U187
g13277 not P1_R1117_U37 ; P1_R1117_U188
g13278 not P1_R1117_U54 ; P1_R1117_U189
g13279 not P1_R1117_U25 ; P1_R1117_U190
g13280 nand P1_R1117_U190 P1_R1117_U26 ; P1_R1117_U191
g13281 nand P1_R1117_U191 P1_R1117_U165 ; P1_R1117_U192
g13282 nand P1_U3078 P1_R1117_U25 ; P1_R1117_U193
g13283 not P1_R1117_U46 ; P1_R1117_U194
g13284 nand P1_U3467 P1_R1117_U30 ; P1_R1117_U195
g13285 nand P1_R1117_U115 P1_R1117_U46 ; P1_R1117_U196
g13286 nand P1_R1117_U30 P1_R1117_U29 ; P1_R1117_U197
g13287 nand P1_R1117_U197 P1_R1117_U27 ; P1_R1117_U198
g13288 nand P1_U3064 P1_R1117_U177 ; P1_R1117_U199
g13289 not P1_R1117_U152 ; P1_R1117_U200
g13290 nand P1_U3476 P1_R1117_U34 ; P1_R1117_U201
g13291 nand P1_U3071 P1_R1117_U31 ; P1_R1117_U202
g13292 nand P1_U3067 P1_R1117_U32 ; P1_R1117_U203
g13293 nand P1_R1117_U188 P1_R1117_U6 ; P1_R1117_U204
g13294 nand P1_R1117_U7 P1_R1117_U204 ; P1_R1117_U205
g13295 nand P1_U3470 P1_R1117_U36 ; P1_R1117_U206
g13296 nand P1_U3476 P1_R1117_U34 ; P1_R1117_U207
g13297 nand P1_R1117_U206 P1_R1117_U152 P1_R1117_U6 ; P1_R1117_U208
g13298 nand P1_R1117_U207 P1_R1117_U205 ; P1_R1117_U209
g13299 not P1_R1117_U44 ; P1_R1117_U210
g13300 nand P1_U3482 P1_R1117_U41 ; P1_R1117_U211
g13301 nand P1_R1117_U117 P1_R1117_U44 ; P1_R1117_U212
g13302 nand P1_R1117_U41 P1_R1117_U40 ; P1_R1117_U213
g13303 nand P1_R1117_U213 P1_R1117_U38 ; P1_R1117_U214
g13304 nand P1_U3084 P1_R1117_U178 ; P1_R1117_U215
g13305 not P1_R1117_U148 ; P1_R1117_U216
g13306 nand P1_U3485 P1_R1117_U43 ; P1_R1117_U217
g13307 nand P1_R1117_U217 P1_R1117_U54 ; P1_R1117_U218
g13308 nand P1_R1117_U210 P1_R1117_U40 ; P1_R1117_U219
g13309 nand P1_R1117_U120 P1_R1117_U219 ; P1_R1117_U220
g13310 nand P1_R1117_U44 P1_R1117_U185 ; P1_R1117_U221
g13311 nand P1_R1117_U119 P1_R1117_U221 ; P1_R1117_U222
g13312 nand P1_R1117_U40 P1_R1117_U185 ; P1_R1117_U223
g13313 nand P1_R1117_U206 P1_R1117_U152 ; P1_R1117_U224
g13314 not P1_R1117_U45 ; P1_R1117_U225
g13315 nand P1_U3067 P1_R1117_U32 ; P1_R1117_U226
g13316 nand P1_R1117_U225 P1_R1117_U226 ; P1_R1117_U227
g13317 nand P1_R1117_U122 P1_R1117_U227 ; P1_R1117_U228
g13318 nand P1_R1117_U45 P1_R1117_U184 ; P1_R1117_U229
g13319 nand P1_U3476 P1_R1117_U34 ; P1_R1117_U230
g13320 nand P1_R1117_U121 P1_R1117_U229 ; P1_R1117_U231
g13321 nand P1_U3067 P1_R1117_U32 ; P1_R1117_U232
g13322 nand P1_R1117_U184 P1_R1117_U232 ; P1_R1117_U233
g13323 nand P1_R1117_U206 P1_R1117_U37 ; P1_R1117_U234
g13324 nand P1_R1117_U194 P1_R1117_U29 ; P1_R1117_U235
g13325 nand P1_R1117_U124 P1_R1117_U235 ; P1_R1117_U236
g13326 nand P1_R1117_U46 P1_R1117_U183 ; P1_R1117_U237
g13327 nand P1_R1117_U123 P1_R1117_U237 ; P1_R1117_U238
g13328 nand P1_R1117_U29 P1_R1117_U183 ; P1_R1117_U239
g13329 nand P1_U3491 P1_R1117_U52 ; P1_R1117_U240
g13330 nand P1_U3063 P1_R1117_U50 ; P1_R1117_U241
g13331 nand P1_U3062 P1_R1117_U51 ; P1_R1117_U242
g13332 nand P1_R1117_U189 P1_R1117_U8 ; P1_R1117_U243
g13333 nand P1_R1117_U9 P1_R1117_U243 ; P1_R1117_U244
g13334 nand P1_U3491 P1_R1117_U52 ; P1_R1117_U245
g13335 nand P1_R1117_U125 P1_R1117_U148 ; P1_R1117_U246
g13336 nand P1_R1117_U245 P1_R1117_U244 ; P1_R1117_U247
g13337 not P1_R1117_U173 ; P1_R1117_U248
g13338 nand P1_U3494 P1_R1117_U56 ; P1_R1117_U249
g13339 nand P1_R1117_U249 P1_R1117_U173 ; P1_R1117_U250
g13340 nand P1_U3072 P1_R1117_U55 ; P1_R1117_U251
g13341 not P1_R1117_U172 ; P1_R1117_U252
g13342 nand P1_U3497 P1_R1117_U58 ; P1_R1117_U253
g13343 nand P1_R1117_U253 P1_R1117_U172 ; P1_R1117_U254
g13344 nand P1_U3080 P1_R1117_U57 ; P1_R1117_U255
g13345 not P1_R1117_U171 ; P1_R1117_U256
g13346 nand P1_U3506 P1_R1117_U61 ; P1_R1117_U257
g13347 nand P1_U3073 P1_R1117_U59 ; P1_R1117_U258
g13348 nand P1_U3074 P1_R1117_U49 ; P1_R1117_U259
g13349 nand P1_R1117_U186 P1_R1117_U180 ; P1_R1117_U260
g13350 nand P1_R1117_U10 P1_R1117_U260 ; P1_R1117_U261
g13351 nand P1_U3500 P1_R1117_U63 ; P1_R1117_U262
g13352 nand P1_U3506 P1_R1117_U61 ; P1_R1117_U263
g13353 nand P1_R1117_U171 P1_R1117_U126 P1_R1117_U257 ; P1_R1117_U264
g13354 nand P1_R1117_U263 P1_R1117_U261 ; P1_R1117_U265
g13355 not P1_R1117_U168 ; P1_R1117_U266
g13356 nand P1_U3509 P1_R1117_U66 ; P1_R1117_U267
g13357 nand P1_R1117_U267 P1_R1117_U168 ; P1_R1117_U268
g13358 nand P1_U3069 P1_R1117_U65 ; P1_R1117_U269
g13359 not P1_R1117_U67 ; P1_R1117_U270
g13360 nand P1_R1117_U270 P1_R1117_U68 ; P1_R1117_U271
g13361 nand P1_R1117_U271 P1_R1117_U167 ; P1_R1117_U272
g13362 nand P1_U3082 P1_R1117_U67 ; P1_R1117_U273
g13363 not P1_R1117_U166 ; P1_R1117_U274
g13364 nand P1_U3514 P1_R1117_U70 ; P1_R1117_U275
g13365 nand P1_R1117_U275 P1_R1117_U166 ; P1_R1117_U276
g13366 nand P1_U3081 P1_R1117_U69 ; P1_R1117_U277
g13367 not P1_R1117_U164 ; P1_R1117_U278
g13368 nand P1_U4025 P1_R1117_U72 ; P1_R1117_U279
g13369 nand P1_R1117_U279 P1_R1117_U164 ; P1_R1117_U280
g13370 nand P1_U3076 P1_R1117_U71 ; P1_R1117_U281
g13371 not P1_R1117_U163 ; P1_R1117_U282
g13372 nand P1_U4022 P1_R1117_U75 ; P1_R1117_U283
g13373 nand P1_U3066 P1_R1117_U73 ; P1_R1117_U284
g13374 nand P1_U3061 P1_R1117_U48 ; P1_R1117_U285
g13375 nand P1_R1117_U187 P1_R1117_U181 ; P1_R1117_U286
g13376 nand P1_R1117_U11 P1_R1117_U286 ; P1_R1117_U287
g13377 nand P1_U4024 P1_R1117_U77 ; P1_R1117_U288
g13378 nand P1_U4022 P1_R1117_U75 ; P1_R1117_U289
g13379 nand P1_R1117_U163 P1_R1117_U127 P1_R1117_U283 ; P1_R1117_U290
g13380 nand P1_R1117_U289 P1_R1117_U287 ; P1_R1117_U291
g13381 not P1_R1117_U160 ; P1_R1117_U292
g13382 nand P1_U4021 P1_R1117_U80 ; P1_R1117_U293
g13383 nand P1_R1117_U293 P1_R1117_U160 ; P1_R1117_U294
g13384 nand P1_U3065 P1_R1117_U79 ; P1_R1117_U295
g13385 not P1_R1117_U159 ; P1_R1117_U296
g13386 nand P1_U4020 P1_R1117_U82 ; P1_R1117_U297
g13387 nand P1_R1117_U297 P1_R1117_U159 ; P1_R1117_U298
g13388 nand P1_U3058 P1_R1117_U81 ; P1_R1117_U299
g13389 not P1_R1117_U89 ; P1_R1117_U300
g13390 nand P1_U4018 P1_R1117_U86 ; P1_R1117_U301
g13391 nand P1_R1117_U89 P1_R1117_U182 P1_R1117_U301 ; P1_R1117_U302
g13392 nand P1_R1117_U86 P1_R1117_U85 ; P1_R1117_U303
g13393 nand P1_R1117_U303 P1_R1117_U83 ; P1_R1117_U304
g13394 nand P1_U3053 P1_R1117_U176 ; P1_R1117_U305
g13395 not P1_R1117_U157 ; P1_R1117_U306
g13396 nand P1_U4017 P1_R1117_U88 ; P1_R1117_U307
g13397 nand P1_U3054 P1_R1117_U87 ; P1_R1117_U308
g13398 nand P1_R1117_U300 P1_R1117_U85 ; P1_R1117_U309
g13399 nand P1_R1117_U133 P1_R1117_U309 ; P1_R1117_U310
g13400 nand P1_R1117_U89 P1_R1117_U182 ; P1_R1117_U311
g13401 nand P1_R1117_U132 P1_R1117_U311 ; P1_R1117_U312
g13402 nand P1_R1117_U85 P1_R1117_U182 ; P1_R1117_U313
g13403 nand P1_R1117_U288 P1_R1117_U163 ; P1_R1117_U314
g13404 not P1_R1117_U90 ; P1_R1117_U315
g13405 nand P1_U3061 P1_R1117_U48 ; P1_R1117_U316
g13406 nand P1_R1117_U315 P1_R1117_U316 ; P1_R1117_U317
g13407 nand P1_R1117_U136 P1_R1117_U317 ; P1_R1117_U318
g13408 nand P1_R1117_U90 P1_R1117_U181 ; P1_R1117_U319
g13409 nand P1_U4022 P1_R1117_U75 ; P1_R1117_U320
g13410 nand P1_R1117_U320 P1_R1117_U319 P1_R1117_U11 ; P1_R1117_U321
g13411 nand P1_U3061 P1_R1117_U48 ; P1_R1117_U322
g13412 nand P1_R1117_U181 P1_R1117_U322 ; P1_R1117_U323
g13413 nand P1_R1117_U288 P1_R1117_U78 ; P1_R1117_U324
g13414 nand P1_R1117_U262 P1_R1117_U171 ; P1_R1117_U325
g13415 not P1_R1117_U91 ; P1_R1117_U326
g13416 nand P1_U3074 P1_R1117_U49 ; P1_R1117_U327
g13417 nand P1_R1117_U326 P1_R1117_U327 ; P1_R1117_U328
g13418 nand P1_R1117_U142 P1_R1117_U328 ; P1_R1117_U329
g13419 nand P1_R1117_U91 P1_R1117_U180 ; P1_R1117_U330
g13420 nand P1_U3506 P1_R1117_U61 ; P1_R1117_U331
g13421 nand P1_R1117_U331 P1_R1117_U330 P1_R1117_U10 ; P1_R1117_U332
g13422 nand P1_U3074 P1_R1117_U49 ; P1_R1117_U333
g13423 nand P1_R1117_U180 P1_R1117_U333 ; P1_R1117_U334
g13424 nand P1_R1117_U262 P1_R1117_U64 ; P1_R1117_U335
g13425 nand P1_R1117_U217 P1_R1117_U148 ; P1_R1117_U336
g13426 not P1_R1117_U92 ; P1_R1117_U337
g13427 nand P1_U3062 P1_R1117_U51 ; P1_R1117_U338
g13428 nand P1_R1117_U337 P1_R1117_U338 ; P1_R1117_U339
g13429 nand P1_R1117_U146 P1_R1117_U339 ; P1_R1117_U340
g13430 nand P1_R1117_U92 P1_R1117_U179 ; P1_R1117_U341
g13431 nand P1_U3491 P1_R1117_U52 ; P1_R1117_U342
g13432 nand P1_R1117_U145 P1_R1117_U341 ; P1_R1117_U343
g13433 nand P1_U3062 P1_R1117_U51 ; P1_R1117_U344
g13434 nand P1_R1117_U179 P1_R1117_U344 ; P1_R1117_U345
g13435 nand P1_U3077 P1_R1117_U24 ; P1_R1117_U346
g13436 nand P1_R1117_U89 P1_R1117_U182 P1_R1117_U301 ; P1_R1117_U347
g13437 nand P1_R1117_U12 P1_R1117_U347 P1_R1117_U130 ; P1_R1117_U348
g13438 nand P1_U3485 P1_R1117_U43 ; P1_R1117_U349
g13439 nand P1_U3083 P1_R1117_U42 ; P1_R1117_U350
g13440 nand P1_R1117_U218 P1_R1117_U148 ; P1_R1117_U351
g13441 nand P1_R1117_U216 P1_R1117_U147 ; P1_R1117_U352
g13442 nand P1_U3482 P1_R1117_U41 ; P1_R1117_U353
g13443 nand P1_U3084 P1_R1117_U38 ; P1_R1117_U354
g13444 nand P1_U3482 P1_R1117_U41 ; P1_R1117_U355
g13445 nand P1_U3084 P1_R1117_U38 ; P1_R1117_U356
g13446 nand P1_R1117_U356 P1_R1117_U355 ; P1_R1117_U357
g13447 nand P1_U3479 P1_R1117_U39 ; P1_R1117_U358
g13448 nand P1_U3070 P1_R1117_U22 ; P1_R1117_U359
g13449 nand P1_R1117_U223 P1_R1117_U44 ; P1_R1117_U360
g13450 nand P1_R1117_U149 P1_R1117_U210 ; P1_R1117_U361
g13451 nand P1_U3476 P1_R1117_U34 ; P1_R1117_U362
g13452 nand P1_U3071 P1_R1117_U31 ; P1_R1117_U363
g13453 nand P1_R1117_U363 P1_R1117_U362 ; P1_R1117_U364
g13454 nand P1_U3473 P1_R1117_U35 ; P1_R1117_U365
g13455 nand P1_U3067 P1_R1117_U32 ; P1_R1117_U366
g13456 nand P1_R1117_U233 P1_R1117_U45 ; P1_R1117_U367
g13457 nand P1_R1117_U150 P1_R1117_U225 ; P1_R1117_U368
g13458 nand P1_U3470 P1_R1117_U36 ; P1_R1117_U369
g13459 nand P1_U3060 P1_R1117_U33 ; P1_R1117_U370
g13460 nand P1_R1117_U234 P1_R1117_U152 ; P1_R1117_U371
g13461 nand P1_R1117_U200 P1_R1117_U151 ; P1_R1117_U372
g13462 nand P1_U3467 P1_R1117_U30 ; P1_R1117_U373
g13463 nand P1_U3064 P1_R1117_U27 ; P1_R1117_U374
g13464 nand P1_U3467 P1_R1117_U30 ; P1_R1117_U375
g13465 nand P1_U3064 P1_R1117_U27 ; P1_R1117_U376
g13466 nand P1_R1117_U376 P1_R1117_U375 ; P1_R1117_U377
g13467 nand P1_U3464 P1_R1117_U28 ; P1_R1117_U378
g13468 nand P1_U3068 P1_R1117_U23 ; P1_R1117_U379
g13469 nand P1_R1117_U239 P1_R1117_U46 ; P1_R1117_U380
g13470 nand P1_R1117_U153 P1_R1117_U194 ; P1_R1117_U381
g13471 nand P1_U4028 P1_R1117_U155 ; P1_R1117_U382
g13472 nand P1_U3055 P1_R1117_U154 ; P1_R1117_U383
g13473 nand P1_U4028 P1_R1117_U155 ; P1_R1117_U384
g13474 nand P1_U3055 P1_R1117_U154 ; P1_R1117_U385
g13475 nand P1_R1117_U385 P1_R1117_U384 ; P1_R1117_U386
g13476 nand P1_U3054 P1_R1117_U386 P1_R1117_U87 ; P1_R1117_U387
g13477 nand P1_R1117_U12 P1_R1117_U88 P1_U4017 ; P1_R1117_U388
g13478 nand P1_U4017 P1_R1117_U88 ; P1_R1117_U389
g13479 nand P1_U3054 P1_R1117_U87 ; P1_R1117_U390
g13480 not P1_R1117_U131 ; P1_R1117_U391
g13481 nand P1_R1117_U306 P1_R1117_U391 ; P1_R1117_U392
g13482 nand P1_R1117_U131 P1_R1117_U157 ; P1_R1117_U393
g13483 nand P1_U4018 P1_R1117_U86 ; P1_R1117_U394
g13484 nand P1_U3053 P1_R1117_U83 ; P1_R1117_U395
g13485 nand P1_U4018 P1_R1117_U86 ; P1_R1117_U396
g13486 nand P1_U3053 P1_R1117_U83 ; P1_R1117_U397
g13487 nand P1_R1117_U397 P1_R1117_U396 ; P1_R1117_U398
g13488 nand P1_U4019 P1_R1117_U84 ; P1_R1117_U399
g13489 nand P1_U3057 P1_R1117_U47 ; P1_R1117_U400
g13490 nand P1_R1117_U313 P1_R1117_U89 ; P1_R1117_U401
g13491 nand P1_R1117_U158 P1_R1117_U300 ; P1_R1117_U402
g13492 nand P1_U4020 P1_R1117_U82 ; P1_R1117_U403
g13493 nand P1_U3058 P1_R1117_U81 ; P1_R1117_U404
g13494 not P1_R1117_U134 ; P1_R1117_U405
g13495 nand P1_R1117_U296 P1_R1117_U405 ; P1_R1117_U406
g13496 nand P1_R1117_U134 P1_R1117_U159 ; P1_R1117_U407
g13497 nand P1_U4021 P1_R1117_U80 ; P1_R1117_U408
g13498 nand P1_U3065 P1_R1117_U79 ; P1_R1117_U409
g13499 not P1_R1117_U135 ; P1_R1117_U410
g13500 nand P1_R1117_U292 P1_R1117_U410 ; P1_R1117_U411
g13501 nand P1_R1117_U135 P1_R1117_U160 ; P1_R1117_U412
g13502 nand P1_U4022 P1_R1117_U75 ; P1_R1117_U413
g13503 nand P1_U3066 P1_R1117_U73 ; P1_R1117_U414
g13504 nand P1_R1117_U414 P1_R1117_U413 ; P1_R1117_U415
g13505 nand P1_U4023 P1_R1117_U76 ; P1_R1117_U416
g13506 nand P1_U3061 P1_R1117_U48 ; P1_R1117_U417
g13507 nand P1_R1117_U323 P1_R1117_U90 ; P1_R1117_U418
g13508 nand P1_R1117_U161 P1_R1117_U315 ; P1_R1117_U419
g13509 nand P1_U4024 P1_R1117_U77 ; P1_R1117_U420
g13510 nand P1_U3075 P1_R1117_U74 ; P1_R1117_U421
g13511 nand P1_R1117_U324 P1_R1117_U163 ; P1_R1117_U422
g13512 nand P1_R1117_U282 P1_R1117_U162 ; P1_R1117_U423
g13513 nand P1_U4025 P1_R1117_U72 ; P1_R1117_U424
g13514 nand P1_U3076 P1_R1117_U71 ; P1_R1117_U425
g13515 not P1_R1117_U137 ; P1_R1117_U426
g13516 nand P1_R1117_U278 P1_R1117_U426 ; P1_R1117_U427
g13517 nand P1_R1117_U137 P1_R1117_U164 ; P1_R1117_U428
g13518 nand P1_U3461 P1_R1117_U26 ; P1_R1117_U429
g13519 nand P1_U3078 P1_R1117_U165 ; P1_R1117_U430
g13520 not P1_R1117_U138 ; P1_R1117_U431
g13521 nand P1_R1117_U431 P1_R1117_U190 ; P1_R1117_U432
g13522 nand P1_R1117_U138 P1_R1117_U25 ; P1_R1117_U433
g13523 nand P1_U3514 P1_R1117_U70 ; P1_R1117_U434
g13524 nand P1_U3081 P1_R1117_U69 ; P1_R1117_U435
g13525 not P1_R1117_U139 ; P1_R1117_U436
g13526 nand P1_R1117_U274 P1_R1117_U436 ; P1_R1117_U437
g13527 nand P1_R1117_U139 P1_R1117_U166 ; P1_R1117_U438
g13528 nand P1_U3512 P1_R1117_U68 ; P1_R1117_U439
g13529 nand P1_U3082 P1_R1117_U167 ; P1_R1117_U440
g13530 not P1_R1117_U140 ; P1_R1117_U441
g13531 nand P1_R1117_U441 P1_R1117_U270 ; P1_R1117_U442
g13532 nand P1_R1117_U140 P1_R1117_U67 ; P1_R1117_U443
g13533 nand P1_U3509 P1_R1117_U66 ; P1_R1117_U444
g13534 nand P1_U3069 P1_R1117_U65 ; P1_R1117_U445
g13535 not P1_R1117_U141 ; P1_R1117_U446
g13536 nand P1_R1117_U266 P1_R1117_U446 ; P1_R1117_U447
g13537 nand P1_R1117_U141 P1_R1117_U168 ; P1_R1117_U448
g13538 nand P1_U3506 P1_R1117_U61 ; P1_R1117_U449
g13539 nand P1_U3073 P1_R1117_U59 ; P1_R1117_U450
g13540 nand P1_R1117_U450 P1_R1117_U449 ; P1_R1117_U451
g13541 nand P1_U3503 P1_R1117_U62 ; P1_R1117_U452
g13542 nand P1_U3074 P1_R1117_U49 ; P1_R1117_U453
g13543 nand P1_R1117_U334 P1_R1117_U91 ; P1_R1117_U454
g13544 nand P1_R1117_U169 P1_R1117_U326 ; P1_R1117_U455
g13545 nand P1_U3500 P1_R1117_U63 ; P1_R1117_U456
g13546 nand P1_U3079 P1_R1117_U60 ; P1_R1117_U457
g13547 nand P1_R1117_U335 P1_R1117_U171 ; P1_R1117_U458
g13548 nand P1_R1117_U256 P1_R1117_U170 ; P1_R1117_U459
g13549 nand P1_U3497 P1_R1117_U58 ; P1_R1117_U460
g13550 nand P1_U3080 P1_R1117_U57 ; P1_R1117_U461
g13551 not P1_R1117_U143 ; P1_R1117_U462
g13552 nand P1_R1117_U252 P1_R1117_U462 ; P1_R1117_U463
g13553 nand P1_R1117_U143 P1_R1117_U172 ; P1_R1117_U464
g13554 nand P1_U3494 P1_R1117_U56 ; P1_R1117_U465
g13555 nand P1_U3072 P1_R1117_U55 ; P1_R1117_U466
g13556 not P1_R1117_U144 ; P1_R1117_U467
g13557 nand P1_R1117_U248 P1_R1117_U467 ; P1_R1117_U468
g13558 nand P1_R1117_U144 P1_R1117_U173 ; P1_R1117_U469
g13559 nand P1_U3491 P1_R1117_U52 ; P1_R1117_U470
g13560 nand P1_U3063 P1_R1117_U50 ; P1_R1117_U471
g13561 nand P1_R1117_U471 P1_R1117_U470 ; P1_R1117_U472
g13562 nand P1_U3488 P1_R1117_U53 ; P1_R1117_U473
g13563 nand P1_U3062 P1_R1117_U51 ; P1_R1117_U474
g13564 nand P1_R1117_U345 P1_R1117_U92 ; P1_R1117_U475
g13565 nand P1_R1117_U174 P1_R1117_U337 ; P1_R1117_U476
g13566 and P1_R1375_U8 P1_R1375_U191 ; P1_R1375_U6
g13567 and P1_R1375_U190 P1_R1375_U100 P1_R1375_U189 ; P1_R1375_U7
g13568 and P1_R1375_U195 P1_R1375_U194 ; P1_R1375_U8
g13569 nand P1_R1375_U7 P1_R1375_U192 ; P1_R1375_U9
g13570 not P1_U3088 ; P1_R1375_U10
g13571 not P1_U3087 ; P1_R1375_U11
g13572 not P1_U3121 ; P1_R1375_U12
g13573 not P1_U3120 ; P1_R1375_U13
g13574 not P1_U3152 ; P1_R1375_U14
g13575 not P1_U3117 ; P1_R1375_U15
g13576 not P1_U3149 ; P1_R1375_U16
g13577 not P1_U3148 ; P1_R1375_U17
g13578 not P1_U3116 ; P1_R1375_U18
g13579 not P1_U3115 ; P1_R1375_U19
g13580 not P1_U3147 ; P1_R1375_U20
g13581 not P1_U3146 ; P1_R1375_U21
g13582 not P1_U3114 ; P1_R1375_U22
g13583 not P1_U3113 ; P1_R1375_U23
g13584 not P1_U3145 ; P1_R1375_U24
g13585 not P1_U3144 ; P1_R1375_U25
g13586 not P1_U3112 ; P1_R1375_U26
g13587 not P1_U3111 ; P1_R1375_U27
g13588 not P1_U3143 ; P1_R1375_U28
g13589 not P1_U3142 ; P1_R1375_U29
g13590 not P1_U3110 ; P1_R1375_U30
g13591 not P1_U3109 ; P1_R1375_U31
g13592 not P1_U3141 ; P1_R1375_U32
g13593 not P1_U3140 ; P1_R1375_U33
g13594 not P1_U3108 ; P1_R1375_U34
g13595 not P1_U3107 ; P1_R1375_U35
g13596 not P1_U3139 ; P1_R1375_U36
g13597 not P1_U3138 ; P1_R1375_U37
g13598 not P1_U3106 ; P1_R1375_U38
g13599 not P1_U3105 ; P1_R1375_U39
g13600 not P1_U3137 ; P1_R1375_U40
g13601 not P1_U3136 ; P1_R1375_U41
g13602 not P1_U3104 ; P1_R1375_U42
g13603 not P1_U3103 ; P1_R1375_U43
g13604 not P1_U3135 ; P1_R1375_U44
g13605 not P1_U3134 ; P1_R1375_U45
g13606 not P1_U3102 ; P1_R1375_U46
g13607 not P1_U3101 ; P1_R1375_U47
g13608 not P1_U3133 ; P1_R1375_U48
g13609 not P1_U3132 ; P1_R1375_U49
g13610 not P1_U3100 ; P1_R1375_U50
g13611 not P1_U3099 ; P1_R1375_U51
g13612 not P1_U3131 ; P1_R1375_U52
g13613 not P1_U3130 ; P1_R1375_U53
g13614 not P1_U3098 ; P1_R1375_U54
g13615 not P1_U3097 ; P1_R1375_U55
g13616 not P1_U3129 ; P1_R1375_U56
g13617 not P1_U3128 ; P1_R1375_U57
g13618 not P1_U3096 ; P1_R1375_U58
g13619 not P1_U3095 ; P1_R1375_U59
g13620 not P1_U3127 ; P1_R1375_U60
g13621 not P1_U3126 ; P1_R1375_U61
g13622 not P1_U3094 ; P1_R1375_U62
g13623 not P1_U3093 ; P1_R1375_U63
g13624 not P1_U3125 ; P1_R1375_U64
g13625 not P1_U3124 ; P1_R1375_U65
g13626 not P1_U3092 ; P1_R1375_U66
g13627 not P1_U3091 ; P1_R1375_U67
g13628 not P1_U3123 ; P1_R1375_U68
g13629 not P1_U3089 ; P1_R1375_U69
g13630 and P1_R1375_U107 P1_R1375_U108 ; P1_R1375_U70
g13631 and P1_R1375_U110 P1_R1375_U111 ; P1_R1375_U71
g13632 and P1_R1375_U113 P1_R1375_U114 ; P1_R1375_U72
g13633 and P1_R1375_U116 P1_R1375_U117 ; P1_R1375_U73
g13634 and P1_R1375_U119 P1_R1375_U120 ; P1_R1375_U74
g13635 and P1_R1375_U122 P1_R1375_U123 ; P1_R1375_U75
g13636 and P1_R1375_U125 P1_R1375_U126 ; P1_R1375_U76
g13637 and P1_R1375_U128 P1_R1375_U129 ; P1_R1375_U77
g13638 and P1_R1375_U131 P1_R1375_U132 ; P1_R1375_U78
g13639 and P1_R1375_U134 P1_R1375_U135 ; P1_R1375_U79
g13640 and P1_R1375_U137 P1_R1375_U138 ; P1_R1375_U80
g13641 and P1_R1375_U140 P1_R1375_U141 ; P1_R1375_U81
g13642 and P1_R1375_U143 P1_R1375_U144 ; P1_R1375_U82
g13643 and P1_R1375_U146 P1_R1375_U147 ; P1_R1375_U83
g13644 and P1_R1375_U149 P1_R1375_U150 ; P1_R1375_U84
g13645 and P1_R1375_U152 P1_R1375_U153 ; P1_R1375_U85
g13646 and P1_R1375_U155 P1_R1375_U156 ; P1_R1375_U86
g13647 and P1_R1375_U158 P1_R1375_U159 ; P1_R1375_U87
g13648 and P1_R1375_U161 P1_R1375_U162 ; P1_R1375_U88
g13649 and P1_R1375_U164 P1_R1375_U165 ; P1_R1375_U89
g13650 and P1_R1375_U167 P1_R1375_U168 ; P1_R1375_U90
g13651 and P1_R1375_U170 P1_R1375_U171 ; P1_R1375_U91
g13652 and P1_R1375_U173 P1_R1375_U174 ; P1_R1375_U92
g13653 and P1_R1375_U176 P1_R1375_U177 ; P1_R1375_U93
g13654 and P1_R1375_U179 P1_R1375_U180 ; P1_R1375_U94
g13655 and P1_R1375_U182 P1_R1375_U183 ; P1_R1375_U95
g13656 and P1_R1375_U186 P1_R1375_U101 ; P1_R1375_U96
g13657 and P1_R1375_U186 P1_U3090 ; P1_R1375_U97
g13658 and P1_R1375_U187 P1_R1375_U188 ; P1_R1375_U98
g13659 not P1_U3119 ; P1_R1375_U99
g13660 and P1_R1375_U197 P1_R1375_U196 ; P1_R1375_U100
g13661 not P1_U3122 ; P1_R1375_U101
g13662 nand P1_U3150 P1_U3151 ; P1_R1375_U102
g13663 nand P1_U3118 P1_R1375_U102 ; P1_R1375_U103
g13664 or P1_U3150 P1_U3151 ; P1_R1375_U104
g13665 nand P1_U3117 P1_R1375_U16 ; P1_R1375_U105
g13666 nand P1_R1375_U104 P1_R1375_U105 P1_R1375_U103 ; P1_R1375_U106
g13667 nand P1_U3149 P1_R1375_U15 ; P1_R1375_U107
g13668 nand P1_U3148 P1_R1375_U18 ; P1_R1375_U108
g13669 nand P1_R1375_U70 P1_R1375_U106 ; P1_R1375_U109
g13670 nand P1_U3116 P1_R1375_U17 ; P1_R1375_U110
g13671 nand P1_U3115 P1_R1375_U20 ; P1_R1375_U111
g13672 nand P1_R1375_U71 P1_R1375_U109 ; P1_R1375_U112
g13673 nand P1_U3147 P1_R1375_U19 ; P1_R1375_U113
g13674 nand P1_U3146 P1_R1375_U22 ; P1_R1375_U114
g13675 nand P1_R1375_U72 P1_R1375_U112 ; P1_R1375_U115
g13676 nand P1_U3114 P1_R1375_U21 ; P1_R1375_U116
g13677 nand P1_U3113 P1_R1375_U24 ; P1_R1375_U117
g13678 nand P1_R1375_U73 P1_R1375_U115 ; P1_R1375_U118
g13679 nand P1_U3145 P1_R1375_U23 ; P1_R1375_U119
g13680 nand P1_U3144 P1_R1375_U26 ; P1_R1375_U120
g13681 nand P1_R1375_U74 P1_R1375_U118 ; P1_R1375_U121
g13682 nand P1_U3112 P1_R1375_U25 ; P1_R1375_U122
g13683 nand P1_U3111 P1_R1375_U28 ; P1_R1375_U123
g13684 nand P1_R1375_U75 P1_R1375_U121 ; P1_R1375_U124
g13685 nand P1_U3143 P1_R1375_U27 ; P1_R1375_U125
g13686 nand P1_U3142 P1_R1375_U30 ; P1_R1375_U126
g13687 nand P1_R1375_U76 P1_R1375_U124 ; P1_R1375_U127
g13688 nand P1_U3110 P1_R1375_U29 ; P1_R1375_U128
g13689 nand P1_U3109 P1_R1375_U32 ; P1_R1375_U129
g13690 nand P1_R1375_U77 P1_R1375_U127 ; P1_R1375_U130
g13691 nand P1_U3141 P1_R1375_U31 ; P1_R1375_U131
g13692 nand P1_U3140 P1_R1375_U34 ; P1_R1375_U132
g13693 nand P1_R1375_U78 P1_R1375_U130 ; P1_R1375_U133
g13694 nand P1_U3108 P1_R1375_U33 ; P1_R1375_U134
g13695 nand P1_U3107 P1_R1375_U36 ; P1_R1375_U135
g13696 nand P1_R1375_U79 P1_R1375_U133 ; P1_R1375_U136
g13697 nand P1_U3139 P1_R1375_U35 ; P1_R1375_U137
g13698 nand P1_U3138 P1_R1375_U38 ; P1_R1375_U138
g13699 nand P1_R1375_U80 P1_R1375_U136 ; P1_R1375_U139
g13700 nand P1_U3106 P1_R1375_U37 ; P1_R1375_U140
g13701 nand P1_U3105 P1_R1375_U40 ; P1_R1375_U141
g13702 nand P1_R1375_U81 P1_R1375_U139 ; P1_R1375_U142
g13703 nand P1_U3137 P1_R1375_U39 ; P1_R1375_U143
g13704 nand P1_U3136 P1_R1375_U42 ; P1_R1375_U144
g13705 nand P1_R1375_U82 P1_R1375_U142 ; P1_R1375_U145
g13706 nand P1_U3104 P1_R1375_U41 ; P1_R1375_U146
g13707 nand P1_U3103 P1_R1375_U44 ; P1_R1375_U147
g13708 nand P1_R1375_U83 P1_R1375_U145 ; P1_R1375_U148
g13709 nand P1_U3135 P1_R1375_U43 ; P1_R1375_U149
g13710 nand P1_U3134 P1_R1375_U46 ; P1_R1375_U150
g13711 nand P1_R1375_U84 P1_R1375_U148 ; P1_R1375_U151
g13712 nand P1_U3102 P1_R1375_U45 ; P1_R1375_U152
g13713 nand P1_U3101 P1_R1375_U48 ; P1_R1375_U153
g13714 nand P1_R1375_U85 P1_R1375_U151 ; P1_R1375_U154
g13715 nand P1_U3133 P1_R1375_U47 ; P1_R1375_U155
g13716 nand P1_U3132 P1_R1375_U50 ; P1_R1375_U156
g13717 nand P1_R1375_U86 P1_R1375_U154 ; P1_R1375_U157
g13718 nand P1_U3100 P1_R1375_U49 ; P1_R1375_U158
g13719 nand P1_U3099 P1_R1375_U52 ; P1_R1375_U159
g13720 nand P1_R1375_U87 P1_R1375_U157 ; P1_R1375_U160
g13721 nand P1_U3131 P1_R1375_U51 ; P1_R1375_U161
g13722 nand P1_U3130 P1_R1375_U54 ; P1_R1375_U162
g13723 nand P1_R1375_U88 P1_R1375_U160 ; P1_R1375_U163
g13724 nand P1_U3098 P1_R1375_U53 ; P1_R1375_U164
g13725 nand P1_U3097 P1_R1375_U56 ; P1_R1375_U165
g13726 nand P1_R1375_U89 P1_R1375_U163 ; P1_R1375_U166
g13727 nand P1_U3129 P1_R1375_U55 ; P1_R1375_U167
g13728 nand P1_U3128 P1_R1375_U58 ; P1_R1375_U168
g13729 nand P1_R1375_U90 P1_R1375_U166 ; P1_R1375_U169
g13730 nand P1_U3096 P1_R1375_U57 ; P1_R1375_U170
g13731 nand P1_U3095 P1_R1375_U60 ; P1_R1375_U171
g13732 nand P1_R1375_U91 P1_R1375_U169 ; P1_R1375_U172
g13733 nand P1_U3127 P1_R1375_U59 ; P1_R1375_U173
g13734 nand P1_U3126 P1_R1375_U62 ; P1_R1375_U174
g13735 nand P1_R1375_U92 P1_R1375_U172 ; P1_R1375_U175
g13736 nand P1_U3094 P1_R1375_U61 ; P1_R1375_U176
g13737 nand P1_U3093 P1_R1375_U64 ; P1_R1375_U177
g13738 nand P1_R1375_U93 P1_R1375_U175 ; P1_R1375_U178
g13739 nand P1_U3125 P1_R1375_U63 ; P1_R1375_U179
g13740 nand P1_U3124 P1_R1375_U66 ; P1_R1375_U180
g13741 nand P1_R1375_U94 P1_R1375_U178 ; P1_R1375_U181
g13742 nand P1_U3092 P1_R1375_U65 ; P1_R1375_U182
g13743 nand P1_U3091 P1_R1375_U68 ; P1_R1375_U183
g13744 nand P1_R1375_U95 P1_R1375_U181 ; P1_R1375_U184
g13745 nand P1_R1375_U96 P1_R1375_U184 ; P1_R1375_U185
g13746 nand P1_U3123 P1_R1375_U67 ; P1_R1375_U186
g13747 nand P1_U3090 P1_R1375_U101 ; P1_R1375_U187
g13748 nand P1_U3089 P1_R1375_U12 ; P1_R1375_U188
g13749 nand P1_R1375_U8 P1_R1375_U191 P1_U3121 P1_R1375_U69 ; P1_R1375_U189
g13750 nand P1_R1375_U8 P1_R1375_U10 P1_U3120 ; P1_R1375_U190
g13751 nand P1_U3088 P1_R1375_U13 ; P1_R1375_U191
g13752 nand P1_R1375_U6 P1_R1375_U193 P1_R1375_U98 P1_R1375_U185 ; P1_R1375_U192
g13753 nand P1_R1375_U97 P1_R1375_U184 ; P1_R1375_U193
g13754 nand P1_U3087 P1_R1375_U99 ; P1_R1375_U194
g13755 nand P1_U3119 P1_R1375_U11 ; P1_R1375_U195
g13756 nand P1_U3152 P1_U3087 P1_R1375_U99 ; P1_R1375_U196
g13757 nand P1_R1375_U14 P1_R1375_U11 P1_U3119 ; P1_R1375_U197
g13758 and P1_U3059 P1_R1352_U7 ; P1_R1352_U6
g13759 not P1_U3056 ; P1_R1352_U7
g13760 and P1_R1207_U184 P1_R1207_U201 ; P1_R1207_U6
g13761 and P1_R1207_U203 P1_R1207_U202 ; P1_R1207_U7
g13762 and P1_R1207_U179 P1_R1207_U240 ; P1_R1207_U8
g13763 and P1_R1207_U242 P1_R1207_U241 ; P1_R1207_U9
g13764 and P1_R1207_U259 P1_R1207_U258 ; P1_R1207_U10
g13765 and P1_R1207_U285 P1_R1207_U284 ; P1_R1207_U11
g13766 and P1_R1207_U383 P1_R1207_U382 ; P1_R1207_U12
g13767 nand P1_R1207_U340 P1_R1207_U343 ; P1_R1207_U13
g13768 nand P1_R1207_U329 P1_R1207_U332 ; P1_R1207_U14
g13769 nand P1_R1207_U318 P1_R1207_U321 ; P1_R1207_U15
g13770 nand P1_R1207_U310 P1_R1207_U312 ; P1_R1207_U16
g13771 nand P1_R1207_U156 P1_R1207_U175 P1_R1207_U348 ; P1_R1207_U17
g13772 nand P1_R1207_U236 P1_R1207_U238 ; P1_R1207_U18
g13773 nand P1_R1207_U228 P1_R1207_U231 ; P1_R1207_U19
g13774 nand P1_R1207_U220 P1_R1207_U222 ; P1_R1207_U20
g13775 nand P1_R1207_U25 P1_R1207_U346 ; P1_R1207_U21
g13776 not P1_U3479 ; P1_R1207_U22
g13777 not P1_U3464 ; P1_R1207_U23
g13778 not P1_U3456 ; P1_R1207_U24
g13779 nand P1_U3456 P1_R1207_U93 ; P1_R1207_U25
g13780 not P1_U3078 ; P1_R1207_U26
g13781 not P1_U3467 ; P1_R1207_U27
g13782 not P1_U3068 ; P1_R1207_U28
g13783 nand P1_U3068 P1_R1207_U23 ; P1_R1207_U29
g13784 not P1_U3064 ; P1_R1207_U30
g13785 not P1_U3476 ; P1_R1207_U31
g13786 not P1_U3473 ; P1_R1207_U32
g13787 not P1_U3470 ; P1_R1207_U33
g13788 not P1_U3071 ; P1_R1207_U34
g13789 not P1_U3067 ; P1_R1207_U35
g13790 not P1_U3060 ; P1_R1207_U36
g13791 nand P1_U3060 P1_R1207_U33 ; P1_R1207_U37
g13792 not P1_U3482 ; P1_R1207_U38
g13793 not P1_U3070 ; P1_R1207_U39
g13794 nand P1_U3070 P1_R1207_U22 ; P1_R1207_U40
g13795 not P1_U3084 ; P1_R1207_U41
g13796 not P1_U3485 ; P1_R1207_U42
g13797 not P1_U3083 ; P1_R1207_U43
g13798 nand P1_R1207_U209 P1_R1207_U208 ; P1_R1207_U44
g13799 nand P1_R1207_U37 P1_R1207_U224 ; P1_R1207_U45
g13800 nand P1_R1207_U193 P1_R1207_U192 ; P1_R1207_U46
g13801 not P1_U4019 ; P1_R1207_U47
g13802 not P1_U4023 ; P1_R1207_U48
g13803 not P1_U3503 ; P1_R1207_U49
g13804 not P1_U3491 ; P1_R1207_U50
g13805 not P1_U3488 ; P1_R1207_U51
g13806 not P1_U3063 ; P1_R1207_U52
g13807 not P1_U3062 ; P1_R1207_U53
g13808 nand P1_U3083 P1_R1207_U42 ; P1_R1207_U54
g13809 not P1_U3494 ; P1_R1207_U55
g13810 not P1_U3072 ; P1_R1207_U56
g13811 not P1_U3497 ; P1_R1207_U57
g13812 not P1_U3080 ; P1_R1207_U58
g13813 not P1_U3506 ; P1_R1207_U59
g13814 not P1_U3500 ; P1_R1207_U60
g13815 not P1_U3073 ; P1_R1207_U61
g13816 not P1_U3074 ; P1_R1207_U62
g13817 not P1_U3079 ; P1_R1207_U63
g13818 nand P1_U3079 P1_R1207_U60 ; P1_R1207_U64
g13819 not P1_U3509 ; P1_R1207_U65
g13820 not P1_U3069 ; P1_R1207_U66
g13821 nand P1_R1207_U269 P1_R1207_U268 ; P1_R1207_U67
g13822 not P1_U3082 ; P1_R1207_U68
g13823 not P1_U3514 ; P1_R1207_U69
g13824 not P1_U3081 ; P1_R1207_U70
g13825 not P1_U4025 ; P1_R1207_U71
g13826 not P1_U3076 ; P1_R1207_U72
g13827 not P1_U4022 ; P1_R1207_U73
g13828 not P1_U4024 ; P1_R1207_U74
g13829 not P1_U3066 ; P1_R1207_U75
g13830 not P1_U3061 ; P1_R1207_U76
g13831 not P1_U3075 ; P1_R1207_U77
g13832 nand P1_U3075 P1_R1207_U74 ; P1_R1207_U78
g13833 not P1_U4021 ; P1_R1207_U79
g13834 not P1_U3065 ; P1_R1207_U80
g13835 not P1_U4020 ; P1_R1207_U81
g13836 not P1_U3058 ; P1_R1207_U82
g13837 not P1_U4018 ; P1_R1207_U83
g13838 not P1_U3057 ; P1_R1207_U84
g13839 nand P1_U3057 P1_R1207_U47 ; P1_R1207_U85
g13840 not P1_U3053 ; P1_R1207_U86
g13841 not P1_U4017 ; P1_R1207_U87
g13842 not P1_U3054 ; P1_R1207_U88
g13843 nand P1_R1207_U299 P1_R1207_U298 ; P1_R1207_U89
g13844 nand P1_R1207_U78 P1_R1207_U314 ; P1_R1207_U90
g13845 nand P1_R1207_U64 P1_R1207_U325 ; P1_R1207_U91
g13846 nand P1_R1207_U54 P1_R1207_U336 ; P1_R1207_U92
g13847 not P1_U3077 ; P1_R1207_U93
g13848 nand P1_R1207_U393 P1_R1207_U392 ; P1_R1207_U94
g13849 nand P1_R1207_U407 P1_R1207_U406 ; P1_R1207_U95
g13850 nand P1_R1207_U412 P1_R1207_U411 ; P1_R1207_U96
g13851 nand P1_R1207_U428 P1_R1207_U427 ; P1_R1207_U97
g13852 nand P1_R1207_U433 P1_R1207_U432 ; P1_R1207_U98
g13853 nand P1_R1207_U438 P1_R1207_U437 ; P1_R1207_U99
g13854 nand P1_R1207_U443 P1_R1207_U442 ; P1_R1207_U100
g13855 nand P1_R1207_U448 P1_R1207_U447 ; P1_R1207_U101
g13856 nand P1_R1207_U464 P1_R1207_U463 ; P1_R1207_U102
g13857 nand P1_R1207_U469 P1_R1207_U468 ; P1_R1207_U103
g13858 nand P1_R1207_U352 P1_R1207_U351 ; P1_R1207_U104
g13859 nand P1_R1207_U361 P1_R1207_U360 ; P1_R1207_U105
g13860 nand P1_R1207_U368 P1_R1207_U367 ; P1_R1207_U106
g13861 nand P1_R1207_U372 P1_R1207_U371 ; P1_R1207_U107
g13862 nand P1_R1207_U381 P1_R1207_U380 ; P1_R1207_U108
g13863 nand P1_R1207_U402 P1_R1207_U401 ; P1_R1207_U109
g13864 nand P1_R1207_U419 P1_R1207_U418 ; P1_R1207_U110
g13865 nand P1_R1207_U423 P1_R1207_U422 ; P1_R1207_U111
g13866 nand P1_R1207_U455 P1_R1207_U454 ; P1_R1207_U112
g13867 nand P1_R1207_U459 P1_R1207_U458 ; P1_R1207_U113
g13868 nand P1_R1207_U476 P1_R1207_U475 ; P1_R1207_U114
g13869 and P1_R1207_U195 P1_R1207_U183 ; P1_R1207_U115
g13870 and P1_R1207_U198 P1_R1207_U199 ; P1_R1207_U116
g13871 and P1_R1207_U211 P1_R1207_U185 ; P1_R1207_U117
g13872 and P1_R1207_U214 P1_R1207_U215 ; P1_R1207_U118
g13873 and P1_R1207_U354 P1_R1207_U353 P1_R1207_U40 ; P1_R1207_U119
g13874 and P1_R1207_U357 P1_R1207_U185 ; P1_R1207_U120
g13875 and P1_R1207_U230 P1_R1207_U7 ; P1_R1207_U121
g13876 and P1_R1207_U364 P1_R1207_U184 ; P1_R1207_U122
g13877 and P1_R1207_U374 P1_R1207_U373 P1_R1207_U29 ; P1_R1207_U123
g13878 and P1_R1207_U377 P1_R1207_U183 ; P1_R1207_U124
g13879 and P1_R1207_U217 P1_R1207_U8 ; P1_R1207_U125
g13880 and P1_R1207_U262 P1_R1207_U180 ; P1_R1207_U126
g13881 and P1_R1207_U288 P1_R1207_U181 ; P1_R1207_U127
g13882 and P1_R1207_U304 P1_R1207_U305 ; P1_R1207_U128
g13883 and P1_R1207_U307 P1_R1207_U386 ; P1_R1207_U129
g13884 and P1_R1207_U305 P1_R1207_U304 P1_R1207_U308 ; P1_R1207_U130
g13885 nand P1_R1207_U390 P1_R1207_U389 ; P1_R1207_U131
g13886 and P1_R1207_U395 P1_R1207_U394 P1_R1207_U85 ; P1_R1207_U132
g13887 and P1_R1207_U398 P1_R1207_U182 ; P1_R1207_U133
g13888 nand P1_R1207_U404 P1_R1207_U403 ; P1_R1207_U134
g13889 nand P1_R1207_U409 P1_R1207_U408 ; P1_R1207_U135
g13890 and P1_R1207_U415 P1_R1207_U181 ; P1_R1207_U136
g13891 nand P1_R1207_U425 P1_R1207_U424 ; P1_R1207_U137
g13892 nand P1_R1207_U430 P1_R1207_U429 ; P1_R1207_U138
g13893 nand P1_R1207_U435 P1_R1207_U434 ; P1_R1207_U139
g13894 nand P1_R1207_U440 P1_R1207_U439 ; P1_R1207_U140
g13895 nand P1_R1207_U445 P1_R1207_U444 ; P1_R1207_U141
g13896 and P1_R1207_U451 P1_R1207_U180 ; P1_R1207_U142
g13897 nand P1_R1207_U461 P1_R1207_U460 ; P1_R1207_U143
g13898 nand P1_R1207_U466 P1_R1207_U465 ; P1_R1207_U144
g13899 and P1_R1207_U342 P1_R1207_U9 ; P1_R1207_U145
g13900 and P1_R1207_U472 P1_R1207_U179 ; P1_R1207_U146
g13901 and P1_R1207_U350 P1_R1207_U349 ; P1_R1207_U147
g13902 nand P1_R1207_U118 P1_R1207_U212 ; P1_R1207_U148
g13903 and P1_R1207_U359 P1_R1207_U358 ; P1_R1207_U149
g13904 and P1_R1207_U366 P1_R1207_U365 ; P1_R1207_U150
g13905 and P1_R1207_U370 P1_R1207_U369 ; P1_R1207_U151
g13906 nand P1_R1207_U116 P1_R1207_U196 ; P1_R1207_U152
g13907 and P1_R1207_U379 P1_R1207_U378 ; P1_R1207_U153
g13908 not P1_U4028 ; P1_R1207_U154
g13909 not P1_U3055 ; P1_R1207_U155
g13910 and P1_R1207_U388 P1_R1207_U387 ; P1_R1207_U156
g13911 nand P1_R1207_U128 P1_R1207_U302 ; P1_R1207_U157
g13912 and P1_R1207_U400 P1_R1207_U399 ; P1_R1207_U158
g13913 nand P1_R1207_U295 P1_R1207_U294 ; P1_R1207_U159
g13914 nand P1_R1207_U291 P1_R1207_U290 ; P1_R1207_U160
g13915 and P1_R1207_U417 P1_R1207_U416 ; P1_R1207_U161
g13916 and P1_R1207_U421 P1_R1207_U420 ; P1_R1207_U162
g13917 nand P1_R1207_U281 P1_R1207_U280 ; P1_R1207_U163
g13918 nand P1_R1207_U277 P1_R1207_U276 ; P1_R1207_U164
g13919 not P1_U3461 ; P1_R1207_U165
g13920 nand P1_R1207_U273 P1_R1207_U272 ; P1_R1207_U166
g13921 not P1_U3512 ; P1_R1207_U167
g13922 nand P1_R1207_U265 P1_R1207_U264 ; P1_R1207_U168
g13923 and P1_R1207_U453 P1_R1207_U452 ; P1_R1207_U169
g13924 and P1_R1207_U457 P1_R1207_U456 ; P1_R1207_U170
g13925 nand P1_R1207_U255 P1_R1207_U254 ; P1_R1207_U171
g13926 nand P1_R1207_U251 P1_R1207_U250 ; P1_R1207_U172
g13927 nand P1_R1207_U247 P1_R1207_U246 ; P1_R1207_U173
g13928 and P1_R1207_U474 P1_R1207_U473 ; P1_R1207_U174
g13929 nand P1_R1207_U129 P1_R1207_U157 ; P1_R1207_U175
g13930 not P1_R1207_U85 ; P1_R1207_U176
g13931 not P1_R1207_U29 ; P1_R1207_U177
g13932 not P1_R1207_U40 ; P1_R1207_U178
g13933 nand P1_U3488 P1_R1207_U53 ; P1_R1207_U179
g13934 nand P1_U3503 P1_R1207_U62 ; P1_R1207_U180
g13935 nand P1_U4023 P1_R1207_U76 ; P1_R1207_U181
g13936 nand P1_U4019 P1_R1207_U84 ; P1_R1207_U182
g13937 nand P1_U3464 P1_R1207_U28 ; P1_R1207_U183
g13938 nand P1_U3473 P1_R1207_U35 ; P1_R1207_U184
g13939 nand P1_U3479 P1_R1207_U39 ; P1_R1207_U185
g13940 not P1_R1207_U64 ; P1_R1207_U186
g13941 not P1_R1207_U78 ; P1_R1207_U187
g13942 not P1_R1207_U37 ; P1_R1207_U188
g13943 not P1_R1207_U54 ; P1_R1207_U189
g13944 not P1_R1207_U25 ; P1_R1207_U190
g13945 nand P1_R1207_U190 P1_R1207_U26 ; P1_R1207_U191
g13946 nand P1_R1207_U191 P1_R1207_U165 ; P1_R1207_U192
g13947 nand P1_U3078 P1_R1207_U25 ; P1_R1207_U193
g13948 not P1_R1207_U46 ; P1_R1207_U194
g13949 nand P1_U3467 P1_R1207_U30 ; P1_R1207_U195
g13950 nand P1_R1207_U115 P1_R1207_U46 ; P1_R1207_U196
g13951 nand P1_R1207_U30 P1_R1207_U29 ; P1_R1207_U197
g13952 nand P1_R1207_U197 P1_R1207_U27 ; P1_R1207_U198
g13953 nand P1_U3064 P1_R1207_U177 ; P1_R1207_U199
g13954 not P1_R1207_U152 ; P1_R1207_U200
g13955 nand P1_U3476 P1_R1207_U34 ; P1_R1207_U201
g13956 nand P1_U3071 P1_R1207_U31 ; P1_R1207_U202
g13957 nand P1_U3067 P1_R1207_U32 ; P1_R1207_U203
g13958 nand P1_R1207_U188 P1_R1207_U6 ; P1_R1207_U204
g13959 nand P1_R1207_U7 P1_R1207_U204 ; P1_R1207_U205
g13960 nand P1_U3470 P1_R1207_U36 ; P1_R1207_U206
g13961 nand P1_U3476 P1_R1207_U34 ; P1_R1207_U207
g13962 nand P1_R1207_U206 P1_R1207_U152 P1_R1207_U6 ; P1_R1207_U208
g13963 nand P1_R1207_U207 P1_R1207_U205 ; P1_R1207_U209
g13964 not P1_R1207_U44 ; P1_R1207_U210
g13965 nand P1_U3482 P1_R1207_U41 ; P1_R1207_U211
g13966 nand P1_R1207_U117 P1_R1207_U44 ; P1_R1207_U212
g13967 nand P1_R1207_U41 P1_R1207_U40 ; P1_R1207_U213
g13968 nand P1_R1207_U213 P1_R1207_U38 ; P1_R1207_U214
g13969 nand P1_U3084 P1_R1207_U178 ; P1_R1207_U215
g13970 not P1_R1207_U148 ; P1_R1207_U216
g13971 nand P1_U3485 P1_R1207_U43 ; P1_R1207_U217
g13972 nand P1_R1207_U217 P1_R1207_U54 ; P1_R1207_U218
g13973 nand P1_R1207_U210 P1_R1207_U40 ; P1_R1207_U219
g13974 nand P1_R1207_U120 P1_R1207_U219 ; P1_R1207_U220
g13975 nand P1_R1207_U44 P1_R1207_U185 ; P1_R1207_U221
g13976 nand P1_R1207_U119 P1_R1207_U221 ; P1_R1207_U222
g13977 nand P1_R1207_U40 P1_R1207_U185 ; P1_R1207_U223
g13978 nand P1_R1207_U206 P1_R1207_U152 ; P1_R1207_U224
g13979 not P1_R1207_U45 ; P1_R1207_U225
g13980 nand P1_U3067 P1_R1207_U32 ; P1_R1207_U226
g13981 nand P1_R1207_U225 P1_R1207_U226 ; P1_R1207_U227
g13982 nand P1_R1207_U122 P1_R1207_U227 ; P1_R1207_U228
g13983 nand P1_R1207_U45 P1_R1207_U184 ; P1_R1207_U229
g13984 nand P1_U3476 P1_R1207_U34 ; P1_R1207_U230
g13985 nand P1_R1207_U121 P1_R1207_U229 ; P1_R1207_U231
g13986 nand P1_U3067 P1_R1207_U32 ; P1_R1207_U232
g13987 nand P1_R1207_U184 P1_R1207_U232 ; P1_R1207_U233
g13988 nand P1_R1207_U206 P1_R1207_U37 ; P1_R1207_U234
g13989 nand P1_R1207_U194 P1_R1207_U29 ; P1_R1207_U235
g13990 nand P1_R1207_U124 P1_R1207_U235 ; P1_R1207_U236
g13991 nand P1_R1207_U46 P1_R1207_U183 ; P1_R1207_U237
g13992 nand P1_R1207_U123 P1_R1207_U237 ; P1_R1207_U238
g13993 nand P1_R1207_U29 P1_R1207_U183 ; P1_R1207_U239
g13994 nand P1_U3491 P1_R1207_U52 ; P1_R1207_U240
g13995 nand P1_U3063 P1_R1207_U50 ; P1_R1207_U241
g13996 nand P1_U3062 P1_R1207_U51 ; P1_R1207_U242
g13997 nand P1_R1207_U189 P1_R1207_U8 ; P1_R1207_U243
g13998 nand P1_R1207_U9 P1_R1207_U243 ; P1_R1207_U244
g13999 nand P1_U3491 P1_R1207_U52 ; P1_R1207_U245
g14000 nand P1_R1207_U125 P1_R1207_U148 ; P1_R1207_U246
g14001 nand P1_R1207_U245 P1_R1207_U244 ; P1_R1207_U247
g14002 not P1_R1207_U173 ; P1_R1207_U248
g14003 nand P1_U3494 P1_R1207_U56 ; P1_R1207_U249
g14004 nand P1_R1207_U249 P1_R1207_U173 ; P1_R1207_U250
g14005 nand P1_U3072 P1_R1207_U55 ; P1_R1207_U251
g14006 not P1_R1207_U172 ; P1_R1207_U252
g14007 nand P1_U3497 P1_R1207_U58 ; P1_R1207_U253
g14008 nand P1_R1207_U253 P1_R1207_U172 ; P1_R1207_U254
g14009 nand P1_U3080 P1_R1207_U57 ; P1_R1207_U255
g14010 not P1_R1207_U171 ; P1_R1207_U256
g14011 nand P1_U3506 P1_R1207_U61 ; P1_R1207_U257
g14012 nand P1_U3073 P1_R1207_U59 ; P1_R1207_U258
g14013 nand P1_U3074 P1_R1207_U49 ; P1_R1207_U259
g14014 nand P1_R1207_U186 P1_R1207_U180 ; P1_R1207_U260
g14015 nand P1_R1207_U10 P1_R1207_U260 ; P1_R1207_U261
g14016 nand P1_U3500 P1_R1207_U63 ; P1_R1207_U262
g14017 nand P1_U3506 P1_R1207_U61 ; P1_R1207_U263
g14018 nand P1_R1207_U171 P1_R1207_U126 P1_R1207_U257 ; P1_R1207_U264
g14019 nand P1_R1207_U263 P1_R1207_U261 ; P1_R1207_U265
g14020 not P1_R1207_U168 ; P1_R1207_U266
g14021 nand P1_U3509 P1_R1207_U66 ; P1_R1207_U267
g14022 nand P1_R1207_U267 P1_R1207_U168 ; P1_R1207_U268
g14023 nand P1_U3069 P1_R1207_U65 ; P1_R1207_U269
g14024 not P1_R1207_U67 ; P1_R1207_U270
g14025 nand P1_R1207_U270 P1_R1207_U68 ; P1_R1207_U271
g14026 nand P1_R1207_U271 P1_R1207_U167 ; P1_R1207_U272
g14027 nand P1_U3082 P1_R1207_U67 ; P1_R1207_U273
g14028 not P1_R1207_U166 ; P1_R1207_U274
g14029 nand P1_U3514 P1_R1207_U70 ; P1_R1207_U275
g14030 nand P1_R1207_U275 P1_R1207_U166 ; P1_R1207_U276
g14031 nand P1_U3081 P1_R1207_U69 ; P1_R1207_U277
g14032 not P1_R1207_U164 ; P1_R1207_U278
g14033 nand P1_U4025 P1_R1207_U72 ; P1_R1207_U279
g14034 nand P1_R1207_U279 P1_R1207_U164 ; P1_R1207_U280
g14035 nand P1_U3076 P1_R1207_U71 ; P1_R1207_U281
g14036 not P1_R1207_U163 ; P1_R1207_U282
g14037 nand P1_U4022 P1_R1207_U75 ; P1_R1207_U283
g14038 nand P1_U3066 P1_R1207_U73 ; P1_R1207_U284
g14039 nand P1_U3061 P1_R1207_U48 ; P1_R1207_U285
g14040 nand P1_R1207_U187 P1_R1207_U181 ; P1_R1207_U286
g14041 nand P1_R1207_U11 P1_R1207_U286 ; P1_R1207_U287
g14042 nand P1_U4024 P1_R1207_U77 ; P1_R1207_U288
g14043 nand P1_U4022 P1_R1207_U75 ; P1_R1207_U289
g14044 nand P1_R1207_U163 P1_R1207_U127 P1_R1207_U283 ; P1_R1207_U290
g14045 nand P1_R1207_U289 P1_R1207_U287 ; P1_R1207_U291
g14046 not P1_R1207_U160 ; P1_R1207_U292
g14047 nand P1_U4021 P1_R1207_U80 ; P1_R1207_U293
g14048 nand P1_R1207_U293 P1_R1207_U160 ; P1_R1207_U294
g14049 nand P1_U3065 P1_R1207_U79 ; P1_R1207_U295
g14050 not P1_R1207_U159 ; P1_R1207_U296
g14051 nand P1_U4020 P1_R1207_U82 ; P1_R1207_U297
g14052 nand P1_R1207_U297 P1_R1207_U159 ; P1_R1207_U298
g14053 nand P1_U3058 P1_R1207_U81 ; P1_R1207_U299
g14054 not P1_R1207_U89 ; P1_R1207_U300
g14055 nand P1_U4018 P1_R1207_U86 ; P1_R1207_U301
g14056 nand P1_R1207_U89 P1_R1207_U182 P1_R1207_U301 ; P1_R1207_U302
g14057 nand P1_R1207_U86 P1_R1207_U85 ; P1_R1207_U303
g14058 nand P1_R1207_U303 P1_R1207_U83 ; P1_R1207_U304
g14059 nand P1_U3053 P1_R1207_U176 ; P1_R1207_U305
g14060 not P1_R1207_U157 ; P1_R1207_U306
g14061 nand P1_U4017 P1_R1207_U88 ; P1_R1207_U307
g14062 nand P1_U3054 P1_R1207_U87 ; P1_R1207_U308
g14063 nand P1_R1207_U300 P1_R1207_U85 ; P1_R1207_U309
g14064 nand P1_R1207_U133 P1_R1207_U309 ; P1_R1207_U310
g14065 nand P1_R1207_U89 P1_R1207_U182 ; P1_R1207_U311
g14066 nand P1_R1207_U132 P1_R1207_U311 ; P1_R1207_U312
g14067 nand P1_R1207_U85 P1_R1207_U182 ; P1_R1207_U313
g14068 nand P1_R1207_U288 P1_R1207_U163 ; P1_R1207_U314
g14069 not P1_R1207_U90 ; P1_R1207_U315
g14070 nand P1_U3061 P1_R1207_U48 ; P1_R1207_U316
g14071 nand P1_R1207_U315 P1_R1207_U316 ; P1_R1207_U317
g14072 nand P1_R1207_U136 P1_R1207_U317 ; P1_R1207_U318
g14073 nand P1_R1207_U90 P1_R1207_U181 ; P1_R1207_U319
g14074 nand P1_U4022 P1_R1207_U75 ; P1_R1207_U320
g14075 nand P1_R1207_U320 P1_R1207_U319 P1_R1207_U11 ; P1_R1207_U321
g14076 nand P1_U3061 P1_R1207_U48 ; P1_R1207_U322
g14077 nand P1_R1207_U181 P1_R1207_U322 ; P1_R1207_U323
g14078 nand P1_R1207_U288 P1_R1207_U78 ; P1_R1207_U324
g14079 nand P1_R1207_U262 P1_R1207_U171 ; P1_R1207_U325
g14080 not P1_R1207_U91 ; P1_R1207_U326
g14081 nand P1_U3074 P1_R1207_U49 ; P1_R1207_U327
g14082 nand P1_R1207_U326 P1_R1207_U327 ; P1_R1207_U328
g14083 nand P1_R1207_U142 P1_R1207_U328 ; P1_R1207_U329
g14084 nand P1_R1207_U91 P1_R1207_U180 ; P1_R1207_U330
g14085 nand P1_U3506 P1_R1207_U61 ; P1_R1207_U331
g14086 nand P1_R1207_U331 P1_R1207_U330 P1_R1207_U10 ; P1_R1207_U332
g14087 nand P1_U3074 P1_R1207_U49 ; P1_R1207_U333
g14088 nand P1_R1207_U180 P1_R1207_U333 ; P1_R1207_U334
g14089 nand P1_R1207_U262 P1_R1207_U64 ; P1_R1207_U335
g14090 nand P1_R1207_U217 P1_R1207_U148 ; P1_R1207_U336
g14091 not P1_R1207_U92 ; P1_R1207_U337
g14092 nand P1_U3062 P1_R1207_U51 ; P1_R1207_U338
g14093 nand P1_R1207_U337 P1_R1207_U338 ; P1_R1207_U339
g14094 nand P1_R1207_U146 P1_R1207_U339 ; P1_R1207_U340
g14095 nand P1_R1207_U92 P1_R1207_U179 ; P1_R1207_U341
g14096 nand P1_U3491 P1_R1207_U52 ; P1_R1207_U342
g14097 nand P1_R1207_U145 P1_R1207_U341 ; P1_R1207_U343
g14098 nand P1_U3062 P1_R1207_U51 ; P1_R1207_U344
g14099 nand P1_R1207_U179 P1_R1207_U344 ; P1_R1207_U345
g14100 nand P1_U3077 P1_R1207_U24 ; P1_R1207_U346
g14101 nand P1_R1207_U89 P1_R1207_U182 P1_R1207_U301 ; P1_R1207_U347
g14102 nand P1_R1207_U12 P1_R1207_U347 P1_R1207_U130 ; P1_R1207_U348
g14103 nand P1_U3485 P1_R1207_U43 ; P1_R1207_U349
g14104 nand P1_U3083 P1_R1207_U42 ; P1_R1207_U350
g14105 nand P1_R1207_U218 P1_R1207_U148 ; P1_R1207_U351
g14106 nand P1_R1207_U216 P1_R1207_U147 ; P1_R1207_U352
g14107 nand P1_U3482 P1_R1207_U41 ; P1_R1207_U353
g14108 nand P1_U3084 P1_R1207_U38 ; P1_R1207_U354
g14109 nand P1_U3482 P1_R1207_U41 ; P1_R1207_U355
g14110 nand P1_U3084 P1_R1207_U38 ; P1_R1207_U356
g14111 nand P1_R1207_U356 P1_R1207_U355 ; P1_R1207_U357
g14112 nand P1_U3479 P1_R1207_U39 ; P1_R1207_U358
g14113 nand P1_U3070 P1_R1207_U22 ; P1_R1207_U359
g14114 nand P1_R1207_U223 P1_R1207_U44 ; P1_R1207_U360
g14115 nand P1_R1207_U149 P1_R1207_U210 ; P1_R1207_U361
g14116 nand P1_U3476 P1_R1207_U34 ; P1_R1207_U362
g14117 nand P1_U3071 P1_R1207_U31 ; P1_R1207_U363
g14118 nand P1_R1207_U363 P1_R1207_U362 ; P1_R1207_U364
g14119 nand P1_U3473 P1_R1207_U35 ; P1_R1207_U365
g14120 nand P1_U3067 P1_R1207_U32 ; P1_R1207_U366
g14121 nand P1_R1207_U233 P1_R1207_U45 ; P1_R1207_U367
g14122 nand P1_R1207_U150 P1_R1207_U225 ; P1_R1207_U368
g14123 nand P1_U3470 P1_R1207_U36 ; P1_R1207_U369
g14124 nand P1_U3060 P1_R1207_U33 ; P1_R1207_U370
g14125 nand P1_R1207_U234 P1_R1207_U152 ; P1_R1207_U371
g14126 nand P1_R1207_U200 P1_R1207_U151 ; P1_R1207_U372
g14127 nand P1_U3467 P1_R1207_U30 ; P1_R1207_U373
g14128 nand P1_U3064 P1_R1207_U27 ; P1_R1207_U374
g14129 nand P1_U3467 P1_R1207_U30 ; P1_R1207_U375
g14130 nand P1_U3064 P1_R1207_U27 ; P1_R1207_U376
g14131 nand P1_R1207_U376 P1_R1207_U375 ; P1_R1207_U377
g14132 nand P1_U3464 P1_R1207_U28 ; P1_R1207_U378
g14133 nand P1_U3068 P1_R1207_U23 ; P1_R1207_U379
g14134 nand P1_R1207_U239 P1_R1207_U46 ; P1_R1207_U380
g14135 nand P1_R1207_U153 P1_R1207_U194 ; P1_R1207_U381
g14136 nand P1_U4028 P1_R1207_U155 ; P1_R1207_U382
g14137 nand P1_U3055 P1_R1207_U154 ; P1_R1207_U383
g14138 nand P1_U4028 P1_R1207_U155 ; P1_R1207_U384
g14139 nand P1_U3055 P1_R1207_U154 ; P1_R1207_U385
g14140 nand P1_R1207_U385 P1_R1207_U384 ; P1_R1207_U386
g14141 nand P1_U3054 P1_R1207_U386 P1_R1207_U87 ; P1_R1207_U387
g14142 nand P1_R1207_U12 P1_R1207_U88 P1_U4017 ; P1_R1207_U388
g14143 nand P1_U4017 P1_R1207_U88 ; P1_R1207_U389
g14144 nand P1_U3054 P1_R1207_U87 ; P1_R1207_U390
g14145 not P1_R1207_U131 ; P1_R1207_U391
g14146 nand P1_R1207_U306 P1_R1207_U391 ; P1_R1207_U392
g14147 nand P1_R1207_U131 P1_R1207_U157 ; P1_R1207_U393
g14148 nand P1_U4018 P1_R1207_U86 ; P1_R1207_U394
g14149 nand P1_U3053 P1_R1207_U83 ; P1_R1207_U395
g14150 nand P1_U4018 P1_R1207_U86 ; P1_R1207_U396
g14151 nand P1_U3053 P1_R1207_U83 ; P1_R1207_U397
g14152 nand P1_R1207_U397 P1_R1207_U396 ; P1_R1207_U398
g14153 nand P1_U4019 P1_R1207_U84 ; P1_R1207_U399
g14154 nand P1_U3057 P1_R1207_U47 ; P1_R1207_U400
g14155 nand P1_R1207_U313 P1_R1207_U89 ; P1_R1207_U401
g14156 nand P1_R1207_U158 P1_R1207_U300 ; P1_R1207_U402
g14157 nand P1_U4020 P1_R1207_U82 ; P1_R1207_U403
g14158 nand P1_U3058 P1_R1207_U81 ; P1_R1207_U404
g14159 not P1_R1207_U134 ; P1_R1207_U405
g14160 nand P1_R1207_U296 P1_R1207_U405 ; P1_R1207_U406
g14161 nand P1_R1207_U134 P1_R1207_U159 ; P1_R1207_U407
g14162 nand P1_U4021 P1_R1207_U80 ; P1_R1207_U408
g14163 nand P1_U3065 P1_R1207_U79 ; P1_R1207_U409
g14164 not P1_R1207_U135 ; P1_R1207_U410
g14165 nand P1_R1207_U292 P1_R1207_U410 ; P1_R1207_U411
g14166 nand P1_R1207_U135 P1_R1207_U160 ; P1_R1207_U412
g14167 nand P1_U4022 P1_R1207_U75 ; P1_R1207_U413
g14168 nand P1_U3066 P1_R1207_U73 ; P1_R1207_U414
g14169 nand P1_R1207_U414 P1_R1207_U413 ; P1_R1207_U415
g14170 nand P1_U4023 P1_R1207_U76 ; P1_R1207_U416
g14171 nand P1_U3061 P1_R1207_U48 ; P1_R1207_U417
g14172 nand P1_R1207_U323 P1_R1207_U90 ; P1_R1207_U418
g14173 nand P1_R1207_U161 P1_R1207_U315 ; P1_R1207_U419
g14174 nand P1_U4024 P1_R1207_U77 ; P1_R1207_U420
g14175 nand P1_U3075 P1_R1207_U74 ; P1_R1207_U421
g14176 nand P1_R1207_U324 P1_R1207_U163 ; P1_R1207_U422
g14177 nand P1_R1207_U282 P1_R1207_U162 ; P1_R1207_U423
g14178 nand P1_U4025 P1_R1207_U72 ; P1_R1207_U424
g14179 nand P1_U3076 P1_R1207_U71 ; P1_R1207_U425
g14180 not P1_R1207_U137 ; P1_R1207_U426
g14181 nand P1_R1207_U278 P1_R1207_U426 ; P1_R1207_U427
g14182 nand P1_R1207_U137 P1_R1207_U164 ; P1_R1207_U428
g14183 nand P1_U3461 P1_R1207_U26 ; P1_R1207_U429
g14184 nand P1_U3078 P1_R1207_U165 ; P1_R1207_U430
g14185 not P1_R1207_U138 ; P1_R1207_U431
g14186 nand P1_R1207_U431 P1_R1207_U190 ; P1_R1207_U432
g14187 nand P1_R1207_U138 P1_R1207_U25 ; P1_R1207_U433
g14188 nand P1_U3514 P1_R1207_U70 ; P1_R1207_U434
g14189 nand P1_U3081 P1_R1207_U69 ; P1_R1207_U435
g14190 not P1_R1207_U139 ; P1_R1207_U436
g14191 nand P1_R1207_U274 P1_R1207_U436 ; P1_R1207_U437
g14192 nand P1_R1207_U139 P1_R1207_U166 ; P1_R1207_U438
g14193 nand P1_U3512 P1_R1207_U68 ; P1_R1207_U439
g14194 nand P1_U3082 P1_R1207_U167 ; P1_R1207_U440
g14195 not P1_R1207_U140 ; P1_R1207_U441
g14196 nand P1_R1207_U441 P1_R1207_U270 ; P1_R1207_U442
g14197 nand P1_R1207_U140 P1_R1207_U67 ; P1_R1207_U443
g14198 nand P1_U3509 P1_R1207_U66 ; P1_R1207_U444
g14199 nand P1_U3069 P1_R1207_U65 ; P1_R1207_U445
g14200 not P1_R1207_U141 ; P1_R1207_U446
g14201 nand P1_R1207_U266 P1_R1207_U446 ; P1_R1207_U447
g14202 nand P1_R1207_U141 P1_R1207_U168 ; P1_R1207_U448
g14203 nand P1_U3506 P1_R1207_U61 ; P1_R1207_U449
g14204 nand P1_U3073 P1_R1207_U59 ; P1_R1207_U450
g14205 nand P1_R1207_U450 P1_R1207_U449 ; P1_R1207_U451
g14206 nand P1_U3503 P1_R1207_U62 ; P1_R1207_U452
g14207 nand P1_U3074 P1_R1207_U49 ; P1_R1207_U453
g14208 nand P1_R1207_U334 P1_R1207_U91 ; P1_R1207_U454
g14209 nand P1_R1207_U169 P1_R1207_U326 ; P1_R1207_U455
g14210 nand P1_U3500 P1_R1207_U63 ; P1_R1207_U456
g14211 nand P1_U3079 P1_R1207_U60 ; P1_R1207_U457
g14212 nand P1_R1207_U335 P1_R1207_U171 ; P1_R1207_U458
g14213 nand P1_R1207_U256 P1_R1207_U170 ; P1_R1207_U459
g14214 nand P1_U3497 P1_R1207_U58 ; P1_R1207_U460
g14215 nand P1_U3080 P1_R1207_U57 ; P1_R1207_U461
g14216 not P1_R1207_U143 ; P1_R1207_U462
g14217 nand P1_R1207_U252 P1_R1207_U462 ; P1_R1207_U463
g14218 nand P1_R1207_U143 P1_R1207_U172 ; P1_R1207_U464
g14219 nand P1_U3494 P1_R1207_U56 ; P1_R1207_U465
g14220 nand P1_U3072 P1_R1207_U55 ; P1_R1207_U466
g14221 not P1_R1207_U144 ; P1_R1207_U467
g14222 nand P1_R1207_U248 P1_R1207_U467 ; P1_R1207_U468
g14223 nand P1_R1207_U144 P1_R1207_U173 ; P1_R1207_U469
g14224 nand P1_U3491 P1_R1207_U52 ; P1_R1207_U470
g14225 nand P1_U3063 P1_R1207_U50 ; P1_R1207_U471
g14226 nand P1_R1207_U471 P1_R1207_U470 ; P1_R1207_U472
g14227 nand P1_U3488 P1_R1207_U53 ; P1_R1207_U473
g14228 nand P1_U3062 P1_R1207_U51 ; P1_R1207_U474
g14229 nand P1_R1207_U345 P1_R1207_U92 ; P1_R1207_U475
g14230 nand P1_R1207_U174 P1_R1207_U337 ; P1_R1207_U476
g14231 and P1_R1165_U202 P1_R1165_U201 ; P1_R1165_U4
g14232 and P1_R1165_U217 P1_R1165_U216 ; P1_R1165_U5
g14233 and P1_R1165_U251 P1_R1165_U250 ; P1_R1165_U6
g14234 and P1_R1165_U269 P1_R1165_U268 ; P1_R1165_U7
g14235 and P1_R1165_U281 P1_R1165_U280 ; P1_R1165_U8
g14236 and P1_R1165_U339 P1_R1165_U336 ; P1_R1165_U9
g14237 and P1_R1165_U330 P1_R1165_U327 ; P1_R1165_U10
g14238 and P1_R1165_U323 P1_R1165_U320 ; P1_R1165_U11
g14239 and P1_R1165_U314 P1_R1165_U311 ; P1_R1165_U12
g14240 and P1_R1165_U240 P1_R1165_U237 ; P1_R1165_U13
g14241 and P1_R1165_U233 P1_R1165_U230 ; P1_R1165_U14
g14242 not P1_U3211 ; P1_R1165_U15
g14243 not P1_U3175 ; P1_R1165_U16
g14244 nand P1_U3175 P1_R1165_U59 ; P1_R1165_U17
g14245 not P1_U3174 ; P1_R1165_U18
g14246 not P1_U3179 ; P1_R1165_U19
g14247 nand P1_U3179 P1_R1165_U61 ; P1_R1165_U20
g14248 not P1_U3178 ; P1_R1165_U21
g14249 not P1_U3181 ; P1_R1165_U22
g14250 not P1_U3180 ; P1_R1165_U23
g14251 nand P1_R1165_U110 P1_R1165_U206 ; P1_R1165_U24
g14252 not P1_U3177 ; P1_R1165_U25
g14253 not P1_U3176 ; P1_R1165_U26
g14254 not P1_U3173 ; P1_R1165_U27
g14255 not P1_U3172 ; P1_R1165_U28
g14256 nand P1_R1165_U226 P1_R1165_U225 ; P1_R1165_U29
g14257 nand P1_R1165_U214 P1_R1165_U213 ; P1_R1165_U30
g14258 nand P1_R1165_U199 P1_R1165_U198 ; P1_R1165_U31
g14259 not P1_U3154 ; P1_R1165_U32
g14260 not P1_U3155 ; P1_R1165_U33
g14261 not P1_U3156 ; P1_R1165_U34
g14262 not P1_U3157 ; P1_R1165_U35
g14263 not P1_U3160 ; P1_R1165_U36
g14264 not P1_U3165 ; P1_R1165_U37
g14265 nand P1_U3165 P1_R1165_U73 ; P1_R1165_U38
g14266 not P1_U3164 ; P1_R1165_U39
g14267 not P1_U3171 ; P1_R1165_U40
g14268 not P1_U3169 ; P1_R1165_U41
g14269 not P1_U3170 ; P1_R1165_U42
g14270 nand P1_U3170 P1_R1165_U76 ; P1_R1165_U43
g14271 not P1_U3168 ; P1_R1165_U44
g14272 not P1_U3167 ; P1_R1165_U45
g14273 not P1_U3166 ; P1_R1165_U46
g14274 not P1_U3163 ; P1_R1165_U47
g14275 not P1_U3162 ; P1_R1165_U48
g14276 nand P1_U3162 P1_R1165_U82 ; P1_R1165_U49
g14277 not P1_U3161 ; P1_R1165_U50
g14278 not P1_U3159 ; P1_R1165_U51
g14279 not P1_U3158 ; P1_R1165_U52
g14280 nand P1_U3155 P1_R1165_U70 ; P1_R1165_U53
g14281 nand P1_R1165_U192 P1_R1165_U307 ; P1_R1165_U54
g14282 nand P1_R1165_U49 P1_R1165_U316 ; P1_R1165_U55
g14283 nand P1_R1165_U266 P1_R1165_U265 ; P1_R1165_U56
g14284 nand P1_R1165_U43 P1_R1165_U332 ; P1_R1165_U57
g14285 nand P1_R1165_U359 P1_R1165_U358 ; P1_R1165_U58
g14286 nand P1_R1165_U388 P1_R1165_U387 ; P1_R1165_U59
g14287 nand P1_R1165_U385 P1_R1165_U384 ; P1_R1165_U60
g14288 nand P1_R1165_U376 P1_R1165_U375 ; P1_R1165_U61
g14289 nand P1_R1165_U373 P1_R1165_U372 ; P1_R1165_U62
g14290 nand P1_R1165_U367 P1_R1165_U366 ; P1_R1165_U63
g14291 nand P1_R1165_U370 P1_R1165_U369 ; P1_R1165_U64
g14292 nand P1_R1165_U379 P1_R1165_U378 ; P1_R1165_U65
g14293 nand P1_R1165_U382 P1_R1165_U381 ; P1_R1165_U66
g14294 nand P1_R1165_U391 P1_R1165_U390 ; P1_R1165_U67
g14295 nand P1_R1165_U431 P1_R1165_U430 ; P1_R1165_U68
g14296 nand P1_R1165_U434 P1_R1165_U433 ; P1_R1165_U69
g14297 nand P1_R1165_U437 P1_R1165_U436 ; P1_R1165_U70
g14298 nand P1_R1165_U440 P1_R1165_U439 ; P1_R1165_U71
g14299 nand P1_R1165_U443 P1_R1165_U442 ; P1_R1165_U72
g14300 nand P1_R1165_U473 P1_R1165_U472 ; P1_R1165_U73
g14301 nand P1_R1165_U470 P1_R1165_U469 ; P1_R1165_U74
g14302 nand P1_R1165_U452 P1_R1165_U451 ; P1_R1165_U75
g14303 nand P1_R1165_U461 P1_R1165_U460 ; P1_R1165_U76
g14304 nand P1_R1165_U455 P1_R1165_U454 ; P1_R1165_U77
g14305 nand P1_R1165_U458 P1_R1165_U457 ; P1_R1165_U78
g14306 nand P1_R1165_U464 P1_R1165_U463 ; P1_R1165_U79
g14307 nand P1_R1165_U467 P1_R1165_U466 ; P1_R1165_U80
g14308 nand P1_R1165_U476 P1_R1165_U475 ; P1_R1165_U81
g14309 nand P1_R1165_U449 P1_R1165_U448 ; P1_R1165_U82
g14310 nand P1_R1165_U446 P1_R1165_U445 ; P1_R1165_U83
g14311 nand P1_R1165_U479 P1_R1165_U478 ; P1_R1165_U84
g14312 nand P1_R1165_U482 P1_R1165_U481 ; P1_R1165_U85
g14313 nand P1_R1165_U488 P1_R1165_U487 ; P1_R1165_U86
g14314 nand P1_R1165_U595 P1_R1165_U594 ; P1_R1165_U87
g14315 nand P1_R1165_U394 P1_R1165_U393 ; P1_R1165_U88
g14316 nand P1_R1165_U401 P1_R1165_U400 ; P1_R1165_U89
g14317 nand P1_R1165_U408 P1_R1165_U407 ; P1_R1165_U90
g14318 nand P1_R1165_U415 P1_R1165_U414 ; P1_R1165_U91
g14319 nand P1_R1165_U422 P1_R1165_U421 ; P1_R1165_U92
g14320 nand P1_R1165_U429 P1_R1165_U428 ; P1_R1165_U93
g14321 nand P1_R1165_U491 P1_R1165_U490 ; P1_R1165_U94
g14322 nand P1_R1165_U498 P1_R1165_U497 ; P1_R1165_U95
g14323 nand P1_R1165_U505 P1_R1165_U504 ; P1_R1165_U96
g14324 nand P1_R1165_U510 P1_R1165_U509 ; P1_R1165_U97
g14325 nand P1_R1165_U517 P1_R1165_U516 ; P1_R1165_U98
g14326 nand P1_R1165_U524 P1_R1165_U523 ; P1_R1165_U99
g14327 nand P1_R1165_U531 P1_R1165_U530 ; P1_R1165_U100
g14328 nand P1_R1165_U538 P1_R1165_U537 ; P1_R1165_U101
g14329 nand P1_R1165_U543 P1_R1165_U542 ; P1_R1165_U102
g14330 nand P1_R1165_U550 P1_R1165_U549 ; P1_R1165_U103
g14331 nand P1_R1165_U557 P1_R1165_U556 ; P1_R1165_U104
g14332 nand P1_R1165_U564 P1_R1165_U563 ; P1_R1165_U105
g14333 nand P1_R1165_U571 P1_R1165_U570 ; P1_R1165_U106
g14334 nand P1_R1165_U578 P1_R1165_U577 ; P1_R1165_U107
g14335 nand P1_R1165_U583 P1_R1165_U582 ; P1_R1165_U108
g14336 nand P1_R1165_U590 P1_R1165_U589 ; P1_R1165_U109
g14337 and P1_R1165_U205 P1_R1165_U204 ; P1_R1165_U110
g14338 and P1_R1165_U221 P1_R1165_U220 ; P1_R1165_U111
g14339 and P1_R1165_U403 P1_R1165_U402 P1_R1165_U17 ; P1_R1165_U112
g14340 and P1_R1165_U232 P1_R1165_U5 ; P1_R1165_U113
g14341 and P1_R1165_U424 P1_R1165_U423 P1_R1165_U20 ; P1_R1165_U114
g14342 and P1_R1165_U239 P1_R1165_U4 ; P1_R1165_U115
g14343 and P1_R1165_U255 P1_R1165_U6 ; P1_R1165_U116
g14344 and P1_R1165_U253 P1_R1165_U187 ; P1_R1165_U117
g14345 and P1_R1165_U273 P1_R1165_U272 ; P1_R1165_U118
g14346 and P1_R1165_U357 P1_R1165_U53 ; P1_R1165_U119
g14347 and P1_R1165_U306 P1_R1165_U301 ; P1_R1165_U120
g14348 and P1_R1165_U354 P1_R1165_U305 ; P1_R1165_U121
g14349 nand P1_R1165_U485 P1_R1165_U484 ; P1_R1165_U122
g14350 and P1_R1165_U500 P1_R1165_U499 P1_R1165_U189 ; P1_R1165_U123
g14351 and P1_R1165_U526 P1_R1165_U525 P1_R1165_U188 ; P1_R1165_U124
g14352 and P1_R1165_U552 P1_R1165_U551 P1_R1165_U38 ; P1_R1165_U125
g14353 and P1_R1165_U329 P1_R1165_U7 ; P1_R1165_U126
g14354 and P1_R1165_U573 P1_R1165_U572 P1_R1165_U187 ; P1_R1165_U127
g14355 and P1_R1165_U338 P1_R1165_U6 ; P1_R1165_U128
g14356 nand P1_R1165_U592 P1_R1165_U591 ; P1_R1165_U129
g14357 not P1_U3201 ; P1_R1165_U130
g14358 and P1_R1165_U362 P1_R1165_U361 ; P1_R1165_U131
g14359 not P1_U3210 ; P1_R1165_U132
g14360 not P1_U3209 ; P1_R1165_U133
g14361 not P1_U3207 ; P1_R1165_U134
g14362 not P1_U3208 ; P1_R1165_U135
g14363 not P1_U3206 ; P1_R1165_U136
g14364 not P1_U3205 ; P1_R1165_U137
g14365 not P1_U3203 ; P1_R1165_U138
g14366 not P1_U3204 ; P1_R1165_U139
g14367 not P1_U3202 ; P1_R1165_U140
g14368 and P1_R1165_U396 P1_R1165_U395 ; P1_R1165_U141
g14369 nand P1_R1165_U111 P1_R1165_U222 ; P1_R1165_U142
g14370 and P1_R1165_U410 P1_R1165_U409 ; P1_R1165_U143
g14371 nand P1_R1165_U210 P1_R1165_U209 ; P1_R1165_U144
g14372 and P1_R1165_U417 P1_R1165_U416 ; P1_R1165_U145
g14373 not P1_U3183 ; P1_R1165_U146
g14374 not P1_U3185 ; P1_R1165_U147
g14375 not P1_U3184 ; P1_R1165_U148
g14376 not P1_U3186 ; P1_R1165_U149
g14377 not P1_U3189 ; P1_R1165_U150
g14378 not P1_U3190 ; P1_R1165_U151
g14379 not P1_U3191 ; P1_R1165_U152
g14380 not P1_U3200 ; P1_R1165_U153
g14381 not P1_U3197 ; P1_R1165_U154
g14382 not P1_U3198 ; P1_R1165_U155
g14383 not P1_U3199 ; P1_R1165_U156
g14384 not P1_U3196 ; P1_R1165_U157
g14385 not P1_U3195 ; P1_R1165_U158
g14386 not P1_U3193 ; P1_R1165_U159
g14387 not P1_U3194 ; P1_R1165_U160
g14388 not P1_U3192 ; P1_R1165_U161
g14389 not P1_U3188 ; P1_R1165_U162
g14390 not P1_U3187 ; P1_R1165_U163
g14391 not P1_U3153 ; P1_R1165_U164
g14392 not P1_U3182 ; P1_R1165_U165
g14393 and P1_R1165_U493 P1_R1165_U492 ; P1_R1165_U166
g14394 nand P1_R1165_U351 P1_R1165_U302 P1_R1165_U53 ; P1_R1165_U167
g14395 nand P1_R1165_U296 P1_R1165_U295 ; P1_R1165_U168
g14396 and P1_R1165_U512 P1_R1165_U511 ; P1_R1165_U169
g14397 nand P1_R1165_U292 P1_R1165_U291 ; P1_R1165_U170
g14398 and P1_R1165_U519 P1_R1165_U518 ; P1_R1165_U171
g14399 nand P1_R1165_U287 P1_R1165_U283 P1_R1165_U288 ; P1_R1165_U172
g14400 and P1_R1165_U533 P1_R1165_U532 ; P1_R1165_U173
g14401 nand P1_R1165_U195 P1_R1165_U194 ; P1_R1165_U174
g14402 nand P1_R1165_U278 P1_R1165_U277 ; P1_R1165_U175
g14403 and P1_R1165_U545 P1_R1165_U544 ; P1_R1165_U176
g14404 nand P1_R1165_U118 P1_R1165_U274 ; P1_R1165_U177
g14405 and P1_R1165_U559 P1_R1165_U558 ; P1_R1165_U178
g14406 nand P1_R1165_U262 P1_R1165_U261 ; P1_R1165_U179
g14407 and P1_R1165_U566 P1_R1165_U565 ; P1_R1165_U180
g14408 nand P1_R1165_U258 P1_R1165_U257 ; P1_R1165_U181
g14409 nand P1_R1165_U248 P1_R1165_U247 ; P1_R1165_U182
g14410 and P1_R1165_U585 P1_R1165_U584 ; P1_R1165_U183
g14411 nand P1_R1165_U244 P1_R1165_U243 ; P1_R1165_U184
g14412 nand P1_R1165_U353 P1_R1165_U352 ; P1_R1165_U185
g14413 not P1_R1165_U20 ; P1_R1165_U186
g14414 nand P1_U3169 P1_R1165_U78 ; P1_R1165_U187
g14415 nand P1_U3161 P1_R1165_U83 ; P1_R1165_U188
g14416 nand P1_U3156 P1_R1165_U69 ; P1_R1165_U189
g14417 not P1_R1165_U43 ; P1_R1165_U190
g14418 not P1_R1165_U49 ; P1_R1165_U191
g14419 nand P1_U3157 P1_R1165_U71 ; P1_R1165_U192
g14420 or P1_U3211 P1_U3181 ; P1_R1165_U193
g14421 nand P1_R1165_U63 P1_R1165_U193 ; P1_R1165_U194
g14422 nand P1_U3181 P1_U3211 ; P1_R1165_U195
g14423 not P1_R1165_U174 ; P1_R1165_U196
g14424 nand P1_R1165_U371 P1_R1165_U23 ; P1_R1165_U197
g14425 nand P1_R1165_U197 P1_R1165_U174 ; P1_R1165_U198
g14426 nand P1_U3180 P1_R1165_U64 ; P1_R1165_U199
g14427 not P1_R1165_U31 ; P1_R1165_U200
g14428 nand P1_R1165_U374 P1_R1165_U21 ; P1_R1165_U201
g14429 nand P1_R1165_U377 P1_R1165_U19 ; P1_R1165_U202
g14430 nand P1_R1165_U21 P1_R1165_U20 ; P1_R1165_U203
g14431 nand P1_R1165_U62 P1_R1165_U203 ; P1_R1165_U204
g14432 nand P1_U3178 P1_R1165_U186 ; P1_R1165_U205
g14433 nand P1_R1165_U4 P1_R1165_U31 ; P1_R1165_U206
g14434 not P1_R1165_U24 ; P1_R1165_U207
g14435 nand P1_R1165_U207 P1_R1165_U25 ; P1_R1165_U208
g14436 nand P1_R1165_U65 P1_R1165_U208 ; P1_R1165_U209
g14437 nand P1_U3177 P1_R1165_U24 ; P1_R1165_U210
g14438 not P1_R1165_U144 ; P1_R1165_U211
g14439 nand P1_R1165_U383 P1_R1165_U26 ; P1_R1165_U212
g14440 nand P1_R1165_U212 P1_R1165_U144 ; P1_R1165_U213
g14441 nand P1_U3176 P1_R1165_U66 ; P1_R1165_U214
g14442 not P1_R1165_U30 ; P1_R1165_U215
g14443 nand P1_R1165_U386 P1_R1165_U18 ; P1_R1165_U216
g14444 nand P1_R1165_U389 P1_R1165_U16 ; P1_R1165_U217
g14445 not P1_R1165_U17 ; P1_R1165_U218
g14446 nand P1_R1165_U18 P1_R1165_U17 ; P1_R1165_U219
g14447 nand P1_R1165_U60 P1_R1165_U219 ; P1_R1165_U220
g14448 nand P1_U3174 P1_R1165_U218 ; P1_R1165_U221
g14449 nand P1_R1165_U5 P1_R1165_U30 ; P1_R1165_U222
g14450 not P1_R1165_U142 ; P1_R1165_U223
g14451 nand P1_R1165_U392 P1_R1165_U27 ; P1_R1165_U224
g14452 nand P1_R1165_U224 P1_R1165_U142 ; P1_R1165_U225
g14453 nand P1_U3173 P1_R1165_U67 ; P1_R1165_U226
g14454 not P1_R1165_U29 ; P1_R1165_U227
g14455 nand P1_R1165_U389 P1_R1165_U16 ; P1_R1165_U228
g14456 nand P1_R1165_U228 P1_R1165_U30 ; P1_R1165_U229
g14457 nand P1_R1165_U112 P1_R1165_U229 ; P1_R1165_U230
g14458 nand P1_R1165_U215 P1_R1165_U17 ; P1_R1165_U231
g14459 nand P1_U3174 P1_R1165_U60 ; P1_R1165_U232
g14460 nand P1_R1165_U113 P1_R1165_U231 ; P1_R1165_U233
g14461 nand P1_R1165_U389 P1_R1165_U16 ; P1_R1165_U234
g14462 nand P1_R1165_U377 P1_R1165_U19 ; P1_R1165_U235
g14463 nand P1_R1165_U235 P1_R1165_U31 ; P1_R1165_U236
g14464 nand P1_R1165_U114 P1_R1165_U236 ; P1_R1165_U237
g14465 nand P1_R1165_U200 P1_R1165_U20 ; P1_R1165_U238
g14466 nand P1_U3178 P1_R1165_U62 ; P1_R1165_U239
g14467 nand P1_R1165_U115 P1_R1165_U238 ; P1_R1165_U240
g14468 nand P1_R1165_U377 P1_R1165_U19 ; P1_R1165_U241
g14469 nand P1_R1165_U227 P1_R1165_U28 ; P1_R1165_U242
g14470 nand P1_R1165_U58 P1_R1165_U242 ; P1_R1165_U243
g14471 nand P1_U3172 P1_R1165_U29 ; P1_R1165_U244
g14472 not P1_R1165_U184 ; P1_R1165_U245
g14473 nand P1_R1165_U453 P1_R1165_U40 ; P1_R1165_U246
g14474 nand P1_R1165_U246 P1_R1165_U184 ; P1_R1165_U247
g14475 nand P1_U3171 P1_R1165_U75 ; P1_R1165_U248
g14476 not P1_R1165_U182 ; P1_R1165_U249
g14477 nand P1_R1165_U456 P1_R1165_U44 ; P1_R1165_U250
g14478 nand P1_R1165_U459 P1_R1165_U41 ; P1_R1165_U251
g14479 nand P1_R1165_U190 P1_R1165_U6 ; P1_R1165_U252
g14480 nand P1_U3168 P1_R1165_U77 ; P1_R1165_U253
g14481 nand P1_R1165_U117 P1_R1165_U252 ; P1_R1165_U254
g14482 nand P1_R1165_U462 P1_R1165_U42 ; P1_R1165_U255
g14483 nand P1_R1165_U456 P1_R1165_U44 ; P1_R1165_U256
g14484 nand P1_R1165_U116 P1_R1165_U182 ; P1_R1165_U257
g14485 nand P1_R1165_U256 P1_R1165_U254 ; P1_R1165_U258
g14486 not P1_R1165_U181 ; P1_R1165_U259
g14487 nand P1_R1165_U465 P1_R1165_U45 ; P1_R1165_U260
g14488 nand P1_R1165_U260 P1_R1165_U181 ; P1_R1165_U261
g14489 nand P1_U3167 P1_R1165_U79 ; P1_R1165_U262
g14490 not P1_R1165_U179 ; P1_R1165_U263
g14491 nand P1_R1165_U468 P1_R1165_U46 ; P1_R1165_U264
g14492 nand P1_R1165_U264 P1_R1165_U179 ; P1_R1165_U265
g14493 nand P1_U3166 P1_R1165_U80 ; P1_R1165_U266
g14494 not P1_R1165_U56 ; P1_R1165_U267
g14495 nand P1_R1165_U471 P1_R1165_U39 ; P1_R1165_U268
g14496 nand P1_R1165_U474 P1_R1165_U37 ; P1_R1165_U269
g14497 not P1_R1165_U38 ; P1_R1165_U270
g14498 nand P1_R1165_U39 P1_R1165_U38 ; P1_R1165_U271
g14499 nand P1_R1165_U74 P1_R1165_U271 ; P1_R1165_U272
g14500 nand P1_U3164 P1_R1165_U270 ; P1_R1165_U273
g14501 nand P1_R1165_U7 P1_R1165_U56 ; P1_R1165_U274
g14502 not P1_R1165_U177 ; P1_R1165_U275
g14503 nand P1_R1165_U477 P1_R1165_U47 ; P1_R1165_U276
g14504 nand P1_R1165_U276 P1_R1165_U177 ; P1_R1165_U277
g14505 nand P1_U3163 P1_R1165_U81 ; P1_R1165_U278
g14506 not P1_R1165_U175 ; P1_R1165_U279
g14507 nand P1_R1165_U444 P1_R1165_U36 ; P1_R1165_U280
g14508 nand P1_R1165_U447 P1_R1165_U50 ; P1_R1165_U281
g14509 nand P1_R1165_U191 P1_R1165_U8 ; P1_R1165_U282
g14510 nand P1_U3160 P1_R1165_U72 ; P1_R1165_U283
g14511 nand P1_R1165_U188 P1_R1165_U282 ; P1_R1165_U284
g14512 nand P1_R1165_U450 P1_R1165_U48 ; P1_R1165_U285
g14513 nand P1_R1165_U444 P1_R1165_U36 ; P1_R1165_U286
g14514 nand P1_R1165_U285 P1_R1165_U175 P1_R1165_U8 ; P1_R1165_U287
g14515 nand P1_R1165_U286 P1_R1165_U284 ; P1_R1165_U288
g14516 not P1_R1165_U172 ; P1_R1165_U289
g14517 nand P1_R1165_U480 P1_R1165_U51 ; P1_R1165_U290
g14518 nand P1_R1165_U290 P1_R1165_U172 ; P1_R1165_U291
g14519 nand P1_U3159 P1_R1165_U84 ; P1_R1165_U292
g14520 not P1_R1165_U170 ; P1_R1165_U293
g14521 nand P1_R1165_U483 P1_R1165_U52 ; P1_R1165_U294
g14522 nand P1_R1165_U294 P1_R1165_U170 ; P1_R1165_U295
g14523 nand P1_U3158 P1_R1165_U85 ; P1_R1165_U296
g14524 not P1_R1165_U168 ; P1_R1165_U297
g14525 nand P1_R1165_U435 P1_R1165_U34 ; P1_R1165_U298
g14526 nand P1_R1165_U192 P1_R1165_U189 ; P1_R1165_U299
g14527 not P1_R1165_U53 ; P1_R1165_U300
g14528 nand P1_R1165_U441 P1_R1165_U35 ; P1_R1165_U301
g14529 nand P1_R1165_U168 P1_R1165_U301 P1_R1165_U185 ; P1_R1165_U302
g14530 not P1_R1165_U167 ; P1_R1165_U303
g14531 nand P1_R1165_U432 P1_R1165_U32 ; P1_R1165_U304
g14532 nand P1_U3154 P1_R1165_U68 ; P1_R1165_U305
g14533 nand P1_R1165_U432 P1_R1165_U32 ; P1_R1165_U306
g14534 nand P1_R1165_U301 P1_R1165_U168 ; P1_R1165_U307
g14535 not P1_R1165_U54 ; P1_R1165_U308
g14536 nand P1_R1165_U435 P1_R1165_U34 ; P1_R1165_U309
g14537 nand P1_R1165_U309 P1_R1165_U54 ; P1_R1165_U310
g14538 nand P1_R1165_U123 P1_R1165_U310 ; P1_R1165_U311
g14539 nand P1_R1165_U308 P1_R1165_U189 ; P1_R1165_U312
g14540 nand P1_U3155 P1_R1165_U70 ; P1_R1165_U313
g14541 nand P1_R1165_U312 P1_R1165_U313 P1_R1165_U185 ; P1_R1165_U314
g14542 nand P1_R1165_U435 P1_R1165_U34 ; P1_R1165_U315
g14543 nand P1_R1165_U285 P1_R1165_U175 ; P1_R1165_U316
g14544 not P1_R1165_U55 ; P1_R1165_U317
g14545 nand P1_R1165_U447 P1_R1165_U50 ; P1_R1165_U318
g14546 nand P1_R1165_U318 P1_R1165_U55 ; P1_R1165_U319
g14547 nand P1_R1165_U124 P1_R1165_U319 ; P1_R1165_U320
g14548 nand P1_R1165_U317 P1_R1165_U188 ; P1_R1165_U321
g14549 nand P1_U3160 P1_R1165_U72 ; P1_R1165_U322
g14550 nand P1_R1165_U322 P1_R1165_U321 P1_R1165_U8 ; P1_R1165_U323
g14551 nand P1_R1165_U447 P1_R1165_U50 ; P1_R1165_U324
g14552 nand P1_R1165_U474 P1_R1165_U37 ; P1_R1165_U325
g14553 nand P1_R1165_U325 P1_R1165_U56 ; P1_R1165_U326
g14554 nand P1_R1165_U125 P1_R1165_U326 ; P1_R1165_U327
g14555 nand P1_R1165_U267 P1_R1165_U38 ; P1_R1165_U328
g14556 nand P1_U3164 P1_R1165_U74 ; P1_R1165_U329
g14557 nand P1_R1165_U126 P1_R1165_U328 ; P1_R1165_U330
g14558 nand P1_R1165_U474 P1_R1165_U37 ; P1_R1165_U331
g14559 nand P1_R1165_U255 P1_R1165_U182 ; P1_R1165_U332
g14560 not P1_R1165_U57 ; P1_R1165_U333
g14561 nand P1_R1165_U459 P1_R1165_U41 ; P1_R1165_U334
g14562 nand P1_R1165_U334 P1_R1165_U57 ; P1_R1165_U335
g14563 nand P1_R1165_U127 P1_R1165_U335 ; P1_R1165_U336
g14564 nand P1_R1165_U333 P1_R1165_U187 ; P1_R1165_U337
g14565 nand P1_U3168 P1_R1165_U77 ; P1_R1165_U338
g14566 nand P1_R1165_U128 P1_R1165_U337 ; P1_R1165_U339
g14567 nand P1_R1165_U459 P1_R1165_U41 ; P1_R1165_U340
g14568 nand P1_R1165_U234 P1_R1165_U17 ; P1_R1165_U341
g14569 nand P1_R1165_U241 P1_R1165_U20 ; P1_R1165_U342
g14570 nand P1_R1165_U315 P1_R1165_U189 ; P1_R1165_U343
g14571 nand P1_R1165_U301 P1_R1165_U192 ; P1_R1165_U344
g14572 nand P1_R1165_U324 P1_R1165_U188 ; P1_R1165_U345
g14573 nand P1_R1165_U285 P1_R1165_U49 ; P1_R1165_U346
g14574 nand P1_R1165_U331 P1_R1165_U38 ; P1_R1165_U347
g14575 nand P1_R1165_U340 P1_R1165_U187 ; P1_R1165_U348
g14576 nand P1_R1165_U255 P1_R1165_U43 ; P1_R1165_U349
g14577 nand P1_R1165_U351 P1_R1165_U302 P1_R1165_U119 ; P1_R1165_U350
g14578 nand P1_R1165_U299 P1_R1165_U185 ; P1_R1165_U351
g14579 nand P1_R1165_U70 P1_R1165_U298 ; P1_R1165_U352
g14580 nand P1_U3155 P1_R1165_U298 ; P1_R1165_U353
g14581 nand P1_R1165_U299 P1_R1165_U185 P1_R1165_U306 ; P1_R1165_U354
g14582 nand P1_R1165_U168 P1_R1165_U185 P1_R1165_U120 ; P1_R1165_U355
g14583 nand P1_R1165_U300 P1_R1165_U306 ; P1_R1165_U356
g14584 nand P1_U3154 P1_R1165_U68 ; P1_R1165_U357
g14585 nand P1_U3211 P1_R1165_U130 ; P1_R1165_U358
g14586 nand P1_U3201 P1_R1165_U15 ; P1_R1165_U359
g14587 not P1_R1165_U58 ; P1_R1165_U360
g14588 nand P1_R1165_U360 P1_U3172 ; P1_R1165_U361
g14589 nand P1_R1165_U58 P1_R1165_U28 ; P1_R1165_U362
g14590 nand P1_R1165_U360 P1_U3172 ; P1_R1165_U363
g14591 nand P1_R1165_U58 P1_R1165_U28 ; P1_R1165_U364
g14592 nand P1_R1165_U364 P1_R1165_U363 ; P1_R1165_U365
g14593 nand P1_U3211 P1_R1165_U132 ; P1_R1165_U366
g14594 nand P1_U3210 P1_R1165_U15 ; P1_R1165_U367
g14595 not P1_R1165_U63 ; P1_R1165_U368
g14596 nand P1_U3211 P1_R1165_U133 ; P1_R1165_U369
g14597 nand P1_U3209 P1_R1165_U15 ; P1_R1165_U370
g14598 not P1_R1165_U64 ; P1_R1165_U371
g14599 nand P1_U3211 P1_R1165_U134 ; P1_R1165_U372
g14600 nand P1_U3207 P1_R1165_U15 ; P1_R1165_U373
g14601 not P1_R1165_U62 ; P1_R1165_U374
g14602 nand P1_U3211 P1_R1165_U135 ; P1_R1165_U375
g14603 nand P1_U3208 P1_R1165_U15 ; P1_R1165_U376
g14604 not P1_R1165_U61 ; P1_R1165_U377
g14605 nand P1_U3211 P1_R1165_U136 ; P1_R1165_U378
g14606 nand P1_U3206 P1_R1165_U15 ; P1_R1165_U379
g14607 not P1_R1165_U65 ; P1_R1165_U380
g14608 nand P1_U3211 P1_R1165_U137 ; P1_R1165_U381
g14609 nand P1_U3205 P1_R1165_U15 ; P1_R1165_U382
g14610 not P1_R1165_U66 ; P1_R1165_U383
g14611 nand P1_U3211 P1_R1165_U138 ; P1_R1165_U384
g14612 nand P1_U3203 P1_R1165_U15 ; P1_R1165_U385
g14613 not P1_R1165_U60 ; P1_R1165_U386
g14614 nand P1_U3211 P1_R1165_U139 ; P1_R1165_U387
g14615 nand P1_U3204 P1_R1165_U15 ; P1_R1165_U388
g14616 not P1_R1165_U59 ; P1_R1165_U389
g14617 nand P1_U3211 P1_R1165_U140 ; P1_R1165_U390
g14618 nand P1_U3202 P1_R1165_U15 ; P1_R1165_U391
g14619 not P1_R1165_U67 ; P1_R1165_U392
g14620 nand P1_R1165_U131 P1_R1165_U29 ; P1_R1165_U393
g14621 nand P1_R1165_U365 P1_R1165_U227 ; P1_R1165_U394
g14622 nand P1_R1165_U392 P1_U3173 ; P1_R1165_U395
g14623 nand P1_R1165_U67 P1_R1165_U27 ; P1_R1165_U396
g14624 nand P1_R1165_U392 P1_U3173 ; P1_R1165_U397
g14625 nand P1_R1165_U67 P1_R1165_U27 ; P1_R1165_U398
g14626 nand P1_R1165_U398 P1_R1165_U397 ; P1_R1165_U399
g14627 nand P1_R1165_U141 P1_R1165_U142 ; P1_R1165_U400
g14628 nand P1_R1165_U223 P1_R1165_U399 ; P1_R1165_U401
g14629 nand P1_R1165_U386 P1_U3174 ; P1_R1165_U402
g14630 nand P1_R1165_U60 P1_R1165_U18 ; P1_R1165_U403
g14631 nand P1_R1165_U389 P1_U3175 ; P1_R1165_U404
g14632 nand P1_R1165_U59 P1_R1165_U16 ; P1_R1165_U405
g14633 nand P1_R1165_U405 P1_R1165_U404 ; P1_R1165_U406
g14634 nand P1_R1165_U341 P1_R1165_U30 ; P1_R1165_U407
g14635 nand P1_R1165_U406 P1_R1165_U215 ; P1_R1165_U408
g14636 nand P1_R1165_U383 P1_U3176 ; P1_R1165_U409
g14637 nand P1_R1165_U66 P1_R1165_U26 ; P1_R1165_U410
g14638 nand P1_R1165_U383 P1_U3176 ; P1_R1165_U411
g14639 nand P1_R1165_U66 P1_R1165_U26 ; P1_R1165_U412
g14640 nand P1_R1165_U412 P1_R1165_U411 ; P1_R1165_U413
g14641 nand P1_R1165_U143 P1_R1165_U144 ; P1_R1165_U414
g14642 nand P1_R1165_U211 P1_R1165_U413 ; P1_R1165_U415
g14643 nand P1_R1165_U380 P1_U3177 ; P1_R1165_U416
g14644 nand P1_R1165_U65 P1_R1165_U25 ; P1_R1165_U417
g14645 nand P1_R1165_U380 P1_U3177 ; P1_R1165_U418
g14646 nand P1_R1165_U65 P1_R1165_U25 ; P1_R1165_U419
g14647 nand P1_R1165_U419 P1_R1165_U418 ; P1_R1165_U420
g14648 nand P1_R1165_U145 P1_R1165_U24 ; P1_R1165_U421
g14649 nand P1_R1165_U420 P1_R1165_U207 ; P1_R1165_U422
g14650 nand P1_R1165_U374 P1_U3178 ; P1_R1165_U423
g14651 nand P1_R1165_U62 P1_R1165_U21 ; P1_R1165_U424
g14652 nand P1_R1165_U377 P1_U3179 ; P1_R1165_U425
g14653 nand P1_R1165_U61 P1_R1165_U19 ; P1_R1165_U426
g14654 nand P1_R1165_U426 P1_R1165_U425 ; P1_R1165_U427
g14655 nand P1_R1165_U342 P1_R1165_U31 ; P1_R1165_U428
g14656 nand P1_R1165_U427 P1_R1165_U200 ; P1_R1165_U429
g14657 nand P1_U3211 P1_R1165_U146 ; P1_R1165_U430
g14658 nand P1_U3183 P1_R1165_U15 ; P1_R1165_U431
g14659 not P1_R1165_U68 ; P1_R1165_U432
g14660 nand P1_U3211 P1_R1165_U147 ; P1_R1165_U433
g14661 nand P1_U3185 P1_R1165_U15 ; P1_R1165_U434
g14662 not P1_R1165_U69 ; P1_R1165_U435
g14663 nand P1_U3211 P1_R1165_U148 ; P1_R1165_U436
g14664 nand P1_U3184 P1_R1165_U15 ; P1_R1165_U437
g14665 not P1_R1165_U70 ; P1_R1165_U438
g14666 nand P1_U3211 P1_R1165_U149 ; P1_R1165_U439
g14667 nand P1_U3186 P1_R1165_U15 ; P1_R1165_U440
g14668 not P1_R1165_U71 ; P1_R1165_U441
g14669 nand P1_U3211 P1_R1165_U150 ; P1_R1165_U442
g14670 nand P1_U3189 P1_R1165_U15 ; P1_R1165_U443
g14671 not P1_R1165_U72 ; P1_R1165_U444
g14672 nand P1_U3211 P1_R1165_U151 ; P1_R1165_U445
g14673 nand P1_U3190 P1_R1165_U15 ; P1_R1165_U446
g14674 not P1_R1165_U83 ; P1_R1165_U447
g14675 nand P1_U3211 P1_R1165_U152 ; P1_R1165_U448
g14676 nand P1_U3191 P1_R1165_U15 ; P1_R1165_U449
g14677 not P1_R1165_U82 ; P1_R1165_U450
g14678 nand P1_U3211 P1_R1165_U153 ; P1_R1165_U451
g14679 nand P1_U3200 P1_R1165_U15 ; P1_R1165_U452
g14680 not P1_R1165_U75 ; P1_R1165_U453
g14681 nand P1_U3211 P1_R1165_U154 ; P1_R1165_U454
g14682 nand P1_U3197 P1_R1165_U15 ; P1_R1165_U455
g14683 not P1_R1165_U77 ; P1_R1165_U456
g14684 nand P1_U3211 P1_R1165_U155 ; P1_R1165_U457
g14685 nand P1_U3198 P1_R1165_U15 ; P1_R1165_U458
g14686 not P1_R1165_U78 ; P1_R1165_U459
g14687 nand P1_U3211 P1_R1165_U156 ; P1_R1165_U460
g14688 nand P1_U3199 P1_R1165_U15 ; P1_R1165_U461
g14689 not P1_R1165_U76 ; P1_R1165_U462
g14690 nand P1_U3211 P1_R1165_U157 ; P1_R1165_U463
g14691 nand P1_U3196 P1_R1165_U15 ; P1_R1165_U464
g14692 not P1_R1165_U79 ; P1_R1165_U465
g14693 nand P1_U3211 P1_R1165_U158 ; P1_R1165_U466
g14694 nand P1_U3195 P1_R1165_U15 ; P1_R1165_U467
g14695 not P1_R1165_U80 ; P1_R1165_U468
g14696 nand P1_U3211 P1_R1165_U159 ; P1_R1165_U469
g14697 nand P1_U3193 P1_R1165_U15 ; P1_R1165_U470
g14698 not P1_R1165_U74 ; P1_R1165_U471
g14699 nand P1_U3211 P1_R1165_U160 ; P1_R1165_U472
g14700 nand P1_U3194 P1_R1165_U15 ; P1_R1165_U473
g14701 not P1_R1165_U73 ; P1_R1165_U474
g14702 nand P1_U3211 P1_R1165_U161 ; P1_R1165_U475
g14703 nand P1_U3192 P1_R1165_U15 ; P1_R1165_U476
g14704 not P1_R1165_U81 ; P1_R1165_U477
g14705 nand P1_U3211 P1_R1165_U162 ; P1_R1165_U478
g14706 nand P1_U3188 P1_R1165_U15 ; P1_R1165_U479
g14707 not P1_R1165_U84 ; P1_R1165_U480
g14708 nand P1_U3211 P1_R1165_U163 ; P1_R1165_U481
g14709 nand P1_U3187 P1_R1165_U15 ; P1_R1165_U482
g14710 not P1_R1165_U85 ; P1_R1165_U483
g14711 nand P1_U3211 P1_R1165_U164 ; P1_R1165_U484
g14712 nand P1_U3153 P1_R1165_U15 ; P1_R1165_U485
g14713 not P1_R1165_U122 ; P1_R1165_U486
g14714 nand P1_U3182 P1_R1165_U486 ; P1_R1165_U487
g14715 nand P1_R1165_U122 P1_R1165_U165 ; P1_R1165_U488
g14716 not P1_R1165_U86 ; P1_R1165_U489
g14717 nand P1_R1165_U350 P1_R1165_U304 P1_R1165_U489 ; P1_R1165_U490
g14718 nand P1_R1165_U356 P1_R1165_U355 P1_R1165_U121 P1_R1165_U86 ; P1_R1165_U491
g14719 nand P1_R1165_U432 P1_U3154 ; P1_R1165_U492
g14720 nand P1_R1165_U68 P1_R1165_U32 ; P1_R1165_U493
g14721 nand P1_R1165_U432 P1_U3154 ; P1_R1165_U494
g14722 nand P1_R1165_U68 P1_R1165_U32 ; P1_R1165_U495
g14723 nand P1_R1165_U495 P1_R1165_U494 ; P1_R1165_U496
g14724 nand P1_R1165_U166 P1_R1165_U167 ; P1_R1165_U497
g14725 nand P1_R1165_U303 P1_R1165_U496 ; P1_R1165_U498
g14726 nand P1_R1165_U438 P1_U3155 ; P1_R1165_U499
g14727 nand P1_R1165_U70 P1_R1165_U33 ; P1_R1165_U500
g14728 nand P1_R1165_U435 P1_U3156 ; P1_R1165_U501
g14729 nand P1_R1165_U69 P1_R1165_U34 ; P1_R1165_U502
g14730 nand P1_R1165_U502 P1_R1165_U501 ; P1_R1165_U503
g14731 nand P1_R1165_U343 P1_R1165_U54 ; P1_R1165_U504
g14732 nand P1_R1165_U503 P1_R1165_U308 ; P1_R1165_U505
g14733 nand P1_R1165_U441 P1_U3157 ; P1_R1165_U506
g14734 nand P1_R1165_U71 P1_R1165_U35 ; P1_R1165_U507
g14735 nand P1_R1165_U507 P1_R1165_U506 ; P1_R1165_U508
g14736 nand P1_R1165_U344 P1_R1165_U168 ; P1_R1165_U509
g14737 nand P1_R1165_U297 P1_R1165_U508 ; P1_R1165_U510
g14738 nand P1_R1165_U483 P1_U3158 ; P1_R1165_U511
g14739 nand P1_R1165_U85 P1_R1165_U52 ; P1_R1165_U512
g14740 nand P1_R1165_U483 P1_U3158 ; P1_R1165_U513
g14741 nand P1_R1165_U85 P1_R1165_U52 ; P1_R1165_U514
g14742 nand P1_R1165_U514 P1_R1165_U513 ; P1_R1165_U515
g14743 nand P1_R1165_U169 P1_R1165_U170 ; P1_R1165_U516
g14744 nand P1_R1165_U293 P1_R1165_U515 ; P1_R1165_U517
g14745 nand P1_R1165_U480 P1_U3159 ; P1_R1165_U518
g14746 nand P1_R1165_U84 P1_R1165_U51 ; P1_R1165_U519
g14747 nand P1_R1165_U480 P1_U3159 ; P1_R1165_U520
g14748 nand P1_R1165_U84 P1_R1165_U51 ; P1_R1165_U521
g14749 nand P1_R1165_U521 P1_R1165_U520 ; P1_R1165_U522
g14750 nand P1_R1165_U171 P1_R1165_U172 ; P1_R1165_U523
g14751 nand P1_R1165_U289 P1_R1165_U522 ; P1_R1165_U524
g14752 nand P1_R1165_U444 P1_U3160 ; P1_R1165_U525
g14753 nand P1_R1165_U72 P1_R1165_U36 ; P1_R1165_U526
g14754 nand P1_R1165_U447 P1_U3161 ; P1_R1165_U527
g14755 nand P1_R1165_U83 P1_R1165_U50 ; P1_R1165_U528
g14756 nand P1_R1165_U528 P1_R1165_U527 ; P1_R1165_U529
g14757 nand P1_R1165_U345 P1_R1165_U55 ; P1_R1165_U530
g14758 nand P1_R1165_U529 P1_R1165_U317 ; P1_R1165_U531
g14759 nand P1_R1165_U371 P1_U3180 ; P1_R1165_U532
g14760 nand P1_R1165_U64 P1_R1165_U23 ; P1_R1165_U533
g14761 nand P1_R1165_U371 P1_U3180 ; P1_R1165_U534
g14762 nand P1_R1165_U64 P1_R1165_U23 ; P1_R1165_U535
g14763 nand P1_R1165_U535 P1_R1165_U534 ; P1_R1165_U536
g14764 nand P1_R1165_U173 P1_R1165_U174 ; P1_R1165_U537
g14765 nand P1_R1165_U196 P1_R1165_U536 ; P1_R1165_U538
g14766 nand P1_R1165_U450 P1_U3162 ; P1_R1165_U539
g14767 nand P1_R1165_U82 P1_R1165_U48 ; P1_R1165_U540
g14768 nand P1_R1165_U540 P1_R1165_U539 ; P1_R1165_U541
g14769 nand P1_R1165_U346 P1_R1165_U175 ; P1_R1165_U542
g14770 nand P1_R1165_U279 P1_R1165_U541 ; P1_R1165_U543
g14771 nand P1_R1165_U477 P1_U3163 ; P1_R1165_U544
g14772 nand P1_R1165_U81 P1_R1165_U47 ; P1_R1165_U545
g14773 nand P1_R1165_U477 P1_U3163 ; P1_R1165_U546
g14774 nand P1_R1165_U81 P1_R1165_U47 ; P1_R1165_U547
g14775 nand P1_R1165_U547 P1_R1165_U546 ; P1_R1165_U548
g14776 nand P1_R1165_U176 P1_R1165_U177 ; P1_R1165_U549
g14777 nand P1_R1165_U275 P1_R1165_U548 ; P1_R1165_U550
g14778 nand P1_R1165_U471 P1_U3164 ; P1_R1165_U551
g14779 nand P1_R1165_U74 P1_R1165_U39 ; P1_R1165_U552
g14780 nand P1_R1165_U474 P1_U3165 ; P1_R1165_U553
g14781 nand P1_R1165_U73 P1_R1165_U37 ; P1_R1165_U554
g14782 nand P1_R1165_U554 P1_R1165_U553 ; P1_R1165_U555
g14783 nand P1_R1165_U347 P1_R1165_U56 ; P1_R1165_U556
g14784 nand P1_R1165_U555 P1_R1165_U267 ; P1_R1165_U557
g14785 nand P1_R1165_U468 P1_U3166 ; P1_R1165_U558
g14786 nand P1_R1165_U80 P1_R1165_U46 ; P1_R1165_U559
g14787 nand P1_R1165_U468 P1_U3166 ; P1_R1165_U560
g14788 nand P1_R1165_U80 P1_R1165_U46 ; P1_R1165_U561
g14789 nand P1_R1165_U561 P1_R1165_U560 ; P1_R1165_U562
g14790 nand P1_R1165_U178 P1_R1165_U179 ; P1_R1165_U563
g14791 nand P1_R1165_U263 P1_R1165_U562 ; P1_R1165_U564
g14792 nand P1_R1165_U465 P1_U3167 ; P1_R1165_U565
g14793 nand P1_R1165_U79 P1_R1165_U45 ; P1_R1165_U566
g14794 nand P1_R1165_U465 P1_U3167 ; P1_R1165_U567
g14795 nand P1_R1165_U79 P1_R1165_U45 ; P1_R1165_U568
g14796 nand P1_R1165_U568 P1_R1165_U567 ; P1_R1165_U569
g14797 nand P1_R1165_U180 P1_R1165_U181 ; P1_R1165_U570
g14798 nand P1_R1165_U259 P1_R1165_U569 ; P1_R1165_U571
g14799 nand P1_R1165_U456 P1_U3168 ; P1_R1165_U572
g14800 nand P1_R1165_U77 P1_R1165_U44 ; P1_R1165_U573
g14801 nand P1_R1165_U459 P1_U3169 ; P1_R1165_U574
g14802 nand P1_R1165_U78 P1_R1165_U41 ; P1_R1165_U575
g14803 nand P1_R1165_U575 P1_R1165_U574 ; P1_R1165_U576
g14804 nand P1_R1165_U348 P1_R1165_U57 ; P1_R1165_U577
g14805 nand P1_R1165_U576 P1_R1165_U333 ; P1_R1165_U578
g14806 nand P1_R1165_U462 P1_U3170 ; P1_R1165_U579
g14807 nand P1_R1165_U76 P1_R1165_U42 ; P1_R1165_U580
g14808 nand P1_R1165_U580 P1_R1165_U579 ; P1_R1165_U581
g14809 nand P1_R1165_U349 P1_R1165_U182 ; P1_R1165_U582
g14810 nand P1_R1165_U249 P1_R1165_U581 ; P1_R1165_U583
g14811 nand P1_R1165_U453 P1_U3171 ; P1_R1165_U584
g14812 nand P1_R1165_U75 P1_R1165_U40 ; P1_R1165_U585
g14813 nand P1_R1165_U453 P1_U3171 ; P1_R1165_U586
g14814 nand P1_R1165_U75 P1_R1165_U40 ; P1_R1165_U587
g14815 nand P1_R1165_U587 P1_R1165_U586 ; P1_R1165_U588
g14816 nand P1_R1165_U183 P1_R1165_U184 ; P1_R1165_U589
g14817 nand P1_R1165_U245 P1_R1165_U588 ; P1_R1165_U590
g14818 nand P1_U3181 P1_R1165_U15 ; P1_R1165_U591
g14819 nand P1_U3211 P1_R1165_U22 ; P1_R1165_U592
g14820 not P1_R1165_U129 ; P1_R1165_U593
g14821 nand P1_R1165_U63 P1_R1165_U593 ; P1_R1165_U594
g14822 nand P1_R1165_U129 P1_R1165_U368 ; P1_R1165_U595
g14823 and P1_R1150_U184 P1_R1150_U201 ; P1_R1150_U6
g14824 and P1_R1150_U203 P1_R1150_U202 ; P1_R1150_U7
g14825 and P1_R1150_U179 P1_R1150_U240 ; P1_R1150_U8
g14826 and P1_R1150_U242 P1_R1150_U241 ; P1_R1150_U9
g14827 and P1_R1150_U259 P1_R1150_U258 ; P1_R1150_U10
g14828 and P1_R1150_U285 P1_R1150_U284 ; P1_R1150_U11
g14829 and P1_R1150_U383 P1_R1150_U382 ; P1_R1150_U12
g14830 nand P1_R1150_U340 P1_R1150_U343 ; P1_R1150_U13
g14831 nand P1_R1150_U329 P1_R1150_U332 ; P1_R1150_U14
g14832 nand P1_R1150_U318 P1_R1150_U321 ; P1_R1150_U15
g14833 nand P1_R1150_U310 P1_R1150_U312 ; P1_R1150_U16
g14834 nand P1_R1150_U156 P1_R1150_U175 P1_R1150_U348 ; P1_R1150_U17
g14835 nand P1_R1150_U236 P1_R1150_U238 ; P1_R1150_U18
g14836 nand P1_R1150_U228 P1_R1150_U231 ; P1_R1150_U19
g14837 nand P1_R1150_U220 P1_R1150_U222 ; P1_R1150_U20
g14838 nand P1_R1150_U25 P1_R1150_U346 ; P1_R1150_U21
g14839 not P1_U3479 ; P1_R1150_U22
g14840 not P1_U3464 ; P1_R1150_U23
g14841 not P1_U3456 ; P1_R1150_U24
g14842 nand P1_U3456 P1_R1150_U93 ; P1_R1150_U25
g14843 not P1_U3078 ; P1_R1150_U26
g14844 not P1_U3467 ; P1_R1150_U27
g14845 not P1_U3068 ; P1_R1150_U28
g14846 nand P1_U3068 P1_R1150_U23 ; P1_R1150_U29
g14847 not P1_U3064 ; P1_R1150_U30
g14848 not P1_U3476 ; P1_R1150_U31
g14849 not P1_U3473 ; P1_R1150_U32
g14850 not P1_U3470 ; P1_R1150_U33
g14851 not P1_U3071 ; P1_R1150_U34
g14852 not P1_U3067 ; P1_R1150_U35
g14853 not P1_U3060 ; P1_R1150_U36
g14854 nand P1_U3060 P1_R1150_U33 ; P1_R1150_U37
g14855 not P1_U3482 ; P1_R1150_U38
g14856 not P1_U3070 ; P1_R1150_U39
g14857 nand P1_U3070 P1_R1150_U22 ; P1_R1150_U40
g14858 not P1_U3084 ; P1_R1150_U41
g14859 not P1_U3485 ; P1_R1150_U42
g14860 not P1_U3083 ; P1_R1150_U43
g14861 nand P1_R1150_U209 P1_R1150_U208 ; P1_R1150_U44
g14862 nand P1_R1150_U37 P1_R1150_U224 ; P1_R1150_U45
g14863 nand P1_R1150_U193 P1_R1150_U192 ; P1_R1150_U46
g14864 not P1_U4019 ; P1_R1150_U47
g14865 not P1_U4023 ; P1_R1150_U48
g14866 not P1_U3503 ; P1_R1150_U49
g14867 not P1_U3491 ; P1_R1150_U50
g14868 not P1_U3488 ; P1_R1150_U51
g14869 not P1_U3063 ; P1_R1150_U52
g14870 not P1_U3062 ; P1_R1150_U53
g14871 nand P1_U3083 P1_R1150_U42 ; P1_R1150_U54
g14872 not P1_U3494 ; P1_R1150_U55
g14873 not P1_U3072 ; P1_R1150_U56
g14874 not P1_U3497 ; P1_R1150_U57
g14875 not P1_U3080 ; P1_R1150_U58
g14876 not P1_U3506 ; P1_R1150_U59
g14877 not P1_U3500 ; P1_R1150_U60
g14878 not P1_U3073 ; P1_R1150_U61
g14879 not P1_U3074 ; P1_R1150_U62
g14880 not P1_U3079 ; P1_R1150_U63
g14881 nand P1_U3079 P1_R1150_U60 ; P1_R1150_U64
g14882 not P1_U3509 ; P1_R1150_U65
g14883 not P1_U3069 ; P1_R1150_U66
g14884 nand P1_R1150_U269 P1_R1150_U268 ; P1_R1150_U67
g14885 not P1_U3082 ; P1_R1150_U68
g14886 not P1_U3514 ; P1_R1150_U69
g14887 not P1_U3081 ; P1_R1150_U70
g14888 not P1_U4025 ; P1_R1150_U71
g14889 not P1_U3076 ; P1_R1150_U72
g14890 not P1_U4022 ; P1_R1150_U73
g14891 not P1_U4024 ; P1_R1150_U74
g14892 not P1_U3066 ; P1_R1150_U75
g14893 not P1_U3061 ; P1_R1150_U76
g14894 not P1_U3075 ; P1_R1150_U77
g14895 nand P1_U3075 P1_R1150_U74 ; P1_R1150_U78
g14896 not P1_U4021 ; P1_R1150_U79
g14897 not P1_U3065 ; P1_R1150_U80
g14898 not P1_U4020 ; P1_R1150_U81
g14899 not P1_U3058 ; P1_R1150_U82
g14900 not P1_U4018 ; P1_R1150_U83
g14901 not P1_U3057 ; P1_R1150_U84
g14902 nand P1_U3057 P1_R1150_U47 ; P1_R1150_U85
g14903 not P1_U3053 ; P1_R1150_U86
g14904 not P1_U4017 ; P1_R1150_U87
g14905 not P1_U3054 ; P1_R1150_U88
g14906 nand P1_R1150_U299 P1_R1150_U298 ; P1_R1150_U89
g14907 nand P1_R1150_U78 P1_R1150_U314 ; P1_R1150_U90
g14908 nand P1_R1150_U64 P1_R1150_U325 ; P1_R1150_U91
g14909 nand P1_R1150_U54 P1_R1150_U336 ; P1_R1150_U92
g14910 not P1_U3077 ; P1_R1150_U93
g14911 nand P1_R1150_U393 P1_R1150_U392 ; P1_R1150_U94
g14912 nand P1_R1150_U407 P1_R1150_U406 ; P1_R1150_U95
g14913 nand P1_R1150_U412 P1_R1150_U411 ; P1_R1150_U96
g14914 nand P1_R1150_U428 P1_R1150_U427 ; P1_R1150_U97
g14915 nand P1_R1150_U433 P1_R1150_U432 ; P1_R1150_U98
g14916 nand P1_R1150_U438 P1_R1150_U437 ; P1_R1150_U99
g14917 nand P1_R1150_U443 P1_R1150_U442 ; P1_R1150_U100
g14918 nand P1_R1150_U448 P1_R1150_U447 ; P1_R1150_U101
g14919 nand P1_R1150_U464 P1_R1150_U463 ; P1_R1150_U102
g14920 nand P1_R1150_U469 P1_R1150_U468 ; P1_R1150_U103
g14921 nand P1_R1150_U352 P1_R1150_U351 ; P1_R1150_U104
g14922 nand P1_R1150_U361 P1_R1150_U360 ; P1_R1150_U105
g14923 nand P1_R1150_U368 P1_R1150_U367 ; P1_R1150_U106
g14924 nand P1_R1150_U372 P1_R1150_U371 ; P1_R1150_U107
g14925 nand P1_R1150_U381 P1_R1150_U380 ; P1_R1150_U108
g14926 nand P1_R1150_U402 P1_R1150_U401 ; P1_R1150_U109
g14927 nand P1_R1150_U419 P1_R1150_U418 ; P1_R1150_U110
g14928 nand P1_R1150_U423 P1_R1150_U422 ; P1_R1150_U111
g14929 nand P1_R1150_U455 P1_R1150_U454 ; P1_R1150_U112
g14930 nand P1_R1150_U459 P1_R1150_U458 ; P1_R1150_U113
g14931 nand P1_R1150_U476 P1_R1150_U475 ; P1_R1150_U114
g14932 and P1_R1150_U195 P1_R1150_U183 ; P1_R1150_U115
g14933 and P1_R1150_U198 P1_R1150_U199 ; P1_R1150_U116
g14934 and P1_R1150_U211 P1_R1150_U185 ; P1_R1150_U117
g14935 and P1_R1150_U214 P1_R1150_U215 ; P1_R1150_U118
g14936 and P1_R1150_U354 P1_R1150_U353 P1_R1150_U40 ; P1_R1150_U119
g14937 and P1_R1150_U357 P1_R1150_U185 ; P1_R1150_U120
g14938 and P1_R1150_U230 P1_R1150_U7 ; P1_R1150_U121
g14939 and P1_R1150_U364 P1_R1150_U184 ; P1_R1150_U122
g14940 and P1_R1150_U374 P1_R1150_U373 P1_R1150_U29 ; P1_R1150_U123
g14941 and P1_R1150_U377 P1_R1150_U183 ; P1_R1150_U124
g14942 and P1_R1150_U217 P1_R1150_U8 ; P1_R1150_U125
g14943 and P1_R1150_U262 P1_R1150_U180 ; P1_R1150_U126
g14944 and P1_R1150_U288 P1_R1150_U181 ; P1_R1150_U127
g14945 and P1_R1150_U304 P1_R1150_U305 ; P1_R1150_U128
g14946 and P1_R1150_U307 P1_R1150_U386 ; P1_R1150_U129
g14947 and P1_R1150_U305 P1_R1150_U304 P1_R1150_U308 ; P1_R1150_U130
g14948 nand P1_R1150_U390 P1_R1150_U389 ; P1_R1150_U131
g14949 and P1_R1150_U395 P1_R1150_U394 P1_R1150_U85 ; P1_R1150_U132
g14950 and P1_R1150_U398 P1_R1150_U182 ; P1_R1150_U133
g14951 nand P1_R1150_U404 P1_R1150_U403 ; P1_R1150_U134
g14952 nand P1_R1150_U409 P1_R1150_U408 ; P1_R1150_U135
g14953 and P1_R1150_U415 P1_R1150_U181 ; P1_R1150_U136
g14954 nand P1_R1150_U425 P1_R1150_U424 ; P1_R1150_U137
g14955 nand P1_R1150_U430 P1_R1150_U429 ; P1_R1150_U138
g14956 nand P1_R1150_U435 P1_R1150_U434 ; P1_R1150_U139
g14957 nand P1_R1150_U440 P1_R1150_U439 ; P1_R1150_U140
g14958 nand P1_R1150_U445 P1_R1150_U444 ; P1_R1150_U141
g14959 and P1_R1150_U451 P1_R1150_U180 ; P1_R1150_U142
g14960 nand P1_R1150_U461 P1_R1150_U460 ; P1_R1150_U143
g14961 nand P1_R1150_U466 P1_R1150_U465 ; P1_R1150_U144
g14962 and P1_R1150_U342 P1_R1150_U9 ; P1_R1150_U145
g14963 and P1_R1150_U472 P1_R1150_U179 ; P1_R1150_U146
g14964 and P1_R1150_U350 P1_R1150_U349 ; P1_R1150_U147
g14965 nand P1_R1150_U118 P1_R1150_U212 ; P1_R1150_U148
g14966 and P1_R1150_U359 P1_R1150_U358 ; P1_R1150_U149
g14967 and P1_R1150_U366 P1_R1150_U365 ; P1_R1150_U150
g14968 and P1_R1150_U370 P1_R1150_U369 ; P1_R1150_U151
g14969 nand P1_R1150_U116 P1_R1150_U196 ; P1_R1150_U152
g14970 and P1_R1150_U379 P1_R1150_U378 ; P1_R1150_U153
g14971 not P1_U4028 ; P1_R1150_U154
g14972 not P1_U3055 ; P1_R1150_U155
g14973 and P1_R1150_U388 P1_R1150_U387 ; P1_R1150_U156
g14974 nand P1_R1150_U128 P1_R1150_U302 ; P1_R1150_U157
g14975 and P1_R1150_U400 P1_R1150_U399 ; P1_R1150_U158
g14976 nand P1_R1150_U295 P1_R1150_U294 ; P1_R1150_U159
g14977 nand P1_R1150_U291 P1_R1150_U290 ; P1_R1150_U160
g14978 and P1_R1150_U417 P1_R1150_U416 ; P1_R1150_U161
g14979 and P1_R1150_U421 P1_R1150_U420 ; P1_R1150_U162
g14980 nand P1_R1150_U281 P1_R1150_U280 ; P1_R1150_U163
g14981 nand P1_R1150_U277 P1_R1150_U276 ; P1_R1150_U164
g14982 not P1_U3461 ; P1_R1150_U165
g14983 nand P1_R1150_U273 P1_R1150_U272 ; P1_R1150_U166
g14984 not P1_U3512 ; P1_R1150_U167
g14985 nand P1_R1150_U265 P1_R1150_U264 ; P1_R1150_U168
g14986 and P1_R1150_U453 P1_R1150_U452 ; P1_R1150_U169
g14987 and P1_R1150_U457 P1_R1150_U456 ; P1_R1150_U170
g14988 nand P1_R1150_U255 P1_R1150_U254 ; P1_R1150_U171
g14989 nand P1_R1150_U251 P1_R1150_U250 ; P1_R1150_U172
g14990 nand P1_R1150_U247 P1_R1150_U246 ; P1_R1150_U173
g14991 and P1_R1150_U474 P1_R1150_U473 ; P1_R1150_U174
g14992 nand P1_R1150_U129 P1_R1150_U157 ; P1_R1150_U175
g14993 not P1_R1150_U85 ; P1_R1150_U176
g14994 not P1_R1150_U29 ; P1_R1150_U177
g14995 not P1_R1150_U40 ; P1_R1150_U178
g14996 nand P1_U3488 P1_R1150_U53 ; P1_R1150_U179
g14997 nand P1_U3503 P1_R1150_U62 ; P1_R1150_U180
g14998 nand P1_U4023 P1_R1150_U76 ; P1_R1150_U181
g14999 nand P1_U4019 P1_R1150_U84 ; P1_R1150_U182
g15000 nand P1_U3464 P1_R1150_U28 ; P1_R1150_U183
g15001 nand P1_U3473 P1_R1150_U35 ; P1_R1150_U184
g15002 nand P1_U3479 P1_R1150_U39 ; P1_R1150_U185
g15003 not P1_R1150_U64 ; P1_R1150_U186
g15004 not P1_R1150_U78 ; P1_R1150_U187
g15005 not P1_R1150_U37 ; P1_R1150_U188
g15006 not P1_R1150_U54 ; P1_R1150_U189
g15007 not P1_R1150_U25 ; P1_R1150_U190
g15008 nand P1_R1150_U190 P1_R1150_U26 ; P1_R1150_U191
g15009 nand P1_R1150_U191 P1_R1150_U165 ; P1_R1150_U192
g15010 nand P1_U3078 P1_R1150_U25 ; P1_R1150_U193
g15011 not P1_R1150_U46 ; P1_R1150_U194
g15012 nand P1_U3467 P1_R1150_U30 ; P1_R1150_U195
g15013 nand P1_R1150_U115 P1_R1150_U46 ; P1_R1150_U196
g15014 nand P1_R1150_U30 P1_R1150_U29 ; P1_R1150_U197
g15015 nand P1_R1150_U197 P1_R1150_U27 ; P1_R1150_U198
g15016 nand P1_U3064 P1_R1150_U177 ; P1_R1150_U199
g15017 not P1_R1150_U152 ; P1_R1150_U200
g15018 nand P1_U3476 P1_R1150_U34 ; P1_R1150_U201
g15019 nand P1_U3071 P1_R1150_U31 ; P1_R1150_U202
g15020 nand P1_U3067 P1_R1150_U32 ; P1_R1150_U203
g15021 nand P1_R1150_U188 P1_R1150_U6 ; P1_R1150_U204
g15022 nand P1_R1150_U7 P1_R1150_U204 ; P1_R1150_U205
g15023 nand P1_U3470 P1_R1150_U36 ; P1_R1150_U206
g15024 nand P1_U3476 P1_R1150_U34 ; P1_R1150_U207
g15025 nand P1_R1150_U206 P1_R1150_U152 P1_R1150_U6 ; P1_R1150_U208
g15026 nand P1_R1150_U207 P1_R1150_U205 ; P1_R1150_U209
g15027 not P1_R1150_U44 ; P1_R1150_U210
g15028 nand P1_U3482 P1_R1150_U41 ; P1_R1150_U211
g15029 nand P1_R1150_U117 P1_R1150_U44 ; P1_R1150_U212
g15030 nand P1_R1150_U41 P1_R1150_U40 ; P1_R1150_U213
g15031 nand P1_R1150_U213 P1_R1150_U38 ; P1_R1150_U214
g15032 nand P1_U3084 P1_R1150_U178 ; P1_R1150_U215
g15033 not P1_R1150_U148 ; P1_R1150_U216
g15034 nand P1_U3485 P1_R1150_U43 ; P1_R1150_U217
g15035 nand P1_R1150_U217 P1_R1150_U54 ; P1_R1150_U218
g15036 nand P1_R1150_U210 P1_R1150_U40 ; P1_R1150_U219
g15037 nand P1_R1150_U120 P1_R1150_U219 ; P1_R1150_U220
g15038 nand P1_R1150_U44 P1_R1150_U185 ; P1_R1150_U221
g15039 nand P1_R1150_U119 P1_R1150_U221 ; P1_R1150_U222
g15040 nand P1_R1150_U40 P1_R1150_U185 ; P1_R1150_U223
g15041 nand P1_R1150_U206 P1_R1150_U152 ; P1_R1150_U224
g15042 not P1_R1150_U45 ; P1_R1150_U225
g15043 nand P1_U3067 P1_R1150_U32 ; P1_R1150_U226
g15044 nand P1_R1150_U225 P1_R1150_U226 ; P1_R1150_U227
g15045 nand P1_R1150_U122 P1_R1150_U227 ; P1_R1150_U228
g15046 nand P1_R1150_U45 P1_R1150_U184 ; P1_R1150_U229
g15047 nand P1_U3476 P1_R1150_U34 ; P1_R1150_U230
g15048 nand P1_R1150_U121 P1_R1150_U229 ; P1_R1150_U231
g15049 nand P1_U3067 P1_R1150_U32 ; P1_R1150_U232
g15050 nand P1_R1150_U184 P1_R1150_U232 ; P1_R1150_U233
g15051 nand P1_R1150_U206 P1_R1150_U37 ; P1_R1150_U234
g15052 nand P1_R1150_U194 P1_R1150_U29 ; P1_R1150_U235
g15053 nand P1_R1150_U124 P1_R1150_U235 ; P1_R1150_U236
g15054 nand P1_R1150_U46 P1_R1150_U183 ; P1_R1150_U237
g15055 nand P1_R1150_U123 P1_R1150_U237 ; P1_R1150_U238
g15056 nand P1_R1150_U29 P1_R1150_U183 ; P1_R1150_U239
g15057 nand P1_U3491 P1_R1150_U52 ; P1_R1150_U240
g15058 nand P1_U3063 P1_R1150_U50 ; P1_R1150_U241
g15059 nand P1_U3062 P1_R1150_U51 ; P1_R1150_U242
g15060 nand P1_R1150_U189 P1_R1150_U8 ; P1_R1150_U243
g15061 nand P1_R1150_U9 P1_R1150_U243 ; P1_R1150_U244
g15062 nand P1_U3491 P1_R1150_U52 ; P1_R1150_U245
g15063 nand P1_R1150_U125 P1_R1150_U148 ; P1_R1150_U246
g15064 nand P1_R1150_U245 P1_R1150_U244 ; P1_R1150_U247
g15065 not P1_R1150_U173 ; P1_R1150_U248
g15066 nand P1_U3494 P1_R1150_U56 ; P1_R1150_U249
g15067 nand P1_R1150_U249 P1_R1150_U173 ; P1_R1150_U250
g15068 nand P1_U3072 P1_R1150_U55 ; P1_R1150_U251
g15069 not P1_R1150_U172 ; P1_R1150_U252
g15070 nand P1_U3497 P1_R1150_U58 ; P1_R1150_U253
g15071 nand P1_R1150_U253 P1_R1150_U172 ; P1_R1150_U254
g15072 nand P1_U3080 P1_R1150_U57 ; P1_R1150_U255
g15073 not P1_R1150_U171 ; P1_R1150_U256
g15074 nand P1_U3506 P1_R1150_U61 ; P1_R1150_U257
g15075 nand P1_U3073 P1_R1150_U59 ; P1_R1150_U258
g15076 nand P1_U3074 P1_R1150_U49 ; P1_R1150_U259
g15077 nand P1_R1150_U186 P1_R1150_U180 ; P1_R1150_U260
g15078 nand P1_R1150_U10 P1_R1150_U260 ; P1_R1150_U261
g15079 nand P1_U3500 P1_R1150_U63 ; P1_R1150_U262
g15080 nand P1_U3506 P1_R1150_U61 ; P1_R1150_U263
g15081 nand P1_R1150_U171 P1_R1150_U126 P1_R1150_U257 ; P1_R1150_U264
g15082 nand P1_R1150_U263 P1_R1150_U261 ; P1_R1150_U265
g15083 not P1_R1150_U168 ; P1_R1150_U266
g15084 nand P1_U3509 P1_R1150_U66 ; P1_R1150_U267
g15085 nand P1_R1150_U267 P1_R1150_U168 ; P1_R1150_U268
g15086 nand P1_U3069 P1_R1150_U65 ; P1_R1150_U269
g15087 not P1_R1150_U67 ; P1_R1150_U270
g15088 nand P1_R1150_U270 P1_R1150_U68 ; P1_R1150_U271
g15089 nand P1_R1150_U271 P1_R1150_U167 ; P1_R1150_U272
g15090 nand P1_U3082 P1_R1150_U67 ; P1_R1150_U273
g15091 not P1_R1150_U166 ; P1_R1150_U274
g15092 nand P1_U3514 P1_R1150_U70 ; P1_R1150_U275
g15093 nand P1_R1150_U275 P1_R1150_U166 ; P1_R1150_U276
g15094 nand P1_U3081 P1_R1150_U69 ; P1_R1150_U277
g15095 not P1_R1150_U164 ; P1_R1150_U278
g15096 nand P1_U4025 P1_R1150_U72 ; P1_R1150_U279
g15097 nand P1_R1150_U279 P1_R1150_U164 ; P1_R1150_U280
g15098 nand P1_U3076 P1_R1150_U71 ; P1_R1150_U281
g15099 not P1_R1150_U163 ; P1_R1150_U282
g15100 nand P1_U4022 P1_R1150_U75 ; P1_R1150_U283
g15101 nand P1_U3066 P1_R1150_U73 ; P1_R1150_U284
g15102 nand P1_U3061 P1_R1150_U48 ; P1_R1150_U285
g15103 nand P1_R1150_U187 P1_R1150_U181 ; P1_R1150_U286
g15104 nand P1_R1150_U11 P1_R1150_U286 ; P1_R1150_U287
g15105 nand P1_U4024 P1_R1150_U77 ; P1_R1150_U288
g15106 nand P1_U4022 P1_R1150_U75 ; P1_R1150_U289
g15107 nand P1_R1150_U163 P1_R1150_U127 P1_R1150_U283 ; P1_R1150_U290
g15108 nand P1_R1150_U289 P1_R1150_U287 ; P1_R1150_U291
g15109 not P1_R1150_U160 ; P1_R1150_U292
g15110 nand P1_U4021 P1_R1150_U80 ; P1_R1150_U293
g15111 nand P1_R1150_U293 P1_R1150_U160 ; P1_R1150_U294
g15112 nand P1_U3065 P1_R1150_U79 ; P1_R1150_U295
g15113 not P1_R1150_U159 ; P1_R1150_U296
g15114 nand P1_U4020 P1_R1150_U82 ; P1_R1150_U297
g15115 nand P1_R1150_U297 P1_R1150_U159 ; P1_R1150_U298
g15116 nand P1_U3058 P1_R1150_U81 ; P1_R1150_U299
g15117 not P1_R1150_U89 ; P1_R1150_U300
g15118 nand P1_U4018 P1_R1150_U86 ; P1_R1150_U301
g15119 nand P1_R1150_U89 P1_R1150_U182 P1_R1150_U301 ; P1_R1150_U302
g15120 nand P1_R1150_U86 P1_R1150_U85 ; P1_R1150_U303
g15121 nand P1_R1150_U303 P1_R1150_U83 ; P1_R1150_U304
g15122 nand P1_U3053 P1_R1150_U176 ; P1_R1150_U305
g15123 not P1_R1150_U157 ; P1_R1150_U306
g15124 nand P1_U4017 P1_R1150_U88 ; P1_R1150_U307
g15125 nand P1_U3054 P1_R1150_U87 ; P1_R1150_U308
g15126 nand P1_R1150_U300 P1_R1150_U85 ; P1_R1150_U309
g15127 nand P1_R1150_U133 P1_R1150_U309 ; P1_R1150_U310
g15128 nand P1_R1150_U89 P1_R1150_U182 ; P1_R1150_U311
g15129 nand P1_R1150_U132 P1_R1150_U311 ; P1_R1150_U312
g15130 nand P1_R1150_U85 P1_R1150_U182 ; P1_R1150_U313
g15131 nand P1_R1150_U288 P1_R1150_U163 ; P1_R1150_U314
g15132 not P1_R1150_U90 ; P1_R1150_U315
g15133 nand P1_U3061 P1_R1150_U48 ; P1_R1150_U316
g15134 nand P1_R1150_U315 P1_R1150_U316 ; P1_R1150_U317
g15135 nand P1_R1150_U136 P1_R1150_U317 ; P1_R1150_U318
g15136 nand P1_R1150_U90 P1_R1150_U181 ; P1_R1150_U319
g15137 nand P1_U4022 P1_R1150_U75 ; P1_R1150_U320
g15138 nand P1_R1150_U320 P1_R1150_U319 P1_R1150_U11 ; P1_R1150_U321
g15139 nand P1_U3061 P1_R1150_U48 ; P1_R1150_U322
g15140 nand P1_R1150_U181 P1_R1150_U322 ; P1_R1150_U323
g15141 nand P1_R1150_U288 P1_R1150_U78 ; P1_R1150_U324
g15142 nand P1_R1150_U262 P1_R1150_U171 ; P1_R1150_U325
g15143 not P1_R1150_U91 ; P1_R1150_U326
g15144 nand P1_U3074 P1_R1150_U49 ; P1_R1150_U327
g15145 nand P1_R1150_U326 P1_R1150_U327 ; P1_R1150_U328
g15146 nand P1_R1150_U142 P1_R1150_U328 ; P1_R1150_U329
g15147 nand P1_R1150_U91 P1_R1150_U180 ; P1_R1150_U330
g15148 nand P1_U3506 P1_R1150_U61 ; P1_R1150_U331
g15149 nand P1_R1150_U331 P1_R1150_U330 P1_R1150_U10 ; P1_R1150_U332
g15150 nand P1_U3074 P1_R1150_U49 ; P1_R1150_U333
g15151 nand P1_R1150_U180 P1_R1150_U333 ; P1_R1150_U334
g15152 nand P1_R1150_U262 P1_R1150_U64 ; P1_R1150_U335
g15153 nand P1_R1150_U217 P1_R1150_U148 ; P1_R1150_U336
g15154 not P1_R1150_U92 ; P1_R1150_U337
g15155 nand P1_U3062 P1_R1150_U51 ; P1_R1150_U338
g15156 nand P1_R1150_U337 P1_R1150_U338 ; P1_R1150_U339
g15157 nand P1_R1150_U146 P1_R1150_U339 ; P1_R1150_U340
g15158 nand P1_R1150_U92 P1_R1150_U179 ; P1_R1150_U341
g15159 nand P1_U3491 P1_R1150_U52 ; P1_R1150_U342
g15160 nand P1_R1150_U145 P1_R1150_U341 ; P1_R1150_U343
g15161 nand P1_U3062 P1_R1150_U51 ; P1_R1150_U344
g15162 nand P1_R1150_U179 P1_R1150_U344 ; P1_R1150_U345
g15163 nand P1_U3077 P1_R1150_U24 ; P1_R1150_U346
g15164 nand P1_R1150_U89 P1_R1150_U182 P1_R1150_U301 ; P1_R1150_U347
g15165 nand P1_R1150_U12 P1_R1150_U347 P1_R1150_U130 ; P1_R1150_U348
g15166 nand P1_U3485 P1_R1150_U43 ; P1_R1150_U349
g15167 nand P1_U3083 P1_R1150_U42 ; P1_R1150_U350
g15168 nand P1_R1150_U218 P1_R1150_U148 ; P1_R1150_U351
g15169 nand P1_R1150_U216 P1_R1150_U147 ; P1_R1150_U352
g15170 nand P1_U3482 P1_R1150_U41 ; P1_R1150_U353
g15171 nand P1_U3084 P1_R1150_U38 ; P1_R1150_U354
g15172 nand P1_U3482 P1_R1150_U41 ; P1_R1150_U355
g15173 nand P1_U3084 P1_R1150_U38 ; P1_R1150_U356
g15174 nand P1_R1150_U356 P1_R1150_U355 ; P1_R1150_U357
g15175 nand P1_U3479 P1_R1150_U39 ; P1_R1150_U358
g15176 nand P1_U3070 P1_R1150_U22 ; P1_R1150_U359
g15177 nand P1_R1150_U223 P1_R1150_U44 ; P1_R1150_U360
g15178 nand P1_R1150_U149 P1_R1150_U210 ; P1_R1150_U361
g15179 nand P1_U3476 P1_R1150_U34 ; P1_R1150_U362
g15180 nand P1_U3071 P1_R1150_U31 ; P1_R1150_U363
g15181 nand P1_R1150_U363 P1_R1150_U362 ; P1_R1150_U364
g15182 nand P1_U3473 P1_R1150_U35 ; P1_R1150_U365
g15183 nand P1_U3067 P1_R1150_U32 ; P1_R1150_U366
g15184 nand P1_R1150_U233 P1_R1150_U45 ; P1_R1150_U367
g15185 nand P1_R1150_U150 P1_R1150_U225 ; P1_R1150_U368
g15186 nand P1_U3470 P1_R1150_U36 ; P1_R1150_U369
g15187 nand P1_U3060 P1_R1150_U33 ; P1_R1150_U370
g15188 nand P1_R1150_U234 P1_R1150_U152 ; P1_R1150_U371
g15189 nand P1_R1150_U200 P1_R1150_U151 ; P1_R1150_U372
g15190 nand P1_U3467 P1_R1150_U30 ; P1_R1150_U373
g15191 nand P1_U3064 P1_R1150_U27 ; P1_R1150_U374
g15192 nand P1_U3467 P1_R1150_U30 ; P1_R1150_U375
g15193 nand P1_U3064 P1_R1150_U27 ; P1_R1150_U376
g15194 nand P1_R1150_U376 P1_R1150_U375 ; P1_R1150_U377
g15195 nand P1_U3464 P1_R1150_U28 ; P1_R1150_U378
g15196 nand P1_U3068 P1_R1150_U23 ; P1_R1150_U379
g15197 nand P1_R1150_U239 P1_R1150_U46 ; P1_R1150_U380
g15198 nand P1_R1150_U153 P1_R1150_U194 ; P1_R1150_U381
g15199 nand P1_U4028 P1_R1150_U155 ; P1_R1150_U382
g15200 nand P1_U3055 P1_R1150_U154 ; P1_R1150_U383
g15201 nand P1_U4028 P1_R1150_U155 ; P1_R1150_U384
g15202 nand P1_U3055 P1_R1150_U154 ; P1_R1150_U385
g15203 nand P1_R1150_U385 P1_R1150_U384 ; P1_R1150_U386
g15204 nand P1_U3054 P1_R1150_U386 P1_R1150_U87 ; P1_R1150_U387
g15205 nand P1_R1150_U12 P1_R1150_U88 P1_U4017 ; P1_R1150_U388
g15206 nand P1_U4017 P1_R1150_U88 ; P1_R1150_U389
g15207 nand P1_U3054 P1_R1150_U87 ; P1_R1150_U390
g15208 not P1_R1150_U131 ; P1_R1150_U391
g15209 nand P1_R1150_U306 P1_R1150_U391 ; P1_R1150_U392
g15210 nand P1_R1150_U131 P1_R1150_U157 ; P1_R1150_U393
g15211 nand P1_U4018 P1_R1150_U86 ; P1_R1150_U394
g15212 nand P1_U3053 P1_R1150_U83 ; P1_R1150_U395
g15213 nand P1_U4018 P1_R1150_U86 ; P1_R1150_U396
g15214 nand P1_U3053 P1_R1150_U83 ; P1_R1150_U397
g15215 nand P1_R1150_U397 P1_R1150_U396 ; P1_R1150_U398
g15216 nand P1_U4019 P1_R1150_U84 ; P1_R1150_U399
g15217 nand P1_U3057 P1_R1150_U47 ; P1_R1150_U400
g15218 nand P1_R1150_U313 P1_R1150_U89 ; P1_R1150_U401
g15219 nand P1_R1150_U158 P1_R1150_U300 ; P1_R1150_U402
g15220 nand P1_U4020 P1_R1150_U82 ; P1_R1150_U403
g15221 nand P1_U3058 P1_R1150_U81 ; P1_R1150_U404
g15222 not P1_R1150_U134 ; P1_R1150_U405
g15223 nand P1_R1150_U296 P1_R1150_U405 ; P1_R1150_U406
g15224 nand P1_R1150_U134 P1_R1150_U159 ; P1_R1150_U407
g15225 nand P1_U4021 P1_R1150_U80 ; P1_R1150_U408
g15226 nand P1_U3065 P1_R1150_U79 ; P1_R1150_U409
g15227 not P1_R1150_U135 ; P1_R1150_U410
g15228 nand P1_R1150_U292 P1_R1150_U410 ; P1_R1150_U411
g15229 nand P1_R1150_U135 P1_R1150_U160 ; P1_R1150_U412
g15230 nand P1_U4022 P1_R1150_U75 ; P1_R1150_U413
g15231 nand P1_U3066 P1_R1150_U73 ; P1_R1150_U414
g15232 nand P1_R1150_U414 P1_R1150_U413 ; P1_R1150_U415
g15233 nand P1_U4023 P1_R1150_U76 ; P1_R1150_U416
g15234 nand P1_U3061 P1_R1150_U48 ; P1_R1150_U417
g15235 nand P1_R1150_U323 P1_R1150_U90 ; P1_R1150_U418
g15236 nand P1_R1150_U161 P1_R1150_U315 ; P1_R1150_U419
g15237 nand P1_U4024 P1_R1150_U77 ; P1_R1150_U420
g15238 nand P1_U3075 P1_R1150_U74 ; P1_R1150_U421
g15239 nand P1_R1150_U324 P1_R1150_U163 ; P1_R1150_U422
g15240 nand P1_R1150_U282 P1_R1150_U162 ; P1_R1150_U423
g15241 nand P1_U4025 P1_R1150_U72 ; P1_R1150_U424
g15242 nand P1_U3076 P1_R1150_U71 ; P1_R1150_U425
g15243 not P1_R1150_U137 ; P1_R1150_U426
g15244 nand P1_R1150_U278 P1_R1150_U426 ; P1_R1150_U427
g15245 nand P1_R1150_U137 P1_R1150_U164 ; P1_R1150_U428
g15246 nand P1_U3461 P1_R1150_U26 ; P1_R1150_U429
g15247 nand P1_U3078 P1_R1150_U165 ; P1_R1150_U430
g15248 not P1_R1150_U138 ; P1_R1150_U431
g15249 nand P1_R1150_U431 P1_R1150_U190 ; P1_R1150_U432
g15250 nand P1_R1150_U138 P1_R1150_U25 ; P1_R1150_U433
g15251 nand P1_U3514 P1_R1150_U70 ; P1_R1150_U434
g15252 nand P1_U3081 P1_R1150_U69 ; P1_R1150_U435
g15253 not P1_R1150_U139 ; P1_R1150_U436
g15254 nand P1_R1150_U274 P1_R1150_U436 ; P1_R1150_U437
g15255 nand P1_R1150_U139 P1_R1150_U166 ; P1_R1150_U438
g15256 nand P1_U3512 P1_R1150_U68 ; P1_R1150_U439
g15257 nand P1_U3082 P1_R1150_U167 ; P1_R1150_U440
g15258 not P1_R1150_U140 ; P1_R1150_U441
g15259 nand P1_R1150_U441 P1_R1150_U270 ; P1_R1150_U442
g15260 nand P1_R1150_U140 P1_R1150_U67 ; P1_R1150_U443
g15261 nand P1_U3509 P1_R1150_U66 ; P1_R1150_U444
g15262 nand P1_U3069 P1_R1150_U65 ; P1_R1150_U445
g15263 not P1_R1150_U141 ; P1_R1150_U446
g15264 nand P1_R1150_U266 P1_R1150_U446 ; P1_R1150_U447
g15265 nand P1_R1150_U141 P1_R1150_U168 ; P1_R1150_U448
g15266 nand P1_U3506 P1_R1150_U61 ; P1_R1150_U449
g15267 nand P1_U3073 P1_R1150_U59 ; P1_R1150_U450
g15268 nand P1_R1150_U450 P1_R1150_U449 ; P1_R1150_U451
g15269 nand P1_U3503 P1_R1150_U62 ; P1_R1150_U452
g15270 nand P1_U3074 P1_R1150_U49 ; P1_R1150_U453
g15271 nand P1_R1150_U334 P1_R1150_U91 ; P1_R1150_U454
g15272 nand P1_R1150_U169 P1_R1150_U326 ; P1_R1150_U455
g15273 nand P1_U3500 P1_R1150_U63 ; P1_R1150_U456
g15274 nand P1_U3079 P1_R1150_U60 ; P1_R1150_U457
g15275 nand P1_R1150_U335 P1_R1150_U171 ; P1_R1150_U458
g15276 nand P1_R1150_U256 P1_R1150_U170 ; P1_R1150_U459
g15277 nand P1_U3497 P1_R1150_U58 ; P1_R1150_U460
g15278 nand P1_U3080 P1_R1150_U57 ; P1_R1150_U461
g15279 not P1_R1150_U143 ; P1_R1150_U462
g15280 nand P1_R1150_U252 P1_R1150_U462 ; P1_R1150_U463
g15281 nand P1_R1150_U143 P1_R1150_U172 ; P1_R1150_U464
g15282 nand P1_U3494 P1_R1150_U56 ; P1_R1150_U465
g15283 nand P1_U3072 P1_R1150_U55 ; P1_R1150_U466
g15284 not P1_R1150_U144 ; P1_R1150_U467
g15285 nand P1_R1150_U248 P1_R1150_U467 ; P1_R1150_U468
g15286 nand P1_R1150_U144 P1_R1150_U173 ; P1_R1150_U469
g15287 nand P1_U3491 P1_R1150_U52 ; P1_R1150_U470
g15288 nand P1_U3063 P1_R1150_U50 ; P1_R1150_U471
g15289 nand P1_R1150_U471 P1_R1150_U470 ; P1_R1150_U472
g15290 nand P1_U3488 P1_R1150_U53 ; P1_R1150_U473
g15291 nand P1_U3062 P1_R1150_U51 ; P1_R1150_U474
g15292 nand P1_R1150_U345 P1_R1150_U92 ; P1_R1150_U475
g15293 nand P1_R1150_U174 P1_R1150_U337 ; P1_R1150_U476
g15294 and P1_R1192_U184 P1_R1192_U201 ; P1_R1192_U6
g15295 and P1_R1192_U203 P1_R1192_U202 ; P1_R1192_U7
g15296 and P1_R1192_U179 P1_R1192_U240 ; P1_R1192_U8
g15297 and P1_R1192_U242 P1_R1192_U241 ; P1_R1192_U9
g15298 and P1_R1192_U259 P1_R1192_U258 ; P1_R1192_U10
g15299 and P1_R1192_U285 P1_R1192_U284 ; P1_R1192_U11
g15300 and P1_R1192_U383 P1_R1192_U382 ; P1_R1192_U12
g15301 nand P1_R1192_U340 P1_R1192_U343 ; P1_R1192_U13
g15302 nand P1_R1192_U329 P1_R1192_U332 ; P1_R1192_U14
g15303 nand P1_R1192_U318 P1_R1192_U321 ; P1_R1192_U15
g15304 nand P1_R1192_U310 P1_R1192_U312 ; P1_R1192_U16
g15305 nand P1_R1192_U156 P1_R1192_U175 P1_R1192_U348 ; P1_R1192_U17
g15306 nand P1_R1192_U236 P1_R1192_U238 ; P1_R1192_U18
g15307 nand P1_R1192_U228 P1_R1192_U231 ; P1_R1192_U19
g15308 nand P1_R1192_U220 P1_R1192_U222 ; P1_R1192_U20
g15309 nand P1_R1192_U25 P1_R1192_U346 ; P1_R1192_U21
g15310 not P1_U3479 ; P1_R1192_U22
g15311 not P1_U3464 ; P1_R1192_U23
g15312 not P1_U3456 ; P1_R1192_U24
g15313 nand P1_U3456 P1_R1192_U93 ; P1_R1192_U25
g15314 not P1_U3078 ; P1_R1192_U26
g15315 not P1_U3467 ; P1_R1192_U27
g15316 not P1_U3068 ; P1_R1192_U28
g15317 nand P1_U3068 P1_R1192_U23 ; P1_R1192_U29
g15318 not P1_U3064 ; P1_R1192_U30
g15319 not P1_U3476 ; P1_R1192_U31
g15320 not P1_U3473 ; P1_R1192_U32
g15321 not P1_U3470 ; P1_R1192_U33
g15322 not P1_U3071 ; P1_R1192_U34
g15323 not P1_U3067 ; P1_R1192_U35
g15324 not P1_U3060 ; P1_R1192_U36
g15325 nand P1_U3060 P1_R1192_U33 ; P1_R1192_U37
g15326 not P1_U3482 ; P1_R1192_U38
g15327 not P1_U3070 ; P1_R1192_U39
g15328 nand P1_U3070 P1_R1192_U22 ; P1_R1192_U40
g15329 not P1_U3084 ; P1_R1192_U41
g15330 not P1_U3485 ; P1_R1192_U42
g15331 not P1_U3083 ; P1_R1192_U43
g15332 nand P1_R1192_U209 P1_R1192_U208 ; P1_R1192_U44
g15333 nand P1_R1192_U37 P1_R1192_U224 ; P1_R1192_U45
g15334 nand P1_R1192_U193 P1_R1192_U192 ; P1_R1192_U46
g15335 not P1_U4019 ; P1_R1192_U47
g15336 not P1_U4023 ; P1_R1192_U48
g15337 not P1_U3503 ; P1_R1192_U49
g15338 not P1_U3491 ; P1_R1192_U50
g15339 not P1_U3488 ; P1_R1192_U51
g15340 not P1_U3063 ; P1_R1192_U52
g15341 not P1_U3062 ; P1_R1192_U53
g15342 nand P1_U3083 P1_R1192_U42 ; P1_R1192_U54
g15343 not P1_U3494 ; P1_R1192_U55
g15344 not P1_U3072 ; P1_R1192_U56
g15345 not P1_U3497 ; P1_R1192_U57
g15346 not P1_U3080 ; P1_R1192_U58
g15347 not P1_U3506 ; P1_R1192_U59
g15348 not P1_U3500 ; P1_R1192_U60
g15349 not P1_U3073 ; P1_R1192_U61
g15350 not P1_U3074 ; P1_R1192_U62
g15351 not P1_U3079 ; P1_R1192_U63
g15352 nand P1_U3079 P1_R1192_U60 ; P1_R1192_U64
g15353 not P1_U3509 ; P1_R1192_U65
g15354 not P1_U3069 ; P1_R1192_U66
g15355 nand P1_R1192_U269 P1_R1192_U268 ; P1_R1192_U67
g15356 not P1_U3082 ; P1_R1192_U68
g15357 not P1_U3514 ; P1_R1192_U69
g15358 not P1_U3081 ; P1_R1192_U70
g15359 not P1_U4025 ; P1_R1192_U71
g15360 not P1_U3076 ; P1_R1192_U72
g15361 not P1_U4022 ; P1_R1192_U73
g15362 not P1_U4024 ; P1_R1192_U74
g15363 not P1_U3066 ; P1_R1192_U75
g15364 not P1_U3061 ; P1_R1192_U76
g15365 not P1_U3075 ; P1_R1192_U77
g15366 nand P1_U3075 P1_R1192_U74 ; P1_R1192_U78
g15367 not P1_U4021 ; P1_R1192_U79
g15368 not P1_U3065 ; P1_R1192_U80
g15369 not P1_U4020 ; P1_R1192_U81
g15370 not P1_U3058 ; P1_R1192_U82
g15371 not P1_U4018 ; P1_R1192_U83
g15372 not P1_U3057 ; P1_R1192_U84
g15373 nand P1_U3057 P1_R1192_U47 ; P1_R1192_U85
g15374 not P1_U3053 ; P1_R1192_U86
g15375 not P1_U4017 ; P1_R1192_U87
g15376 not P1_U3054 ; P1_R1192_U88
g15377 nand P1_R1192_U299 P1_R1192_U298 ; P1_R1192_U89
g15378 nand P1_R1192_U78 P1_R1192_U314 ; P1_R1192_U90
g15379 nand P1_R1192_U64 P1_R1192_U325 ; P1_R1192_U91
g15380 nand P1_R1192_U54 P1_R1192_U336 ; P1_R1192_U92
g15381 not P1_U3077 ; P1_R1192_U93
g15382 nand P1_R1192_U393 P1_R1192_U392 ; P1_R1192_U94
g15383 nand P1_R1192_U407 P1_R1192_U406 ; P1_R1192_U95
g15384 nand P1_R1192_U412 P1_R1192_U411 ; P1_R1192_U96
g15385 nand P1_R1192_U428 P1_R1192_U427 ; P1_R1192_U97
g15386 nand P1_R1192_U433 P1_R1192_U432 ; P1_R1192_U98
g15387 nand P1_R1192_U438 P1_R1192_U437 ; P1_R1192_U99
g15388 nand P1_R1192_U443 P1_R1192_U442 ; P1_R1192_U100
g15389 nand P1_R1192_U448 P1_R1192_U447 ; P1_R1192_U101
g15390 nand P1_R1192_U464 P1_R1192_U463 ; P1_R1192_U102
g15391 nand P1_R1192_U469 P1_R1192_U468 ; P1_R1192_U103
g15392 nand P1_R1192_U352 P1_R1192_U351 ; P1_R1192_U104
g15393 nand P1_R1192_U361 P1_R1192_U360 ; P1_R1192_U105
g15394 nand P1_R1192_U368 P1_R1192_U367 ; P1_R1192_U106
g15395 nand P1_R1192_U372 P1_R1192_U371 ; P1_R1192_U107
g15396 nand P1_R1192_U381 P1_R1192_U380 ; P1_R1192_U108
g15397 nand P1_R1192_U402 P1_R1192_U401 ; P1_R1192_U109
g15398 nand P1_R1192_U419 P1_R1192_U418 ; P1_R1192_U110
g15399 nand P1_R1192_U423 P1_R1192_U422 ; P1_R1192_U111
g15400 nand P1_R1192_U455 P1_R1192_U454 ; P1_R1192_U112
g15401 nand P1_R1192_U459 P1_R1192_U458 ; P1_R1192_U113
g15402 nand P1_R1192_U476 P1_R1192_U475 ; P1_R1192_U114
g15403 and P1_R1192_U195 P1_R1192_U183 ; P1_R1192_U115
g15404 and P1_R1192_U198 P1_R1192_U199 ; P1_R1192_U116
g15405 and P1_R1192_U211 P1_R1192_U185 ; P1_R1192_U117
g15406 and P1_R1192_U214 P1_R1192_U215 ; P1_R1192_U118
g15407 and P1_R1192_U354 P1_R1192_U353 P1_R1192_U40 ; P1_R1192_U119
g15408 and P1_R1192_U357 P1_R1192_U185 ; P1_R1192_U120
g15409 and P1_R1192_U230 P1_R1192_U7 ; P1_R1192_U121
g15410 and P1_R1192_U364 P1_R1192_U184 ; P1_R1192_U122
g15411 and P1_R1192_U374 P1_R1192_U373 P1_R1192_U29 ; P1_R1192_U123
g15412 and P1_R1192_U377 P1_R1192_U183 ; P1_R1192_U124
g15413 and P1_R1192_U217 P1_R1192_U8 ; P1_R1192_U125
g15414 and P1_R1192_U262 P1_R1192_U180 ; P1_R1192_U126
g15415 and P1_R1192_U288 P1_R1192_U181 ; P1_R1192_U127
g15416 and P1_R1192_U304 P1_R1192_U305 ; P1_R1192_U128
g15417 and P1_R1192_U307 P1_R1192_U386 ; P1_R1192_U129
g15418 and P1_R1192_U305 P1_R1192_U304 P1_R1192_U308 ; P1_R1192_U130
g15419 nand P1_R1192_U390 P1_R1192_U389 ; P1_R1192_U131
g15420 and P1_R1192_U395 P1_R1192_U394 P1_R1192_U85 ; P1_R1192_U132
g15421 and P1_R1192_U398 P1_R1192_U182 ; P1_R1192_U133
g15422 nand P1_R1192_U404 P1_R1192_U403 ; P1_R1192_U134
g15423 nand P1_R1192_U409 P1_R1192_U408 ; P1_R1192_U135
g15424 and P1_R1192_U415 P1_R1192_U181 ; P1_R1192_U136
g15425 nand P1_R1192_U425 P1_R1192_U424 ; P1_R1192_U137
g15426 nand P1_R1192_U430 P1_R1192_U429 ; P1_R1192_U138
g15427 nand P1_R1192_U435 P1_R1192_U434 ; P1_R1192_U139
g15428 nand P1_R1192_U440 P1_R1192_U439 ; P1_R1192_U140
g15429 nand P1_R1192_U445 P1_R1192_U444 ; P1_R1192_U141
g15430 and P1_R1192_U451 P1_R1192_U180 ; P1_R1192_U142
g15431 nand P1_R1192_U461 P1_R1192_U460 ; P1_R1192_U143
g15432 nand P1_R1192_U466 P1_R1192_U465 ; P1_R1192_U144
g15433 and P1_R1192_U342 P1_R1192_U9 ; P1_R1192_U145
g15434 and P1_R1192_U472 P1_R1192_U179 ; P1_R1192_U146
g15435 and P1_R1192_U350 P1_R1192_U349 ; P1_R1192_U147
g15436 nand P1_R1192_U118 P1_R1192_U212 ; P1_R1192_U148
g15437 and P1_R1192_U359 P1_R1192_U358 ; P1_R1192_U149
g15438 and P1_R1192_U366 P1_R1192_U365 ; P1_R1192_U150
g15439 and P1_R1192_U370 P1_R1192_U369 ; P1_R1192_U151
g15440 nand P1_R1192_U116 P1_R1192_U196 ; P1_R1192_U152
g15441 and P1_R1192_U379 P1_R1192_U378 ; P1_R1192_U153
g15442 not P1_U4028 ; P1_R1192_U154
g15443 not P1_U3055 ; P1_R1192_U155
g15444 and P1_R1192_U388 P1_R1192_U387 ; P1_R1192_U156
g15445 nand P1_R1192_U128 P1_R1192_U302 ; P1_R1192_U157
g15446 and P1_R1192_U400 P1_R1192_U399 ; P1_R1192_U158
g15447 nand P1_R1192_U295 P1_R1192_U294 ; P1_R1192_U159
g15448 nand P1_R1192_U291 P1_R1192_U290 ; P1_R1192_U160
g15449 and P1_R1192_U417 P1_R1192_U416 ; P1_R1192_U161
g15450 and P1_R1192_U421 P1_R1192_U420 ; P1_R1192_U162
g15451 nand P1_R1192_U281 P1_R1192_U280 ; P1_R1192_U163
g15452 nand P1_R1192_U277 P1_R1192_U276 ; P1_R1192_U164
g15453 not P1_U3461 ; P1_R1192_U165
g15454 nand P1_R1192_U273 P1_R1192_U272 ; P1_R1192_U166
g15455 not P1_U3512 ; P1_R1192_U167
g15456 nand P1_R1192_U265 P1_R1192_U264 ; P1_R1192_U168
g15457 and P1_R1192_U453 P1_R1192_U452 ; P1_R1192_U169
g15458 and P1_R1192_U457 P1_R1192_U456 ; P1_R1192_U170
g15459 nand P1_R1192_U255 P1_R1192_U254 ; P1_R1192_U171
g15460 nand P1_R1192_U251 P1_R1192_U250 ; P1_R1192_U172
g15461 nand P1_R1192_U247 P1_R1192_U246 ; P1_R1192_U173
g15462 and P1_R1192_U474 P1_R1192_U473 ; P1_R1192_U174
g15463 nand P1_R1192_U129 P1_R1192_U157 ; P1_R1192_U175
g15464 not P1_R1192_U85 ; P1_R1192_U176
g15465 not P1_R1192_U29 ; P1_R1192_U177
g15466 not P1_R1192_U40 ; P1_R1192_U178
g15467 nand P1_U3488 P1_R1192_U53 ; P1_R1192_U179
g15468 nand P1_U3503 P1_R1192_U62 ; P1_R1192_U180
g15469 nand P1_U4023 P1_R1192_U76 ; P1_R1192_U181
g15470 nand P1_U4019 P1_R1192_U84 ; P1_R1192_U182
g15471 nand P1_U3464 P1_R1192_U28 ; P1_R1192_U183
g15472 nand P1_U3473 P1_R1192_U35 ; P1_R1192_U184
g15473 nand P1_U3479 P1_R1192_U39 ; P1_R1192_U185
g15474 not P1_R1192_U64 ; P1_R1192_U186
g15475 not P1_R1192_U78 ; P1_R1192_U187
g15476 not P1_R1192_U37 ; P1_R1192_U188
g15477 not P1_R1192_U54 ; P1_R1192_U189
g15478 not P1_R1192_U25 ; P1_R1192_U190
g15479 nand P1_R1192_U190 P1_R1192_U26 ; P1_R1192_U191
g15480 nand P1_R1192_U191 P1_R1192_U165 ; P1_R1192_U192
g15481 nand P1_U3078 P1_R1192_U25 ; P1_R1192_U193
g15482 not P1_R1192_U46 ; P1_R1192_U194
g15483 nand P1_U3467 P1_R1192_U30 ; P1_R1192_U195
g15484 nand P1_R1192_U115 P1_R1192_U46 ; P1_R1192_U196
g15485 nand P1_R1192_U30 P1_R1192_U29 ; P1_R1192_U197
g15486 nand P1_R1192_U197 P1_R1192_U27 ; P1_R1192_U198
g15487 nand P1_U3064 P1_R1192_U177 ; P1_R1192_U199
g15488 not P1_R1192_U152 ; P1_R1192_U200
g15489 nand P1_U3476 P1_R1192_U34 ; P1_R1192_U201
g15490 nand P1_U3071 P1_R1192_U31 ; P1_R1192_U202
g15491 nand P1_U3067 P1_R1192_U32 ; P1_R1192_U203
g15492 nand P1_R1192_U188 P1_R1192_U6 ; P1_R1192_U204
g15493 nand P1_R1192_U7 P1_R1192_U204 ; P1_R1192_U205
g15494 nand P1_U3470 P1_R1192_U36 ; P1_R1192_U206
g15495 nand P1_U3476 P1_R1192_U34 ; P1_R1192_U207
g15496 nand P1_R1192_U206 P1_R1192_U152 P1_R1192_U6 ; P1_R1192_U208
g15497 nand P1_R1192_U207 P1_R1192_U205 ; P1_R1192_U209
g15498 not P1_R1192_U44 ; P1_R1192_U210
g15499 nand P1_U3482 P1_R1192_U41 ; P1_R1192_U211
g15500 nand P1_R1192_U117 P1_R1192_U44 ; P1_R1192_U212
g15501 nand P1_R1192_U41 P1_R1192_U40 ; P1_R1192_U213
g15502 nand P1_R1192_U213 P1_R1192_U38 ; P1_R1192_U214
g15503 nand P1_U3084 P1_R1192_U178 ; P1_R1192_U215
g15504 not P1_R1192_U148 ; P1_R1192_U216
g15505 nand P1_U3485 P1_R1192_U43 ; P1_R1192_U217
g15506 nand P1_R1192_U217 P1_R1192_U54 ; P1_R1192_U218
g15507 nand P1_R1192_U210 P1_R1192_U40 ; P1_R1192_U219
g15508 nand P1_R1192_U120 P1_R1192_U219 ; P1_R1192_U220
g15509 nand P1_R1192_U44 P1_R1192_U185 ; P1_R1192_U221
g15510 nand P1_R1192_U119 P1_R1192_U221 ; P1_R1192_U222
g15511 nand P1_R1192_U40 P1_R1192_U185 ; P1_R1192_U223
g15512 nand P1_R1192_U206 P1_R1192_U152 ; P1_R1192_U224
g15513 not P1_R1192_U45 ; P1_R1192_U225
g15514 nand P1_U3067 P1_R1192_U32 ; P1_R1192_U226
g15515 nand P1_R1192_U225 P1_R1192_U226 ; P1_R1192_U227
g15516 nand P1_R1192_U122 P1_R1192_U227 ; P1_R1192_U228
g15517 nand P1_R1192_U45 P1_R1192_U184 ; P1_R1192_U229
g15518 nand P1_U3476 P1_R1192_U34 ; P1_R1192_U230
g15519 nand P1_R1192_U121 P1_R1192_U229 ; P1_R1192_U231
g15520 nand P1_U3067 P1_R1192_U32 ; P1_R1192_U232
g15521 nand P1_R1192_U184 P1_R1192_U232 ; P1_R1192_U233
g15522 nand P1_R1192_U206 P1_R1192_U37 ; P1_R1192_U234
g15523 nand P1_R1192_U194 P1_R1192_U29 ; P1_R1192_U235
g15524 nand P1_R1192_U124 P1_R1192_U235 ; P1_R1192_U236
g15525 nand P1_R1192_U46 P1_R1192_U183 ; P1_R1192_U237
g15526 nand P1_R1192_U123 P1_R1192_U237 ; P1_R1192_U238
g15527 nand P1_R1192_U29 P1_R1192_U183 ; P1_R1192_U239
g15528 nand P1_U3491 P1_R1192_U52 ; P1_R1192_U240
g15529 nand P1_U3063 P1_R1192_U50 ; P1_R1192_U241
g15530 nand P1_U3062 P1_R1192_U51 ; P1_R1192_U242
g15531 nand P1_R1192_U189 P1_R1192_U8 ; P1_R1192_U243
g15532 nand P1_R1192_U9 P1_R1192_U243 ; P1_R1192_U244
g15533 nand P1_U3491 P1_R1192_U52 ; P1_R1192_U245
g15534 nand P1_R1192_U125 P1_R1192_U148 ; P1_R1192_U246
g15535 nand P1_R1192_U245 P1_R1192_U244 ; P1_R1192_U247
g15536 not P1_R1192_U173 ; P1_R1192_U248
g15537 nand P1_U3494 P1_R1192_U56 ; P1_R1192_U249
g15538 nand P1_R1192_U249 P1_R1192_U173 ; P1_R1192_U250
g15539 nand P1_U3072 P1_R1192_U55 ; P1_R1192_U251
g15540 not P1_R1192_U172 ; P1_R1192_U252
g15541 nand P1_U3497 P1_R1192_U58 ; P1_R1192_U253
g15542 nand P1_R1192_U253 P1_R1192_U172 ; P1_R1192_U254
g15543 nand P1_U3080 P1_R1192_U57 ; P1_R1192_U255
g15544 not P1_R1192_U171 ; P1_R1192_U256
g15545 nand P1_U3506 P1_R1192_U61 ; P1_R1192_U257
g15546 nand P1_U3073 P1_R1192_U59 ; P1_R1192_U258
g15547 nand P1_U3074 P1_R1192_U49 ; P1_R1192_U259
g15548 nand P1_R1192_U186 P1_R1192_U180 ; P1_R1192_U260
g15549 nand P1_R1192_U10 P1_R1192_U260 ; P1_R1192_U261
g15550 nand P1_U3500 P1_R1192_U63 ; P1_R1192_U262
g15551 nand P1_U3506 P1_R1192_U61 ; P1_R1192_U263
g15552 nand P1_R1192_U171 P1_R1192_U126 P1_R1192_U257 ; P1_R1192_U264
g15553 nand P1_R1192_U263 P1_R1192_U261 ; P1_R1192_U265
g15554 not P1_R1192_U168 ; P1_R1192_U266
g15555 nand P1_U3509 P1_R1192_U66 ; P1_R1192_U267
g15556 nand P1_R1192_U267 P1_R1192_U168 ; P1_R1192_U268
g15557 nand P1_U3069 P1_R1192_U65 ; P1_R1192_U269
g15558 not P1_R1192_U67 ; P1_R1192_U270
g15559 nand P1_R1192_U270 P1_R1192_U68 ; P1_R1192_U271
g15560 nand P1_R1192_U271 P1_R1192_U167 ; P1_R1192_U272
g15561 nand P1_U3082 P1_R1192_U67 ; P1_R1192_U273
g15562 not P1_R1192_U166 ; P1_R1192_U274
g15563 nand P1_U3514 P1_R1192_U70 ; P1_R1192_U275
g15564 nand P1_R1192_U275 P1_R1192_U166 ; P1_R1192_U276
g15565 nand P1_U3081 P1_R1192_U69 ; P1_R1192_U277
g15566 not P1_R1192_U164 ; P1_R1192_U278
g15567 nand P1_U4025 P1_R1192_U72 ; P1_R1192_U279
g15568 nand P1_R1192_U279 P1_R1192_U164 ; P1_R1192_U280
g15569 nand P1_U3076 P1_R1192_U71 ; P1_R1192_U281
g15570 not P1_R1192_U163 ; P1_R1192_U282
g15571 nand P1_U4022 P1_R1192_U75 ; P1_R1192_U283
g15572 nand P1_U3066 P1_R1192_U73 ; P1_R1192_U284
g15573 nand P1_U3061 P1_R1192_U48 ; P1_R1192_U285
g15574 nand P1_R1192_U187 P1_R1192_U181 ; P1_R1192_U286
g15575 nand P1_R1192_U11 P1_R1192_U286 ; P1_R1192_U287
g15576 nand P1_U4024 P1_R1192_U77 ; P1_R1192_U288
g15577 nand P1_U4022 P1_R1192_U75 ; P1_R1192_U289
g15578 nand P1_R1192_U163 P1_R1192_U127 P1_R1192_U283 ; P1_R1192_U290
g15579 nand P1_R1192_U289 P1_R1192_U287 ; P1_R1192_U291
g15580 not P1_R1192_U160 ; P1_R1192_U292
g15581 nand P1_U4021 P1_R1192_U80 ; P1_R1192_U293
g15582 nand P1_R1192_U293 P1_R1192_U160 ; P1_R1192_U294
g15583 nand P1_U3065 P1_R1192_U79 ; P1_R1192_U295
g15584 not P1_R1192_U159 ; P1_R1192_U296
g15585 nand P1_U4020 P1_R1192_U82 ; P1_R1192_U297
g15586 nand P1_R1192_U297 P1_R1192_U159 ; P1_R1192_U298
g15587 nand P1_U3058 P1_R1192_U81 ; P1_R1192_U299
g15588 not P1_R1192_U89 ; P1_R1192_U300
g15589 nand P1_U4018 P1_R1192_U86 ; P1_R1192_U301
g15590 nand P1_R1192_U89 P1_R1192_U182 P1_R1192_U301 ; P1_R1192_U302
g15591 nand P1_R1192_U86 P1_R1192_U85 ; P1_R1192_U303
g15592 nand P1_R1192_U303 P1_R1192_U83 ; P1_R1192_U304
g15593 nand P1_U3053 P1_R1192_U176 ; P1_R1192_U305
g15594 not P1_R1192_U157 ; P1_R1192_U306
g15595 nand P1_U4017 P1_R1192_U88 ; P1_R1192_U307
g15596 nand P1_U3054 P1_R1192_U87 ; P1_R1192_U308
g15597 nand P1_R1192_U300 P1_R1192_U85 ; P1_R1192_U309
g15598 nand P1_R1192_U133 P1_R1192_U309 ; P1_R1192_U310
g15599 nand P1_R1192_U89 P1_R1192_U182 ; P1_R1192_U311
g15600 nand P1_R1192_U132 P1_R1192_U311 ; P1_R1192_U312
g15601 nand P1_R1192_U85 P1_R1192_U182 ; P1_R1192_U313
g15602 nand P1_R1192_U288 P1_R1192_U163 ; P1_R1192_U314
g15603 not P1_R1192_U90 ; P1_R1192_U315
g15604 nand P1_U3061 P1_R1192_U48 ; P1_R1192_U316
g15605 nand P1_R1192_U315 P1_R1192_U316 ; P1_R1192_U317
g15606 nand P1_R1192_U136 P1_R1192_U317 ; P1_R1192_U318
g15607 nand P1_R1192_U90 P1_R1192_U181 ; P1_R1192_U319
g15608 nand P1_U4022 P1_R1192_U75 ; P1_R1192_U320
g15609 nand P1_R1192_U320 P1_R1192_U319 P1_R1192_U11 ; P1_R1192_U321
g15610 nand P1_U3061 P1_R1192_U48 ; P1_R1192_U322
g15611 nand P1_R1192_U181 P1_R1192_U322 ; P1_R1192_U323
g15612 nand P1_R1192_U288 P1_R1192_U78 ; P1_R1192_U324
g15613 nand P1_R1192_U262 P1_R1192_U171 ; P1_R1192_U325
g15614 not P1_R1192_U91 ; P1_R1192_U326
g15615 nand P1_U3074 P1_R1192_U49 ; P1_R1192_U327
g15616 nand P1_R1192_U326 P1_R1192_U327 ; P1_R1192_U328
g15617 nand P1_R1192_U142 P1_R1192_U328 ; P1_R1192_U329
g15618 nand P1_R1192_U91 P1_R1192_U180 ; P1_R1192_U330
g15619 nand P1_U3506 P1_R1192_U61 ; P1_R1192_U331
g15620 nand P1_R1192_U331 P1_R1192_U330 P1_R1192_U10 ; P1_R1192_U332
g15621 nand P1_U3074 P1_R1192_U49 ; P1_R1192_U333
g15622 nand P1_R1192_U180 P1_R1192_U333 ; P1_R1192_U334
g15623 nand P1_R1192_U262 P1_R1192_U64 ; P1_R1192_U335
g15624 nand P1_R1192_U217 P1_R1192_U148 ; P1_R1192_U336
g15625 not P1_R1192_U92 ; P1_R1192_U337
g15626 nand P1_U3062 P1_R1192_U51 ; P1_R1192_U338
g15627 nand P1_R1192_U337 P1_R1192_U338 ; P1_R1192_U339
g15628 nand P1_R1192_U146 P1_R1192_U339 ; P1_R1192_U340
g15629 nand P1_R1192_U92 P1_R1192_U179 ; P1_R1192_U341
g15630 nand P1_U3491 P1_R1192_U52 ; P1_R1192_U342
g15631 nand P1_R1192_U145 P1_R1192_U341 ; P1_R1192_U343
g15632 nand P1_U3062 P1_R1192_U51 ; P1_R1192_U344
g15633 nand P1_R1192_U179 P1_R1192_U344 ; P1_R1192_U345
g15634 nand P1_U3077 P1_R1192_U24 ; P1_R1192_U346
g15635 nand P1_R1192_U89 P1_R1192_U182 P1_R1192_U301 ; P1_R1192_U347
g15636 nand P1_R1192_U12 P1_R1192_U347 P1_R1192_U130 ; P1_R1192_U348
g15637 nand P1_U3485 P1_R1192_U43 ; P1_R1192_U349
g15638 nand P1_U3083 P1_R1192_U42 ; P1_R1192_U350
g15639 nand P1_R1192_U218 P1_R1192_U148 ; P1_R1192_U351
g15640 nand P1_R1192_U216 P1_R1192_U147 ; P1_R1192_U352
g15641 nand P1_U3482 P1_R1192_U41 ; P1_R1192_U353
g15642 nand P1_U3084 P1_R1192_U38 ; P1_R1192_U354
g15643 nand P1_U3482 P1_R1192_U41 ; P1_R1192_U355
g15644 nand P1_U3084 P1_R1192_U38 ; P1_R1192_U356
g15645 nand P1_R1192_U356 P1_R1192_U355 ; P1_R1192_U357
g15646 nand P1_U3479 P1_R1192_U39 ; P1_R1192_U358
g15647 nand P1_U3070 P1_R1192_U22 ; P1_R1192_U359
g15648 nand P1_R1192_U223 P1_R1192_U44 ; P1_R1192_U360
g15649 nand P1_R1192_U149 P1_R1192_U210 ; P1_R1192_U361
g15650 nand P1_U3476 P1_R1192_U34 ; P1_R1192_U362
g15651 nand P1_U3071 P1_R1192_U31 ; P1_R1192_U363
g15652 nand P1_R1192_U363 P1_R1192_U362 ; P1_R1192_U364
g15653 nand P1_U3473 P1_R1192_U35 ; P1_R1192_U365
g15654 nand P1_U3067 P1_R1192_U32 ; P1_R1192_U366
g15655 nand P1_R1192_U233 P1_R1192_U45 ; P1_R1192_U367
g15656 nand P1_R1192_U150 P1_R1192_U225 ; P1_R1192_U368
g15657 nand P1_U3470 P1_R1192_U36 ; P1_R1192_U369
g15658 nand P1_U3060 P1_R1192_U33 ; P1_R1192_U370
g15659 nand P1_R1192_U234 P1_R1192_U152 ; P1_R1192_U371
g15660 nand P1_R1192_U200 P1_R1192_U151 ; P1_R1192_U372
g15661 nand P1_U3467 P1_R1192_U30 ; P1_R1192_U373
g15662 nand P1_U3064 P1_R1192_U27 ; P1_R1192_U374
g15663 nand P1_U3467 P1_R1192_U30 ; P1_R1192_U375
g15664 nand P1_U3064 P1_R1192_U27 ; P1_R1192_U376
g15665 nand P1_R1192_U376 P1_R1192_U375 ; P1_R1192_U377
g15666 nand P1_U3464 P1_R1192_U28 ; P1_R1192_U378
g15667 nand P1_U3068 P1_R1192_U23 ; P1_R1192_U379
g15668 nand P1_R1192_U239 P1_R1192_U46 ; P1_R1192_U380
g15669 nand P1_R1192_U153 P1_R1192_U194 ; P1_R1192_U381
g15670 nand P1_U4028 P1_R1192_U155 ; P1_R1192_U382
g15671 nand P1_U3055 P1_R1192_U154 ; P1_R1192_U383
g15672 nand P1_U4028 P1_R1192_U155 ; P1_R1192_U384
g15673 nand P1_U3055 P1_R1192_U154 ; P1_R1192_U385
g15674 nand P1_R1192_U385 P1_R1192_U384 ; P1_R1192_U386
g15675 nand P1_U3054 P1_R1192_U386 P1_R1192_U87 ; P1_R1192_U387
g15676 nand P1_R1192_U12 P1_R1192_U88 P1_U4017 ; P1_R1192_U388
g15677 nand P1_U4017 P1_R1192_U88 ; P1_R1192_U389
g15678 nand P1_U3054 P1_R1192_U87 ; P1_R1192_U390
g15679 not P1_R1192_U131 ; P1_R1192_U391
g15680 nand P1_R1192_U306 P1_R1192_U391 ; P1_R1192_U392
g15681 nand P1_R1192_U131 P1_R1192_U157 ; P1_R1192_U393
g15682 nand P1_U4018 P1_R1192_U86 ; P1_R1192_U394
g15683 nand P1_U3053 P1_R1192_U83 ; P1_R1192_U395
g15684 nand P1_U4018 P1_R1192_U86 ; P1_R1192_U396
g15685 nand P1_U3053 P1_R1192_U83 ; P1_R1192_U397
g15686 nand P1_R1192_U397 P1_R1192_U396 ; P1_R1192_U398
g15687 nand P1_U4019 P1_R1192_U84 ; P1_R1192_U399
g15688 nand P1_U3057 P1_R1192_U47 ; P1_R1192_U400
g15689 nand P1_R1192_U313 P1_R1192_U89 ; P1_R1192_U401
g15690 nand P1_R1192_U158 P1_R1192_U300 ; P1_R1192_U402
g15691 nand P1_U4020 P1_R1192_U82 ; P1_R1192_U403
g15692 nand P1_U3058 P1_R1192_U81 ; P1_R1192_U404
g15693 not P1_R1192_U134 ; P1_R1192_U405
g15694 nand P1_R1192_U296 P1_R1192_U405 ; P1_R1192_U406
g15695 nand P1_R1192_U134 P1_R1192_U159 ; P1_R1192_U407
g15696 nand P1_U4021 P1_R1192_U80 ; P1_R1192_U408
g15697 nand P1_U3065 P1_R1192_U79 ; P1_R1192_U409
g15698 not P1_R1192_U135 ; P1_R1192_U410
g15699 nand P1_R1192_U292 P1_R1192_U410 ; P1_R1192_U411
g15700 nand P1_R1192_U135 P1_R1192_U160 ; P1_R1192_U412
g15701 nand P1_U4022 P1_R1192_U75 ; P1_R1192_U413
g15702 nand P1_U3066 P1_R1192_U73 ; P1_R1192_U414
g15703 nand P1_R1192_U414 P1_R1192_U413 ; P1_R1192_U415
g15704 nand P1_U4023 P1_R1192_U76 ; P1_R1192_U416
g15705 nand P1_U3061 P1_R1192_U48 ; P1_R1192_U417
g15706 nand P1_R1192_U323 P1_R1192_U90 ; P1_R1192_U418
g15707 nand P1_R1192_U161 P1_R1192_U315 ; P1_R1192_U419
g15708 nand P1_U4024 P1_R1192_U77 ; P1_R1192_U420
g15709 nand P1_U3075 P1_R1192_U74 ; P1_R1192_U421
g15710 nand P1_R1192_U324 P1_R1192_U163 ; P1_R1192_U422
g15711 nand P1_R1192_U282 P1_R1192_U162 ; P1_R1192_U423
g15712 nand P1_U4025 P1_R1192_U72 ; P1_R1192_U424
g15713 nand P1_U3076 P1_R1192_U71 ; P1_R1192_U425
g15714 not P1_R1192_U137 ; P1_R1192_U426
g15715 nand P1_R1192_U278 P1_R1192_U426 ; P1_R1192_U427
g15716 nand P1_R1192_U137 P1_R1192_U164 ; P1_R1192_U428
g15717 nand P1_U3461 P1_R1192_U26 ; P1_R1192_U429
g15718 nand P1_U3078 P1_R1192_U165 ; P1_R1192_U430
g15719 not P1_R1192_U138 ; P1_R1192_U431
g15720 nand P1_R1192_U431 P1_R1192_U190 ; P1_R1192_U432
g15721 nand P1_R1192_U138 P1_R1192_U25 ; P1_R1192_U433
g15722 nand P1_U3514 P1_R1192_U70 ; P1_R1192_U434
g15723 nand P1_U3081 P1_R1192_U69 ; P1_R1192_U435
g15724 not P1_R1192_U139 ; P1_R1192_U436
g15725 nand P1_R1192_U274 P1_R1192_U436 ; P1_R1192_U437
g15726 nand P1_R1192_U139 P1_R1192_U166 ; P1_R1192_U438
g15727 nand P1_U3512 P1_R1192_U68 ; P1_R1192_U439
g15728 nand P1_U3082 P1_R1192_U167 ; P1_R1192_U440
g15729 not P1_R1192_U140 ; P1_R1192_U441
g15730 nand P1_R1192_U441 P1_R1192_U270 ; P1_R1192_U442
g15731 nand P1_R1192_U140 P1_R1192_U67 ; P1_R1192_U443
g15732 nand P1_U3509 P1_R1192_U66 ; P1_R1192_U444
g15733 nand P1_U3069 P1_R1192_U65 ; P1_R1192_U445
g15734 not P1_R1192_U141 ; P1_R1192_U446
g15735 nand P1_R1192_U266 P1_R1192_U446 ; P1_R1192_U447
g15736 nand P1_R1192_U141 P1_R1192_U168 ; P1_R1192_U448
g15737 nand P1_U3506 P1_R1192_U61 ; P1_R1192_U449
g15738 nand P1_U3073 P1_R1192_U59 ; P1_R1192_U450
g15739 nand P1_R1192_U450 P1_R1192_U449 ; P1_R1192_U451
g15740 nand P1_U3503 P1_R1192_U62 ; P1_R1192_U452
g15741 nand P1_U3074 P1_R1192_U49 ; P1_R1192_U453
g15742 nand P1_R1192_U334 P1_R1192_U91 ; P1_R1192_U454
g15743 nand P1_R1192_U169 P1_R1192_U326 ; P1_R1192_U455
g15744 nand P1_U3500 P1_R1192_U63 ; P1_R1192_U456
g15745 nand P1_U3079 P1_R1192_U60 ; P1_R1192_U457
g15746 nand P1_R1192_U335 P1_R1192_U171 ; P1_R1192_U458
g15747 nand P1_R1192_U256 P1_R1192_U170 ; P1_R1192_U459
g15748 nand P1_U3497 P1_R1192_U58 ; P1_R1192_U460
g15749 nand P1_U3080 P1_R1192_U57 ; P1_R1192_U461
g15750 not P1_R1192_U143 ; P1_R1192_U462
g15751 nand P1_R1192_U252 P1_R1192_U462 ; P1_R1192_U463
g15752 nand P1_R1192_U143 P1_R1192_U172 ; P1_R1192_U464
g15753 nand P1_U3494 P1_R1192_U56 ; P1_R1192_U465
g15754 nand P1_U3072 P1_R1192_U55 ; P1_R1192_U466
g15755 not P1_R1192_U144 ; P1_R1192_U467
g15756 nand P1_R1192_U248 P1_R1192_U467 ; P1_R1192_U468
g15757 nand P1_R1192_U144 P1_R1192_U173 ; P1_R1192_U469
g15758 nand P1_U3491 P1_R1192_U52 ; P1_R1192_U470
g15759 nand P1_U3063 P1_R1192_U50 ; P1_R1192_U471
g15760 nand P1_R1192_U471 P1_R1192_U470 ; P1_R1192_U472
g15761 nand P1_U3488 P1_R1192_U53 ; P1_R1192_U473
g15762 nand P1_U3062 P1_R1192_U51 ; P1_R1192_U474
g15763 nand P1_R1192_U345 P1_R1192_U92 ; P1_R1192_U475
g15764 nand P1_R1192_U174 P1_R1192_U337 ; P1_R1192_U476
g15765 and P1_R1171_U176 P1_R1171_U175 ; P1_R1171_U4
g15766 and P1_R1171_U177 P1_R1171_U178 ; P1_R1171_U5
g15767 and P1_R1171_U194 P1_R1171_U193 ; P1_R1171_U6
g15768 and P1_R1171_U234 P1_R1171_U233 ; P1_R1171_U7
g15769 and P1_R1171_U243 P1_R1171_U242 ; P1_R1171_U8
g15770 and P1_R1171_U261 P1_R1171_U260 ; P1_R1171_U9
g15771 and P1_R1171_U269 P1_R1171_U268 ; P1_R1171_U10
g15772 and P1_R1171_U348 P1_R1171_U345 ; P1_R1171_U11
g15773 and P1_R1171_U341 P1_R1171_U338 ; P1_R1171_U12
g15774 and P1_R1171_U332 P1_R1171_U329 ; P1_R1171_U13
g15775 and P1_R1171_U323 P1_R1171_U320 ; P1_R1171_U14
g15776 and P1_R1171_U317 P1_R1171_U315 ; P1_R1171_U15
g15777 and P1_R1171_U310 P1_R1171_U307 ; P1_R1171_U16
g15778 and P1_R1171_U232 P1_R1171_U229 ; P1_R1171_U17
g15779 and P1_R1171_U224 P1_R1171_U221 ; P1_R1171_U18
g15780 and P1_R1171_U210 P1_R1171_U207 ; P1_R1171_U19
g15781 not P1_U3476 ; P1_R1171_U20
g15782 not P1_U3071 ; P1_R1171_U21
g15783 not P1_U3070 ; P1_R1171_U22
g15784 nand P1_U3071 P1_U3476 ; P1_R1171_U23
g15785 not P1_U3479 ; P1_R1171_U24
g15786 not P1_U3470 ; P1_R1171_U25
g15787 not P1_U3060 ; P1_R1171_U26
g15788 not P1_U3067 ; P1_R1171_U27
g15789 not P1_U3464 ; P1_R1171_U28
g15790 not P1_U3068 ; P1_R1171_U29
g15791 not P1_U3456 ; P1_R1171_U30
g15792 not P1_U3077 ; P1_R1171_U31
g15793 nand P1_U3077 P1_U3456 ; P1_R1171_U32
g15794 not P1_U3467 ; P1_R1171_U33
g15795 not P1_U3064 ; P1_R1171_U34
g15796 nand P1_U3060 P1_U3470 ; P1_R1171_U35
g15797 not P1_U3473 ; P1_R1171_U36
g15798 not P1_U3482 ; P1_R1171_U37
g15799 not P1_U3084 ; P1_R1171_U38
g15800 not P1_U3083 ; P1_R1171_U39
g15801 not P1_U3485 ; P1_R1171_U40
g15802 nand P1_R1171_U62 P1_R1171_U202 ; P1_R1171_U41
g15803 nand P1_R1171_U118 P1_R1171_U190 ; P1_R1171_U42
g15804 nand P1_R1171_U179 P1_R1171_U180 ; P1_R1171_U43
g15805 nand P1_U3461 P1_U3078 ; P1_R1171_U44
g15806 nand P1_R1171_U122 P1_R1171_U216 ; P1_R1171_U45
g15807 nand P1_R1171_U213 P1_R1171_U212 ; P1_R1171_U46
g15808 not P1_U4018 ; P1_R1171_U47
g15809 not P1_U3053 ; P1_R1171_U48
g15810 not P1_U3057 ; P1_R1171_U49
g15811 not P1_U4019 ; P1_R1171_U50
g15812 not P1_U4020 ; P1_R1171_U51
g15813 not P1_U3058 ; P1_R1171_U52
g15814 not P1_U4021 ; P1_R1171_U53
g15815 not P1_U3065 ; P1_R1171_U54
g15816 not P1_U4024 ; P1_R1171_U55
g15817 not P1_U3075 ; P1_R1171_U56
g15818 not P1_U3506 ; P1_R1171_U57
g15819 not P1_U3073 ; P1_R1171_U58
g15820 not P1_U3069 ; P1_R1171_U59
g15821 nand P1_U3073 P1_U3506 ; P1_R1171_U60
g15822 not P1_U3509 ; P1_R1171_U61
g15823 nand P1_U3084 P1_U3482 ; P1_R1171_U62
g15824 not P1_U3488 ; P1_R1171_U63
g15825 not P1_U3062 ; P1_R1171_U64
g15826 not P1_U3494 ; P1_R1171_U65
g15827 not P1_U3072 ; P1_R1171_U66
g15828 not P1_U3491 ; P1_R1171_U67
g15829 not P1_U3063 ; P1_R1171_U68
g15830 nand P1_U3063 P1_U3491 ; P1_R1171_U69
g15831 not P1_U3497 ; P1_R1171_U70
g15832 not P1_U3080 ; P1_R1171_U71
g15833 not P1_U3500 ; P1_R1171_U72
g15834 not P1_U3079 ; P1_R1171_U73
g15835 not P1_U3503 ; P1_R1171_U74
g15836 not P1_U3074 ; P1_R1171_U75
g15837 not P1_U3512 ; P1_R1171_U76
g15838 not P1_U3082 ; P1_R1171_U77
g15839 nand P1_U3082 P1_U3512 ; P1_R1171_U78
g15840 not P1_U3514 ; P1_R1171_U79
g15841 not P1_U3081 ; P1_R1171_U80
g15842 nand P1_U3081 P1_U3514 ; P1_R1171_U81
g15843 not P1_U4025 ; P1_R1171_U82
g15844 not P1_U4023 ; P1_R1171_U83
g15845 not P1_U3061 ; P1_R1171_U84
g15846 not P1_U4022 ; P1_R1171_U85
g15847 not P1_U3066 ; P1_R1171_U86
g15848 nand P1_U4019 P1_U3057 ; P1_R1171_U87
g15849 not P1_U3054 ; P1_R1171_U88
g15850 not P1_U4017 ; P1_R1171_U89
g15851 nand P1_R1171_U303 P1_R1171_U173 ; P1_R1171_U90
g15852 not P1_U3076 ; P1_R1171_U91
g15853 nand P1_R1171_U78 P1_R1171_U312 ; P1_R1171_U92
g15854 nand P1_R1171_U258 P1_R1171_U257 ; P1_R1171_U93
g15855 nand P1_R1171_U69 P1_R1171_U334 ; P1_R1171_U94
g15856 nand P1_R1171_U454 P1_R1171_U453 ; P1_R1171_U95
g15857 nand P1_R1171_U501 P1_R1171_U500 ; P1_R1171_U96
g15858 nand P1_R1171_U372 P1_R1171_U371 ; P1_R1171_U97
g15859 nand P1_R1171_U377 P1_R1171_U376 ; P1_R1171_U98
g15860 nand P1_R1171_U384 P1_R1171_U383 ; P1_R1171_U99
g15861 nand P1_R1171_U391 P1_R1171_U390 ; P1_R1171_U100
g15862 nand P1_R1171_U396 P1_R1171_U395 ; P1_R1171_U101
g15863 nand P1_R1171_U405 P1_R1171_U404 ; P1_R1171_U102
g15864 nand P1_R1171_U412 P1_R1171_U411 ; P1_R1171_U103
g15865 nand P1_R1171_U419 P1_R1171_U418 ; P1_R1171_U104
g15866 nand P1_R1171_U426 P1_R1171_U425 ; P1_R1171_U105
g15867 nand P1_R1171_U431 P1_R1171_U430 ; P1_R1171_U106
g15868 nand P1_R1171_U438 P1_R1171_U437 ; P1_R1171_U107
g15869 nand P1_R1171_U445 P1_R1171_U444 ; P1_R1171_U108
g15870 nand P1_R1171_U459 P1_R1171_U458 ; P1_R1171_U109
g15871 nand P1_R1171_U464 P1_R1171_U463 ; P1_R1171_U110
g15872 nand P1_R1171_U471 P1_R1171_U470 ; P1_R1171_U111
g15873 nand P1_R1171_U478 P1_R1171_U477 ; P1_R1171_U112
g15874 nand P1_R1171_U485 P1_R1171_U484 ; P1_R1171_U113
g15875 nand P1_R1171_U492 P1_R1171_U491 ; P1_R1171_U114
g15876 nand P1_R1171_U497 P1_R1171_U496 ; P1_R1171_U115
g15877 and P1_U3464 P1_U3068 ; P1_R1171_U116
g15878 and P1_R1171_U186 P1_R1171_U184 ; P1_R1171_U117
g15879 and P1_R1171_U191 P1_R1171_U189 ; P1_R1171_U118
g15880 and P1_R1171_U198 P1_R1171_U197 ; P1_R1171_U119
g15881 and P1_R1171_U379 P1_R1171_U378 P1_R1171_U23 ; P1_R1171_U120
g15882 and P1_R1171_U209 P1_R1171_U6 ; P1_R1171_U121
g15883 and P1_R1171_U217 P1_R1171_U215 ; P1_R1171_U122
g15884 and P1_R1171_U386 P1_R1171_U385 P1_R1171_U35 ; P1_R1171_U123
g15885 and P1_R1171_U223 P1_R1171_U4 ; P1_R1171_U124
g15886 and P1_R1171_U231 P1_R1171_U178 ; P1_R1171_U125
g15887 and P1_R1171_U201 P1_R1171_U7 ; P1_R1171_U126
g15888 and P1_R1171_U236 P1_R1171_U168 ; P1_R1171_U127
g15889 and P1_R1171_U245 P1_R1171_U169 ; P1_R1171_U128
g15890 and P1_R1171_U265 P1_R1171_U264 ; P1_R1171_U129
g15891 and P1_R1171_U10 P1_R1171_U279 ; P1_R1171_U130
g15892 and P1_R1171_U282 P1_R1171_U277 ; P1_R1171_U131
g15893 and P1_R1171_U298 P1_R1171_U295 ; P1_R1171_U132
g15894 and P1_R1171_U365 P1_R1171_U299 ; P1_R1171_U133
g15895 and P1_R1171_U156 P1_R1171_U275 ; P1_R1171_U134
g15896 and P1_R1171_U466 P1_R1171_U465 P1_R1171_U60 ; P1_R1171_U135
g15897 and P1_R1171_U487 P1_R1171_U486 P1_R1171_U169 ; P1_R1171_U136
g15898 and P1_R1171_U340 P1_R1171_U8 ; P1_R1171_U137
g15899 and P1_R1171_U499 P1_R1171_U498 P1_R1171_U168 ; P1_R1171_U138
g15900 and P1_R1171_U347 P1_R1171_U7 ; P1_R1171_U139
g15901 nand P1_R1171_U119 P1_R1171_U199 ; P1_R1171_U140
g15902 nand P1_R1171_U214 P1_R1171_U226 ; P1_R1171_U141
g15903 not P1_U3055 ; P1_R1171_U142
g15904 not P1_U4028 ; P1_R1171_U143
g15905 and P1_R1171_U400 P1_R1171_U399 ; P1_R1171_U144
g15906 nand P1_R1171_U301 P1_R1171_U166 P1_R1171_U361 ; P1_R1171_U145
g15907 and P1_R1171_U407 P1_R1171_U406 ; P1_R1171_U146
g15908 nand P1_R1171_U367 P1_R1171_U366 P1_R1171_U133 ; P1_R1171_U147
g15909 and P1_R1171_U414 P1_R1171_U413 ; P1_R1171_U148
g15910 nand P1_R1171_U362 P1_R1171_U296 P1_R1171_U87 ; P1_R1171_U149
g15911 and P1_R1171_U421 P1_R1171_U420 ; P1_R1171_U150
g15912 nand P1_R1171_U290 P1_R1171_U289 ; P1_R1171_U151
g15913 and P1_R1171_U433 P1_R1171_U432 ; P1_R1171_U152
g15914 nand P1_R1171_U286 P1_R1171_U285 ; P1_R1171_U153
g15915 and P1_R1171_U440 P1_R1171_U439 ; P1_R1171_U154
g15916 nand P1_R1171_U131 P1_R1171_U281 ; P1_R1171_U155
g15917 and P1_R1171_U447 P1_R1171_U446 ; P1_R1171_U156
g15918 and P1_R1171_U452 P1_R1171_U451 ; P1_R1171_U157
g15919 nand P1_R1171_U44 P1_R1171_U324 ; P1_R1171_U158
g15920 nand P1_R1171_U129 P1_R1171_U266 ; P1_R1171_U159
g15921 and P1_R1171_U473 P1_R1171_U472 ; P1_R1171_U160
g15922 nand P1_R1171_U254 P1_R1171_U253 ; P1_R1171_U161
g15923 and P1_R1171_U480 P1_R1171_U479 ; P1_R1171_U162
g15924 nand P1_R1171_U250 P1_R1171_U249 ; P1_R1171_U163
g15925 nand P1_R1171_U240 P1_R1171_U239 ; P1_R1171_U164
g15926 nand P1_R1171_U364 P1_R1171_U363 ; P1_R1171_U165
g15927 nand P1_U3054 P1_R1171_U147 ; P1_R1171_U166
g15928 not P1_R1171_U35 ; P1_R1171_U167
g15929 nand P1_U3485 P1_U3083 ; P1_R1171_U168
g15930 nand P1_U3072 P1_U3494 ; P1_R1171_U169
g15931 nand P1_U3058 P1_U4020 ; P1_R1171_U170
g15932 not P1_R1171_U69 ; P1_R1171_U171
g15933 not P1_R1171_U78 ; P1_R1171_U172
g15934 nand P1_U3065 P1_U4021 ; P1_R1171_U173
g15935 not P1_R1171_U62 ; P1_R1171_U174
g15936 or P1_U3067 P1_U3473 ; P1_R1171_U175
g15937 or P1_U3060 P1_U3470 ; P1_R1171_U176
g15938 or P1_U3467 P1_U3064 ; P1_R1171_U177
g15939 or P1_U3464 P1_U3068 ; P1_R1171_U178
g15940 not P1_R1171_U32 ; P1_R1171_U179
g15941 or P1_U3461 P1_U3078 ; P1_R1171_U180
g15942 not P1_R1171_U43 ; P1_R1171_U181
g15943 not P1_R1171_U44 ; P1_R1171_U182
g15944 nand P1_R1171_U43 P1_R1171_U44 ; P1_R1171_U183
g15945 nand P1_R1171_U116 P1_R1171_U177 ; P1_R1171_U184
g15946 nand P1_R1171_U5 P1_R1171_U183 ; P1_R1171_U185
g15947 nand P1_U3064 P1_U3467 ; P1_R1171_U186
g15948 nand P1_R1171_U117 P1_R1171_U185 ; P1_R1171_U187
g15949 nand P1_R1171_U36 P1_R1171_U35 ; P1_R1171_U188
g15950 nand P1_U3067 P1_R1171_U188 ; P1_R1171_U189
g15951 nand P1_R1171_U4 P1_R1171_U187 ; P1_R1171_U190
g15952 nand P1_U3473 P1_R1171_U167 ; P1_R1171_U191
g15953 not P1_R1171_U42 ; P1_R1171_U192
g15954 or P1_U3070 P1_U3479 ; P1_R1171_U193
g15955 or P1_U3071 P1_U3476 ; P1_R1171_U194
g15956 not P1_R1171_U23 ; P1_R1171_U195
g15957 nand P1_R1171_U24 P1_R1171_U23 ; P1_R1171_U196
g15958 nand P1_U3070 P1_R1171_U196 ; P1_R1171_U197
g15959 nand P1_U3479 P1_R1171_U195 ; P1_R1171_U198
g15960 nand P1_R1171_U6 P1_R1171_U42 ; P1_R1171_U199
g15961 not P1_R1171_U140 ; P1_R1171_U200
g15962 or P1_U3482 P1_U3084 ; P1_R1171_U201
g15963 nand P1_R1171_U201 P1_R1171_U140 ; P1_R1171_U202
g15964 not P1_R1171_U41 ; P1_R1171_U203
g15965 or P1_U3083 P1_U3485 ; P1_R1171_U204
g15966 or P1_U3476 P1_U3071 ; P1_R1171_U205
g15967 nand P1_R1171_U205 P1_R1171_U42 ; P1_R1171_U206
g15968 nand P1_R1171_U120 P1_R1171_U206 ; P1_R1171_U207
g15969 nand P1_R1171_U192 P1_R1171_U23 ; P1_R1171_U208
g15970 nand P1_U3479 P1_U3070 ; P1_R1171_U209
g15971 nand P1_R1171_U121 P1_R1171_U208 ; P1_R1171_U210
g15972 or P1_U3071 P1_U3476 ; P1_R1171_U211
g15973 nand P1_R1171_U182 P1_R1171_U178 ; P1_R1171_U212
g15974 nand P1_U3068 P1_U3464 ; P1_R1171_U213
g15975 not P1_R1171_U46 ; P1_R1171_U214
g15976 nand P1_R1171_U181 P1_R1171_U5 ; P1_R1171_U215
g15977 nand P1_R1171_U46 P1_R1171_U177 ; P1_R1171_U216
g15978 nand P1_U3064 P1_U3467 ; P1_R1171_U217
g15979 not P1_R1171_U45 ; P1_R1171_U218
g15980 or P1_U3470 P1_U3060 ; P1_R1171_U219
g15981 nand P1_R1171_U219 P1_R1171_U45 ; P1_R1171_U220
g15982 nand P1_R1171_U123 P1_R1171_U220 ; P1_R1171_U221
g15983 nand P1_R1171_U218 P1_R1171_U35 ; P1_R1171_U222
g15984 nand P1_U3473 P1_U3067 ; P1_R1171_U223
g15985 nand P1_R1171_U124 P1_R1171_U222 ; P1_R1171_U224
g15986 or P1_U3060 P1_U3470 ; P1_R1171_U225
g15987 nand P1_R1171_U181 P1_R1171_U178 ; P1_R1171_U226
g15988 not P1_R1171_U141 ; P1_R1171_U227
g15989 nand P1_U3064 P1_U3467 ; P1_R1171_U228
g15990 nand P1_R1171_U398 P1_R1171_U397 P1_R1171_U44 P1_R1171_U43 ; P1_R1171_U229
g15991 nand P1_R1171_U44 P1_R1171_U43 ; P1_R1171_U230
g15992 nand P1_U3068 P1_U3464 ; P1_R1171_U231
g15993 nand P1_R1171_U125 P1_R1171_U230 ; P1_R1171_U232
g15994 or P1_U3083 P1_U3485 ; P1_R1171_U233
g15995 or P1_U3062 P1_U3488 ; P1_R1171_U234
g15996 nand P1_R1171_U174 P1_R1171_U7 ; P1_R1171_U235
g15997 nand P1_U3062 P1_U3488 ; P1_R1171_U236
g15998 nand P1_R1171_U127 P1_R1171_U235 ; P1_R1171_U237
g15999 or P1_U3488 P1_U3062 ; P1_R1171_U238
g16000 nand P1_R1171_U126 P1_R1171_U140 ; P1_R1171_U239
g16001 nand P1_R1171_U238 P1_R1171_U237 ; P1_R1171_U240
g16002 not P1_R1171_U164 ; P1_R1171_U241
g16003 or P1_U3080 P1_U3497 ; P1_R1171_U242
g16004 or P1_U3072 P1_U3494 ; P1_R1171_U243
g16005 nand P1_R1171_U171 P1_R1171_U8 ; P1_R1171_U244
g16006 nand P1_U3080 P1_U3497 ; P1_R1171_U245
g16007 nand P1_R1171_U128 P1_R1171_U244 ; P1_R1171_U246
g16008 or P1_U3491 P1_U3063 ; P1_R1171_U247
g16009 or P1_U3497 P1_U3080 ; P1_R1171_U248
g16010 nand P1_R1171_U247 P1_R1171_U164 P1_R1171_U8 ; P1_R1171_U249
g16011 nand P1_R1171_U248 P1_R1171_U246 ; P1_R1171_U250
g16012 not P1_R1171_U163 ; P1_R1171_U251
g16013 or P1_U3500 P1_U3079 ; P1_R1171_U252
g16014 nand P1_R1171_U252 P1_R1171_U163 ; P1_R1171_U253
g16015 nand P1_U3079 P1_U3500 ; P1_R1171_U254
g16016 not P1_R1171_U161 ; P1_R1171_U255
g16017 or P1_U3503 P1_U3074 ; P1_R1171_U256
g16018 nand P1_R1171_U256 P1_R1171_U161 ; P1_R1171_U257
g16019 nand P1_U3074 P1_U3503 ; P1_R1171_U258
g16020 not P1_R1171_U93 ; P1_R1171_U259
g16021 or P1_U3069 P1_U3509 ; P1_R1171_U260
g16022 or P1_U3073 P1_U3506 ; P1_R1171_U261
g16023 not P1_R1171_U60 ; P1_R1171_U262
g16024 nand P1_R1171_U61 P1_R1171_U60 ; P1_R1171_U263
g16025 nand P1_U3069 P1_R1171_U263 ; P1_R1171_U264
g16026 nand P1_U3509 P1_R1171_U262 ; P1_R1171_U265
g16027 nand P1_R1171_U9 P1_R1171_U93 ; P1_R1171_U266
g16028 not P1_R1171_U159 ; P1_R1171_U267
g16029 or P1_U3076 P1_U4025 ; P1_R1171_U268
g16030 or P1_U3081 P1_U3514 ; P1_R1171_U269
g16031 or P1_U3075 P1_U4024 ; P1_R1171_U270
g16032 not P1_R1171_U81 ; P1_R1171_U271
g16033 nand P1_U4025 P1_R1171_U271 ; P1_R1171_U272
g16034 nand P1_R1171_U272 P1_R1171_U91 ; P1_R1171_U273
g16035 nand P1_R1171_U81 P1_R1171_U82 ; P1_R1171_U274
g16036 nand P1_R1171_U274 P1_R1171_U273 ; P1_R1171_U275
g16037 nand P1_R1171_U172 P1_R1171_U10 ; P1_R1171_U276
g16038 nand P1_U3075 P1_U4024 ; P1_R1171_U277
g16039 nand P1_R1171_U275 P1_R1171_U276 ; P1_R1171_U278
g16040 or P1_U3512 P1_U3082 ; P1_R1171_U279
g16041 or P1_U4024 P1_U3075 ; P1_R1171_U280
g16042 nand P1_R1171_U270 P1_R1171_U159 P1_R1171_U130 ; P1_R1171_U281
g16043 nand P1_R1171_U280 P1_R1171_U278 ; P1_R1171_U282
g16044 not P1_R1171_U155 ; P1_R1171_U283
g16045 or P1_U4023 P1_U3061 ; P1_R1171_U284
g16046 nand P1_R1171_U284 P1_R1171_U155 ; P1_R1171_U285
g16047 nand P1_U3061 P1_U4023 ; P1_R1171_U286
g16048 not P1_R1171_U153 ; P1_R1171_U287
g16049 or P1_U4022 P1_U3066 ; P1_R1171_U288
g16050 nand P1_R1171_U288 P1_R1171_U153 ; P1_R1171_U289
g16051 nand P1_U3066 P1_U4022 ; P1_R1171_U290
g16052 not P1_R1171_U151 ; P1_R1171_U291
g16053 or P1_U3058 P1_U4020 ; P1_R1171_U292
g16054 nand P1_R1171_U173 P1_R1171_U170 ; P1_R1171_U293
g16055 not P1_R1171_U87 ; P1_R1171_U294
g16056 or P1_U4021 P1_U3065 ; P1_R1171_U295
g16057 nand P1_R1171_U151 P1_R1171_U295 P1_R1171_U165 ; P1_R1171_U296
g16058 not P1_R1171_U149 ; P1_R1171_U297
g16059 or P1_U4018 P1_U3053 ; P1_R1171_U298
g16060 nand P1_U3053 P1_U4018 ; P1_R1171_U299
g16061 not P1_R1171_U147 ; P1_R1171_U300
g16062 nand P1_U4017 P1_R1171_U147 ; P1_R1171_U301
g16063 not P1_R1171_U145 ; P1_R1171_U302
g16064 nand P1_R1171_U295 P1_R1171_U151 ; P1_R1171_U303
g16065 not P1_R1171_U90 ; P1_R1171_U304
g16066 or P1_U4020 P1_U3058 ; P1_R1171_U305
g16067 nand P1_R1171_U305 P1_R1171_U90 ; P1_R1171_U306
g16068 nand P1_R1171_U306 P1_R1171_U170 P1_R1171_U150 ; P1_R1171_U307
g16069 nand P1_R1171_U304 P1_R1171_U170 ; P1_R1171_U308
g16070 nand P1_U4019 P1_U3057 ; P1_R1171_U309
g16071 nand P1_R1171_U308 P1_R1171_U309 P1_R1171_U165 ; P1_R1171_U310
g16072 or P1_U3058 P1_U4020 ; P1_R1171_U311
g16073 nand P1_R1171_U279 P1_R1171_U159 ; P1_R1171_U312
g16074 not P1_R1171_U92 ; P1_R1171_U313
g16075 nand P1_R1171_U10 P1_R1171_U92 ; P1_R1171_U314
g16076 nand P1_R1171_U134 P1_R1171_U314 ; P1_R1171_U315
g16077 nand P1_R1171_U314 P1_R1171_U275 ; P1_R1171_U316
g16078 nand P1_R1171_U450 P1_R1171_U316 ; P1_R1171_U317
g16079 or P1_U3514 P1_U3081 ; P1_R1171_U318
g16080 nand P1_R1171_U318 P1_R1171_U92 ; P1_R1171_U319
g16081 nand P1_R1171_U319 P1_R1171_U81 P1_R1171_U157 ; P1_R1171_U320
g16082 nand P1_R1171_U313 P1_R1171_U81 ; P1_R1171_U321
g16083 nand P1_U3076 P1_U4025 ; P1_R1171_U322
g16084 nand P1_R1171_U322 P1_R1171_U321 P1_R1171_U10 ; P1_R1171_U323
g16085 or P1_U3461 P1_U3078 ; P1_R1171_U324
g16086 not P1_R1171_U158 ; P1_R1171_U325
g16087 or P1_U3081 P1_U3514 ; P1_R1171_U326
g16088 or P1_U3506 P1_U3073 ; P1_R1171_U327
g16089 nand P1_R1171_U327 P1_R1171_U93 ; P1_R1171_U328
g16090 nand P1_R1171_U135 P1_R1171_U328 ; P1_R1171_U329
g16091 nand P1_R1171_U259 P1_R1171_U60 ; P1_R1171_U330
g16092 nand P1_U3509 P1_U3069 ; P1_R1171_U331
g16093 nand P1_R1171_U331 P1_R1171_U330 P1_R1171_U9 ; P1_R1171_U332
g16094 or P1_U3073 P1_U3506 ; P1_R1171_U333
g16095 nand P1_R1171_U247 P1_R1171_U164 ; P1_R1171_U334
g16096 not P1_R1171_U94 ; P1_R1171_U335
g16097 or P1_U3494 P1_U3072 ; P1_R1171_U336
g16098 nand P1_R1171_U336 P1_R1171_U94 ; P1_R1171_U337
g16099 nand P1_R1171_U136 P1_R1171_U337 ; P1_R1171_U338
g16100 nand P1_R1171_U335 P1_R1171_U169 ; P1_R1171_U339
g16101 nand P1_U3080 P1_U3497 ; P1_R1171_U340
g16102 nand P1_R1171_U137 P1_R1171_U339 ; P1_R1171_U341
g16103 or P1_U3072 P1_U3494 ; P1_R1171_U342
g16104 or P1_U3485 P1_U3083 ; P1_R1171_U343
g16105 nand P1_R1171_U343 P1_R1171_U41 ; P1_R1171_U344
g16106 nand P1_R1171_U138 P1_R1171_U344 ; P1_R1171_U345
g16107 nand P1_R1171_U203 P1_R1171_U168 ; P1_R1171_U346
g16108 nand P1_U3062 P1_U3488 ; P1_R1171_U347
g16109 nand P1_R1171_U139 P1_R1171_U346 ; P1_R1171_U348
g16110 nand P1_R1171_U204 P1_R1171_U168 ; P1_R1171_U349
g16111 nand P1_R1171_U201 P1_R1171_U62 ; P1_R1171_U350
g16112 nand P1_R1171_U211 P1_R1171_U23 ; P1_R1171_U351
g16113 nand P1_R1171_U225 P1_R1171_U35 ; P1_R1171_U352
g16114 nand P1_R1171_U228 P1_R1171_U177 ; P1_R1171_U353
g16115 nand P1_R1171_U311 P1_R1171_U170 ; P1_R1171_U354
g16116 nand P1_R1171_U295 P1_R1171_U173 ; P1_R1171_U355
g16117 nand P1_R1171_U326 P1_R1171_U81 ; P1_R1171_U356
g16118 nand P1_R1171_U279 P1_R1171_U78 ; P1_R1171_U357
g16119 nand P1_R1171_U333 P1_R1171_U60 ; P1_R1171_U358
g16120 nand P1_R1171_U342 P1_R1171_U169 ; P1_R1171_U359
g16121 nand P1_R1171_U247 P1_R1171_U69 ; P1_R1171_U360
g16122 nand P1_U4017 P1_U3054 ; P1_R1171_U361
g16123 nand P1_R1171_U293 P1_R1171_U165 ; P1_R1171_U362
g16124 nand P1_U3057 P1_R1171_U292 ; P1_R1171_U363
g16125 nand P1_U4019 P1_R1171_U292 ; P1_R1171_U364
g16126 nand P1_R1171_U293 P1_R1171_U165 P1_R1171_U298 ; P1_R1171_U365
g16127 nand P1_R1171_U151 P1_R1171_U165 P1_R1171_U132 ; P1_R1171_U366
g16128 nand P1_R1171_U294 P1_R1171_U298 ; P1_R1171_U367
g16129 nand P1_U3083 P1_R1171_U40 ; P1_R1171_U368
g16130 nand P1_U3485 P1_R1171_U39 ; P1_R1171_U369
g16131 nand P1_R1171_U369 P1_R1171_U368 ; P1_R1171_U370
g16132 nand P1_R1171_U349 P1_R1171_U41 ; P1_R1171_U371
g16133 nand P1_R1171_U370 P1_R1171_U203 ; P1_R1171_U372
g16134 nand P1_U3084 P1_R1171_U37 ; P1_R1171_U373
g16135 nand P1_U3482 P1_R1171_U38 ; P1_R1171_U374
g16136 nand P1_R1171_U374 P1_R1171_U373 ; P1_R1171_U375
g16137 nand P1_R1171_U350 P1_R1171_U140 ; P1_R1171_U376
g16138 nand P1_R1171_U200 P1_R1171_U375 ; P1_R1171_U377
g16139 nand P1_U3070 P1_R1171_U24 ; P1_R1171_U378
g16140 nand P1_U3479 P1_R1171_U22 ; P1_R1171_U379
g16141 nand P1_U3071 P1_R1171_U20 ; P1_R1171_U380
g16142 nand P1_U3476 P1_R1171_U21 ; P1_R1171_U381
g16143 nand P1_R1171_U381 P1_R1171_U380 ; P1_R1171_U382
g16144 nand P1_R1171_U351 P1_R1171_U42 ; P1_R1171_U383
g16145 nand P1_R1171_U382 P1_R1171_U192 ; P1_R1171_U384
g16146 nand P1_U3067 P1_R1171_U36 ; P1_R1171_U385
g16147 nand P1_U3473 P1_R1171_U27 ; P1_R1171_U386
g16148 nand P1_U3060 P1_R1171_U25 ; P1_R1171_U387
g16149 nand P1_U3470 P1_R1171_U26 ; P1_R1171_U388
g16150 nand P1_R1171_U388 P1_R1171_U387 ; P1_R1171_U389
g16151 nand P1_R1171_U352 P1_R1171_U45 ; P1_R1171_U390
g16152 nand P1_R1171_U389 P1_R1171_U218 ; P1_R1171_U391
g16153 nand P1_U3064 P1_R1171_U33 ; P1_R1171_U392
g16154 nand P1_U3467 P1_R1171_U34 ; P1_R1171_U393
g16155 nand P1_R1171_U393 P1_R1171_U392 ; P1_R1171_U394
g16156 nand P1_R1171_U353 P1_R1171_U141 ; P1_R1171_U395
g16157 nand P1_R1171_U227 P1_R1171_U394 ; P1_R1171_U396
g16158 nand P1_U3068 P1_R1171_U28 ; P1_R1171_U397
g16159 nand P1_U3464 P1_R1171_U29 ; P1_R1171_U398
g16160 nand P1_U3055 P1_R1171_U143 ; P1_R1171_U399
g16161 nand P1_U4028 P1_R1171_U142 ; P1_R1171_U400
g16162 nand P1_U3055 P1_R1171_U143 ; P1_R1171_U401
g16163 nand P1_U4028 P1_R1171_U142 ; P1_R1171_U402
g16164 nand P1_R1171_U402 P1_R1171_U401 ; P1_R1171_U403
g16165 nand P1_R1171_U144 P1_R1171_U145 ; P1_R1171_U404
g16166 nand P1_R1171_U302 P1_R1171_U403 ; P1_R1171_U405
g16167 nand P1_U3054 P1_R1171_U89 ; P1_R1171_U406
g16168 nand P1_U4017 P1_R1171_U88 ; P1_R1171_U407
g16169 nand P1_U3054 P1_R1171_U89 ; P1_R1171_U408
g16170 nand P1_U4017 P1_R1171_U88 ; P1_R1171_U409
g16171 nand P1_R1171_U409 P1_R1171_U408 ; P1_R1171_U410
g16172 nand P1_R1171_U146 P1_R1171_U147 ; P1_R1171_U411
g16173 nand P1_R1171_U300 P1_R1171_U410 ; P1_R1171_U412
g16174 nand P1_U3053 P1_R1171_U47 ; P1_R1171_U413
g16175 nand P1_U4018 P1_R1171_U48 ; P1_R1171_U414
g16176 nand P1_U3053 P1_R1171_U47 ; P1_R1171_U415
g16177 nand P1_U4018 P1_R1171_U48 ; P1_R1171_U416
g16178 nand P1_R1171_U416 P1_R1171_U415 ; P1_R1171_U417
g16179 nand P1_R1171_U148 P1_R1171_U149 ; P1_R1171_U418
g16180 nand P1_R1171_U297 P1_R1171_U417 ; P1_R1171_U419
g16181 nand P1_U3057 P1_R1171_U50 ; P1_R1171_U420
g16182 nand P1_U4019 P1_R1171_U49 ; P1_R1171_U421
g16183 nand P1_U3058 P1_R1171_U51 ; P1_R1171_U422
g16184 nand P1_U4020 P1_R1171_U52 ; P1_R1171_U423
g16185 nand P1_R1171_U423 P1_R1171_U422 ; P1_R1171_U424
g16186 nand P1_R1171_U354 P1_R1171_U90 ; P1_R1171_U425
g16187 nand P1_R1171_U424 P1_R1171_U304 ; P1_R1171_U426
g16188 nand P1_U3065 P1_R1171_U53 ; P1_R1171_U427
g16189 nand P1_U4021 P1_R1171_U54 ; P1_R1171_U428
g16190 nand P1_R1171_U428 P1_R1171_U427 ; P1_R1171_U429
g16191 nand P1_R1171_U355 P1_R1171_U151 ; P1_R1171_U430
g16192 nand P1_R1171_U291 P1_R1171_U429 ; P1_R1171_U431
g16193 nand P1_U3066 P1_R1171_U85 ; P1_R1171_U432
g16194 nand P1_U4022 P1_R1171_U86 ; P1_R1171_U433
g16195 nand P1_U3066 P1_R1171_U85 ; P1_R1171_U434
g16196 nand P1_U4022 P1_R1171_U86 ; P1_R1171_U435
g16197 nand P1_R1171_U435 P1_R1171_U434 ; P1_R1171_U436
g16198 nand P1_R1171_U152 P1_R1171_U153 ; P1_R1171_U437
g16199 nand P1_R1171_U287 P1_R1171_U436 ; P1_R1171_U438
g16200 nand P1_U3061 P1_R1171_U83 ; P1_R1171_U439
g16201 nand P1_U4023 P1_R1171_U84 ; P1_R1171_U440
g16202 nand P1_U3061 P1_R1171_U83 ; P1_R1171_U441
g16203 nand P1_U4023 P1_R1171_U84 ; P1_R1171_U442
g16204 nand P1_R1171_U442 P1_R1171_U441 ; P1_R1171_U443
g16205 nand P1_R1171_U154 P1_R1171_U155 ; P1_R1171_U444
g16206 nand P1_R1171_U283 P1_R1171_U443 ; P1_R1171_U445
g16207 nand P1_U3075 P1_R1171_U55 ; P1_R1171_U446
g16208 nand P1_U4024 P1_R1171_U56 ; P1_R1171_U447
g16209 nand P1_U3075 P1_R1171_U55 ; P1_R1171_U448
g16210 nand P1_U4024 P1_R1171_U56 ; P1_R1171_U449
g16211 nand P1_R1171_U449 P1_R1171_U448 ; P1_R1171_U450
g16212 nand P1_U3076 P1_R1171_U82 ; P1_R1171_U451
g16213 nand P1_U4025 P1_R1171_U91 ; P1_R1171_U452
g16214 nand P1_R1171_U179 P1_R1171_U158 ; P1_R1171_U453
g16215 nand P1_R1171_U325 P1_R1171_U32 ; P1_R1171_U454
g16216 nand P1_U3081 P1_R1171_U79 ; P1_R1171_U455
g16217 nand P1_U3514 P1_R1171_U80 ; P1_R1171_U456
g16218 nand P1_R1171_U456 P1_R1171_U455 ; P1_R1171_U457
g16219 nand P1_R1171_U356 P1_R1171_U92 ; P1_R1171_U458
g16220 nand P1_R1171_U457 P1_R1171_U313 ; P1_R1171_U459
g16221 nand P1_U3082 P1_R1171_U76 ; P1_R1171_U460
g16222 nand P1_U3512 P1_R1171_U77 ; P1_R1171_U461
g16223 nand P1_R1171_U461 P1_R1171_U460 ; P1_R1171_U462
g16224 nand P1_R1171_U357 P1_R1171_U159 ; P1_R1171_U463
g16225 nand P1_R1171_U267 P1_R1171_U462 ; P1_R1171_U464
g16226 nand P1_U3069 P1_R1171_U61 ; P1_R1171_U465
g16227 nand P1_U3509 P1_R1171_U59 ; P1_R1171_U466
g16228 nand P1_U3073 P1_R1171_U57 ; P1_R1171_U467
g16229 nand P1_U3506 P1_R1171_U58 ; P1_R1171_U468
g16230 nand P1_R1171_U468 P1_R1171_U467 ; P1_R1171_U469
g16231 nand P1_R1171_U358 P1_R1171_U93 ; P1_R1171_U470
g16232 nand P1_R1171_U469 P1_R1171_U259 ; P1_R1171_U471
g16233 nand P1_U3074 P1_R1171_U74 ; P1_R1171_U472
g16234 nand P1_U3503 P1_R1171_U75 ; P1_R1171_U473
g16235 nand P1_U3074 P1_R1171_U74 ; P1_R1171_U474
g16236 nand P1_U3503 P1_R1171_U75 ; P1_R1171_U475
g16237 nand P1_R1171_U475 P1_R1171_U474 ; P1_R1171_U476
g16238 nand P1_R1171_U160 P1_R1171_U161 ; P1_R1171_U477
g16239 nand P1_R1171_U255 P1_R1171_U476 ; P1_R1171_U478
g16240 nand P1_U3079 P1_R1171_U72 ; P1_R1171_U479
g16241 nand P1_U3500 P1_R1171_U73 ; P1_R1171_U480
g16242 nand P1_U3079 P1_R1171_U72 ; P1_R1171_U481
g16243 nand P1_U3500 P1_R1171_U73 ; P1_R1171_U482
g16244 nand P1_R1171_U482 P1_R1171_U481 ; P1_R1171_U483
g16245 nand P1_R1171_U162 P1_R1171_U163 ; P1_R1171_U484
g16246 nand P1_R1171_U251 P1_R1171_U483 ; P1_R1171_U485
g16247 nand P1_U3080 P1_R1171_U70 ; P1_R1171_U486
g16248 nand P1_U3497 P1_R1171_U71 ; P1_R1171_U487
g16249 nand P1_U3072 P1_R1171_U65 ; P1_R1171_U488
g16250 nand P1_U3494 P1_R1171_U66 ; P1_R1171_U489
g16251 nand P1_R1171_U489 P1_R1171_U488 ; P1_R1171_U490
g16252 nand P1_R1171_U359 P1_R1171_U94 ; P1_R1171_U491
g16253 nand P1_R1171_U490 P1_R1171_U335 ; P1_R1171_U492
g16254 nand P1_U3063 P1_R1171_U67 ; P1_R1171_U493
g16255 nand P1_U3491 P1_R1171_U68 ; P1_R1171_U494
g16256 nand P1_R1171_U494 P1_R1171_U493 ; P1_R1171_U495
g16257 nand P1_R1171_U360 P1_R1171_U164 ; P1_R1171_U496
g16258 nand P1_R1171_U241 P1_R1171_U495 ; P1_R1171_U497
g16259 nand P1_U3062 P1_R1171_U63 ; P1_R1171_U498
g16260 nand P1_U3488 P1_R1171_U64 ; P1_R1171_U499
g16261 nand P1_U3077 P1_R1171_U30 ; P1_R1171_U500
g16262 nand P1_U3456 P1_R1171_U31 ; P1_R1171_U501
g16263 and P1_R1138_U176 P1_R1138_U175 ; P1_R1138_U4
g16264 and P1_R1138_U177 P1_R1138_U178 ; P1_R1138_U5
g16265 and P1_R1138_U194 P1_R1138_U193 ; P1_R1138_U6
g16266 and P1_R1138_U234 P1_R1138_U233 ; P1_R1138_U7
g16267 and P1_R1138_U243 P1_R1138_U242 ; P1_R1138_U8
g16268 and P1_R1138_U261 P1_R1138_U260 ; P1_R1138_U9
g16269 and P1_R1138_U269 P1_R1138_U268 ; P1_R1138_U10
g16270 and P1_R1138_U348 P1_R1138_U345 ; P1_R1138_U11
g16271 and P1_R1138_U341 P1_R1138_U338 ; P1_R1138_U12
g16272 and P1_R1138_U332 P1_R1138_U329 ; P1_R1138_U13
g16273 and P1_R1138_U323 P1_R1138_U320 ; P1_R1138_U14
g16274 and P1_R1138_U317 P1_R1138_U315 ; P1_R1138_U15
g16275 and P1_R1138_U310 P1_R1138_U307 ; P1_R1138_U16
g16276 and P1_R1138_U232 P1_R1138_U229 ; P1_R1138_U17
g16277 and P1_R1138_U224 P1_R1138_U221 ; P1_R1138_U18
g16278 and P1_R1138_U210 P1_R1138_U207 ; P1_R1138_U19
g16279 not P1_U3476 ; P1_R1138_U20
g16280 not P1_U3071 ; P1_R1138_U21
g16281 not P1_U3070 ; P1_R1138_U22
g16282 nand P1_U3071 P1_U3476 ; P1_R1138_U23
g16283 not P1_U3479 ; P1_R1138_U24
g16284 not P1_U3470 ; P1_R1138_U25
g16285 not P1_U3060 ; P1_R1138_U26
g16286 not P1_U3067 ; P1_R1138_U27
g16287 not P1_U3464 ; P1_R1138_U28
g16288 not P1_U3068 ; P1_R1138_U29
g16289 not P1_U3456 ; P1_R1138_U30
g16290 not P1_U3077 ; P1_R1138_U31
g16291 nand P1_U3077 P1_U3456 ; P1_R1138_U32
g16292 not P1_U3467 ; P1_R1138_U33
g16293 not P1_U3064 ; P1_R1138_U34
g16294 nand P1_U3060 P1_U3470 ; P1_R1138_U35
g16295 not P1_U3473 ; P1_R1138_U36
g16296 not P1_U3482 ; P1_R1138_U37
g16297 not P1_U3084 ; P1_R1138_U38
g16298 not P1_U3083 ; P1_R1138_U39
g16299 not P1_U3485 ; P1_R1138_U40
g16300 nand P1_R1138_U62 P1_R1138_U202 ; P1_R1138_U41
g16301 nand P1_R1138_U118 P1_R1138_U190 ; P1_R1138_U42
g16302 nand P1_R1138_U179 P1_R1138_U180 ; P1_R1138_U43
g16303 nand P1_U3461 P1_U3078 ; P1_R1138_U44
g16304 nand P1_R1138_U122 P1_R1138_U216 ; P1_R1138_U45
g16305 nand P1_R1138_U213 P1_R1138_U212 ; P1_R1138_U46
g16306 not P1_U4018 ; P1_R1138_U47
g16307 not P1_U3053 ; P1_R1138_U48
g16308 not P1_U3057 ; P1_R1138_U49
g16309 not P1_U4019 ; P1_R1138_U50
g16310 not P1_U4020 ; P1_R1138_U51
g16311 not P1_U3058 ; P1_R1138_U52
g16312 not P1_U4021 ; P1_R1138_U53
g16313 not P1_U3065 ; P1_R1138_U54
g16314 not P1_U4024 ; P1_R1138_U55
g16315 not P1_U3075 ; P1_R1138_U56
g16316 not P1_U3506 ; P1_R1138_U57
g16317 not P1_U3073 ; P1_R1138_U58
g16318 not P1_U3069 ; P1_R1138_U59
g16319 nand P1_U3073 P1_U3506 ; P1_R1138_U60
g16320 not P1_U3509 ; P1_R1138_U61
g16321 nand P1_U3084 P1_U3482 ; P1_R1138_U62
g16322 not P1_U3488 ; P1_R1138_U63
g16323 not P1_U3062 ; P1_R1138_U64
g16324 not P1_U3494 ; P1_R1138_U65
g16325 not P1_U3072 ; P1_R1138_U66
g16326 not P1_U3491 ; P1_R1138_U67
g16327 not P1_U3063 ; P1_R1138_U68
g16328 nand P1_U3063 P1_U3491 ; P1_R1138_U69
g16329 not P1_U3497 ; P1_R1138_U70
g16330 not P1_U3080 ; P1_R1138_U71
g16331 not P1_U3500 ; P1_R1138_U72
g16332 not P1_U3079 ; P1_R1138_U73
g16333 not P1_U3503 ; P1_R1138_U74
g16334 not P1_U3074 ; P1_R1138_U75
g16335 not P1_U3512 ; P1_R1138_U76
g16336 not P1_U3082 ; P1_R1138_U77
g16337 nand P1_U3082 P1_U3512 ; P1_R1138_U78
g16338 not P1_U3514 ; P1_R1138_U79
g16339 not P1_U3081 ; P1_R1138_U80
g16340 nand P1_U3081 P1_U3514 ; P1_R1138_U81
g16341 not P1_U4025 ; P1_R1138_U82
g16342 not P1_U4023 ; P1_R1138_U83
g16343 not P1_U3061 ; P1_R1138_U84
g16344 not P1_U4022 ; P1_R1138_U85
g16345 not P1_U3066 ; P1_R1138_U86
g16346 nand P1_U4019 P1_U3057 ; P1_R1138_U87
g16347 not P1_U3054 ; P1_R1138_U88
g16348 not P1_U4017 ; P1_R1138_U89
g16349 nand P1_R1138_U303 P1_R1138_U173 ; P1_R1138_U90
g16350 not P1_U3076 ; P1_R1138_U91
g16351 nand P1_R1138_U78 P1_R1138_U312 ; P1_R1138_U92
g16352 nand P1_R1138_U258 P1_R1138_U257 ; P1_R1138_U93
g16353 nand P1_R1138_U69 P1_R1138_U334 ; P1_R1138_U94
g16354 nand P1_R1138_U454 P1_R1138_U453 ; P1_R1138_U95
g16355 nand P1_R1138_U501 P1_R1138_U500 ; P1_R1138_U96
g16356 nand P1_R1138_U372 P1_R1138_U371 ; P1_R1138_U97
g16357 nand P1_R1138_U377 P1_R1138_U376 ; P1_R1138_U98
g16358 nand P1_R1138_U384 P1_R1138_U383 ; P1_R1138_U99
g16359 nand P1_R1138_U391 P1_R1138_U390 ; P1_R1138_U100
g16360 nand P1_R1138_U396 P1_R1138_U395 ; P1_R1138_U101
g16361 nand P1_R1138_U405 P1_R1138_U404 ; P1_R1138_U102
g16362 nand P1_R1138_U412 P1_R1138_U411 ; P1_R1138_U103
g16363 nand P1_R1138_U419 P1_R1138_U418 ; P1_R1138_U104
g16364 nand P1_R1138_U426 P1_R1138_U425 ; P1_R1138_U105
g16365 nand P1_R1138_U431 P1_R1138_U430 ; P1_R1138_U106
g16366 nand P1_R1138_U438 P1_R1138_U437 ; P1_R1138_U107
g16367 nand P1_R1138_U445 P1_R1138_U444 ; P1_R1138_U108
g16368 nand P1_R1138_U459 P1_R1138_U458 ; P1_R1138_U109
g16369 nand P1_R1138_U464 P1_R1138_U463 ; P1_R1138_U110
g16370 nand P1_R1138_U471 P1_R1138_U470 ; P1_R1138_U111
g16371 nand P1_R1138_U478 P1_R1138_U477 ; P1_R1138_U112
g16372 nand P1_R1138_U485 P1_R1138_U484 ; P1_R1138_U113
g16373 nand P1_R1138_U492 P1_R1138_U491 ; P1_R1138_U114
g16374 nand P1_R1138_U497 P1_R1138_U496 ; P1_R1138_U115
g16375 and P1_U3464 P1_U3068 ; P1_R1138_U116
g16376 and P1_R1138_U186 P1_R1138_U184 ; P1_R1138_U117
g16377 and P1_R1138_U191 P1_R1138_U189 ; P1_R1138_U118
g16378 and P1_R1138_U198 P1_R1138_U197 ; P1_R1138_U119
g16379 and P1_R1138_U379 P1_R1138_U378 P1_R1138_U23 ; P1_R1138_U120
g16380 and P1_R1138_U209 P1_R1138_U6 ; P1_R1138_U121
g16381 and P1_R1138_U217 P1_R1138_U215 ; P1_R1138_U122
g16382 and P1_R1138_U386 P1_R1138_U385 P1_R1138_U35 ; P1_R1138_U123
g16383 and P1_R1138_U223 P1_R1138_U4 ; P1_R1138_U124
g16384 and P1_R1138_U231 P1_R1138_U178 ; P1_R1138_U125
g16385 and P1_R1138_U201 P1_R1138_U7 ; P1_R1138_U126
g16386 and P1_R1138_U236 P1_R1138_U168 ; P1_R1138_U127
g16387 and P1_R1138_U245 P1_R1138_U169 ; P1_R1138_U128
g16388 and P1_R1138_U265 P1_R1138_U264 ; P1_R1138_U129
g16389 and P1_R1138_U10 P1_R1138_U279 ; P1_R1138_U130
g16390 and P1_R1138_U282 P1_R1138_U277 ; P1_R1138_U131
g16391 and P1_R1138_U298 P1_R1138_U295 ; P1_R1138_U132
g16392 and P1_R1138_U365 P1_R1138_U299 ; P1_R1138_U133
g16393 and P1_R1138_U156 P1_R1138_U275 ; P1_R1138_U134
g16394 and P1_R1138_U466 P1_R1138_U465 P1_R1138_U60 ; P1_R1138_U135
g16395 and P1_R1138_U487 P1_R1138_U486 P1_R1138_U169 ; P1_R1138_U136
g16396 and P1_R1138_U340 P1_R1138_U8 ; P1_R1138_U137
g16397 and P1_R1138_U499 P1_R1138_U498 P1_R1138_U168 ; P1_R1138_U138
g16398 and P1_R1138_U347 P1_R1138_U7 ; P1_R1138_U139
g16399 nand P1_R1138_U119 P1_R1138_U199 ; P1_R1138_U140
g16400 nand P1_R1138_U214 P1_R1138_U226 ; P1_R1138_U141
g16401 not P1_U3055 ; P1_R1138_U142
g16402 not P1_U4028 ; P1_R1138_U143
g16403 and P1_R1138_U400 P1_R1138_U399 ; P1_R1138_U144
g16404 nand P1_R1138_U301 P1_R1138_U166 P1_R1138_U361 ; P1_R1138_U145
g16405 and P1_R1138_U407 P1_R1138_U406 ; P1_R1138_U146
g16406 nand P1_R1138_U367 P1_R1138_U366 P1_R1138_U133 ; P1_R1138_U147
g16407 and P1_R1138_U414 P1_R1138_U413 ; P1_R1138_U148
g16408 nand P1_R1138_U362 P1_R1138_U296 P1_R1138_U87 ; P1_R1138_U149
g16409 and P1_R1138_U421 P1_R1138_U420 ; P1_R1138_U150
g16410 nand P1_R1138_U290 P1_R1138_U289 ; P1_R1138_U151
g16411 and P1_R1138_U433 P1_R1138_U432 ; P1_R1138_U152
g16412 nand P1_R1138_U286 P1_R1138_U285 ; P1_R1138_U153
g16413 and P1_R1138_U440 P1_R1138_U439 ; P1_R1138_U154
g16414 nand P1_R1138_U131 P1_R1138_U281 ; P1_R1138_U155
g16415 and P1_R1138_U447 P1_R1138_U446 ; P1_R1138_U156
g16416 and P1_R1138_U452 P1_R1138_U451 ; P1_R1138_U157
g16417 nand P1_R1138_U44 P1_R1138_U324 ; P1_R1138_U158
g16418 nand P1_R1138_U129 P1_R1138_U266 ; P1_R1138_U159
g16419 and P1_R1138_U473 P1_R1138_U472 ; P1_R1138_U160
g16420 nand P1_R1138_U254 P1_R1138_U253 ; P1_R1138_U161
g16421 and P1_R1138_U480 P1_R1138_U479 ; P1_R1138_U162
g16422 nand P1_R1138_U250 P1_R1138_U249 ; P1_R1138_U163
g16423 nand P1_R1138_U240 P1_R1138_U239 ; P1_R1138_U164
g16424 nand P1_R1138_U364 P1_R1138_U363 ; P1_R1138_U165
g16425 nand P1_U3054 P1_R1138_U147 ; P1_R1138_U166
g16426 not P1_R1138_U35 ; P1_R1138_U167
g16427 nand P1_U3485 P1_U3083 ; P1_R1138_U168
g16428 nand P1_U3072 P1_U3494 ; P1_R1138_U169
g16429 nand P1_U3058 P1_U4020 ; P1_R1138_U170
g16430 not P1_R1138_U69 ; P1_R1138_U171
g16431 not P1_R1138_U78 ; P1_R1138_U172
g16432 nand P1_U3065 P1_U4021 ; P1_R1138_U173
g16433 not P1_R1138_U62 ; P1_R1138_U174
g16434 or P1_U3067 P1_U3473 ; P1_R1138_U175
g16435 or P1_U3060 P1_U3470 ; P1_R1138_U176
g16436 or P1_U3467 P1_U3064 ; P1_R1138_U177
g16437 or P1_U3464 P1_U3068 ; P1_R1138_U178
g16438 not P1_R1138_U32 ; P1_R1138_U179
g16439 or P1_U3461 P1_U3078 ; P1_R1138_U180
g16440 not P1_R1138_U43 ; P1_R1138_U181
g16441 not P1_R1138_U44 ; P1_R1138_U182
g16442 nand P1_R1138_U43 P1_R1138_U44 ; P1_R1138_U183
g16443 nand P1_R1138_U116 P1_R1138_U177 ; P1_R1138_U184
g16444 nand P1_R1138_U5 P1_R1138_U183 ; P1_R1138_U185
g16445 nand P1_U3064 P1_U3467 ; P1_R1138_U186
g16446 nand P1_R1138_U117 P1_R1138_U185 ; P1_R1138_U187
g16447 nand P1_R1138_U36 P1_R1138_U35 ; P1_R1138_U188
g16448 nand P1_U3067 P1_R1138_U188 ; P1_R1138_U189
g16449 nand P1_R1138_U4 P1_R1138_U187 ; P1_R1138_U190
g16450 nand P1_U3473 P1_R1138_U167 ; P1_R1138_U191
g16451 not P1_R1138_U42 ; P1_R1138_U192
g16452 or P1_U3070 P1_U3479 ; P1_R1138_U193
g16453 or P1_U3071 P1_U3476 ; P1_R1138_U194
g16454 not P1_R1138_U23 ; P1_R1138_U195
g16455 nand P1_R1138_U24 P1_R1138_U23 ; P1_R1138_U196
g16456 nand P1_U3070 P1_R1138_U196 ; P1_R1138_U197
g16457 nand P1_U3479 P1_R1138_U195 ; P1_R1138_U198
g16458 nand P1_R1138_U6 P1_R1138_U42 ; P1_R1138_U199
g16459 not P1_R1138_U140 ; P1_R1138_U200
g16460 or P1_U3482 P1_U3084 ; P1_R1138_U201
g16461 nand P1_R1138_U201 P1_R1138_U140 ; P1_R1138_U202
g16462 not P1_R1138_U41 ; P1_R1138_U203
g16463 or P1_U3083 P1_U3485 ; P1_R1138_U204
g16464 or P1_U3476 P1_U3071 ; P1_R1138_U205
g16465 nand P1_R1138_U205 P1_R1138_U42 ; P1_R1138_U206
g16466 nand P1_R1138_U120 P1_R1138_U206 ; P1_R1138_U207
g16467 nand P1_R1138_U192 P1_R1138_U23 ; P1_R1138_U208
g16468 nand P1_U3479 P1_U3070 ; P1_R1138_U209
g16469 nand P1_R1138_U121 P1_R1138_U208 ; P1_R1138_U210
g16470 or P1_U3071 P1_U3476 ; P1_R1138_U211
g16471 nand P1_R1138_U182 P1_R1138_U178 ; P1_R1138_U212
g16472 nand P1_U3068 P1_U3464 ; P1_R1138_U213
g16473 not P1_R1138_U46 ; P1_R1138_U214
g16474 nand P1_R1138_U181 P1_R1138_U5 ; P1_R1138_U215
g16475 nand P1_R1138_U46 P1_R1138_U177 ; P1_R1138_U216
g16476 nand P1_U3064 P1_U3467 ; P1_R1138_U217
g16477 not P1_R1138_U45 ; P1_R1138_U218
g16478 or P1_U3470 P1_U3060 ; P1_R1138_U219
g16479 nand P1_R1138_U219 P1_R1138_U45 ; P1_R1138_U220
g16480 nand P1_R1138_U123 P1_R1138_U220 ; P1_R1138_U221
g16481 nand P1_R1138_U218 P1_R1138_U35 ; P1_R1138_U222
g16482 nand P1_U3473 P1_U3067 ; P1_R1138_U223
g16483 nand P1_R1138_U124 P1_R1138_U222 ; P1_R1138_U224
g16484 or P1_U3060 P1_U3470 ; P1_R1138_U225
g16485 nand P1_R1138_U181 P1_R1138_U178 ; P1_R1138_U226
g16486 not P1_R1138_U141 ; P1_R1138_U227
g16487 nand P1_U3064 P1_U3467 ; P1_R1138_U228
g16488 nand P1_R1138_U398 P1_R1138_U397 P1_R1138_U44 P1_R1138_U43 ; P1_R1138_U229
g16489 nand P1_R1138_U44 P1_R1138_U43 ; P1_R1138_U230
g16490 nand P1_U3068 P1_U3464 ; P1_R1138_U231
g16491 nand P1_R1138_U125 P1_R1138_U230 ; P1_R1138_U232
g16492 or P1_U3083 P1_U3485 ; P1_R1138_U233
g16493 or P1_U3062 P1_U3488 ; P1_R1138_U234
g16494 nand P1_R1138_U174 P1_R1138_U7 ; P1_R1138_U235
g16495 nand P1_U3062 P1_U3488 ; P1_R1138_U236
g16496 nand P1_R1138_U127 P1_R1138_U235 ; P1_R1138_U237
g16497 or P1_U3488 P1_U3062 ; P1_R1138_U238
g16498 nand P1_R1138_U126 P1_R1138_U140 ; P1_R1138_U239
g16499 nand P1_R1138_U238 P1_R1138_U237 ; P1_R1138_U240
g16500 not P1_R1138_U164 ; P1_R1138_U241
g16501 or P1_U3080 P1_U3497 ; P1_R1138_U242
g16502 or P1_U3072 P1_U3494 ; P1_R1138_U243
g16503 nand P1_R1138_U171 P1_R1138_U8 ; P1_R1138_U244
g16504 nand P1_U3080 P1_U3497 ; P1_R1138_U245
g16505 nand P1_R1138_U128 P1_R1138_U244 ; P1_R1138_U246
g16506 or P1_U3491 P1_U3063 ; P1_R1138_U247
g16507 or P1_U3497 P1_U3080 ; P1_R1138_U248
g16508 nand P1_R1138_U247 P1_R1138_U164 P1_R1138_U8 ; P1_R1138_U249
g16509 nand P1_R1138_U248 P1_R1138_U246 ; P1_R1138_U250
g16510 not P1_R1138_U163 ; P1_R1138_U251
g16511 or P1_U3500 P1_U3079 ; P1_R1138_U252
g16512 nand P1_R1138_U252 P1_R1138_U163 ; P1_R1138_U253
g16513 nand P1_U3079 P1_U3500 ; P1_R1138_U254
g16514 not P1_R1138_U161 ; P1_R1138_U255
g16515 or P1_U3503 P1_U3074 ; P1_R1138_U256
g16516 nand P1_R1138_U256 P1_R1138_U161 ; P1_R1138_U257
g16517 nand P1_U3074 P1_U3503 ; P1_R1138_U258
g16518 not P1_R1138_U93 ; P1_R1138_U259
g16519 or P1_U3069 P1_U3509 ; P1_R1138_U260
g16520 or P1_U3073 P1_U3506 ; P1_R1138_U261
g16521 not P1_R1138_U60 ; P1_R1138_U262
g16522 nand P1_R1138_U61 P1_R1138_U60 ; P1_R1138_U263
g16523 nand P1_U3069 P1_R1138_U263 ; P1_R1138_U264
g16524 nand P1_U3509 P1_R1138_U262 ; P1_R1138_U265
g16525 nand P1_R1138_U9 P1_R1138_U93 ; P1_R1138_U266
g16526 not P1_R1138_U159 ; P1_R1138_U267
g16527 or P1_U3076 P1_U4025 ; P1_R1138_U268
g16528 or P1_U3081 P1_U3514 ; P1_R1138_U269
g16529 or P1_U3075 P1_U4024 ; P1_R1138_U270
g16530 not P1_R1138_U81 ; P1_R1138_U271
g16531 nand P1_U4025 P1_R1138_U271 ; P1_R1138_U272
g16532 nand P1_R1138_U272 P1_R1138_U91 ; P1_R1138_U273
g16533 nand P1_R1138_U81 P1_R1138_U82 ; P1_R1138_U274
g16534 nand P1_R1138_U274 P1_R1138_U273 ; P1_R1138_U275
g16535 nand P1_R1138_U172 P1_R1138_U10 ; P1_R1138_U276
g16536 nand P1_U3075 P1_U4024 ; P1_R1138_U277
g16537 nand P1_R1138_U275 P1_R1138_U276 ; P1_R1138_U278
g16538 or P1_U3512 P1_U3082 ; P1_R1138_U279
g16539 or P1_U4024 P1_U3075 ; P1_R1138_U280
g16540 nand P1_R1138_U270 P1_R1138_U159 P1_R1138_U130 ; P1_R1138_U281
g16541 nand P1_R1138_U280 P1_R1138_U278 ; P1_R1138_U282
g16542 not P1_R1138_U155 ; P1_R1138_U283
g16543 or P1_U4023 P1_U3061 ; P1_R1138_U284
g16544 nand P1_R1138_U284 P1_R1138_U155 ; P1_R1138_U285
g16545 nand P1_U3061 P1_U4023 ; P1_R1138_U286
g16546 not P1_R1138_U153 ; P1_R1138_U287
g16547 or P1_U4022 P1_U3066 ; P1_R1138_U288
g16548 nand P1_R1138_U288 P1_R1138_U153 ; P1_R1138_U289
g16549 nand P1_U3066 P1_U4022 ; P1_R1138_U290
g16550 not P1_R1138_U151 ; P1_R1138_U291
g16551 or P1_U3058 P1_U4020 ; P1_R1138_U292
g16552 nand P1_R1138_U173 P1_R1138_U170 ; P1_R1138_U293
g16553 not P1_R1138_U87 ; P1_R1138_U294
g16554 or P1_U4021 P1_U3065 ; P1_R1138_U295
g16555 nand P1_R1138_U151 P1_R1138_U295 P1_R1138_U165 ; P1_R1138_U296
g16556 not P1_R1138_U149 ; P1_R1138_U297
g16557 or P1_U4018 P1_U3053 ; P1_R1138_U298
g16558 nand P1_U3053 P1_U4018 ; P1_R1138_U299
g16559 not P1_R1138_U147 ; P1_R1138_U300
g16560 nand P1_U4017 P1_R1138_U147 ; P1_R1138_U301
g16561 not P1_R1138_U145 ; P1_R1138_U302
g16562 nand P1_R1138_U295 P1_R1138_U151 ; P1_R1138_U303
g16563 not P1_R1138_U90 ; P1_R1138_U304
g16564 or P1_U4020 P1_U3058 ; P1_R1138_U305
g16565 nand P1_R1138_U305 P1_R1138_U90 ; P1_R1138_U306
g16566 nand P1_R1138_U306 P1_R1138_U170 P1_R1138_U150 ; P1_R1138_U307
g16567 nand P1_R1138_U304 P1_R1138_U170 ; P1_R1138_U308
g16568 nand P1_U4019 P1_U3057 ; P1_R1138_U309
g16569 nand P1_R1138_U308 P1_R1138_U309 P1_R1138_U165 ; P1_R1138_U310
g16570 or P1_U3058 P1_U4020 ; P1_R1138_U311
g16571 nand P1_R1138_U279 P1_R1138_U159 ; P1_R1138_U312
g16572 not P1_R1138_U92 ; P1_R1138_U313
g16573 nand P1_R1138_U10 P1_R1138_U92 ; P1_R1138_U314
g16574 nand P1_R1138_U134 P1_R1138_U314 ; P1_R1138_U315
g16575 nand P1_R1138_U314 P1_R1138_U275 ; P1_R1138_U316
g16576 nand P1_R1138_U450 P1_R1138_U316 ; P1_R1138_U317
g16577 or P1_U3514 P1_U3081 ; P1_R1138_U318
g16578 nand P1_R1138_U318 P1_R1138_U92 ; P1_R1138_U319
g16579 nand P1_R1138_U319 P1_R1138_U81 P1_R1138_U157 ; P1_R1138_U320
g16580 nand P1_R1138_U313 P1_R1138_U81 ; P1_R1138_U321
g16581 nand P1_U3076 P1_U4025 ; P1_R1138_U322
g16582 nand P1_R1138_U322 P1_R1138_U321 P1_R1138_U10 ; P1_R1138_U323
g16583 or P1_U3461 P1_U3078 ; P1_R1138_U324
g16584 not P1_R1138_U158 ; P1_R1138_U325
g16585 or P1_U3081 P1_U3514 ; P1_R1138_U326
g16586 or P1_U3506 P1_U3073 ; P1_R1138_U327
g16587 nand P1_R1138_U327 P1_R1138_U93 ; P1_R1138_U328
g16588 nand P1_R1138_U135 P1_R1138_U328 ; P1_R1138_U329
g16589 nand P1_R1138_U259 P1_R1138_U60 ; P1_R1138_U330
g16590 nand P1_U3509 P1_U3069 ; P1_R1138_U331
g16591 nand P1_R1138_U331 P1_R1138_U330 P1_R1138_U9 ; P1_R1138_U332
g16592 or P1_U3073 P1_U3506 ; P1_R1138_U333
g16593 nand P1_R1138_U247 P1_R1138_U164 ; P1_R1138_U334
g16594 not P1_R1138_U94 ; P1_R1138_U335
g16595 or P1_U3494 P1_U3072 ; P1_R1138_U336
g16596 nand P1_R1138_U336 P1_R1138_U94 ; P1_R1138_U337
g16597 nand P1_R1138_U136 P1_R1138_U337 ; P1_R1138_U338
g16598 nand P1_R1138_U335 P1_R1138_U169 ; P1_R1138_U339
g16599 nand P1_U3080 P1_U3497 ; P1_R1138_U340
g16600 nand P1_R1138_U137 P1_R1138_U339 ; P1_R1138_U341
g16601 or P1_U3072 P1_U3494 ; P1_R1138_U342
g16602 or P1_U3485 P1_U3083 ; P1_R1138_U343
g16603 nand P1_R1138_U343 P1_R1138_U41 ; P1_R1138_U344
g16604 nand P1_R1138_U138 P1_R1138_U344 ; P1_R1138_U345
g16605 nand P1_R1138_U203 P1_R1138_U168 ; P1_R1138_U346
g16606 nand P1_U3062 P1_U3488 ; P1_R1138_U347
g16607 nand P1_R1138_U139 P1_R1138_U346 ; P1_R1138_U348
g16608 nand P1_R1138_U204 P1_R1138_U168 ; P1_R1138_U349
g16609 nand P1_R1138_U201 P1_R1138_U62 ; P1_R1138_U350
g16610 nand P1_R1138_U211 P1_R1138_U23 ; P1_R1138_U351
g16611 nand P1_R1138_U225 P1_R1138_U35 ; P1_R1138_U352
g16612 nand P1_R1138_U228 P1_R1138_U177 ; P1_R1138_U353
g16613 nand P1_R1138_U311 P1_R1138_U170 ; P1_R1138_U354
g16614 nand P1_R1138_U295 P1_R1138_U173 ; P1_R1138_U355
g16615 nand P1_R1138_U326 P1_R1138_U81 ; P1_R1138_U356
g16616 nand P1_R1138_U279 P1_R1138_U78 ; P1_R1138_U357
g16617 nand P1_R1138_U333 P1_R1138_U60 ; P1_R1138_U358
g16618 nand P1_R1138_U342 P1_R1138_U169 ; P1_R1138_U359
g16619 nand P1_R1138_U247 P1_R1138_U69 ; P1_R1138_U360
g16620 nand P1_U4017 P1_U3054 ; P1_R1138_U361
g16621 nand P1_R1138_U293 P1_R1138_U165 ; P1_R1138_U362
g16622 nand P1_U3057 P1_R1138_U292 ; P1_R1138_U363
g16623 nand P1_U4019 P1_R1138_U292 ; P1_R1138_U364
g16624 nand P1_R1138_U293 P1_R1138_U165 P1_R1138_U298 ; P1_R1138_U365
g16625 nand P1_R1138_U151 P1_R1138_U165 P1_R1138_U132 ; P1_R1138_U366
g16626 nand P1_R1138_U294 P1_R1138_U298 ; P1_R1138_U367
g16627 nand P1_U3083 P1_R1138_U40 ; P1_R1138_U368
g16628 nand P1_U3485 P1_R1138_U39 ; P1_R1138_U369
g16629 nand P1_R1138_U369 P1_R1138_U368 ; P1_R1138_U370
g16630 nand P1_R1138_U349 P1_R1138_U41 ; P1_R1138_U371
g16631 nand P1_R1138_U370 P1_R1138_U203 ; P1_R1138_U372
g16632 nand P1_U3084 P1_R1138_U37 ; P1_R1138_U373
g16633 nand P1_U3482 P1_R1138_U38 ; P1_R1138_U374
g16634 nand P1_R1138_U374 P1_R1138_U373 ; P1_R1138_U375
g16635 nand P1_R1138_U350 P1_R1138_U140 ; P1_R1138_U376
g16636 nand P1_R1138_U200 P1_R1138_U375 ; P1_R1138_U377
g16637 nand P1_U3070 P1_R1138_U24 ; P1_R1138_U378
g16638 nand P1_U3479 P1_R1138_U22 ; P1_R1138_U379
g16639 nand P1_U3071 P1_R1138_U20 ; P1_R1138_U380
g16640 nand P1_U3476 P1_R1138_U21 ; P1_R1138_U381
g16641 nand P1_R1138_U381 P1_R1138_U380 ; P1_R1138_U382
g16642 nand P1_R1138_U351 P1_R1138_U42 ; P1_R1138_U383
g16643 nand P1_R1138_U382 P1_R1138_U192 ; P1_R1138_U384
g16644 nand P1_U3067 P1_R1138_U36 ; P1_R1138_U385
g16645 nand P1_U3473 P1_R1138_U27 ; P1_R1138_U386
g16646 nand P1_U3060 P1_R1138_U25 ; P1_R1138_U387
g16647 nand P1_U3470 P1_R1138_U26 ; P1_R1138_U388
g16648 nand P1_R1138_U388 P1_R1138_U387 ; P1_R1138_U389
g16649 nand P1_R1138_U352 P1_R1138_U45 ; P1_R1138_U390
g16650 nand P1_R1138_U389 P1_R1138_U218 ; P1_R1138_U391
g16651 nand P1_U3064 P1_R1138_U33 ; P1_R1138_U392
g16652 nand P1_U3467 P1_R1138_U34 ; P1_R1138_U393
g16653 nand P1_R1138_U393 P1_R1138_U392 ; P1_R1138_U394
g16654 nand P1_R1138_U353 P1_R1138_U141 ; P1_R1138_U395
g16655 nand P1_R1138_U227 P1_R1138_U394 ; P1_R1138_U396
g16656 nand P1_U3068 P1_R1138_U28 ; P1_R1138_U397
g16657 nand P1_U3464 P1_R1138_U29 ; P1_R1138_U398
g16658 nand P1_U3055 P1_R1138_U143 ; P1_R1138_U399
g16659 nand P1_U4028 P1_R1138_U142 ; P1_R1138_U400
g16660 nand P1_U3055 P1_R1138_U143 ; P1_R1138_U401
g16661 nand P1_U4028 P1_R1138_U142 ; P1_R1138_U402
g16662 nand P1_R1138_U402 P1_R1138_U401 ; P1_R1138_U403
g16663 nand P1_R1138_U144 P1_R1138_U145 ; P1_R1138_U404
g16664 nand P1_R1138_U302 P1_R1138_U403 ; P1_R1138_U405
g16665 nand P1_U3054 P1_R1138_U89 ; P1_R1138_U406
g16666 nand P1_U4017 P1_R1138_U88 ; P1_R1138_U407
g16667 nand P1_U3054 P1_R1138_U89 ; P1_R1138_U408
g16668 nand P1_U4017 P1_R1138_U88 ; P1_R1138_U409
g16669 nand P1_R1138_U409 P1_R1138_U408 ; P1_R1138_U410
g16670 nand P1_R1138_U146 P1_R1138_U147 ; P1_R1138_U411
g16671 nand P1_R1138_U300 P1_R1138_U410 ; P1_R1138_U412
g16672 nand P1_U3053 P1_R1138_U47 ; P1_R1138_U413
g16673 nand P1_U4018 P1_R1138_U48 ; P1_R1138_U414
g16674 nand P1_U3053 P1_R1138_U47 ; P1_R1138_U415
g16675 nand P1_U4018 P1_R1138_U48 ; P1_R1138_U416
g16676 nand P1_R1138_U416 P1_R1138_U415 ; P1_R1138_U417
g16677 nand P1_R1138_U148 P1_R1138_U149 ; P1_R1138_U418
g16678 nand P1_R1138_U297 P1_R1138_U417 ; P1_R1138_U419
g16679 nand P1_U3057 P1_R1138_U50 ; P1_R1138_U420
g16680 nand P1_U4019 P1_R1138_U49 ; P1_R1138_U421
g16681 nand P1_U3058 P1_R1138_U51 ; P1_R1138_U422
g16682 nand P1_U4020 P1_R1138_U52 ; P1_R1138_U423
g16683 nand P1_R1138_U423 P1_R1138_U422 ; P1_R1138_U424
g16684 nand P1_R1138_U354 P1_R1138_U90 ; P1_R1138_U425
g16685 nand P1_R1138_U424 P1_R1138_U304 ; P1_R1138_U426
g16686 nand P1_U3065 P1_R1138_U53 ; P1_R1138_U427
g16687 nand P1_U4021 P1_R1138_U54 ; P1_R1138_U428
g16688 nand P1_R1138_U428 P1_R1138_U427 ; P1_R1138_U429
g16689 nand P1_R1138_U355 P1_R1138_U151 ; P1_R1138_U430
g16690 nand P1_R1138_U291 P1_R1138_U429 ; P1_R1138_U431
g16691 nand P1_U3066 P1_R1138_U85 ; P1_R1138_U432
g16692 nand P1_U4022 P1_R1138_U86 ; P1_R1138_U433
g16693 nand P1_U3066 P1_R1138_U85 ; P1_R1138_U434
g16694 nand P1_U4022 P1_R1138_U86 ; P1_R1138_U435
g16695 nand P1_R1138_U435 P1_R1138_U434 ; P1_R1138_U436
g16696 nand P1_R1138_U152 P1_R1138_U153 ; P1_R1138_U437
g16697 nand P1_R1138_U287 P1_R1138_U436 ; P1_R1138_U438
g16698 nand P1_U3061 P1_R1138_U83 ; P1_R1138_U439
g16699 nand P1_U4023 P1_R1138_U84 ; P1_R1138_U440
g16700 nand P1_U3061 P1_R1138_U83 ; P1_R1138_U441
g16701 nand P1_U4023 P1_R1138_U84 ; P1_R1138_U442
g16702 nand P1_R1138_U442 P1_R1138_U441 ; P1_R1138_U443
g16703 nand P1_R1138_U154 P1_R1138_U155 ; P1_R1138_U444
g16704 nand P1_R1138_U283 P1_R1138_U443 ; P1_R1138_U445
g16705 nand P1_U3075 P1_R1138_U55 ; P1_R1138_U446
g16706 nand P1_U4024 P1_R1138_U56 ; P1_R1138_U447
g16707 nand P1_U3075 P1_R1138_U55 ; P1_R1138_U448
g16708 nand P1_U4024 P1_R1138_U56 ; P1_R1138_U449
g16709 nand P1_R1138_U449 P1_R1138_U448 ; P1_R1138_U450
g16710 nand P1_U3076 P1_R1138_U82 ; P1_R1138_U451
g16711 nand P1_U4025 P1_R1138_U91 ; P1_R1138_U452
g16712 nand P1_R1138_U179 P1_R1138_U158 ; P1_R1138_U453
g16713 nand P1_R1138_U325 P1_R1138_U32 ; P1_R1138_U454
g16714 nand P1_U3081 P1_R1138_U79 ; P1_R1138_U455
g16715 nand P1_U3514 P1_R1138_U80 ; P1_R1138_U456
g16716 nand P1_R1138_U456 P1_R1138_U455 ; P1_R1138_U457
g16717 nand P1_R1138_U356 P1_R1138_U92 ; P1_R1138_U458
g16718 nand P1_R1138_U457 P1_R1138_U313 ; P1_R1138_U459
g16719 nand P1_U3082 P1_R1138_U76 ; P1_R1138_U460
g16720 nand P1_U3512 P1_R1138_U77 ; P1_R1138_U461
g16721 nand P1_R1138_U461 P1_R1138_U460 ; P1_R1138_U462
g16722 nand P1_R1138_U357 P1_R1138_U159 ; P1_R1138_U463
g16723 nand P1_R1138_U267 P1_R1138_U462 ; P1_R1138_U464
g16724 nand P1_U3069 P1_R1138_U61 ; P1_R1138_U465
g16725 nand P1_U3509 P1_R1138_U59 ; P1_R1138_U466
g16726 nand P1_U3073 P1_R1138_U57 ; P1_R1138_U467
g16727 nand P1_U3506 P1_R1138_U58 ; P1_R1138_U468
g16728 nand P1_R1138_U468 P1_R1138_U467 ; P1_R1138_U469
g16729 nand P1_R1138_U358 P1_R1138_U93 ; P1_R1138_U470
g16730 nand P1_R1138_U469 P1_R1138_U259 ; P1_R1138_U471
g16731 nand P1_U3074 P1_R1138_U74 ; P1_R1138_U472
g16732 nand P1_U3503 P1_R1138_U75 ; P1_R1138_U473
g16733 nand P1_U3074 P1_R1138_U74 ; P1_R1138_U474
g16734 nand P1_U3503 P1_R1138_U75 ; P1_R1138_U475
g16735 nand P1_R1138_U475 P1_R1138_U474 ; P1_R1138_U476
g16736 nand P1_R1138_U160 P1_R1138_U161 ; P1_R1138_U477
g16737 nand P1_R1138_U255 P1_R1138_U476 ; P1_R1138_U478
g16738 nand P1_U3079 P1_R1138_U72 ; P1_R1138_U479
g16739 nand P1_U3500 P1_R1138_U73 ; P1_R1138_U480
g16740 nand P1_U3079 P1_R1138_U72 ; P1_R1138_U481
g16741 nand P1_U3500 P1_R1138_U73 ; P1_R1138_U482
g16742 nand P1_R1138_U482 P1_R1138_U481 ; P1_R1138_U483
g16743 nand P1_R1138_U162 P1_R1138_U163 ; P1_R1138_U484
g16744 nand P1_R1138_U251 P1_R1138_U483 ; P1_R1138_U485
g16745 nand P1_U3080 P1_R1138_U70 ; P1_R1138_U486
g16746 nand P1_U3497 P1_R1138_U71 ; P1_R1138_U487
g16747 nand P1_U3072 P1_R1138_U65 ; P1_R1138_U488
g16748 nand P1_U3494 P1_R1138_U66 ; P1_R1138_U489
g16749 nand P1_R1138_U489 P1_R1138_U488 ; P1_R1138_U490
g16750 nand P1_R1138_U359 P1_R1138_U94 ; P1_R1138_U491
g16751 nand P1_R1138_U490 P1_R1138_U335 ; P1_R1138_U492
g16752 nand P1_U3063 P1_R1138_U67 ; P1_R1138_U493
g16753 nand P1_U3491 P1_R1138_U68 ; P1_R1138_U494
g16754 nand P1_R1138_U494 P1_R1138_U493 ; P1_R1138_U495
g16755 nand P1_R1138_U360 P1_R1138_U164 ; P1_R1138_U496
g16756 nand P1_R1138_U241 P1_R1138_U495 ; P1_R1138_U497
g16757 nand P1_U3062 P1_R1138_U63 ; P1_R1138_U498
g16758 nand P1_U3488 P1_R1138_U64 ; P1_R1138_U499
g16759 nand P1_U3077 P1_R1138_U30 ; P1_R1138_U500
g16760 nand P1_U3456 P1_R1138_U31 ; P1_R1138_U501
g16761 and P1_R1222_U176 P1_R1222_U175 ; P1_R1222_U4
g16762 and P1_R1222_U177 P1_R1222_U178 ; P1_R1222_U5
g16763 and P1_R1222_U194 P1_R1222_U193 ; P1_R1222_U6
g16764 and P1_R1222_U234 P1_R1222_U233 ; P1_R1222_U7
g16765 and P1_R1222_U243 P1_R1222_U242 ; P1_R1222_U8
g16766 and P1_R1222_U261 P1_R1222_U260 ; P1_R1222_U9
g16767 and P1_R1222_U269 P1_R1222_U268 ; P1_R1222_U10
g16768 and P1_R1222_U348 P1_R1222_U345 ; P1_R1222_U11
g16769 and P1_R1222_U341 P1_R1222_U338 ; P1_R1222_U12
g16770 and P1_R1222_U332 P1_R1222_U329 ; P1_R1222_U13
g16771 and P1_R1222_U323 P1_R1222_U320 ; P1_R1222_U14
g16772 and P1_R1222_U317 P1_R1222_U315 ; P1_R1222_U15
g16773 and P1_R1222_U310 P1_R1222_U307 ; P1_R1222_U16
g16774 and P1_R1222_U232 P1_R1222_U229 ; P1_R1222_U17
g16775 and P1_R1222_U224 P1_R1222_U221 ; P1_R1222_U18
g16776 and P1_R1222_U210 P1_R1222_U207 ; P1_R1222_U19
g16777 not P1_U3476 ; P1_R1222_U20
g16778 not P1_U3071 ; P1_R1222_U21
g16779 not P1_U3070 ; P1_R1222_U22
g16780 nand P1_U3071 P1_U3476 ; P1_R1222_U23
g16781 not P1_U3479 ; P1_R1222_U24
g16782 not P1_U3470 ; P1_R1222_U25
g16783 not P1_U3060 ; P1_R1222_U26
g16784 not P1_U3067 ; P1_R1222_U27
g16785 not P1_U3464 ; P1_R1222_U28
g16786 not P1_U3068 ; P1_R1222_U29
g16787 not P1_U3456 ; P1_R1222_U30
g16788 not P1_U3077 ; P1_R1222_U31
g16789 nand P1_U3077 P1_U3456 ; P1_R1222_U32
g16790 not P1_U3467 ; P1_R1222_U33
g16791 not P1_U3064 ; P1_R1222_U34
g16792 nand P1_U3060 P1_U3470 ; P1_R1222_U35
g16793 not P1_U3473 ; P1_R1222_U36
g16794 not P1_U3482 ; P1_R1222_U37
g16795 not P1_U3084 ; P1_R1222_U38
g16796 not P1_U3083 ; P1_R1222_U39
g16797 not P1_U3485 ; P1_R1222_U40
g16798 nand P1_R1222_U62 P1_R1222_U202 ; P1_R1222_U41
g16799 nand P1_R1222_U118 P1_R1222_U190 ; P1_R1222_U42
g16800 nand P1_R1222_U179 P1_R1222_U180 ; P1_R1222_U43
g16801 nand P1_U3461 P1_U3078 ; P1_R1222_U44
g16802 nand P1_R1222_U122 P1_R1222_U216 ; P1_R1222_U45
g16803 nand P1_R1222_U213 P1_R1222_U212 ; P1_R1222_U46
g16804 not P1_U4018 ; P1_R1222_U47
g16805 not P1_U3053 ; P1_R1222_U48
g16806 not P1_U3057 ; P1_R1222_U49
g16807 not P1_U4019 ; P1_R1222_U50
g16808 not P1_U4020 ; P1_R1222_U51
g16809 not P1_U3058 ; P1_R1222_U52
g16810 not P1_U4021 ; P1_R1222_U53
g16811 not P1_U3065 ; P1_R1222_U54
g16812 not P1_U4024 ; P1_R1222_U55
g16813 not P1_U3075 ; P1_R1222_U56
g16814 not P1_U3506 ; P1_R1222_U57
g16815 not P1_U3073 ; P1_R1222_U58
g16816 not P1_U3069 ; P1_R1222_U59
g16817 nand P1_U3073 P1_U3506 ; P1_R1222_U60
g16818 not P1_U3509 ; P1_R1222_U61
g16819 nand P1_U3084 P1_U3482 ; P1_R1222_U62
g16820 not P1_U3488 ; P1_R1222_U63
g16821 not P1_U3062 ; P1_R1222_U64
g16822 not P1_U3494 ; P1_R1222_U65
g16823 not P1_U3072 ; P1_R1222_U66
g16824 not P1_U3491 ; P1_R1222_U67
g16825 not P1_U3063 ; P1_R1222_U68
g16826 nand P1_U3063 P1_U3491 ; P1_R1222_U69
g16827 not P1_U3497 ; P1_R1222_U70
g16828 not P1_U3080 ; P1_R1222_U71
g16829 not P1_U3500 ; P1_R1222_U72
g16830 not P1_U3079 ; P1_R1222_U73
g16831 not P1_U3503 ; P1_R1222_U74
g16832 not P1_U3074 ; P1_R1222_U75
g16833 not P1_U3512 ; P1_R1222_U76
g16834 not P1_U3082 ; P1_R1222_U77
g16835 nand P1_U3082 P1_U3512 ; P1_R1222_U78
g16836 not P1_U3514 ; P1_R1222_U79
g16837 not P1_U3081 ; P1_R1222_U80
g16838 nand P1_U3081 P1_U3514 ; P1_R1222_U81
g16839 not P1_U4025 ; P1_R1222_U82
g16840 not P1_U4023 ; P1_R1222_U83
g16841 not P1_U3061 ; P1_R1222_U84
g16842 not P1_U4022 ; P1_R1222_U85
g16843 not P1_U3066 ; P1_R1222_U86
g16844 nand P1_U4019 P1_U3057 ; P1_R1222_U87
g16845 not P1_U3054 ; P1_R1222_U88
g16846 not P1_U4017 ; P1_R1222_U89
g16847 nand P1_R1222_U303 P1_R1222_U173 ; P1_R1222_U90
g16848 not P1_U3076 ; P1_R1222_U91
g16849 nand P1_R1222_U78 P1_R1222_U312 ; P1_R1222_U92
g16850 nand P1_R1222_U258 P1_R1222_U257 ; P1_R1222_U93
g16851 nand P1_R1222_U69 P1_R1222_U334 ; P1_R1222_U94
g16852 nand P1_R1222_U454 P1_R1222_U453 ; P1_R1222_U95
g16853 nand P1_R1222_U501 P1_R1222_U500 ; P1_R1222_U96
g16854 nand P1_R1222_U372 P1_R1222_U371 ; P1_R1222_U97
g16855 nand P1_R1222_U377 P1_R1222_U376 ; P1_R1222_U98
g16856 nand P1_R1222_U384 P1_R1222_U383 ; P1_R1222_U99
g16857 nand P1_R1222_U391 P1_R1222_U390 ; P1_R1222_U100
g16858 nand P1_R1222_U396 P1_R1222_U395 ; P1_R1222_U101
g16859 nand P1_R1222_U405 P1_R1222_U404 ; P1_R1222_U102
g16860 nand P1_R1222_U412 P1_R1222_U411 ; P1_R1222_U103
g16861 nand P1_R1222_U419 P1_R1222_U418 ; P1_R1222_U104
g16862 nand P1_R1222_U426 P1_R1222_U425 ; P1_R1222_U105
g16863 nand P1_R1222_U431 P1_R1222_U430 ; P1_R1222_U106
g16864 nand P1_R1222_U438 P1_R1222_U437 ; P1_R1222_U107
g16865 nand P1_R1222_U445 P1_R1222_U444 ; P1_R1222_U108
g16866 nand P1_R1222_U459 P1_R1222_U458 ; P1_R1222_U109
g16867 nand P1_R1222_U464 P1_R1222_U463 ; P1_R1222_U110
g16868 nand P1_R1222_U471 P1_R1222_U470 ; P1_R1222_U111
g16869 nand P1_R1222_U478 P1_R1222_U477 ; P1_R1222_U112
g16870 nand P1_R1222_U485 P1_R1222_U484 ; P1_R1222_U113
g16871 nand P1_R1222_U492 P1_R1222_U491 ; P1_R1222_U114
g16872 nand P1_R1222_U497 P1_R1222_U496 ; P1_R1222_U115
g16873 and P1_U3464 P1_U3068 ; P1_R1222_U116
g16874 and P1_R1222_U186 P1_R1222_U184 ; P1_R1222_U117
g16875 and P1_R1222_U191 P1_R1222_U189 ; P1_R1222_U118
g16876 and P1_R1222_U198 P1_R1222_U197 ; P1_R1222_U119
g16877 and P1_R1222_U379 P1_R1222_U378 P1_R1222_U23 ; P1_R1222_U120
g16878 and P1_R1222_U209 P1_R1222_U6 ; P1_R1222_U121
g16879 and P1_R1222_U217 P1_R1222_U215 ; P1_R1222_U122
g16880 and P1_R1222_U386 P1_R1222_U385 P1_R1222_U35 ; P1_R1222_U123
g16881 and P1_R1222_U223 P1_R1222_U4 ; P1_R1222_U124
g16882 and P1_R1222_U231 P1_R1222_U178 ; P1_R1222_U125
g16883 and P1_R1222_U201 P1_R1222_U7 ; P1_R1222_U126
g16884 and P1_R1222_U236 P1_R1222_U168 ; P1_R1222_U127
g16885 and P1_R1222_U245 P1_R1222_U169 ; P1_R1222_U128
g16886 and P1_R1222_U265 P1_R1222_U264 ; P1_R1222_U129
g16887 and P1_R1222_U10 P1_R1222_U279 ; P1_R1222_U130
g16888 and P1_R1222_U282 P1_R1222_U277 ; P1_R1222_U131
g16889 and P1_R1222_U298 P1_R1222_U295 ; P1_R1222_U132
g16890 and P1_R1222_U365 P1_R1222_U299 ; P1_R1222_U133
g16891 and P1_R1222_U156 P1_R1222_U275 ; P1_R1222_U134
g16892 and P1_R1222_U466 P1_R1222_U465 P1_R1222_U60 ; P1_R1222_U135
g16893 and P1_R1222_U487 P1_R1222_U486 P1_R1222_U169 ; P1_R1222_U136
g16894 and P1_R1222_U340 P1_R1222_U8 ; P1_R1222_U137
g16895 and P1_R1222_U499 P1_R1222_U498 P1_R1222_U168 ; P1_R1222_U138
g16896 and P1_R1222_U347 P1_R1222_U7 ; P1_R1222_U139
g16897 nand P1_R1222_U119 P1_R1222_U199 ; P1_R1222_U140
g16898 nand P1_R1222_U214 P1_R1222_U226 ; P1_R1222_U141
g16899 not P1_U3055 ; P1_R1222_U142
g16900 not P1_U4028 ; P1_R1222_U143
g16901 and P1_R1222_U400 P1_R1222_U399 ; P1_R1222_U144
g16902 nand P1_R1222_U301 P1_R1222_U166 P1_R1222_U361 ; P1_R1222_U145
g16903 and P1_R1222_U407 P1_R1222_U406 ; P1_R1222_U146
g16904 nand P1_R1222_U367 P1_R1222_U366 P1_R1222_U133 ; P1_R1222_U147
g16905 and P1_R1222_U414 P1_R1222_U413 ; P1_R1222_U148
g16906 nand P1_R1222_U362 P1_R1222_U296 P1_R1222_U87 ; P1_R1222_U149
g16907 and P1_R1222_U421 P1_R1222_U420 ; P1_R1222_U150
g16908 nand P1_R1222_U290 P1_R1222_U289 ; P1_R1222_U151
g16909 and P1_R1222_U433 P1_R1222_U432 ; P1_R1222_U152
g16910 nand P1_R1222_U286 P1_R1222_U285 ; P1_R1222_U153
g16911 and P1_R1222_U440 P1_R1222_U439 ; P1_R1222_U154
g16912 nand P1_R1222_U131 P1_R1222_U281 ; P1_R1222_U155
g16913 and P1_R1222_U447 P1_R1222_U446 ; P1_R1222_U156
g16914 and P1_R1222_U452 P1_R1222_U451 ; P1_R1222_U157
g16915 nand P1_R1222_U44 P1_R1222_U324 ; P1_R1222_U158
g16916 nand P1_R1222_U129 P1_R1222_U266 ; P1_R1222_U159
g16917 and P1_R1222_U473 P1_R1222_U472 ; P1_R1222_U160
g16918 nand P1_R1222_U254 P1_R1222_U253 ; P1_R1222_U161
g16919 and P1_R1222_U480 P1_R1222_U479 ; P1_R1222_U162
g16920 nand P1_R1222_U250 P1_R1222_U249 ; P1_R1222_U163
g16921 nand P1_R1222_U240 P1_R1222_U239 ; P1_R1222_U164
g16922 nand P1_R1222_U364 P1_R1222_U363 ; P1_R1222_U165
g16923 nand P1_U3054 P1_R1222_U147 ; P1_R1222_U166
g16924 not P1_R1222_U35 ; P1_R1222_U167
g16925 nand P1_U3485 P1_U3083 ; P1_R1222_U168
g16926 nand P1_U3072 P1_U3494 ; P1_R1222_U169
g16927 nand P1_U3058 P1_U4020 ; P1_R1222_U170
g16928 not P1_R1222_U69 ; P1_R1222_U171
g16929 not P1_R1222_U78 ; P1_R1222_U172
g16930 nand P1_U3065 P1_U4021 ; P1_R1222_U173
g16931 not P1_R1222_U62 ; P1_R1222_U174
g16932 or P1_U3067 P1_U3473 ; P1_R1222_U175
g16933 or P1_U3060 P1_U3470 ; P1_R1222_U176
g16934 or P1_U3467 P1_U3064 ; P1_R1222_U177
g16935 or P1_U3464 P1_U3068 ; P1_R1222_U178
g16936 not P1_R1222_U32 ; P1_R1222_U179
g16937 or P1_U3461 P1_U3078 ; P1_R1222_U180
g16938 not P1_R1222_U43 ; P1_R1222_U181
g16939 not P1_R1222_U44 ; P1_R1222_U182
g16940 nand P1_R1222_U43 P1_R1222_U44 ; P1_R1222_U183
g16941 nand P1_R1222_U116 P1_R1222_U177 ; P1_R1222_U184
g16942 nand P1_R1222_U5 P1_R1222_U183 ; P1_R1222_U185
g16943 nand P1_U3064 P1_U3467 ; P1_R1222_U186
g16944 nand P1_R1222_U117 P1_R1222_U185 ; P1_R1222_U187
g16945 nand P1_R1222_U36 P1_R1222_U35 ; P1_R1222_U188
g16946 nand P1_U3067 P1_R1222_U188 ; P1_R1222_U189
g16947 nand P1_R1222_U4 P1_R1222_U187 ; P1_R1222_U190
g16948 nand P1_U3473 P1_R1222_U167 ; P1_R1222_U191
g16949 not P1_R1222_U42 ; P1_R1222_U192
g16950 or P1_U3070 P1_U3479 ; P1_R1222_U193
g16951 or P1_U3071 P1_U3476 ; P1_R1222_U194
g16952 not P1_R1222_U23 ; P1_R1222_U195
g16953 nand P1_R1222_U24 P1_R1222_U23 ; P1_R1222_U196
g16954 nand P1_U3070 P1_R1222_U196 ; P1_R1222_U197
g16955 nand P1_U3479 P1_R1222_U195 ; P1_R1222_U198
g16956 nand P1_R1222_U6 P1_R1222_U42 ; P1_R1222_U199
g16957 not P1_R1222_U140 ; P1_R1222_U200
g16958 or P1_U3482 P1_U3084 ; P1_R1222_U201
g16959 nand P1_R1222_U201 P1_R1222_U140 ; P1_R1222_U202
g16960 not P1_R1222_U41 ; P1_R1222_U203
g16961 or P1_U3083 P1_U3485 ; P1_R1222_U204
g16962 or P1_U3476 P1_U3071 ; P1_R1222_U205
g16963 nand P1_R1222_U205 P1_R1222_U42 ; P1_R1222_U206
g16964 nand P1_R1222_U120 P1_R1222_U206 ; P1_R1222_U207
g16965 nand P1_R1222_U192 P1_R1222_U23 ; P1_R1222_U208
g16966 nand P1_U3479 P1_U3070 ; P1_R1222_U209
g16967 nand P1_R1222_U121 P1_R1222_U208 ; P1_R1222_U210
g16968 or P1_U3071 P1_U3476 ; P1_R1222_U211
g16969 nand P1_R1222_U182 P1_R1222_U178 ; P1_R1222_U212
g16970 nand P1_U3068 P1_U3464 ; P1_R1222_U213
g16971 not P1_R1222_U46 ; P1_R1222_U214
g16972 nand P1_R1222_U181 P1_R1222_U5 ; P1_R1222_U215
g16973 nand P1_R1222_U46 P1_R1222_U177 ; P1_R1222_U216
g16974 nand P1_U3064 P1_U3467 ; P1_R1222_U217
g16975 not P1_R1222_U45 ; P1_R1222_U218
g16976 or P1_U3470 P1_U3060 ; P1_R1222_U219
g16977 nand P1_R1222_U219 P1_R1222_U45 ; P1_R1222_U220
g16978 nand P1_R1222_U123 P1_R1222_U220 ; P1_R1222_U221
g16979 nand P1_R1222_U218 P1_R1222_U35 ; P1_R1222_U222
g16980 nand P1_U3473 P1_U3067 ; P1_R1222_U223
g16981 nand P1_R1222_U124 P1_R1222_U222 ; P1_R1222_U224
g16982 or P1_U3060 P1_U3470 ; P1_R1222_U225
g16983 nand P1_R1222_U181 P1_R1222_U178 ; P1_R1222_U226
g16984 not P1_R1222_U141 ; P1_R1222_U227
g16985 nand P1_U3064 P1_U3467 ; P1_R1222_U228
g16986 nand P1_R1222_U398 P1_R1222_U397 P1_R1222_U44 P1_R1222_U43 ; P1_R1222_U229
g16987 nand P1_R1222_U44 P1_R1222_U43 ; P1_R1222_U230
g16988 nand P1_U3068 P1_U3464 ; P1_R1222_U231
g16989 nand P1_R1222_U125 P1_R1222_U230 ; P1_R1222_U232
g16990 or P1_U3083 P1_U3485 ; P1_R1222_U233
g16991 or P1_U3062 P1_U3488 ; P1_R1222_U234
g16992 nand P1_R1222_U174 P1_R1222_U7 ; P1_R1222_U235
g16993 nand P1_U3062 P1_U3488 ; P1_R1222_U236
g16994 nand P1_R1222_U127 P1_R1222_U235 ; P1_R1222_U237
g16995 or P1_U3488 P1_U3062 ; P1_R1222_U238
g16996 nand P1_R1222_U126 P1_R1222_U140 ; P1_R1222_U239
g16997 nand P1_R1222_U238 P1_R1222_U237 ; P1_R1222_U240
g16998 not P1_R1222_U164 ; P1_R1222_U241
g16999 or P1_U3080 P1_U3497 ; P1_R1222_U242
g17000 or P1_U3072 P1_U3494 ; P1_R1222_U243
g17001 nand P1_R1222_U171 P1_R1222_U8 ; P1_R1222_U244
g17002 nand P1_U3080 P1_U3497 ; P1_R1222_U245
g17003 nand P1_R1222_U128 P1_R1222_U244 ; P1_R1222_U246
g17004 or P1_U3491 P1_U3063 ; P1_R1222_U247
g17005 or P1_U3497 P1_U3080 ; P1_R1222_U248
g17006 nand P1_R1222_U247 P1_R1222_U164 P1_R1222_U8 ; P1_R1222_U249
g17007 nand P1_R1222_U248 P1_R1222_U246 ; P1_R1222_U250
g17008 not P1_R1222_U163 ; P1_R1222_U251
g17009 or P1_U3500 P1_U3079 ; P1_R1222_U252
g17010 nand P1_R1222_U252 P1_R1222_U163 ; P1_R1222_U253
g17011 nand P1_U3079 P1_U3500 ; P1_R1222_U254
g17012 not P1_R1222_U161 ; P1_R1222_U255
g17013 or P1_U3503 P1_U3074 ; P1_R1222_U256
g17014 nand P1_R1222_U256 P1_R1222_U161 ; P1_R1222_U257
g17015 nand P1_U3074 P1_U3503 ; P1_R1222_U258
g17016 not P1_R1222_U93 ; P1_R1222_U259
g17017 or P1_U3069 P1_U3509 ; P1_R1222_U260
g17018 or P1_U3073 P1_U3506 ; P1_R1222_U261
g17019 not P1_R1222_U60 ; P1_R1222_U262
g17020 nand P1_R1222_U61 P1_R1222_U60 ; P1_R1222_U263
g17021 nand P1_U3069 P1_R1222_U263 ; P1_R1222_U264
g17022 nand P1_U3509 P1_R1222_U262 ; P1_R1222_U265
g17023 nand P1_R1222_U9 P1_R1222_U93 ; P1_R1222_U266
g17024 not P1_R1222_U159 ; P1_R1222_U267
g17025 or P1_U3076 P1_U4025 ; P1_R1222_U268
g17026 or P1_U3081 P1_U3514 ; P1_R1222_U269
g17027 or P1_U3075 P1_U4024 ; P1_R1222_U270
g17028 not P1_R1222_U81 ; P1_R1222_U271
g17029 nand P1_U4025 P1_R1222_U271 ; P1_R1222_U272
g17030 nand P1_R1222_U272 P1_R1222_U91 ; P1_R1222_U273
g17031 nand P1_R1222_U81 P1_R1222_U82 ; P1_R1222_U274
g17032 nand P1_R1222_U274 P1_R1222_U273 ; P1_R1222_U275
g17033 nand P1_R1222_U172 P1_R1222_U10 ; P1_R1222_U276
g17034 nand P1_U3075 P1_U4024 ; P1_R1222_U277
g17035 nand P1_R1222_U275 P1_R1222_U276 ; P1_R1222_U278
g17036 or P1_U3512 P1_U3082 ; P1_R1222_U279
g17037 or P1_U4024 P1_U3075 ; P1_R1222_U280
g17038 nand P1_R1222_U270 P1_R1222_U159 P1_R1222_U130 ; P1_R1222_U281
g17039 nand P1_R1222_U280 P1_R1222_U278 ; P1_R1222_U282
g17040 not P1_R1222_U155 ; P1_R1222_U283
g17041 or P1_U4023 P1_U3061 ; P1_R1222_U284
g17042 nand P1_R1222_U284 P1_R1222_U155 ; P1_R1222_U285
g17043 nand P1_U3061 P1_U4023 ; P1_R1222_U286
g17044 not P1_R1222_U153 ; P1_R1222_U287
g17045 or P1_U4022 P1_U3066 ; P1_R1222_U288
g17046 nand P1_R1222_U288 P1_R1222_U153 ; P1_R1222_U289
g17047 nand P1_U3066 P1_U4022 ; P1_R1222_U290
g17048 not P1_R1222_U151 ; P1_R1222_U291
g17049 or P1_U3058 P1_U4020 ; P1_R1222_U292
g17050 nand P1_R1222_U173 P1_R1222_U170 ; P1_R1222_U293
g17051 not P1_R1222_U87 ; P1_R1222_U294
g17052 or P1_U4021 P1_U3065 ; P1_R1222_U295
g17053 nand P1_R1222_U151 P1_R1222_U295 P1_R1222_U165 ; P1_R1222_U296
g17054 not P1_R1222_U149 ; P1_R1222_U297
g17055 or P1_U4018 P1_U3053 ; P1_R1222_U298
g17056 nand P1_U3053 P1_U4018 ; P1_R1222_U299
g17057 not P1_R1222_U147 ; P1_R1222_U300
g17058 nand P1_U4017 P1_R1222_U147 ; P1_R1222_U301
g17059 not P1_R1222_U145 ; P1_R1222_U302
g17060 nand P1_R1222_U295 P1_R1222_U151 ; P1_R1222_U303
g17061 not P1_R1222_U90 ; P1_R1222_U304
g17062 or P1_U4020 P1_U3058 ; P1_R1222_U305
g17063 nand P1_R1222_U305 P1_R1222_U90 ; P1_R1222_U306
g17064 nand P1_R1222_U306 P1_R1222_U170 P1_R1222_U150 ; P1_R1222_U307
g17065 nand P1_R1222_U304 P1_R1222_U170 ; P1_R1222_U308
g17066 nand P1_U4019 P1_U3057 ; P1_R1222_U309
g17067 nand P1_R1222_U308 P1_R1222_U309 P1_R1222_U165 ; P1_R1222_U310
g17068 or P1_U3058 P1_U4020 ; P1_R1222_U311
g17069 nand P1_R1222_U279 P1_R1222_U159 ; P1_R1222_U312
g17070 not P1_R1222_U92 ; P1_R1222_U313
g17071 nand P1_R1222_U10 P1_R1222_U92 ; P1_R1222_U314
g17072 nand P1_R1222_U134 P1_R1222_U314 ; P1_R1222_U315
g17073 nand P1_R1222_U314 P1_R1222_U275 ; P1_R1222_U316
g17074 nand P1_R1222_U450 P1_R1222_U316 ; P1_R1222_U317
g17075 or P1_U3514 P1_U3081 ; P1_R1222_U318
g17076 nand P1_R1222_U318 P1_R1222_U92 ; P1_R1222_U319
g17077 nand P1_R1222_U319 P1_R1222_U81 P1_R1222_U157 ; P1_R1222_U320
g17078 nand P1_R1222_U313 P1_R1222_U81 ; P1_R1222_U321
g17079 nand P1_U3076 P1_U4025 ; P1_R1222_U322
g17080 nand P1_R1222_U322 P1_R1222_U321 P1_R1222_U10 ; P1_R1222_U323
g17081 or P1_U3461 P1_U3078 ; P1_R1222_U324
g17082 not P1_R1222_U158 ; P1_R1222_U325
g17083 or P1_U3081 P1_U3514 ; P1_R1222_U326
g17084 or P1_U3506 P1_U3073 ; P1_R1222_U327
g17085 nand P1_R1222_U327 P1_R1222_U93 ; P1_R1222_U328
g17086 nand P1_R1222_U135 P1_R1222_U328 ; P1_R1222_U329
g17087 nand P1_R1222_U259 P1_R1222_U60 ; P1_R1222_U330
g17088 nand P1_U3509 P1_U3069 ; P1_R1222_U331
g17089 nand P1_R1222_U331 P1_R1222_U330 P1_R1222_U9 ; P1_R1222_U332
g17090 or P1_U3073 P1_U3506 ; P1_R1222_U333
g17091 nand P1_R1222_U247 P1_R1222_U164 ; P1_R1222_U334
g17092 not P1_R1222_U94 ; P1_R1222_U335
g17093 or P1_U3494 P1_U3072 ; P1_R1222_U336
g17094 nand P1_R1222_U336 P1_R1222_U94 ; P1_R1222_U337
g17095 nand P1_R1222_U136 P1_R1222_U337 ; P1_R1222_U338
g17096 nand P1_R1222_U335 P1_R1222_U169 ; P1_R1222_U339
g17097 nand P1_U3080 P1_U3497 ; P1_R1222_U340
g17098 nand P1_R1222_U137 P1_R1222_U339 ; P1_R1222_U341
g17099 or P1_U3072 P1_U3494 ; P1_R1222_U342
g17100 or P1_U3485 P1_U3083 ; P1_R1222_U343
g17101 nand P1_R1222_U343 P1_R1222_U41 ; P1_R1222_U344
g17102 nand P1_R1222_U138 P1_R1222_U344 ; P1_R1222_U345
g17103 nand P1_R1222_U203 P1_R1222_U168 ; P1_R1222_U346
g17104 nand P1_U3062 P1_U3488 ; P1_R1222_U347
g17105 nand P1_R1222_U139 P1_R1222_U346 ; P1_R1222_U348
g17106 nand P1_R1222_U204 P1_R1222_U168 ; P1_R1222_U349
g17107 nand P1_R1222_U201 P1_R1222_U62 ; P1_R1222_U350
g17108 nand P1_R1222_U211 P1_R1222_U23 ; P1_R1222_U351
g17109 nand P1_R1222_U225 P1_R1222_U35 ; P1_R1222_U352
g17110 nand P1_R1222_U228 P1_R1222_U177 ; P1_R1222_U353
g17111 nand P1_R1222_U311 P1_R1222_U170 ; P1_R1222_U354
g17112 nand P1_R1222_U295 P1_R1222_U173 ; P1_R1222_U355
g17113 nand P1_R1222_U326 P1_R1222_U81 ; P1_R1222_U356
g17114 nand P1_R1222_U279 P1_R1222_U78 ; P1_R1222_U357
g17115 nand P1_R1222_U333 P1_R1222_U60 ; P1_R1222_U358
g17116 nand P1_R1222_U342 P1_R1222_U169 ; P1_R1222_U359
g17117 nand P1_R1222_U247 P1_R1222_U69 ; P1_R1222_U360
g17118 nand P1_U4017 P1_U3054 ; P1_R1222_U361
g17119 nand P1_R1222_U293 P1_R1222_U165 ; P1_R1222_U362
g17120 nand P1_U3057 P1_R1222_U292 ; P1_R1222_U363
g17121 nand P1_U4019 P1_R1222_U292 ; P1_R1222_U364
g17122 nand P1_R1222_U293 P1_R1222_U165 P1_R1222_U298 ; P1_R1222_U365
g17123 nand P1_R1222_U151 P1_R1222_U165 P1_R1222_U132 ; P1_R1222_U366
g17124 nand P1_R1222_U294 P1_R1222_U298 ; P1_R1222_U367
g17125 nand P1_U3083 P1_R1222_U40 ; P1_R1222_U368
g17126 nand P1_U3485 P1_R1222_U39 ; P1_R1222_U369
g17127 nand P1_R1222_U369 P1_R1222_U368 ; P1_R1222_U370
g17128 nand P1_R1222_U349 P1_R1222_U41 ; P1_R1222_U371
g17129 nand P1_R1222_U370 P1_R1222_U203 ; P1_R1222_U372
g17130 nand P1_U3084 P1_R1222_U37 ; P1_R1222_U373
g17131 nand P1_U3482 P1_R1222_U38 ; P1_R1222_U374
g17132 nand P1_R1222_U374 P1_R1222_U373 ; P1_R1222_U375
g17133 nand P1_R1222_U350 P1_R1222_U140 ; P1_R1222_U376
g17134 nand P1_R1222_U200 P1_R1222_U375 ; P1_R1222_U377
g17135 nand P1_U3070 P1_R1222_U24 ; P1_R1222_U378
g17136 nand P1_U3479 P1_R1222_U22 ; P1_R1222_U379
g17137 nand P1_U3071 P1_R1222_U20 ; P1_R1222_U380
g17138 nand P1_U3476 P1_R1222_U21 ; P1_R1222_U381
g17139 nand P1_R1222_U381 P1_R1222_U380 ; P1_R1222_U382
g17140 nand P1_R1222_U351 P1_R1222_U42 ; P1_R1222_U383
g17141 nand P1_R1222_U382 P1_R1222_U192 ; P1_R1222_U384
g17142 nand P1_U3067 P1_R1222_U36 ; P1_R1222_U385
g17143 nand P1_U3473 P1_R1222_U27 ; P1_R1222_U386
g17144 nand P1_U3060 P1_R1222_U25 ; P1_R1222_U387
g17145 nand P1_U3470 P1_R1222_U26 ; P1_R1222_U388
g17146 nand P1_R1222_U388 P1_R1222_U387 ; P1_R1222_U389
g17147 nand P1_R1222_U352 P1_R1222_U45 ; P1_R1222_U390
g17148 nand P1_R1222_U389 P1_R1222_U218 ; P1_R1222_U391
g17149 nand P1_U3064 P1_R1222_U33 ; P1_R1222_U392
g17150 nand P1_U3467 P1_R1222_U34 ; P1_R1222_U393
g17151 nand P1_R1222_U393 P1_R1222_U392 ; P1_R1222_U394
g17152 nand P1_R1222_U353 P1_R1222_U141 ; P1_R1222_U395
g17153 nand P1_R1222_U227 P1_R1222_U394 ; P1_R1222_U396
g17154 nand P1_U3068 P1_R1222_U28 ; P1_R1222_U397
g17155 nand P1_U3464 P1_R1222_U29 ; P1_R1222_U398
g17156 nand P1_U3055 P1_R1222_U143 ; P1_R1222_U399
g17157 nand P1_U4028 P1_R1222_U142 ; P1_R1222_U400
g17158 nand P1_U3055 P1_R1222_U143 ; P1_R1222_U401
g17159 nand P1_U4028 P1_R1222_U142 ; P1_R1222_U402
g17160 nand P1_R1222_U402 P1_R1222_U401 ; P1_R1222_U403
g17161 nand P1_R1222_U144 P1_R1222_U145 ; P1_R1222_U404
g17162 nand P1_R1222_U302 P1_R1222_U403 ; P1_R1222_U405
g17163 nand P1_U3054 P1_R1222_U89 ; P1_R1222_U406
g17164 nand P1_U4017 P1_R1222_U88 ; P1_R1222_U407
g17165 nand P1_U3054 P1_R1222_U89 ; P1_R1222_U408
g17166 nand P1_U4017 P1_R1222_U88 ; P1_R1222_U409
g17167 nand P1_R1222_U409 P1_R1222_U408 ; P1_R1222_U410
g17168 nand P1_R1222_U146 P1_R1222_U147 ; P1_R1222_U411
g17169 nand P1_R1222_U300 P1_R1222_U410 ; P1_R1222_U412
g17170 nand P1_U3053 P1_R1222_U47 ; P1_R1222_U413
g17171 nand P1_U4018 P1_R1222_U48 ; P1_R1222_U414
g17172 nand P1_U3053 P1_R1222_U47 ; P1_R1222_U415
g17173 nand P1_U4018 P1_R1222_U48 ; P1_R1222_U416
g17174 nand P1_R1222_U416 P1_R1222_U415 ; P1_R1222_U417
g17175 nand P1_R1222_U148 P1_R1222_U149 ; P1_R1222_U418
g17176 nand P1_R1222_U297 P1_R1222_U417 ; P1_R1222_U419
g17177 nand P1_U3057 P1_R1222_U50 ; P1_R1222_U420
g17178 nand P1_U4019 P1_R1222_U49 ; P1_R1222_U421
g17179 nand P1_U3058 P1_R1222_U51 ; P1_R1222_U422
g17180 nand P1_U4020 P1_R1222_U52 ; P1_R1222_U423
g17181 nand P1_R1222_U423 P1_R1222_U422 ; P1_R1222_U424
g17182 nand P1_R1222_U354 P1_R1222_U90 ; P1_R1222_U425
g17183 nand P1_R1222_U424 P1_R1222_U304 ; P1_R1222_U426
g17184 nand P1_U3065 P1_R1222_U53 ; P1_R1222_U427
g17185 nand P1_U4021 P1_R1222_U54 ; P1_R1222_U428
g17186 nand P1_R1222_U428 P1_R1222_U427 ; P1_R1222_U429
g17187 nand P1_R1222_U355 P1_R1222_U151 ; P1_R1222_U430
g17188 nand P1_R1222_U291 P1_R1222_U429 ; P1_R1222_U431
g17189 nand P1_U3066 P1_R1222_U85 ; P1_R1222_U432
g17190 nand P1_U4022 P1_R1222_U86 ; P1_R1222_U433
g17191 nand P1_U3066 P1_R1222_U85 ; P1_R1222_U434
g17192 nand P1_U4022 P1_R1222_U86 ; P1_R1222_U435
g17193 nand P1_R1222_U435 P1_R1222_U434 ; P1_R1222_U436
g17194 nand P1_R1222_U152 P1_R1222_U153 ; P1_R1222_U437
g17195 nand P1_R1222_U287 P1_R1222_U436 ; P1_R1222_U438
g17196 nand P1_U3061 P1_R1222_U83 ; P1_R1222_U439
g17197 nand P1_U4023 P1_R1222_U84 ; P1_R1222_U440
g17198 nand P1_U3061 P1_R1222_U83 ; P1_R1222_U441
g17199 nand P1_U4023 P1_R1222_U84 ; P1_R1222_U442
g17200 nand P1_R1222_U442 P1_R1222_U441 ; P1_R1222_U443
g17201 nand P1_R1222_U154 P1_R1222_U155 ; P1_R1222_U444
g17202 nand P1_R1222_U283 P1_R1222_U443 ; P1_R1222_U445
g17203 nand P1_U3075 P1_R1222_U55 ; P1_R1222_U446
g17204 nand P1_U4024 P1_R1222_U56 ; P1_R1222_U447
g17205 nand P1_U3075 P1_R1222_U55 ; P1_R1222_U448
g17206 nand P1_U4024 P1_R1222_U56 ; P1_R1222_U449
g17207 nand P1_R1222_U449 P1_R1222_U448 ; P1_R1222_U450
g17208 nand P1_U3076 P1_R1222_U82 ; P1_R1222_U451
g17209 nand P1_U4025 P1_R1222_U91 ; P1_R1222_U452
g17210 nand P1_R1222_U179 P1_R1222_U158 ; P1_R1222_U453
g17211 nand P1_R1222_U325 P1_R1222_U32 ; P1_R1222_U454
g17212 nand P1_U3081 P1_R1222_U79 ; P1_R1222_U455
g17213 nand P1_U3514 P1_R1222_U80 ; P1_R1222_U456
g17214 nand P1_R1222_U456 P1_R1222_U455 ; P1_R1222_U457
g17215 nand P1_R1222_U356 P1_R1222_U92 ; P1_R1222_U458
g17216 nand P1_R1222_U457 P1_R1222_U313 ; P1_R1222_U459
g17217 nand P1_U3082 P1_R1222_U76 ; P1_R1222_U460
g17218 nand P1_U3512 P1_R1222_U77 ; P1_R1222_U461
g17219 nand P1_R1222_U461 P1_R1222_U460 ; P1_R1222_U462
g17220 nand P1_R1222_U357 P1_R1222_U159 ; P1_R1222_U463
g17221 nand P1_R1222_U267 P1_R1222_U462 ; P1_R1222_U464
g17222 nand P1_U3069 P1_R1222_U61 ; P1_R1222_U465
g17223 nand P1_U3509 P1_R1222_U59 ; P1_R1222_U466
g17224 nand P1_U3073 P1_R1222_U57 ; P1_R1222_U467
g17225 nand P1_U3506 P1_R1222_U58 ; P1_R1222_U468
g17226 nand P1_R1222_U468 P1_R1222_U467 ; P1_R1222_U469
g17227 nand P1_R1222_U358 P1_R1222_U93 ; P1_R1222_U470
g17228 nand P1_R1222_U469 P1_R1222_U259 ; P1_R1222_U471
g17229 nand P1_U3074 P1_R1222_U74 ; P1_R1222_U472
g17230 nand P1_U3503 P1_R1222_U75 ; P1_R1222_U473
g17231 nand P1_U3074 P1_R1222_U74 ; P1_R1222_U474
g17232 nand P1_U3503 P1_R1222_U75 ; P1_R1222_U475
g17233 nand P1_R1222_U475 P1_R1222_U474 ; P1_R1222_U476
g17234 nand P1_R1222_U160 P1_R1222_U161 ; P1_R1222_U477
g17235 nand P1_R1222_U255 P1_R1222_U476 ; P1_R1222_U478
g17236 nand P1_U3079 P1_R1222_U72 ; P1_R1222_U479
g17237 nand P1_U3500 P1_R1222_U73 ; P1_R1222_U480
g17238 nand P1_U3079 P1_R1222_U72 ; P1_R1222_U481
g17239 nand P1_U3500 P1_R1222_U73 ; P1_R1222_U482
g17240 nand P1_R1222_U482 P1_R1222_U481 ; P1_R1222_U483
g17241 nand P1_R1222_U162 P1_R1222_U163 ; P1_R1222_U484
g17242 nand P1_R1222_U251 P1_R1222_U483 ; P1_R1222_U485
g17243 nand P1_U3080 P1_R1222_U70 ; P1_R1222_U486
g17244 nand P1_U3497 P1_R1222_U71 ; P1_R1222_U487
g17245 nand P1_U3072 P1_R1222_U65 ; P1_R1222_U488
g17246 nand P1_U3494 P1_R1222_U66 ; P1_R1222_U489
g17247 nand P1_R1222_U489 P1_R1222_U488 ; P1_R1222_U490
g17248 nand P1_R1222_U359 P1_R1222_U94 ; P1_R1222_U491
g17249 nand P1_R1222_U490 P1_R1222_U335 ; P1_R1222_U492
g17250 nand P1_U3063 P1_R1222_U67 ; P1_R1222_U493
g17251 nand P1_U3491 P1_R1222_U68 ; P1_R1222_U494
g17252 nand P1_R1222_U494 P1_R1222_U493 ; P1_R1222_U495
g17253 nand P1_R1222_U360 P1_R1222_U164 ; P1_R1222_U496
g17254 nand P1_R1222_U241 P1_R1222_U495 ; P1_R1222_U497
g17255 nand P1_U3062 P1_R1222_U63 ; P1_R1222_U498
g17256 nand P1_U3488 P1_R1222_U64 ; P1_R1222_U499
g17257 nand P1_U3077 P1_R1222_U30 ; P1_R1222_U500
g17258 nand P1_U3456 P1_R1222_U31 ; P1_R1222_U501
g17259 not P2_REG3_REG_3__SCAN_IN ; P2_ADD_1119_U4
g17260 and P2_ADD_1119_U78 P2_ADD_1119_U106 ; P2_ADD_1119_U5
g17261 not P2_REG3_REG_5__SCAN_IN ; P2_ADD_1119_U6
g17262 not P2_REG3_REG_4__SCAN_IN ; P2_ADD_1119_U7
g17263 nand P2_REG3_REG_4__SCAN_IN P2_REG3_REG_5__SCAN_IN P2_REG3_REG_3__SCAN_IN ; P2_ADD_1119_U8
g17264 not P2_REG3_REG_7__SCAN_IN ; P2_ADD_1119_U9
g17265 not P2_REG3_REG_6__SCAN_IN ; P2_ADD_1119_U10
g17266 nand P2_ADD_1119_U75 P2_ADD_1119_U85 ; P2_ADD_1119_U11
g17267 not P2_REG3_REG_8__SCAN_IN ; P2_ADD_1119_U12
g17268 not P2_REG3_REG_9__SCAN_IN ; P2_ADD_1119_U13
g17269 nand P2_ADD_1119_U76 P2_ADD_1119_U87 ; P2_ADD_1119_U14
g17270 not P2_REG3_REG_11__SCAN_IN ; P2_ADD_1119_U15
g17271 not P2_REG3_REG_10__SCAN_IN ; P2_ADD_1119_U16
g17272 nand P2_ADD_1119_U77 P2_ADD_1119_U89 ; P2_ADD_1119_U17
g17273 not P2_REG3_REG_12__SCAN_IN ; P2_ADD_1119_U18
g17274 nand P2_ADD_1119_U91 P2_REG3_REG_12__SCAN_IN ; P2_ADD_1119_U19
g17275 not P2_REG3_REG_13__SCAN_IN ; P2_ADD_1119_U20
g17276 nand P2_ADD_1119_U92 P2_REG3_REG_13__SCAN_IN ; P2_ADD_1119_U21
g17277 not P2_REG3_REG_14__SCAN_IN ; P2_ADD_1119_U22
g17278 nand P2_ADD_1119_U93 P2_REG3_REG_14__SCAN_IN ; P2_ADD_1119_U23
g17279 not P2_REG3_REG_15__SCAN_IN ; P2_ADD_1119_U24
g17280 nand P2_ADD_1119_U94 P2_REG3_REG_15__SCAN_IN ; P2_ADD_1119_U25
g17281 not P2_REG3_REG_16__SCAN_IN ; P2_ADD_1119_U26
g17282 nand P2_ADD_1119_U95 P2_REG3_REG_16__SCAN_IN ; P2_ADD_1119_U27
g17283 not P2_REG3_REG_17__SCAN_IN ; P2_ADD_1119_U28
g17284 nand P2_ADD_1119_U96 P2_REG3_REG_17__SCAN_IN ; P2_ADD_1119_U29
g17285 not P2_REG3_REG_18__SCAN_IN ; P2_ADD_1119_U30
g17286 nand P2_ADD_1119_U97 P2_REG3_REG_18__SCAN_IN ; P2_ADD_1119_U31
g17287 not P2_REG3_REG_19__SCAN_IN ; P2_ADD_1119_U32
g17288 nand P2_ADD_1119_U98 P2_REG3_REG_19__SCAN_IN ; P2_ADD_1119_U33
g17289 not P2_REG3_REG_20__SCAN_IN ; P2_ADD_1119_U34
g17290 nand P2_ADD_1119_U99 P2_REG3_REG_20__SCAN_IN ; P2_ADD_1119_U35
g17291 not P2_REG3_REG_21__SCAN_IN ; P2_ADD_1119_U36
g17292 nand P2_ADD_1119_U100 P2_REG3_REG_21__SCAN_IN ; P2_ADD_1119_U37
g17293 not P2_REG3_REG_22__SCAN_IN ; P2_ADD_1119_U38
g17294 nand P2_ADD_1119_U101 P2_REG3_REG_22__SCAN_IN ; P2_ADD_1119_U39
g17295 not P2_REG3_REG_23__SCAN_IN ; P2_ADD_1119_U40
g17296 nand P2_ADD_1119_U102 P2_REG3_REG_23__SCAN_IN ; P2_ADD_1119_U41
g17297 not P2_REG3_REG_24__SCAN_IN ; P2_ADD_1119_U42
g17298 nand P2_ADD_1119_U103 P2_REG3_REG_24__SCAN_IN ; P2_ADD_1119_U43
g17299 not P2_REG3_REG_25__SCAN_IN ; P2_ADD_1119_U44
g17300 nand P2_ADD_1119_U104 P2_REG3_REG_25__SCAN_IN ; P2_ADD_1119_U45
g17301 not P2_REG3_REG_26__SCAN_IN ; P2_ADD_1119_U46
g17302 nand P2_ADD_1119_U105 P2_REG3_REG_26__SCAN_IN ; P2_ADD_1119_U47
g17303 not P2_REG3_REG_28__SCAN_IN ; P2_ADD_1119_U48
g17304 not P2_REG3_REG_27__SCAN_IN ; P2_ADD_1119_U49
g17305 nand P2_ADD_1119_U109 P2_ADD_1119_U108 ; P2_ADD_1119_U50
g17306 nand P2_ADD_1119_U111 P2_ADD_1119_U110 ; P2_ADD_1119_U51
g17307 nand P2_ADD_1119_U113 P2_ADD_1119_U112 ; P2_ADD_1119_U52
g17308 nand P2_ADD_1119_U115 P2_ADD_1119_U114 ; P2_ADD_1119_U53
g17309 nand P2_ADD_1119_U117 P2_ADD_1119_U116 ; P2_ADD_1119_U54
g17310 nand P2_ADD_1119_U119 P2_ADD_1119_U118 ; P2_ADD_1119_U55
g17311 nand P2_ADD_1119_U121 P2_ADD_1119_U120 ; P2_ADD_1119_U56
g17312 nand P2_ADD_1119_U123 P2_ADD_1119_U122 ; P2_ADD_1119_U57
g17313 nand P2_ADD_1119_U125 P2_ADD_1119_U124 ; P2_ADD_1119_U58
g17314 nand P2_ADD_1119_U127 P2_ADD_1119_U126 ; P2_ADD_1119_U59
g17315 nand P2_ADD_1119_U129 P2_ADD_1119_U128 ; P2_ADD_1119_U60
g17316 nand P2_ADD_1119_U131 P2_ADD_1119_U130 ; P2_ADD_1119_U61
g17317 nand P2_ADD_1119_U133 P2_ADD_1119_U132 ; P2_ADD_1119_U62
g17318 nand P2_ADD_1119_U135 P2_ADD_1119_U134 ; P2_ADD_1119_U63
g17319 nand P2_ADD_1119_U137 P2_ADD_1119_U136 ; P2_ADD_1119_U64
g17320 nand P2_ADD_1119_U139 P2_ADD_1119_U138 ; P2_ADD_1119_U65
g17321 nand P2_ADD_1119_U141 P2_ADD_1119_U140 ; P2_ADD_1119_U66
g17322 nand P2_ADD_1119_U143 P2_ADD_1119_U142 ; P2_ADD_1119_U67
g17323 nand P2_ADD_1119_U145 P2_ADD_1119_U144 ; P2_ADD_1119_U68
g17324 nand P2_ADD_1119_U147 P2_ADD_1119_U146 ; P2_ADD_1119_U69
g17325 nand P2_ADD_1119_U149 P2_ADD_1119_U148 ; P2_ADD_1119_U70
g17326 nand P2_ADD_1119_U151 P2_ADD_1119_U150 ; P2_ADD_1119_U71
g17327 nand P2_ADD_1119_U153 P2_ADD_1119_U152 ; P2_ADD_1119_U72
g17328 nand P2_ADD_1119_U155 P2_ADD_1119_U154 ; P2_ADD_1119_U73
g17329 nand P2_ADD_1119_U157 P2_ADD_1119_U156 ; P2_ADD_1119_U74
g17330 and P2_REG3_REG_6__SCAN_IN P2_REG3_REG_7__SCAN_IN ; P2_ADD_1119_U75
g17331 and P2_REG3_REG_9__SCAN_IN P2_REG3_REG_8__SCAN_IN ; P2_ADD_1119_U76
g17332 and P2_REG3_REG_11__SCAN_IN P2_REG3_REG_10__SCAN_IN ; P2_ADD_1119_U77
g17333 and P2_REG3_REG_28__SCAN_IN P2_REG3_REG_27__SCAN_IN ; P2_ADD_1119_U78
g17334 nand P2_ADD_1119_U87 P2_REG3_REG_8__SCAN_IN ; P2_ADD_1119_U79
g17335 nand P2_ADD_1119_U85 P2_REG3_REG_6__SCAN_IN ; P2_ADD_1119_U80
g17336 nand P2_REG3_REG_4__SCAN_IN P2_REG3_REG_3__SCAN_IN ; P2_ADD_1119_U81
g17337 nand P2_ADD_1119_U106 P2_REG3_REG_27__SCAN_IN ; P2_ADD_1119_U82
g17338 nand P2_ADD_1119_U89 P2_REG3_REG_10__SCAN_IN ; P2_ADD_1119_U83
g17339 not P2_ADD_1119_U81 ; P2_ADD_1119_U84
g17340 not P2_ADD_1119_U8 ; P2_ADD_1119_U85
g17341 not P2_ADD_1119_U80 ; P2_ADD_1119_U86
g17342 not P2_ADD_1119_U11 ; P2_ADD_1119_U87
g17343 not P2_ADD_1119_U79 ; P2_ADD_1119_U88
g17344 not P2_ADD_1119_U14 ; P2_ADD_1119_U89
g17345 not P2_ADD_1119_U83 ; P2_ADD_1119_U90
g17346 not P2_ADD_1119_U17 ; P2_ADD_1119_U91
g17347 not P2_ADD_1119_U19 ; P2_ADD_1119_U92
g17348 not P2_ADD_1119_U21 ; P2_ADD_1119_U93
g17349 not P2_ADD_1119_U23 ; P2_ADD_1119_U94
g17350 not P2_ADD_1119_U25 ; P2_ADD_1119_U95
g17351 not P2_ADD_1119_U27 ; P2_ADD_1119_U96
g17352 not P2_ADD_1119_U29 ; P2_ADD_1119_U97
g17353 not P2_ADD_1119_U31 ; P2_ADD_1119_U98
g17354 not P2_ADD_1119_U33 ; P2_ADD_1119_U99
g17355 not P2_ADD_1119_U35 ; P2_ADD_1119_U100
g17356 not P2_ADD_1119_U37 ; P2_ADD_1119_U101
g17357 not P2_ADD_1119_U39 ; P2_ADD_1119_U102
g17358 not P2_ADD_1119_U41 ; P2_ADD_1119_U103
g17359 not P2_ADD_1119_U43 ; P2_ADD_1119_U104
g17360 not P2_ADD_1119_U45 ; P2_ADD_1119_U105
g17361 not P2_ADD_1119_U47 ; P2_ADD_1119_U106
g17362 not P2_ADD_1119_U82 ; P2_ADD_1119_U107
g17363 nand P2_ADD_1119_U79 P2_REG3_REG_9__SCAN_IN ; P2_ADD_1119_U108
g17364 nand P2_ADD_1119_U88 P2_ADD_1119_U13 ; P2_ADD_1119_U109
g17365 nand P2_ADD_1119_U11 P2_REG3_REG_8__SCAN_IN ; P2_ADD_1119_U110
g17366 nand P2_ADD_1119_U87 P2_ADD_1119_U12 ; P2_ADD_1119_U111
g17367 nand P2_ADD_1119_U80 P2_REG3_REG_7__SCAN_IN ; P2_ADD_1119_U112
g17368 nand P2_ADD_1119_U86 P2_ADD_1119_U9 ; P2_ADD_1119_U113
g17369 nand P2_ADD_1119_U8 P2_REG3_REG_6__SCAN_IN ; P2_ADD_1119_U114
g17370 nand P2_ADD_1119_U85 P2_ADD_1119_U10 ; P2_ADD_1119_U115
g17371 nand P2_ADD_1119_U81 P2_REG3_REG_5__SCAN_IN ; P2_ADD_1119_U116
g17372 nand P2_ADD_1119_U84 P2_ADD_1119_U6 ; P2_ADD_1119_U117
g17373 nand P2_ADD_1119_U4 P2_REG3_REG_4__SCAN_IN ; P2_ADD_1119_U118
g17374 nand P2_ADD_1119_U7 P2_REG3_REG_3__SCAN_IN ; P2_ADD_1119_U119
g17375 nand P2_ADD_1119_U82 P2_REG3_REG_28__SCAN_IN ; P2_ADD_1119_U120
g17376 nand P2_ADD_1119_U107 P2_ADD_1119_U48 ; P2_ADD_1119_U121
g17377 nand P2_ADD_1119_U47 P2_REG3_REG_27__SCAN_IN ; P2_ADD_1119_U122
g17378 nand P2_ADD_1119_U106 P2_ADD_1119_U49 ; P2_ADD_1119_U123
g17379 nand P2_ADD_1119_U45 P2_REG3_REG_26__SCAN_IN ; P2_ADD_1119_U124
g17380 nand P2_ADD_1119_U105 P2_ADD_1119_U46 ; P2_ADD_1119_U125
g17381 nand P2_ADD_1119_U43 P2_REG3_REG_25__SCAN_IN ; P2_ADD_1119_U126
g17382 nand P2_ADD_1119_U104 P2_ADD_1119_U44 ; P2_ADD_1119_U127
g17383 nand P2_ADD_1119_U41 P2_REG3_REG_24__SCAN_IN ; P2_ADD_1119_U128
g17384 nand P2_ADD_1119_U103 P2_ADD_1119_U42 ; P2_ADD_1119_U129
g17385 nand P2_ADD_1119_U39 P2_REG3_REG_23__SCAN_IN ; P2_ADD_1119_U130
g17386 nand P2_ADD_1119_U102 P2_ADD_1119_U40 ; P2_ADD_1119_U131
g17387 nand P2_ADD_1119_U37 P2_REG3_REG_22__SCAN_IN ; P2_ADD_1119_U132
g17388 nand P2_ADD_1119_U101 P2_ADD_1119_U38 ; P2_ADD_1119_U133
g17389 nand P2_ADD_1119_U35 P2_REG3_REG_21__SCAN_IN ; P2_ADD_1119_U134
g17390 nand P2_ADD_1119_U100 P2_ADD_1119_U36 ; P2_ADD_1119_U135
g17391 nand P2_ADD_1119_U33 P2_REG3_REG_20__SCAN_IN ; P2_ADD_1119_U136
g17392 nand P2_ADD_1119_U99 P2_ADD_1119_U34 ; P2_ADD_1119_U137
g17393 nand P2_ADD_1119_U31 P2_REG3_REG_19__SCAN_IN ; P2_ADD_1119_U138
g17394 nand P2_ADD_1119_U98 P2_ADD_1119_U32 ; P2_ADD_1119_U139
g17395 nand P2_ADD_1119_U29 P2_REG3_REG_18__SCAN_IN ; P2_ADD_1119_U140
g17396 nand P2_ADD_1119_U97 P2_ADD_1119_U30 ; P2_ADD_1119_U141
g17397 nand P2_ADD_1119_U27 P2_REG3_REG_17__SCAN_IN ; P2_ADD_1119_U142
g17398 nand P2_ADD_1119_U96 P2_ADD_1119_U28 ; P2_ADD_1119_U143
g17399 nand P2_ADD_1119_U25 P2_REG3_REG_16__SCAN_IN ; P2_ADD_1119_U144
g17400 nand P2_ADD_1119_U95 P2_ADD_1119_U26 ; P2_ADD_1119_U145
g17401 nand P2_ADD_1119_U23 P2_REG3_REG_15__SCAN_IN ; P2_ADD_1119_U146
g17402 nand P2_ADD_1119_U94 P2_ADD_1119_U24 ; P2_ADD_1119_U147
g17403 nand P2_ADD_1119_U21 P2_REG3_REG_14__SCAN_IN ; P2_ADD_1119_U148
g17404 nand P2_ADD_1119_U93 P2_ADD_1119_U22 ; P2_ADD_1119_U149
g17405 nand P2_ADD_1119_U19 P2_REG3_REG_13__SCAN_IN ; P2_ADD_1119_U150
g17406 nand P2_ADD_1119_U92 P2_ADD_1119_U20 ; P2_ADD_1119_U151
g17407 nand P2_ADD_1119_U17 P2_REG3_REG_12__SCAN_IN ; P2_ADD_1119_U152
g17408 nand P2_ADD_1119_U91 P2_ADD_1119_U18 ; P2_ADD_1119_U153
g17409 nand P2_ADD_1119_U83 P2_REG3_REG_11__SCAN_IN ; P2_ADD_1119_U154
g17410 nand P2_ADD_1119_U90 P2_ADD_1119_U15 ; P2_ADD_1119_U155
g17411 nand P2_ADD_1119_U14 P2_REG3_REG_10__SCAN_IN ; P2_ADD_1119_U156
g17412 nand P2_ADD_1119_U89 P2_ADD_1119_U16 ; P2_ADD_1119_U157
g17413 and P2_SUB_1108_U172 P2_SUB_1108_U40 ; P2_SUB_1108_U6
g17414 and P2_SUB_1108_U170 P2_SUB_1108_U140 ; P2_SUB_1108_U7
g17415 and P2_SUB_1108_U169 P2_SUB_1108_U37 ; P2_SUB_1108_U8
g17416 and P2_SUB_1108_U168 P2_SUB_1108_U38 ; P2_SUB_1108_U9
g17417 and P2_SUB_1108_U166 P2_SUB_1108_U143 ; P2_SUB_1108_U10
g17418 and P2_SUB_1108_U165 P2_SUB_1108_U30 ; P2_SUB_1108_U11
g17419 and P2_SUB_1108_U164 P2_SUB_1108_U36 ; P2_SUB_1108_U12
g17420 and P2_SUB_1108_U162 P2_SUB_1108_U32 ; P2_SUB_1108_U13
g17421 and P2_SUB_1108_U160 P2_SUB_1108_U33 ; P2_SUB_1108_U14
g17422 and P2_SUB_1108_U159 P2_SUB_1108_U109 ; P2_SUB_1108_U15
g17423 and P2_SUB_1108_U157 P2_SUB_1108_U29 ; P2_SUB_1108_U16
g17424 and P2_SUB_1108_U155 P2_SUB_1108_U23 ; P2_SUB_1108_U17
g17425 and P2_SUB_1108_U138 P2_SUB_1108_U128 ; P2_SUB_1108_U18
g17426 and P2_SUB_1108_U137 P2_SUB_1108_U25 ; P2_SUB_1108_U19
g17427 and P2_SUB_1108_U136 P2_SUB_1108_U26 ; P2_SUB_1108_U20
g17428 and P2_SUB_1108_U134 P2_SUB_1108_U131 ; P2_SUB_1108_U21
g17429 and P2_SUB_1108_U133 P2_SUB_1108_U24 ; P2_SUB_1108_U22
g17430 or P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_2__SCAN_IN ; P2_SUB_1108_U23
g17431 nand P2_SUB_1108_U45 P2_SUB_1108_U174 P2_SUB_1108_U44 ; P2_SUB_1108_U24
g17432 nand P2_SUB_1108_U46 P2_SUB_1108_U174 ; P2_SUB_1108_U25
g17433 nand P2_SUB_1108_U47 P2_SUB_1108_U129 ; P2_SUB_1108_U26
g17434 not P2_IR_REG_7__SCAN_IN ; P2_SUB_1108_U27
g17435 not P2_IR_REG_3__SCAN_IN ; P2_SUB_1108_U28
g17436 nand P2_SUB_1108_U57 P2_SUB_1108_U52 ; P2_SUB_1108_U29
g17437 nand P2_SUB_1108_U91 P2_SUB_1108_U90 P2_SUB_1108_U89 P2_SUB_1108_U88 ; P2_SUB_1108_U30
g17438 nand P2_SUB_1108_U92 P2_SUB_1108_U144 ; P2_SUB_1108_U31
g17439 nand P2_SUB_1108_U93 P2_SUB_1108_U147 ; P2_SUB_1108_U32
g17440 nand P2_SUB_1108_U149 P2_SUB_1108_U34 ; P2_SUB_1108_U33
g17441 not P2_IR_REG_24__SCAN_IN ; P2_SUB_1108_U34
g17442 nand P2_SUB_1108_U147 P2_SUB_1108_U115 ; P2_SUB_1108_U35
g17443 nand P2_SUB_1108_U94 P2_SUB_1108_U144 ; P2_SUB_1108_U36
g17444 nand P2_SUB_1108_U95 P2_SUB_1108_U132 ; P2_SUB_1108_U37
g17445 nand P2_SUB_1108_U96 P2_SUB_1108_U141 ; P2_SUB_1108_U38
g17446 not P2_IR_REG_15__SCAN_IN ; P2_SUB_1108_U39
g17447 nand P2_SUB_1108_U97 P2_SUB_1108_U132 ; P2_SUB_1108_U40
g17448 not P2_IR_REG_11__SCAN_IN ; P2_SUB_1108_U41
g17449 nand P2_SUB_1108_U196 P2_SUB_1108_U195 ; P2_SUB_1108_U42
g17450 nand P2_SUB_1108_U180 P2_SUB_1108_U179 ; P2_SUB_1108_U43
g17451 nor P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U44
g17452 nor P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN ; P2_SUB_1108_U45
g17453 nor P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN ; P2_SUB_1108_U46
g17454 nor P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U47
g17455 nor P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN P2_IR_REG_13__SCAN_IN ; P2_SUB_1108_U48
g17456 nor P2_IR_REG_14__SCAN_IN P2_IR_REG_15__SCAN_IN P2_IR_REG_16__SCAN_IN P2_IR_REG_17__SCAN_IN ; P2_SUB_1108_U49
g17457 nor P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN ; P2_SUB_1108_U50
g17458 nor P2_IR_REG_20__SCAN_IN P2_IR_REG_21__SCAN_IN P2_IR_REG_22__SCAN_IN ; P2_SUB_1108_U51
g17459 and P2_SUB_1108_U51 P2_SUB_1108_U50 P2_SUB_1108_U49 P2_SUB_1108_U48 ; P2_SUB_1108_U52
g17460 nor P2_IR_REG_23__SCAN_IN P2_IR_REG_24__SCAN_IN P2_IR_REG_25__SCAN_IN P2_IR_REG_26__SCAN_IN ; P2_SUB_1108_U53
g17461 nor P2_IR_REG_2__SCAN_IN P2_IR_REG_27__SCAN_IN P2_IR_REG_28__SCAN_IN P2_IR_REG_29__SCAN_IN ; P2_SUB_1108_U54
g17462 nor P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U55
g17463 nor P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U56
g17464 and P2_SUB_1108_U56 P2_SUB_1108_U55 P2_SUB_1108_U54 P2_SUB_1108_U53 ; P2_SUB_1108_U57
g17465 nor P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN P2_IR_REG_13__SCAN_IN ; P2_SUB_1108_U58
g17466 nor P2_IR_REG_14__SCAN_IN P2_IR_REG_15__SCAN_IN P2_IR_REG_16__SCAN_IN P2_IR_REG_17__SCAN_IN ; P2_SUB_1108_U59
g17467 nor P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN ; P2_SUB_1108_U60
g17468 nor P2_IR_REG_20__SCAN_IN P2_IR_REG_21__SCAN_IN P2_IR_REG_22__SCAN_IN ; P2_SUB_1108_U61
g17469 and P2_SUB_1108_U61 P2_SUB_1108_U60 P2_SUB_1108_U59 P2_SUB_1108_U58 ; P2_SUB_1108_U62
g17470 nor P2_IR_REG_23__SCAN_IN P2_IR_REG_24__SCAN_IN P2_IR_REG_25__SCAN_IN P2_IR_REG_26__SCAN_IN ; P2_SUB_1108_U63
g17471 nor P2_IR_REG_2__SCAN_IN P2_IR_REG_27__SCAN_IN P2_IR_REG_28__SCAN_IN ; P2_SUB_1108_U64
g17472 nor P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U65
g17473 nor P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U66
g17474 and P2_SUB_1108_U66 P2_SUB_1108_U65 P2_SUB_1108_U64 P2_SUB_1108_U63 ; P2_SUB_1108_U67
g17475 nor P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN P2_IR_REG_13__SCAN_IN ; P2_SUB_1108_U68
g17476 nor P2_IR_REG_14__SCAN_IN P2_IR_REG_15__SCAN_IN P2_IR_REG_16__SCAN_IN ; P2_SUB_1108_U69
g17477 nor P2_IR_REG_1__SCAN_IN P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN ; P2_SUB_1108_U70
g17478 nor P2_IR_REG_0__SCAN_IN P2_IR_REG_20__SCAN_IN P2_IR_REG_21__SCAN_IN ; P2_SUB_1108_U71
g17479 and P2_SUB_1108_U71 P2_SUB_1108_U70 P2_SUB_1108_U69 P2_SUB_1108_U68 ; P2_SUB_1108_U72
g17480 nor P2_IR_REG_22__SCAN_IN P2_IR_REG_23__SCAN_IN P2_IR_REG_24__SCAN_IN P2_IR_REG_25__SCAN_IN ; P2_SUB_1108_U73
g17481 nor P2_IR_REG_2__SCAN_IN P2_IR_REG_26__SCAN_IN P2_IR_REG_27__SCAN_IN ; P2_SUB_1108_U74
g17482 nor P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U75
g17483 nor P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U76
g17484 and P2_SUB_1108_U76 P2_SUB_1108_U75 P2_SUB_1108_U74 P2_SUB_1108_U73 ; P2_SUB_1108_U77
g17485 nor P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN P2_IR_REG_13__SCAN_IN ; P2_SUB_1108_U78
g17486 nor P2_IR_REG_14__SCAN_IN P2_IR_REG_15__SCAN_IN P2_IR_REG_16__SCAN_IN ; P2_SUB_1108_U79
g17487 nor P2_IR_REG_1__SCAN_IN P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN ; P2_SUB_1108_U80
g17488 nor P2_IR_REG_0__SCAN_IN P2_IR_REG_20__SCAN_IN P2_IR_REG_21__SCAN_IN ; P2_SUB_1108_U81
g17489 and P2_SUB_1108_U81 P2_SUB_1108_U80 P2_SUB_1108_U79 P2_SUB_1108_U78 ; P2_SUB_1108_U82
g17490 nor P2_IR_REG_22__SCAN_IN P2_IR_REG_23__SCAN_IN P2_IR_REG_24__SCAN_IN P2_IR_REG_25__SCAN_IN ; P2_SUB_1108_U83
g17491 nor P2_IR_REG_2__SCAN_IN P2_IR_REG_3__SCAN_IN P2_IR_REG_26__SCAN_IN ; P2_SUB_1108_U84
g17492 nor P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U85
g17493 nor P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U86
g17494 and P2_SUB_1108_U86 P2_SUB_1108_U85 P2_SUB_1108_U84 P2_SUB_1108_U83 ; P2_SUB_1108_U87
g17495 nor P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN P2_IR_REG_13__SCAN_IN P2_IR_REG_14__SCAN_IN ; P2_SUB_1108_U88
g17496 nor P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN P2_IR_REG_15__SCAN_IN P2_IR_REG_16__SCAN_IN ; P2_SUB_1108_U89
g17497 nor P2_IR_REG_2__SCAN_IN P2_IR_REG_3__SCAN_IN P2_IR_REG_4__SCAN_IN P2_IR_REG_5__SCAN_IN ; P2_SUB_1108_U90
g17498 nor P2_IR_REG_6__SCAN_IN P2_IR_REG_7__SCAN_IN P2_IR_REG_8__SCAN_IN P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U91
g17499 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN P2_IR_REG_19__SCAN_IN P2_IR_REG_20__SCAN_IN ; P2_SUB_1108_U92
g17500 nor P2_IR_REG_21__SCAN_IN P2_IR_REG_22__SCAN_IN P2_IR_REG_23__SCAN_IN ; P2_SUB_1108_U93
g17501 nor P2_IR_REG_17__SCAN_IN P2_IR_REG_18__SCAN_IN ; P2_SUB_1108_U94
g17502 nor P2_IR_REG_9__SCAN_IN P2_IR_REG_10__SCAN_IN P2_IR_REG_11__SCAN_IN P2_IR_REG_12__SCAN_IN ; P2_SUB_1108_U95
g17503 nor P2_IR_REG_13__SCAN_IN P2_IR_REG_14__SCAN_IN ; P2_SUB_1108_U96
g17504 nor P2_IR_REG_9__SCAN_IN P2_IR_REG_10__SCAN_IN ; P2_SUB_1108_U97
g17505 not P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U98
g17506 and P2_SUB_1108_U176 P2_SUB_1108_U175 ; P2_SUB_1108_U99
g17507 not P2_IR_REG_5__SCAN_IN ; P2_SUB_1108_U100
g17508 and P2_SUB_1108_U178 P2_SUB_1108_U177 ; P2_SUB_1108_U101
g17509 not P2_IR_REG_31__SCAN_IN ; P2_SUB_1108_U102
g17510 not P2_IR_REG_30__SCAN_IN ; P2_SUB_1108_U103
g17511 and P2_SUB_1108_U182 P2_SUB_1108_U181 ; P2_SUB_1108_U104
g17512 not P2_IR_REG_28__SCAN_IN ; P2_SUB_1108_U105
g17513 nand P2_SUB_1108_U77 P2_SUB_1108_U72 ; P2_SUB_1108_U106
g17514 and P2_SUB_1108_U184 P2_SUB_1108_U183 ; P2_SUB_1108_U107
g17515 not P2_IR_REG_27__SCAN_IN ; P2_SUB_1108_U108
g17516 nand P2_SUB_1108_U87 P2_SUB_1108_U82 ; P2_SUB_1108_U109
g17517 and P2_SUB_1108_U186 P2_SUB_1108_U185 ; P2_SUB_1108_U110
g17518 not P2_IR_REG_25__SCAN_IN ; P2_SUB_1108_U111
g17519 and P2_SUB_1108_U188 P2_SUB_1108_U187 ; P2_SUB_1108_U112
g17520 not P2_IR_REG_22__SCAN_IN ; P2_SUB_1108_U113
g17521 and P2_SUB_1108_U190 P2_SUB_1108_U189 ; P2_SUB_1108_U114
g17522 not P2_IR_REG_21__SCAN_IN ; P2_SUB_1108_U115
g17523 and P2_SUB_1108_U192 P2_SUB_1108_U191 ; P2_SUB_1108_U116
g17524 not P2_IR_REG_20__SCAN_IN ; P2_SUB_1108_U117
g17525 nand P2_SUB_1108_U145 P2_SUB_1108_U122 ; P2_SUB_1108_U118
g17526 and P2_SUB_1108_U194 P2_SUB_1108_U193 ; P2_SUB_1108_U119
g17527 not P2_IR_REG_1__SCAN_IN ; P2_SUB_1108_U120
g17528 not P2_IR_REG_0__SCAN_IN ; P2_SUB_1108_U121
g17529 not P2_IR_REG_19__SCAN_IN ; P2_SUB_1108_U122
g17530 and P2_SUB_1108_U198 P2_SUB_1108_U197 ; P2_SUB_1108_U123
g17531 not P2_IR_REG_17__SCAN_IN ; P2_SUB_1108_U124
g17532 and P2_SUB_1108_U200 P2_SUB_1108_U199 ; P2_SUB_1108_U125
g17533 not P2_IR_REG_13__SCAN_IN ; P2_SUB_1108_U126
g17534 and P2_SUB_1108_U202 P2_SUB_1108_U201 ; P2_SUB_1108_U127
g17535 nand P2_SUB_1108_U174 P2_SUB_1108_U28 ; P2_SUB_1108_U128
g17536 not P2_SUB_1108_U25 ; P2_SUB_1108_U129
g17537 not P2_SUB_1108_U26 ; P2_SUB_1108_U130
g17538 nand P2_SUB_1108_U130 P2_SUB_1108_U27 ; P2_SUB_1108_U131
g17539 not P2_SUB_1108_U24 ; P2_SUB_1108_U132
g17540 nand P2_SUB_1108_U131 P2_IR_REG_8__SCAN_IN ; P2_SUB_1108_U133
g17541 nand P2_SUB_1108_U26 P2_IR_REG_7__SCAN_IN ; P2_SUB_1108_U134
g17542 nand P2_SUB_1108_U129 P2_SUB_1108_U100 ; P2_SUB_1108_U135
g17543 nand P2_SUB_1108_U135 P2_IR_REG_6__SCAN_IN ; P2_SUB_1108_U136
g17544 nand P2_SUB_1108_U128 P2_IR_REG_4__SCAN_IN ; P2_SUB_1108_U137
g17545 nand P2_SUB_1108_U23 P2_IR_REG_3__SCAN_IN ; P2_SUB_1108_U138
g17546 not P2_SUB_1108_U40 ; P2_SUB_1108_U139
g17547 nand P2_SUB_1108_U139 P2_SUB_1108_U41 ; P2_SUB_1108_U140
g17548 not P2_SUB_1108_U37 ; P2_SUB_1108_U141
g17549 not P2_SUB_1108_U38 ; P2_SUB_1108_U142
g17550 nand P2_SUB_1108_U142 P2_SUB_1108_U39 ; P2_SUB_1108_U143
g17551 not P2_SUB_1108_U30 ; P2_SUB_1108_U144
g17552 not P2_SUB_1108_U36 ; P2_SUB_1108_U145
g17553 not P2_SUB_1108_U118 ; P2_SUB_1108_U146
g17554 not P2_SUB_1108_U31 ; P2_SUB_1108_U147
g17555 not P2_SUB_1108_U35 ; P2_SUB_1108_U148
g17556 not P2_SUB_1108_U32 ; P2_SUB_1108_U149
g17557 not P2_SUB_1108_U33 ; P2_SUB_1108_U150
g17558 not P2_SUB_1108_U109 ; P2_SUB_1108_U151
g17559 not P2_SUB_1108_U106 ; P2_SUB_1108_U152
g17560 not P2_SUB_1108_U29 ; P2_SUB_1108_U153
g17561 or P2_IR_REG_0__SCAN_IN P2_IR_REG_1__SCAN_IN ; P2_SUB_1108_U154
g17562 nand P2_SUB_1108_U154 P2_IR_REG_2__SCAN_IN ; P2_SUB_1108_U155
g17563 nand P2_SUB_1108_U67 P2_SUB_1108_U62 ; P2_SUB_1108_U156
g17564 nand P2_SUB_1108_U156 P2_IR_REG_29__SCAN_IN ; P2_SUB_1108_U157
g17565 nand P2_SUB_1108_U150 P2_SUB_1108_U111 ; P2_SUB_1108_U158
g17566 nand P2_SUB_1108_U158 P2_IR_REG_26__SCAN_IN ; P2_SUB_1108_U159
g17567 nand P2_SUB_1108_U32 P2_IR_REG_24__SCAN_IN ; P2_SUB_1108_U160
g17568 nand P2_SUB_1108_U148 P2_SUB_1108_U113 ; P2_SUB_1108_U161
g17569 nand P2_SUB_1108_U161 P2_IR_REG_23__SCAN_IN ; P2_SUB_1108_U162
g17570 nand P2_SUB_1108_U144 P2_SUB_1108_U124 ; P2_SUB_1108_U163
g17571 nand P2_SUB_1108_U163 P2_IR_REG_18__SCAN_IN ; P2_SUB_1108_U164
g17572 nand P2_SUB_1108_U143 P2_IR_REG_16__SCAN_IN ; P2_SUB_1108_U165
g17573 nand P2_SUB_1108_U38 P2_IR_REG_15__SCAN_IN ; P2_SUB_1108_U166
g17574 nand P2_SUB_1108_U141 P2_SUB_1108_U126 ; P2_SUB_1108_U167
g17575 nand P2_SUB_1108_U167 P2_IR_REG_14__SCAN_IN ; P2_SUB_1108_U168
g17576 nand P2_SUB_1108_U140 P2_IR_REG_12__SCAN_IN ; P2_SUB_1108_U169
g17577 nand P2_SUB_1108_U40 P2_IR_REG_11__SCAN_IN ; P2_SUB_1108_U170
g17578 nand P2_SUB_1108_U132 P2_SUB_1108_U98 ; P2_SUB_1108_U171
g17579 nand P2_SUB_1108_U171 P2_IR_REG_10__SCAN_IN ; P2_SUB_1108_U172
g17580 nand P2_SUB_1108_U153 P2_SUB_1108_U103 ; P2_SUB_1108_U173
g17581 not P2_SUB_1108_U23 ; P2_SUB_1108_U174
g17582 nand P2_SUB_1108_U24 P2_IR_REG_9__SCAN_IN ; P2_SUB_1108_U175
g17583 nand P2_SUB_1108_U132 P2_SUB_1108_U98 ; P2_SUB_1108_U176
g17584 nand P2_SUB_1108_U25 P2_IR_REG_5__SCAN_IN ; P2_SUB_1108_U177
g17585 nand P2_SUB_1108_U129 P2_SUB_1108_U100 ; P2_SUB_1108_U178
g17586 nand P2_SUB_1108_U173 P2_SUB_1108_U102 ; P2_SUB_1108_U179
g17587 nand P2_SUB_1108_U153 P2_SUB_1108_U103 P2_IR_REG_31__SCAN_IN ; P2_SUB_1108_U180
g17588 nand P2_SUB_1108_U29 P2_IR_REG_30__SCAN_IN ; P2_SUB_1108_U181
g17589 nand P2_SUB_1108_U153 P2_SUB_1108_U103 ; P2_SUB_1108_U182
g17590 nand P2_SUB_1108_U106 P2_IR_REG_28__SCAN_IN ; P2_SUB_1108_U183
g17591 nand P2_SUB_1108_U152 P2_SUB_1108_U105 ; P2_SUB_1108_U184
g17592 nand P2_SUB_1108_U109 P2_IR_REG_27__SCAN_IN ; P2_SUB_1108_U185
g17593 nand P2_SUB_1108_U151 P2_SUB_1108_U108 ; P2_SUB_1108_U186
g17594 nand P2_SUB_1108_U33 P2_IR_REG_25__SCAN_IN ; P2_SUB_1108_U187
g17595 nand P2_SUB_1108_U150 P2_SUB_1108_U111 ; P2_SUB_1108_U188
g17596 nand P2_SUB_1108_U35 P2_IR_REG_22__SCAN_IN ; P2_SUB_1108_U189
g17597 nand P2_SUB_1108_U148 P2_SUB_1108_U113 ; P2_SUB_1108_U190
g17598 nand P2_SUB_1108_U31 P2_IR_REG_21__SCAN_IN ; P2_SUB_1108_U191
g17599 nand P2_SUB_1108_U147 P2_SUB_1108_U115 ; P2_SUB_1108_U192
g17600 nand P2_SUB_1108_U118 P2_IR_REG_20__SCAN_IN ; P2_SUB_1108_U193
g17601 nand P2_SUB_1108_U146 P2_SUB_1108_U117 ; P2_SUB_1108_U194
g17602 nand P2_SUB_1108_U121 P2_IR_REG_1__SCAN_IN ; P2_SUB_1108_U195
g17603 nand P2_SUB_1108_U120 P2_IR_REG_0__SCAN_IN ; P2_SUB_1108_U196
g17604 nand P2_SUB_1108_U36 P2_IR_REG_19__SCAN_IN ; P2_SUB_1108_U197
g17605 nand P2_SUB_1108_U145 P2_SUB_1108_U122 ; P2_SUB_1108_U198
g17606 nand P2_SUB_1108_U30 P2_IR_REG_17__SCAN_IN ; P2_SUB_1108_U199
g17607 nand P2_SUB_1108_U144 P2_SUB_1108_U124 ; P2_SUB_1108_U200
g17608 nand P2_SUB_1108_U37 P2_IR_REG_13__SCAN_IN ; P2_SUB_1108_U201
g17609 nand P2_SUB_1108_U141 P2_SUB_1108_U126 ; P2_SUB_1108_U202
g17610 and P2_U3061 P2_R1299_U7 ; P2_R1299_U6
g17611 not P2_U3058 ; P2_R1299_U7
g17612 and P2_R1312_U172 P2_R1312_U170 P2_R1312_U171 ; P2_R1312_U6
g17613 and P2_R1312_U85 P2_R1312_U84 ; P2_R1312_U7
g17614 and P2_R1312_U7 P2_R1312_U173 ; P2_R1312_U8
g17615 and P2_R1312_U183 P2_R1312_U182 ; P2_R1312_U9
g17616 and P2_R1312_U213 P2_R1312_U212 ; P2_R1312_U10
g17617 and P2_R1312_U14 P2_R1312_U82 P2_R1312_U169 ; P2_R1312_U11
g17618 and P2_R1312_U157 P2_R1312_U156 P2_R1312_U155 P2_R1312_U154 ; P2_R1312_U12
g17619 and P2_R1312_U176 P2_R1312_U175 P2_R1312_U174 P2_R1312_U173 ; P2_R1312_U13
g17620 and P2_R1312_U162 P2_R1312_U161 P2_R1312_U164 ; P2_R1312_U14
g17621 and P2_R1312_U6 P2_R1312_U11 P2_R1312_U83 P2_R1312_U165 P2_R1312_U17 ; P2_R1312_U15
g17622 and P2_R1312_U165 P2_R1312_U163 ; P2_R1312_U16
g17623 and P2_R1312_U225 P2_R1312_U224 ; P2_R1312_U17
g17624 nand P2_R1312_U152 P2_R1312_U151 P2_R1312_U150 P2_R1312_U147 P2_R1312_U144 ; P2_R1312_U18
g17625 not P2_U3090 ; P2_R1312_U19
g17626 not P2_U3093 ; P2_R1312_U20
g17627 not P2_U3091 ; P2_R1312_U21
g17628 not P2_U3092 ; P2_R1312_U22
g17629 not P2_U3126 ; P2_R1312_U23
g17630 not P2_U3123 ; P2_R1312_U24
g17631 not P2_U3089 ; P2_R1312_U25
g17632 not P2_U3121 ; P2_R1312_U26
g17633 not P2_U3105 ; P2_R1312_U27
g17634 not P2_U3106 ; P2_R1312_U28
g17635 not P2_U3108 ; P2_R1312_U29
g17636 not P2_U3107 ; P2_R1312_U30
g17637 not P2_U3109 ; P2_R1312_U31
g17638 not P2_U3110 ; P2_R1312_U32
g17639 not P2_U3111 ; P2_R1312_U33
g17640 not P2_U3112 ; P2_R1312_U34
g17641 not P2_U3115 ; P2_R1312_U35
g17642 not P2_U3116 ; P2_R1312_U36
g17643 not P2_U3114 ; P2_R1312_U37
g17644 not P2_U3113 ; P2_R1312_U38
g17645 not P2_U3104 ; P2_R1312_U39
g17646 not P2_U3094 ; P2_R1312_U40
g17647 not P2_U3102 ; P2_R1312_U41
g17648 not P2_U3101 ; P2_R1312_U42
g17649 not P2_U3103 ; P2_R1312_U43
g17650 not P2_U3100 ; P2_R1312_U44
g17651 not P2_U3099 ; P2_R1312_U45
g17652 not P2_U3095 ; P2_R1312_U46
g17653 not P2_U3097 ; P2_R1312_U47
g17654 not P2_U3098 ; P2_R1312_U48
g17655 not P2_U3096 ; P2_R1312_U49
g17656 not P2_U3149 ; P2_R1312_U50
g17657 not P2_U3117 ; P2_R1312_U51
g17658 not P2_U3118 ; P2_R1312_U52
g17659 not P2_U3119 ; P2_R1312_U53
g17660 not P2_U3151 ; P2_R1312_U54
g17661 not P2_U3127 ; P2_R1312_U55
g17662 not P2_U3125 ; P2_R1312_U56
g17663 not P2_U3124 ; P2_R1312_U57
g17664 not P2_U3140 ; P2_R1312_U58
g17665 not P2_U3141 ; P2_R1312_U59
g17666 not P2_U3143 ; P2_R1312_U60
g17667 not P2_U3128 ; P2_R1312_U61
g17668 not P2_U3129 ; P2_R1312_U62
g17669 not P2_U3131 ; P2_R1312_U63
g17670 not P2_U3134 ; P2_R1312_U64
g17671 not P2_U3135 ; P2_R1312_U65
g17672 not P2_U3137 ; P2_R1312_U66
g17673 not P2_U3146 ; P2_R1312_U67
g17674 not P2_U3147 ; P2_R1312_U68
g17675 not P2_U3133 ; P2_R1312_U69
g17676 not P2_U3139 ; P2_R1312_U70
g17677 not P2_U3145 ; P2_R1312_U71
g17678 not P2_U3130 ; P2_R1312_U72
g17679 not P2_U3132 ; P2_R1312_U73
g17680 not P2_U3136 ; P2_R1312_U74
g17681 not P2_U3138 ; P2_R1312_U75
g17682 not P2_U3142 ; P2_R1312_U76
g17683 not P2_U3144 ; P2_R1312_U77
g17684 not P2_U3148 ; P2_R1312_U78
g17685 not P2_U3150 ; P2_R1312_U79
g17686 not P2_U3122 ; P2_R1312_U80
g17687 and P2_R1312_U17 P2_R1312_U166 ; P2_R1312_U81
g17688 and P2_R1312_U160 P2_R1312_U159 ; P2_R1312_U82
g17689 and P2_R1312_U163 P2_R1312_U158 ; P2_R1312_U83
g17690 and P2_R1312_U177 P2_R1312_U176 P2_R1312_U175 P2_R1312_U174 ; P2_R1312_U84
g17691 and P2_R1312_U179 P2_R1312_U178 P2_R1312_U180 ; P2_R1312_U85
g17692 and P2_R1312_U168 P2_R1312_U51 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U86
g17693 and P2_U3149 P2_R1312_U12 ; P2_R1312_U87
g17694 and P2_R1312_U186 P2_R1312_U173 ; P2_R1312_U88
g17695 and P2_R1312_U88 P2_R1312_U185 P2_R1312_U168 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U89
g17696 and P2_R1312_U7 P2_R1312_U187 P2_R1312_U91 ; P2_R1312_U90
g17697 and P2_R1312_U9 P2_R1312_U12 ; P2_R1312_U91
g17698 and P2_R1312_U167 P2_R1312_U53 P2_R1312_U166 ; P2_R1312_U92
g17699 and P2_U3151 P2_R1312_U9 P2_R1312_U12 ; P2_R1312_U93
g17700 and P2_U3127 P2_R1312_U46 ; P2_R1312_U94
g17701 and P2_R1312_U194 P2_R1312_U195 ; P2_R1312_U95
g17702 and P2_R1312_U167 P2_R1312_U168 P2_R1312_U166 ; P2_R1312_U96
g17703 and P2_R1312_U167 P2_R1312_U29 P2_R1312_U173 P2_R1312_U168 ; P2_R1312_U97
g17704 and P2_R1312_U176 P2_R1312_U174 P2_U3140 ; P2_R1312_U98
g17705 and P2_R1312_U168 P2_R1312_U31 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U99
g17706 and P2_R1312_U13 P2_U3141 ; P2_R1312_U100
g17707 and P2_R1312_U167 P2_R1312_U33 P2_R1312_U177 P2_R1312_U168 ; P2_R1312_U101
g17708 and P2_R1312_U103 P2_R1312_U13 ; P2_R1312_U102
g17709 and P2_U3143 P2_R1312_U178 ; P2_R1312_U103
g17710 and P2_R1312_U168 P2_R1312_U49 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U104
g17711 and P2_R1312_U164 P2_R1312_U47 P2_R1312_U168 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U105
g17712 and P2_R1312_U167 P2_R1312_U45 P2_R1312_U169 P2_R1312_U168 ; P2_R1312_U106
g17713 and P2_U3131 P2_R1312_U16 ; P2_R1312_U107
g17714 and P2_R1312_U167 P2_R1312_U41 P2_R1312_U171 P2_R1312_U168 ; P2_R1312_U108
g17715 and P2_U3134 P2_R1312_U16 ; P2_R1312_U109
g17716 and P2_R1312_U167 P2_R1312_U43 P2_R1312_U170 P2_R1312_U168 ; P2_R1312_U110
g17717 and P2_R1312_U11 P2_R1312_U171 P2_R1312_U17 P2_R1312_U112 P2_R1312_U166 ; P2_R1312_U111
g17718 and P2_U3135 P2_R1312_U16 ; P2_R1312_U112
g17719 and P2_R1312_U167 P2_R1312_U27 P2_R1312_U166 ; P2_R1312_U113
g17720 and P2_U3137 P2_R1312_U168 ; P2_R1312_U114
g17721 and P2_R1312_U157 P2_R1312_U37 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U115
g17722 and P2_R1312_U156 P2_R1312_U35 P2_R1312_U157 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U116
g17723 and P2_R1312_U168 P2_R1312_U42 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U117
g17724 and P2_U3133 P2_R1312_U16 ; P2_R1312_U118
g17725 and P2_R1312_U168 P2_R1312_U30 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U119
g17726 and P2_R1312_U174 P2_R1312_U173 P2_U3139 ; P2_R1312_U120
g17727 and P2_R1312_U168 P2_R1312_U38 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U121
g17728 and P2_R1312_U161 P2_R1312_U48 P2_R1312_U164 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U122
g17729 and P2_R1312_U169 P2_R1312_U168 ; P2_R1312_U123
g17730 and P2_R1312_U160 P2_R1312_U44 P2_R1312_U168 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U124
g17731 and P2_U3132 P2_R1312_U16 ; P2_R1312_U125
g17732 and P2_R1312_U167 P2_R1312_U39 ; P2_R1312_U126
g17733 and P2_R1312_U17 P2_R1312_U168 P2_R1312_U126 ; P2_R1312_U127
g17734 and P2_R1312_U6 P2_U3136 ; P2_R1312_U128
g17735 and P2_R1312_U168 P2_R1312_U28 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U129
g17736 and P2_U3138 P2_R1312_U173 ; P2_R1312_U130
g17737 and P2_R1312_U168 P2_R1312_U32 P2_R1312_U167 P2_R1312_U166 ; P2_R1312_U131
g17738 and P2_R1312_U133 P2_R1312_U13 ; P2_R1312_U132
g17739 and P2_U3142 P2_R1312_U177 ; P2_R1312_U133
g17740 and P2_R1312_U167 P2_R1312_U34 P2_R1312_U177 P2_R1312_U168 ; P2_R1312_U134
g17741 and P2_R1312_U13 P2_R1312_U136 ; P2_R1312_U135
g17742 and P2_R1312_U179 P2_R1312_U178 P2_U3144 ; P2_R1312_U136
g17743 and P2_R1312_U157 P2_R1312_U156 P2_R1312_U154 P2_R1312_U36 P2_R1312_U166 ; P2_R1312_U137
g17744 and P2_U3148 P2_R1312_U8 P2_R1312_U168 P2_R1312_U167 ; P2_R1312_U138
g17745 and P2_R1312_U167 P2_R1312_U52 P2_R1312_U221 P2_R1312_U168 ; P2_R1312_U139
g17746 and P2_U3150 P2_R1312_U12 ; P2_R1312_U140
g17747 and P2_R1312_U181 P2_R1312_U153 ; P2_R1312_U141
g17748 and P2_R1312_U192 P2_R1312_U188 ; P2_R1312_U142
g17749 and P2_R1312_U199 P2_R1312_U197 P2_R1312_U198 ; P2_R1312_U143
g17750 and P2_R1312_U142 P2_R1312_U141 P2_R1312_U143 ; P2_R1312_U144
g17751 and P2_R1312_U203 P2_R1312_U202 ; P2_R1312_U145
g17752 and P2_R1312_U205 P2_R1312_U204 ; P2_R1312_U146
g17753 and P2_R1312_U201 P2_R1312_U200 P2_R1312_U145 P2_R1312_U146 P2_R1312_U206 ; P2_R1312_U147
g17754 and P2_R1312_U210 P2_R1312_U209 ; P2_R1312_U148
g17755 and P2_R1312_U214 P2_R1312_U215 ; P2_R1312_U149
g17756 and P2_R1312_U208 P2_R1312_U207 P2_R1312_U148 P2_R1312_U149 P2_R1312_U211 ; P2_R1312_U150
g17757 and P2_R1312_U219 P2_R1312_U218 P2_R1312_U217 P2_R1312_U216 ; P2_R1312_U151
g17758 and P2_R1312_U10 P2_R1312_U220 P2_R1312_U222 ; P2_R1312_U152
g17759 nand P2_R1312_U81 P2_R1312_U191 ; P2_R1312_U153
g17760 nand P2_U3115 P2_R1312_U68 ; P2_R1312_U154
g17761 nand P2_U3116 P2_R1312_U78 ; P2_R1312_U155
g17762 nand P2_U3114 P2_R1312_U67 ; P2_R1312_U156
g17763 nand P2_U3113 P2_R1312_U71 ; P2_R1312_U157
g17764 nand P2_U3104 P2_R1312_U74 ; P2_R1312_U158
g17765 nand P2_U3100 P2_R1312_U73 ; P2_R1312_U159
g17766 nand P2_U3099 P2_R1312_U63 ; P2_R1312_U160
g17767 nand P2_U3097 P2_R1312_U62 ; P2_R1312_U161
g17768 nand P2_U3098 P2_R1312_U72 ; P2_R1312_U162
g17769 nand P2_U3094 P2_R1312_U23 ; P2_R1312_U163
g17770 nand P2_U3096 P2_R1312_U61 ; P2_R1312_U164
g17771 nand P2_U3093 P2_R1312_U56 ; P2_R1312_U165
g17772 nand P2_U3090 P2_R1312_U80 ; P2_R1312_U166
g17773 nand P2_U3091 P2_R1312_U24 ; P2_R1312_U167
g17774 nand P2_U3092 P2_R1312_U57 ; P2_R1312_U168
g17775 nand P2_U3095 P2_R1312_U55 ; P2_R1312_U169
g17776 nand P2_U3102 P2_R1312_U64 ; P2_R1312_U170
g17777 nand P2_U3101 P2_R1312_U69 ; P2_R1312_U171
g17778 nand P2_U3103 P2_R1312_U65 ; P2_R1312_U172
g17779 nand P2_U3105 P2_R1312_U66 ; P2_R1312_U173
g17780 nand P2_U3106 P2_R1312_U75 ; P2_R1312_U174
g17781 nand P2_U3108 P2_R1312_U58 ; P2_R1312_U175
g17782 nand P2_U3107 P2_R1312_U70 ; P2_R1312_U176
g17783 nand P2_U3109 P2_R1312_U59 ; P2_R1312_U177
g17784 nand P2_U3110 P2_R1312_U76 ; P2_R1312_U178
g17785 nand P2_U3111 P2_R1312_U60 ; P2_R1312_U179
g17786 nand P2_U3112 P2_R1312_U77 ; P2_R1312_U180
g17787 nand P2_R1312_U8 P2_R1312_U87 P2_R1312_U15 P2_R1312_U86 ; P2_R1312_U181
g17788 nand P2_U3117 P2_R1312_U50 ; P2_R1312_U182
g17789 nand P2_U3118 P2_R1312_U79 ; P2_R1312_U183
g17790 nand P2_U3152 P2_U3153 ; P2_R1312_U184
g17791 nand P2_U3120 P2_R1312_U184 ; P2_R1312_U185
g17792 nand P2_U3119 P2_R1312_U54 ; P2_R1312_U186
g17793 or P2_U3152 P2_U3153 ; P2_R1312_U187
g17794 nand P2_R1312_U15 P2_R1312_U90 P2_R1312_U89 ; P2_R1312_U188
g17795 nand P2_R1312_U165 P2_R1312_U40 P2_R1312_U167 P2_U3126 P2_R1312_U168 ; P2_R1312_U189
g17796 nand P2_U3123 P2_R1312_U21 ; P2_R1312_U190
g17797 nand P2_R1312_U190 P2_R1312_U189 ; P2_R1312_U191
g17798 nand P2_R1312_U8 P2_R1312_U93 P2_R1312_U168 P2_R1312_U15 P2_R1312_U92 ; P2_R1312_U192
g17799 nand P2_R1312_U94 P2_R1312_U16 ; P2_R1312_U193
g17800 nand P2_U3125 P2_R1312_U20 ; P2_R1312_U194
g17801 nand P2_U3124 P2_R1312_U22 ; P2_R1312_U195
g17802 nand P2_R1312_U95 P2_R1312_U193 ; P2_R1312_U196
g17803 nand P2_R1312_U17 P2_R1312_U196 P2_R1312_U96 ; P2_R1312_U197
g17804 nand P2_R1312_U98 P2_R1312_U15 P2_R1312_U166 P2_R1312_U97 ; P2_R1312_U198
g17805 nand P2_R1312_U100 P2_R1312_U15 P2_R1312_U99 ; P2_R1312_U199
g17806 nand P2_R1312_U15 P2_R1312_U102 P2_R1312_U166 P2_R1312_U101 ; P2_R1312_U200
g17807 nand P2_U3128 P2_R1312_U16 P2_R1312_U17 P2_R1312_U169 P2_R1312_U104 ; P2_R1312_U201
g17808 nand P2_U3129 P2_R1312_U16 P2_R1312_U17 P2_R1312_U169 P2_R1312_U105 ; P2_R1312_U202
g17809 nand P2_R1312_U17 P2_R1312_U14 P2_R1312_U107 P2_R1312_U166 P2_R1312_U106 ; P2_R1312_U203
g17810 nand P2_R1312_U17 P2_R1312_U11 P2_R1312_U109 P2_R1312_U166 P2_R1312_U108 ; P2_R1312_U204
g17811 nand P2_R1312_U110 P2_R1312_U111 ; P2_R1312_U205
g17812 nand P2_R1312_U114 P2_R1312_U15 P2_R1312_U113 ; P2_R1312_U206
g17813 nand P2_U3146 P2_R1312_U8 P2_R1312_U168 P2_R1312_U15 P2_R1312_U115 ; P2_R1312_U207
g17814 nand P2_U3147 P2_R1312_U8 P2_R1312_U168 P2_R1312_U15 P2_R1312_U116 ; P2_R1312_U208
g17815 nand P2_R1312_U17 P2_R1312_U11 P2_R1312_U118 P2_R1312_U117 ; P2_R1312_U209
g17816 nand P2_R1312_U120 P2_R1312_U15 P2_R1312_U119 ; P2_R1312_U210
g17817 nand P2_R1312_U8 P2_U3145 P2_R1312_U15 P2_R1312_U121 ; P2_R1312_U211
g17818 nand P2_R1312_U227 P2_R1312_U226 P2_R1312_U223 ; P2_R1312_U212
g17819 nand P2_R1312_U17 P2_U3122 P2_R1312_U19 ; P2_R1312_U213
g17820 nand P2_U3130 P2_R1312_U16 P2_R1312_U17 P2_R1312_U123 P2_R1312_U122 ; P2_R1312_U214
g17821 nand P2_R1312_U14 P2_R1312_U169 P2_R1312_U17 P2_R1312_U125 P2_R1312_U124 ; P2_R1312_U215
g17822 nand P2_R1312_U11 P2_R1312_U128 P2_R1312_U16 P2_R1312_U166 P2_R1312_U127 ; P2_R1312_U216
g17823 nand P2_R1312_U130 P2_R1312_U15 P2_R1312_U129 ; P2_R1312_U217
g17824 nand P2_R1312_U15 P2_R1312_U132 P2_R1312_U131 ; P2_R1312_U218
g17825 nand P2_R1312_U15 P2_R1312_U135 P2_R1312_U166 P2_R1312_U134 ; P2_R1312_U219
g17826 nand P2_R1312_U15 P2_R1312_U138 P2_R1312_U137 ; P2_R1312_U220
g17827 nand P2_U3117 P2_R1312_U50 ; P2_R1312_U221
g17828 nand P2_R1312_U8 P2_R1312_U140 P2_R1312_U15 P2_R1312_U166 P2_R1312_U139 ; P2_R1312_U222
g17829 nand P2_U3121 P2_U3089 ; P2_R1312_U223
g17830 nand P2_U3089 P2_R1312_U26 ; P2_R1312_U224
g17831 nand P2_U3121 P2_R1312_U25 ; P2_R1312_U225
g17832 or P2_U3154 P2_U3121 ; P2_R1312_U226
g17833 nand P2_U3154 P2_R1312_U25 ; P2_R1312_U227
g17834 not P2_U3061 ; P2_R1335_U6
g17835 not P2_U3058 ; P2_R1335_U7
g17836 and P2_R1335_U10 P2_R1335_U9 ; P2_R1335_U8
g17837 nand P2_U3058 P2_R1335_U6 ; P2_R1335_U9
g17838 nand P2_U3061 P2_R1335_U7 ; P2_R1335_U10
g17839 and P2_R1209_U95 P2_R1209_U94 ; P2_R1209_U4
g17840 and P2_R1209_U96 P2_R1209_U97 ; P2_R1209_U5
g17841 and P2_R1209_U113 P2_R1209_U112 ; P2_R1209_U6
g17842 and P2_R1209_U155 P2_R1209_U154 ; P2_R1209_U7
g17843 and P2_R1209_U164 P2_R1209_U163 ; P2_R1209_U8
g17844 and P2_R1209_U182 P2_R1209_U181 ; P2_R1209_U9
g17845 and P2_R1209_U218 P2_R1209_U215 ; P2_R1209_U10
g17846 and P2_R1209_U211 P2_R1209_U208 ; P2_R1209_U11
g17847 and P2_R1209_U202 P2_R1209_U199 ; P2_R1209_U12
g17848 and P2_R1209_U196 P2_R1209_U192 ; P2_R1209_U13
g17849 and P2_R1209_U151 P2_R1209_U148 ; P2_R1209_U14
g17850 and P2_R1209_U143 P2_R1209_U140 ; P2_R1209_U15
g17851 and P2_R1209_U129 P2_R1209_U126 ; P2_R1209_U16
g17852 not P2_REG1_REG_6__SCAN_IN ; P2_R1209_U17
g17853 not P2_U3446 ; P2_R1209_U18
g17854 not P2_U3449 ; P2_R1209_U19
g17855 nand P2_U3446 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U20
g17856 not P2_REG1_REG_7__SCAN_IN ; P2_R1209_U21
g17857 not P2_REG1_REG_4__SCAN_IN ; P2_R1209_U22
g17858 not P2_U3440 ; P2_R1209_U23
g17859 not P2_U3443 ; P2_R1209_U24
g17860 not P2_REG1_REG_2__SCAN_IN ; P2_R1209_U25
g17861 not P2_U3434 ; P2_R1209_U26
g17862 not P2_REG1_REG_0__SCAN_IN ; P2_R1209_U27
g17863 not P2_U3425 ; P2_R1209_U28
g17864 nand P2_U3425 P2_REG1_REG_0__SCAN_IN ; P2_R1209_U29
g17865 not P2_REG1_REG_3__SCAN_IN ; P2_R1209_U30
g17866 not P2_U3437 ; P2_R1209_U31
g17867 nand P2_U3440 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U32
g17868 not P2_REG1_REG_5__SCAN_IN ; P2_R1209_U33
g17869 not P2_REG1_REG_8__SCAN_IN ; P2_R1209_U34
g17870 not P2_U3452 ; P2_R1209_U35
g17871 not P2_U3455 ; P2_R1209_U36
g17872 not P2_REG1_REG_9__SCAN_IN ; P2_R1209_U37
g17873 nand P2_R1209_U49 P2_R1209_U121 ; P2_R1209_U38
g17874 nand P2_R1209_U110 P2_R1209_U108 P2_R1209_U109 ; P2_R1209_U39
g17875 nand P2_R1209_U98 P2_R1209_U99 ; P2_R1209_U40
g17876 nand P2_U3431 P2_REG1_REG_1__SCAN_IN ; P2_R1209_U41
g17877 nand P2_R1209_U136 P2_R1209_U134 P2_R1209_U135 ; P2_R1209_U42
g17878 nand P2_R1209_U132 P2_R1209_U131 ; P2_R1209_U43
g17879 not P2_REG1_REG_16__SCAN_IN ; P2_R1209_U44
g17880 not P2_U3476 ; P2_R1209_U45
g17881 not P2_U3479 ; P2_R1209_U46
g17882 nand P2_U3476 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U47
g17883 not P2_REG1_REG_17__SCAN_IN ; P2_R1209_U48
g17884 nand P2_U3452 P2_REG1_REG_8__SCAN_IN ; P2_R1209_U49
g17885 not P2_REG1_REG_10__SCAN_IN ; P2_R1209_U50
g17886 not P2_U3458 ; P2_R1209_U51
g17887 not P2_REG1_REG_12__SCAN_IN ; P2_R1209_U52
g17888 not P2_U3464 ; P2_R1209_U53
g17889 not P2_REG1_REG_11__SCAN_IN ; P2_R1209_U54
g17890 not P2_U3461 ; P2_R1209_U55
g17891 nand P2_U3461 P2_REG1_REG_11__SCAN_IN ; P2_R1209_U56
g17892 not P2_REG1_REG_13__SCAN_IN ; P2_R1209_U57
g17893 not P2_U3467 ; P2_R1209_U58
g17894 not P2_REG1_REG_14__SCAN_IN ; P2_R1209_U59
g17895 not P2_U3470 ; P2_R1209_U60
g17896 not P2_REG1_REG_15__SCAN_IN ; P2_R1209_U61
g17897 not P2_U3473 ; P2_R1209_U62
g17898 not P2_REG1_REG_18__SCAN_IN ; P2_R1209_U63
g17899 not P2_U3482 ; P2_R1209_U64
g17900 nand P2_R1209_U186 P2_R1209_U185 P2_R1209_U187 ; P2_R1209_U65
g17901 nand P2_R1209_U179 P2_R1209_U178 ; P2_R1209_U66
g17902 nand P2_R1209_U56 P2_R1209_U204 ; P2_R1209_U67
g17903 nand P2_R1209_U259 P2_R1209_U258 ; P2_R1209_U68
g17904 nand P2_R1209_U308 P2_R1209_U307 ; P2_R1209_U69
g17905 nand P2_R1209_U231 P2_R1209_U230 ; P2_R1209_U70
g17906 nand P2_R1209_U236 P2_R1209_U235 ; P2_R1209_U71
g17907 nand P2_R1209_U243 P2_R1209_U242 ; P2_R1209_U72
g17908 nand P2_R1209_U250 P2_R1209_U249 ; P2_R1209_U73
g17909 nand P2_R1209_U255 P2_R1209_U254 ; P2_R1209_U74
g17910 nand P2_R1209_U271 P2_R1209_U270 ; P2_R1209_U75
g17911 nand P2_R1209_U278 P2_R1209_U277 ; P2_R1209_U76
g17912 nand P2_R1209_U285 P2_R1209_U284 ; P2_R1209_U77
g17913 nand P2_R1209_U292 P2_R1209_U291 ; P2_R1209_U78
g17914 nand P2_R1209_U299 P2_R1209_U298 ; P2_R1209_U79
g17915 nand P2_R1209_U304 P2_R1209_U303 ; P2_R1209_U80
g17916 nand P2_R1209_U117 P2_R1209_U116 P2_R1209_U118 ; P2_R1209_U81
g17917 nand P2_R1209_U133 P2_R1209_U145 ; P2_R1209_U82
g17918 nand P2_R1209_U41 P2_R1209_U152 ; P2_R1209_U83
g17919 not P2_U3424 ; P2_R1209_U84
g17920 not P2_REG1_REG_19__SCAN_IN ; P2_R1209_U85
g17921 nand P2_R1209_U175 P2_R1209_U174 ; P2_R1209_U86
g17922 nand P2_R1209_U171 P2_R1209_U170 ; P2_R1209_U87
g17923 nand P2_R1209_U161 P2_R1209_U160 ; P2_R1209_U88
g17924 not P2_R1209_U32 ; P2_R1209_U89
g17925 nand P2_U3455 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U90
g17926 nand P2_U3464 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U91
g17927 not P2_R1209_U56 ; P2_R1209_U92
g17928 not P2_R1209_U49 ; P2_R1209_U93
g17929 or P2_U3443 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U94
g17930 or P2_U3440 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U95
g17931 or P2_U3437 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U96
g17932 or P2_U3434 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U97
g17933 not P2_R1209_U29 ; P2_R1209_U98
g17934 or P2_U3431 P2_REG1_REG_1__SCAN_IN ; P2_R1209_U99
g17935 not P2_R1209_U40 ; P2_R1209_U100
g17936 not P2_R1209_U41 ; P2_R1209_U101
g17937 nand P2_R1209_U40 P2_R1209_U41 ; P2_R1209_U102
g17938 nand P2_U3434 P2_R1209_U96 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U103
g17939 nand P2_R1209_U5 P2_R1209_U102 ; P2_R1209_U104
g17940 nand P2_U3437 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U105
g17941 nand P2_R1209_U105 P2_R1209_U103 P2_R1209_U104 ; P2_R1209_U106
g17942 nand P2_R1209_U33 P2_R1209_U32 ; P2_R1209_U107
g17943 nand P2_U3443 P2_R1209_U107 ; P2_R1209_U108
g17944 nand P2_R1209_U4 P2_R1209_U106 ; P2_R1209_U109
g17945 nand P2_R1209_U89 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U110
g17946 not P2_R1209_U39 ; P2_R1209_U111
g17947 or P2_U3449 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U112
g17948 or P2_U3446 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U113
g17949 not P2_R1209_U20 ; P2_R1209_U114
g17950 nand P2_R1209_U21 P2_R1209_U20 ; P2_R1209_U115
g17951 nand P2_U3449 P2_R1209_U115 ; P2_R1209_U116
g17952 nand P2_R1209_U114 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U117
g17953 nand P2_R1209_U6 P2_R1209_U39 ; P2_R1209_U118
g17954 not P2_R1209_U81 ; P2_R1209_U119
g17955 or P2_U3452 P2_REG1_REG_8__SCAN_IN ; P2_R1209_U120
g17956 nand P2_R1209_U120 P2_R1209_U81 ; P2_R1209_U121
g17957 not P2_R1209_U38 ; P2_R1209_U122
g17958 or P2_U3455 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U123
g17959 or P2_U3446 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U124
g17960 nand P2_R1209_U124 P2_R1209_U39 ; P2_R1209_U125
g17961 nand P2_R1209_U238 P2_R1209_U237 P2_R1209_U20 P2_R1209_U125 ; P2_R1209_U126
g17962 nand P2_R1209_U111 P2_R1209_U20 ; P2_R1209_U127
g17963 nand P2_U3449 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U128
g17964 nand P2_R1209_U128 P2_R1209_U6 P2_R1209_U127 ; P2_R1209_U129
g17965 or P2_U3446 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U130
g17966 nand P2_R1209_U101 P2_R1209_U97 ; P2_R1209_U131
g17967 nand P2_U3434 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U132
g17968 not P2_R1209_U43 ; P2_R1209_U133
g17969 nand P2_R1209_U100 P2_R1209_U5 ; P2_R1209_U134
g17970 nand P2_R1209_U43 P2_R1209_U96 ; P2_R1209_U135
g17971 nand P2_U3437 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U136
g17972 not P2_R1209_U42 ; P2_R1209_U137
g17973 or P2_U3440 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U138
g17974 nand P2_R1209_U138 P2_R1209_U42 ; P2_R1209_U139
g17975 nand P2_R1209_U245 P2_R1209_U244 P2_R1209_U32 P2_R1209_U139 ; P2_R1209_U140
g17976 nand P2_R1209_U137 P2_R1209_U32 ; P2_R1209_U141
g17977 nand P2_U3443 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U142
g17978 nand P2_R1209_U142 P2_R1209_U4 P2_R1209_U141 ; P2_R1209_U143
g17979 or P2_U3440 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U144
g17980 nand P2_R1209_U100 P2_R1209_U97 ; P2_R1209_U145
g17981 not P2_R1209_U82 ; P2_R1209_U146
g17982 nand P2_U3437 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U147
g17983 nand P2_R1209_U257 P2_R1209_U256 P2_R1209_U41 P2_R1209_U40 ; P2_R1209_U148
g17984 nand P2_R1209_U41 P2_R1209_U40 ; P2_R1209_U149
g17985 nand P2_U3434 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U150
g17986 nand P2_R1209_U150 P2_R1209_U97 P2_R1209_U149 ; P2_R1209_U151
g17987 or P2_U3431 P2_REG1_REG_1__SCAN_IN ; P2_R1209_U152
g17988 not P2_R1209_U83 ; P2_R1209_U153
g17989 or P2_U3455 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U154
g17990 or P2_U3458 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U155
g17991 nand P2_R1209_U93 P2_R1209_U7 ; P2_R1209_U156
g17992 nand P2_U3458 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U157
g17993 nand P2_R1209_U157 P2_R1209_U90 P2_R1209_U156 ; P2_R1209_U158
g17994 or P2_U3458 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U159
g17995 nand P2_R1209_U120 P2_R1209_U7 P2_R1209_U81 ; P2_R1209_U160
g17996 nand P2_R1209_U159 P2_R1209_U158 ; P2_R1209_U161
g17997 not P2_R1209_U88 ; P2_R1209_U162
g17998 or P2_U3467 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U163
g17999 or P2_U3464 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U164
g18000 nand P2_R1209_U92 P2_R1209_U8 ; P2_R1209_U165
g18001 nand P2_U3467 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U166
g18002 nand P2_R1209_U166 P2_R1209_U91 P2_R1209_U165 ; P2_R1209_U167
g18003 or P2_U3461 P2_REG1_REG_11__SCAN_IN ; P2_R1209_U168
g18004 or P2_U3467 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U169
g18005 nand P2_R1209_U168 P2_R1209_U8 P2_R1209_U88 ; P2_R1209_U170
g18006 nand P2_R1209_U169 P2_R1209_U167 ; P2_R1209_U171
g18007 not P2_R1209_U87 ; P2_R1209_U172
g18008 or P2_U3470 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U173
g18009 nand P2_R1209_U173 P2_R1209_U87 ; P2_R1209_U174
g18010 nand P2_U3470 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U175
g18011 not P2_R1209_U86 ; P2_R1209_U176
g18012 or P2_U3473 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U177
g18013 nand P2_R1209_U177 P2_R1209_U86 ; P2_R1209_U178
g18014 nand P2_U3473 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U179
g18015 not P2_R1209_U66 ; P2_R1209_U180
g18016 or P2_U3479 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U181
g18017 or P2_U3476 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U182
g18018 not P2_R1209_U47 ; P2_R1209_U183
g18019 nand P2_R1209_U48 P2_R1209_U47 ; P2_R1209_U184
g18020 nand P2_U3479 P2_R1209_U184 ; P2_R1209_U185
g18021 nand P2_R1209_U183 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U186
g18022 nand P2_R1209_U9 P2_R1209_U66 ; P2_R1209_U187
g18023 not P2_R1209_U65 ; P2_R1209_U188
g18024 or P2_U3482 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U189
g18025 nand P2_R1209_U189 P2_R1209_U65 ; P2_R1209_U190
g18026 nand P2_U3482 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U191
g18027 nand P2_R1209_U261 P2_R1209_U260 P2_R1209_U191 P2_R1209_U190 ; P2_R1209_U192
g18028 nand P2_U3482 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U193
g18029 nand P2_R1209_U188 P2_R1209_U193 ; P2_R1209_U194
g18030 or P2_U3482 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U195
g18031 nand P2_R1209_U195 P2_R1209_U264 P2_R1209_U194 ; P2_R1209_U196
g18032 or P2_U3476 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U197
g18033 nand P2_R1209_U197 P2_R1209_U66 ; P2_R1209_U198
g18034 nand P2_R1209_U273 P2_R1209_U272 P2_R1209_U47 P2_R1209_U198 ; P2_R1209_U199
g18035 nand P2_R1209_U180 P2_R1209_U47 ; P2_R1209_U200
g18036 nand P2_U3479 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U201
g18037 nand P2_R1209_U201 P2_R1209_U9 P2_R1209_U200 ; P2_R1209_U202
g18038 or P2_U3476 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U203
g18039 nand P2_R1209_U168 P2_R1209_U88 ; P2_R1209_U204
g18040 not P2_R1209_U67 ; P2_R1209_U205
g18041 or P2_U3464 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U206
g18042 nand P2_R1209_U206 P2_R1209_U67 ; P2_R1209_U207
g18043 nand P2_R1209_U294 P2_R1209_U293 P2_R1209_U91 P2_R1209_U207 ; P2_R1209_U208
g18044 nand P2_R1209_U205 P2_R1209_U91 ; P2_R1209_U209
g18045 nand P2_U3467 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U210
g18046 nand P2_R1209_U210 P2_R1209_U8 P2_R1209_U209 ; P2_R1209_U211
g18047 or P2_U3464 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U212
g18048 or P2_U3455 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U213
g18049 nand P2_R1209_U213 P2_R1209_U38 ; P2_R1209_U214
g18050 nand P2_R1209_U306 P2_R1209_U305 P2_R1209_U90 P2_R1209_U214 ; P2_R1209_U215
g18051 nand P2_R1209_U122 P2_R1209_U90 ; P2_R1209_U216
g18052 nand P2_U3458 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U217
g18053 nand P2_R1209_U217 P2_R1209_U7 P2_R1209_U216 ; P2_R1209_U218
g18054 nand P2_R1209_U123 P2_R1209_U90 ; P2_R1209_U219
g18055 nand P2_R1209_U120 P2_R1209_U49 ; P2_R1209_U220
g18056 nand P2_R1209_U130 P2_R1209_U20 ; P2_R1209_U221
g18057 nand P2_R1209_U144 P2_R1209_U32 ; P2_R1209_U222
g18058 nand P2_R1209_U147 P2_R1209_U96 ; P2_R1209_U223
g18059 nand P2_R1209_U203 P2_R1209_U47 ; P2_R1209_U224
g18060 nand P2_R1209_U212 P2_R1209_U91 ; P2_R1209_U225
g18061 nand P2_R1209_U168 P2_R1209_U56 ; P2_R1209_U226
g18062 nand P2_U3455 P2_R1209_U37 ; P2_R1209_U227
g18063 nand P2_R1209_U36 P2_REG1_REG_9__SCAN_IN ; P2_R1209_U228
g18064 nand P2_R1209_U228 P2_R1209_U227 ; P2_R1209_U229
g18065 nand P2_R1209_U219 P2_R1209_U38 ; P2_R1209_U230
g18066 nand P2_R1209_U229 P2_R1209_U122 ; P2_R1209_U231
g18067 nand P2_U3452 P2_R1209_U34 ; P2_R1209_U232
g18068 nand P2_R1209_U35 P2_REG1_REG_8__SCAN_IN ; P2_R1209_U233
g18069 nand P2_R1209_U233 P2_R1209_U232 ; P2_R1209_U234
g18070 nand P2_R1209_U220 P2_R1209_U81 ; P2_R1209_U235
g18071 nand P2_R1209_U119 P2_R1209_U234 ; P2_R1209_U236
g18072 nand P2_U3449 P2_R1209_U21 ; P2_R1209_U237
g18073 nand P2_R1209_U19 P2_REG1_REG_7__SCAN_IN ; P2_R1209_U238
g18074 nand P2_U3446 P2_R1209_U17 ; P2_R1209_U239
g18075 nand P2_R1209_U18 P2_REG1_REG_6__SCAN_IN ; P2_R1209_U240
g18076 nand P2_R1209_U240 P2_R1209_U239 ; P2_R1209_U241
g18077 nand P2_R1209_U221 P2_R1209_U39 ; P2_R1209_U242
g18078 nand P2_R1209_U241 P2_R1209_U111 ; P2_R1209_U243
g18079 nand P2_U3443 P2_R1209_U33 ; P2_R1209_U244
g18080 nand P2_R1209_U24 P2_REG1_REG_5__SCAN_IN ; P2_R1209_U245
g18081 nand P2_U3440 P2_R1209_U22 ; P2_R1209_U246
g18082 nand P2_R1209_U23 P2_REG1_REG_4__SCAN_IN ; P2_R1209_U247
g18083 nand P2_R1209_U247 P2_R1209_U246 ; P2_R1209_U248
g18084 nand P2_R1209_U222 P2_R1209_U42 ; P2_R1209_U249
g18085 nand P2_R1209_U248 P2_R1209_U137 ; P2_R1209_U250
g18086 nand P2_U3437 P2_R1209_U30 ; P2_R1209_U251
g18087 nand P2_R1209_U31 P2_REG1_REG_3__SCAN_IN ; P2_R1209_U252
g18088 nand P2_R1209_U252 P2_R1209_U251 ; P2_R1209_U253
g18089 nand P2_R1209_U223 P2_R1209_U82 ; P2_R1209_U254
g18090 nand P2_R1209_U146 P2_R1209_U253 ; P2_R1209_U255
g18091 nand P2_U3434 P2_R1209_U25 ; P2_R1209_U256
g18092 nand P2_R1209_U26 P2_REG1_REG_2__SCAN_IN ; P2_R1209_U257
g18093 nand P2_R1209_U98 P2_R1209_U83 ; P2_R1209_U258
g18094 nand P2_R1209_U153 P2_R1209_U29 ; P2_R1209_U259
g18095 nand P2_U3424 P2_R1209_U85 ; P2_R1209_U260
g18096 nand P2_R1209_U84 P2_REG1_REG_19__SCAN_IN ; P2_R1209_U261
g18097 nand P2_U3424 P2_R1209_U85 ; P2_R1209_U262
g18098 nand P2_R1209_U84 P2_REG1_REG_19__SCAN_IN ; P2_R1209_U263
g18099 nand P2_R1209_U263 P2_R1209_U262 ; P2_R1209_U264
g18100 nand P2_U3482 P2_R1209_U63 ; P2_R1209_U265
g18101 nand P2_R1209_U64 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U266
g18102 nand P2_U3482 P2_R1209_U63 ; P2_R1209_U267
g18103 nand P2_R1209_U64 P2_REG1_REG_18__SCAN_IN ; P2_R1209_U268
g18104 nand P2_R1209_U268 P2_R1209_U267 ; P2_R1209_U269
g18105 nand P2_R1209_U266 P2_R1209_U265 P2_R1209_U65 ; P2_R1209_U270
g18106 nand P2_R1209_U269 P2_R1209_U188 ; P2_R1209_U271
g18107 nand P2_U3479 P2_R1209_U48 ; P2_R1209_U272
g18108 nand P2_R1209_U46 P2_REG1_REG_17__SCAN_IN ; P2_R1209_U273
g18109 nand P2_U3476 P2_R1209_U44 ; P2_R1209_U274
g18110 nand P2_R1209_U45 P2_REG1_REG_16__SCAN_IN ; P2_R1209_U275
g18111 nand P2_R1209_U275 P2_R1209_U274 ; P2_R1209_U276
g18112 nand P2_R1209_U224 P2_R1209_U66 ; P2_R1209_U277
g18113 nand P2_R1209_U276 P2_R1209_U180 ; P2_R1209_U278
g18114 nand P2_U3473 P2_R1209_U61 ; P2_R1209_U279
g18115 nand P2_R1209_U62 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U280
g18116 nand P2_U3473 P2_R1209_U61 ; P2_R1209_U281
g18117 nand P2_R1209_U62 P2_REG1_REG_15__SCAN_IN ; P2_R1209_U282
g18118 nand P2_R1209_U282 P2_R1209_U281 ; P2_R1209_U283
g18119 nand P2_R1209_U280 P2_R1209_U279 P2_R1209_U86 ; P2_R1209_U284
g18120 nand P2_R1209_U176 P2_R1209_U283 ; P2_R1209_U285
g18121 nand P2_U3470 P2_R1209_U59 ; P2_R1209_U286
g18122 nand P2_R1209_U60 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U287
g18123 nand P2_U3470 P2_R1209_U59 ; P2_R1209_U288
g18124 nand P2_R1209_U60 P2_REG1_REG_14__SCAN_IN ; P2_R1209_U289
g18125 nand P2_R1209_U289 P2_R1209_U288 ; P2_R1209_U290
g18126 nand P2_R1209_U287 P2_R1209_U286 P2_R1209_U87 ; P2_R1209_U291
g18127 nand P2_R1209_U172 P2_R1209_U290 ; P2_R1209_U292
g18128 nand P2_U3467 P2_R1209_U57 ; P2_R1209_U293
g18129 nand P2_R1209_U58 P2_REG1_REG_13__SCAN_IN ; P2_R1209_U294
g18130 nand P2_U3464 P2_R1209_U52 ; P2_R1209_U295
g18131 nand P2_R1209_U53 P2_REG1_REG_12__SCAN_IN ; P2_R1209_U296
g18132 nand P2_R1209_U296 P2_R1209_U295 ; P2_R1209_U297
g18133 nand P2_R1209_U225 P2_R1209_U67 ; P2_R1209_U298
g18134 nand P2_R1209_U297 P2_R1209_U205 ; P2_R1209_U299
g18135 nand P2_U3461 P2_R1209_U54 ; P2_R1209_U300
g18136 nand P2_R1209_U55 P2_REG1_REG_11__SCAN_IN ; P2_R1209_U301
g18137 nand P2_R1209_U301 P2_R1209_U300 ; P2_R1209_U302
g18138 nand P2_R1209_U226 P2_R1209_U88 ; P2_R1209_U303
g18139 nand P2_R1209_U162 P2_R1209_U302 ; P2_R1209_U304
g18140 nand P2_U3458 P2_R1209_U50 ; P2_R1209_U305
g18141 nand P2_R1209_U51 P2_REG1_REG_10__SCAN_IN ; P2_R1209_U306
g18142 nand P2_U3425 P2_R1209_U27 ; P2_R1209_U307
g18143 nand P2_R1209_U28 P2_REG1_REG_0__SCAN_IN ; P2_R1209_U308
g18144 and P2_R1170_U95 P2_R1170_U94 ; P2_R1170_U4
g18145 and P2_R1170_U96 P2_R1170_U97 ; P2_R1170_U5
g18146 and P2_R1170_U113 P2_R1170_U112 ; P2_R1170_U6
g18147 and P2_R1170_U155 P2_R1170_U154 ; P2_R1170_U7
g18148 and P2_R1170_U164 P2_R1170_U163 ; P2_R1170_U8
g18149 and P2_R1170_U182 P2_R1170_U181 ; P2_R1170_U9
g18150 and P2_R1170_U218 P2_R1170_U215 ; P2_R1170_U10
g18151 and P2_R1170_U211 P2_R1170_U208 ; P2_R1170_U11
g18152 and P2_R1170_U202 P2_R1170_U199 ; P2_R1170_U12
g18153 and P2_R1170_U196 P2_R1170_U192 ; P2_R1170_U13
g18154 and P2_R1170_U151 P2_R1170_U148 ; P2_R1170_U14
g18155 and P2_R1170_U143 P2_R1170_U140 ; P2_R1170_U15
g18156 and P2_R1170_U129 P2_R1170_U126 ; P2_R1170_U16
g18157 not P2_REG2_REG_6__SCAN_IN ; P2_R1170_U17
g18158 not P2_U3446 ; P2_R1170_U18
g18159 not P2_U3449 ; P2_R1170_U19
g18160 nand P2_U3446 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U20
g18161 not P2_REG2_REG_7__SCAN_IN ; P2_R1170_U21
g18162 not P2_REG2_REG_4__SCAN_IN ; P2_R1170_U22
g18163 not P2_U3440 ; P2_R1170_U23
g18164 not P2_U3443 ; P2_R1170_U24
g18165 not P2_REG2_REG_2__SCAN_IN ; P2_R1170_U25
g18166 not P2_U3434 ; P2_R1170_U26
g18167 not P2_REG2_REG_0__SCAN_IN ; P2_R1170_U27
g18168 not P2_U3425 ; P2_R1170_U28
g18169 nand P2_U3425 P2_REG2_REG_0__SCAN_IN ; P2_R1170_U29
g18170 not P2_REG2_REG_3__SCAN_IN ; P2_R1170_U30
g18171 not P2_U3437 ; P2_R1170_U31
g18172 nand P2_U3440 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U32
g18173 not P2_REG2_REG_5__SCAN_IN ; P2_R1170_U33
g18174 not P2_REG2_REG_8__SCAN_IN ; P2_R1170_U34
g18175 not P2_U3452 ; P2_R1170_U35
g18176 not P2_U3455 ; P2_R1170_U36
g18177 not P2_REG2_REG_9__SCAN_IN ; P2_R1170_U37
g18178 nand P2_R1170_U49 P2_R1170_U121 ; P2_R1170_U38
g18179 nand P2_R1170_U110 P2_R1170_U108 P2_R1170_U109 ; P2_R1170_U39
g18180 nand P2_R1170_U98 P2_R1170_U99 ; P2_R1170_U40
g18181 nand P2_U3431 P2_REG2_REG_1__SCAN_IN ; P2_R1170_U41
g18182 nand P2_R1170_U136 P2_R1170_U134 P2_R1170_U135 ; P2_R1170_U42
g18183 nand P2_R1170_U132 P2_R1170_U131 ; P2_R1170_U43
g18184 not P2_REG2_REG_16__SCAN_IN ; P2_R1170_U44
g18185 not P2_U3476 ; P2_R1170_U45
g18186 not P2_U3479 ; P2_R1170_U46
g18187 nand P2_U3476 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U47
g18188 not P2_REG2_REG_17__SCAN_IN ; P2_R1170_U48
g18189 nand P2_U3452 P2_REG2_REG_8__SCAN_IN ; P2_R1170_U49
g18190 not P2_REG2_REG_10__SCAN_IN ; P2_R1170_U50
g18191 not P2_U3458 ; P2_R1170_U51
g18192 not P2_REG2_REG_12__SCAN_IN ; P2_R1170_U52
g18193 not P2_U3464 ; P2_R1170_U53
g18194 not P2_REG2_REG_11__SCAN_IN ; P2_R1170_U54
g18195 not P2_U3461 ; P2_R1170_U55
g18196 nand P2_U3461 P2_REG2_REG_11__SCAN_IN ; P2_R1170_U56
g18197 not P2_REG2_REG_13__SCAN_IN ; P2_R1170_U57
g18198 not P2_U3467 ; P2_R1170_U58
g18199 not P2_REG2_REG_14__SCAN_IN ; P2_R1170_U59
g18200 not P2_U3470 ; P2_R1170_U60
g18201 not P2_REG2_REG_15__SCAN_IN ; P2_R1170_U61
g18202 not P2_U3473 ; P2_R1170_U62
g18203 not P2_REG2_REG_18__SCAN_IN ; P2_R1170_U63
g18204 not P2_U3482 ; P2_R1170_U64
g18205 nand P2_R1170_U186 P2_R1170_U185 P2_R1170_U187 ; P2_R1170_U65
g18206 nand P2_R1170_U179 P2_R1170_U178 ; P2_R1170_U66
g18207 nand P2_R1170_U56 P2_R1170_U204 ; P2_R1170_U67
g18208 nand P2_R1170_U259 P2_R1170_U258 ; P2_R1170_U68
g18209 nand P2_R1170_U308 P2_R1170_U307 ; P2_R1170_U69
g18210 nand P2_R1170_U231 P2_R1170_U230 ; P2_R1170_U70
g18211 nand P2_R1170_U236 P2_R1170_U235 ; P2_R1170_U71
g18212 nand P2_R1170_U243 P2_R1170_U242 ; P2_R1170_U72
g18213 nand P2_R1170_U250 P2_R1170_U249 ; P2_R1170_U73
g18214 nand P2_R1170_U255 P2_R1170_U254 ; P2_R1170_U74
g18215 nand P2_R1170_U271 P2_R1170_U270 ; P2_R1170_U75
g18216 nand P2_R1170_U278 P2_R1170_U277 ; P2_R1170_U76
g18217 nand P2_R1170_U285 P2_R1170_U284 ; P2_R1170_U77
g18218 nand P2_R1170_U292 P2_R1170_U291 ; P2_R1170_U78
g18219 nand P2_R1170_U299 P2_R1170_U298 ; P2_R1170_U79
g18220 nand P2_R1170_U304 P2_R1170_U303 ; P2_R1170_U80
g18221 nand P2_R1170_U117 P2_R1170_U116 P2_R1170_U118 ; P2_R1170_U81
g18222 nand P2_R1170_U133 P2_R1170_U145 ; P2_R1170_U82
g18223 nand P2_R1170_U41 P2_R1170_U152 ; P2_R1170_U83
g18224 not P2_U3424 ; P2_R1170_U84
g18225 not P2_REG2_REG_19__SCAN_IN ; P2_R1170_U85
g18226 nand P2_R1170_U175 P2_R1170_U174 ; P2_R1170_U86
g18227 nand P2_R1170_U171 P2_R1170_U170 ; P2_R1170_U87
g18228 nand P2_R1170_U161 P2_R1170_U160 ; P2_R1170_U88
g18229 not P2_R1170_U32 ; P2_R1170_U89
g18230 nand P2_U3455 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U90
g18231 nand P2_U3464 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U91
g18232 not P2_R1170_U56 ; P2_R1170_U92
g18233 not P2_R1170_U49 ; P2_R1170_U93
g18234 or P2_U3443 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U94
g18235 or P2_U3440 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U95
g18236 or P2_U3437 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U96
g18237 or P2_U3434 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U97
g18238 not P2_R1170_U29 ; P2_R1170_U98
g18239 or P2_U3431 P2_REG2_REG_1__SCAN_IN ; P2_R1170_U99
g18240 not P2_R1170_U40 ; P2_R1170_U100
g18241 not P2_R1170_U41 ; P2_R1170_U101
g18242 nand P2_R1170_U40 P2_R1170_U41 ; P2_R1170_U102
g18243 nand P2_U3434 P2_R1170_U96 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U103
g18244 nand P2_R1170_U5 P2_R1170_U102 ; P2_R1170_U104
g18245 nand P2_U3437 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U105
g18246 nand P2_R1170_U105 P2_R1170_U103 P2_R1170_U104 ; P2_R1170_U106
g18247 nand P2_R1170_U33 P2_R1170_U32 ; P2_R1170_U107
g18248 nand P2_U3443 P2_R1170_U107 ; P2_R1170_U108
g18249 nand P2_R1170_U4 P2_R1170_U106 ; P2_R1170_U109
g18250 nand P2_R1170_U89 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U110
g18251 not P2_R1170_U39 ; P2_R1170_U111
g18252 or P2_U3449 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U112
g18253 or P2_U3446 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U113
g18254 not P2_R1170_U20 ; P2_R1170_U114
g18255 nand P2_R1170_U21 P2_R1170_U20 ; P2_R1170_U115
g18256 nand P2_U3449 P2_R1170_U115 ; P2_R1170_U116
g18257 nand P2_R1170_U114 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U117
g18258 nand P2_R1170_U6 P2_R1170_U39 ; P2_R1170_U118
g18259 not P2_R1170_U81 ; P2_R1170_U119
g18260 or P2_U3452 P2_REG2_REG_8__SCAN_IN ; P2_R1170_U120
g18261 nand P2_R1170_U120 P2_R1170_U81 ; P2_R1170_U121
g18262 not P2_R1170_U38 ; P2_R1170_U122
g18263 or P2_U3455 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U123
g18264 or P2_U3446 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U124
g18265 nand P2_R1170_U124 P2_R1170_U39 ; P2_R1170_U125
g18266 nand P2_R1170_U238 P2_R1170_U237 P2_R1170_U20 P2_R1170_U125 ; P2_R1170_U126
g18267 nand P2_R1170_U111 P2_R1170_U20 ; P2_R1170_U127
g18268 nand P2_U3449 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U128
g18269 nand P2_R1170_U128 P2_R1170_U6 P2_R1170_U127 ; P2_R1170_U129
g18270 or P2_U3446 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U130
g18271 nand P2_R1170_U101 P2_R1170_U97 ; P2_R1170_U131
g18272 nand P2_U3434 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U132
g18273 not P2_R1170_U43 ; P2_R1170_U133
g18274 nand P2_R1170_U100 P2_R1170_U5 ; P2_R1170_U134
g18275 nand P2_R1170_U43 P2_R1170_U96 ; P2_R1170_U135
g18276 nand P2_U3437 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U136
g18277 not P2_R1170_U42 ; P2_R1170_U137
g18278 or P2_U3440 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U138
g18279 nand P2_R1170_U138 P2_R1170_U42 ; P2_R1170_U139
g18280 nand P2_R1170_U245 P2_R1170_U244 P2_R1170_U32 P2_R1170_U139 ; P2_R1170_U140
g18281 nand P2_R1170_U137 P2_R1170_U32 ; P2_R1170_U141
g18282 nand P2_U3443 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U142
g18283 nand P2_R1170_U142 P2_R1170_U4 P2_R1170_U141 ; P2_R1170_U143
g18284 or P2_U3440 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U144
g18285 nand P2_R1170_U100 P2_R1170_U97 ; P2_R1170_U145
g18286 not P2_R1170_U82 ; P2_R1170_U146
g18287 nand P2_U3437 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U147
g18288 nand P2_R1170_U257 P2_R1170_U256 P2_R1170_U41 P2_R1170_U40 ; P2_R1170_U148
g18289 nand P2_R1170_U41 P2_R1170_U40 ; P2_R1170_U149
g18290 nand P2_U3434 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U150
g18291 nand P2_R1170_U150 P2_R1170_U97 P2_R1170_U149 ; P2_R1170_U151
g18292 or P2_U3431 P2_REG2_REG_1__SCAN_IN ; P2_R1170_U152
g18293 not P2_R1170_U83 ; P2_R1170_U153
g18294 or P2_U3455 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U154
g18295 or P2_U3458 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U155
g18296 nand P2_R1170_U93 P2_R1170_U7 ; P2_R1170_U156
g18297 nand P2_U3458 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U157
g18298 nand P2_R1170_U157 P2_R1170_U90 P2_R1170_U156 ; P2_R1170_U158
g18299 or P2_U3458 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U159
g18300 nand P2_R1170_U120 P2_R1170_U7 P2_R1170_U81 ; P2_R1170_U160
g18301 nand P2_R1170_U159 P2_R1170_U158 ; P2_R1170_U161
g18302 not P2_R1170_U88 ; P2_R1170_U162
g18303 or P2_U3467 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U163
g18304 or P2_U3464 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U164
g18305 nand P2_R1170_U92 P2_R1170_U8 ; P2_R1170_U165
g18306 nand P2_U3467 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U166
g18307 nand P2_R1170_U166 P2_R1170_U91 P2_R1170_U165 ; P2_R1170_U167
g18308 or P2_U3461 P2_REG2_REG_11__SCAN_IN ; P2_R1170_U168
g18309 or P2_U3467 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U169
g18310 nand P2_R1170_U168 P2_R1170_U8 P2_R1170_U88 ; P2_R1170_U170
g18311 nand P2_R1170_U169 P2_R1170_U167 ; P2_R1170_U171
g18312 not P2_R1170_U87 ; P2_R1170_U172
g18313 or P2_U3470 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U173
g18314 nand P2_R1170_U173 P2_R1170_U87 ; P2_R1170_U174
g18315 nand P2_U3470 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U175
g18316 not P2_R1170_U86 ; P2_R1170_U176
g18317 or P2_U3473 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U177
g18318 nand P2_R1170_U177 P2_R1170_U86 ; P2_R1170_U178
g18319 nand P2_U3473 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U179
g18320 not P2_R1170_U66 ; P2_R1170_U180
g18321 or P2_U3479 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U181
g18322 or P2_U3476 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U182
g18323 not P2_R1170_U47 ; P2_R1170_U183
g18324 nand P2_R1170_U48 P2_R1170_U47 ; P2_R1170_U184
g18325 nand P2_U3479 P2_R1170_U184 ; P2_R1170_U185
g18326 nand P2_R1170_U183 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U186
g18327 nand P2_R1170_U9 P2_R1170_U66 ; P2_R1170_U187
g18328 not P2_R1170_U65 ; P2_R1170_U188
g18329 or P2_U3482 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U189
g18330 nand P2_R1170_U189 P2_R1170_U65 ; P2_R1170_U190
g18331 nand P2_U3482 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U191
g18332 nand P2_R1170_U261 P2_R1170_U260 P2_R1170_U191 P2_R1170_U190 ; P2_R1170_U192
g18333 nand P2_U3482 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U193
g18334 nand P2_R1170_U188 P2_R1170_U193 ; P2_R1170_U194
g18335 or P2_U3482 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U195
g18336 nand P2_R1170_U195 P2_R1170_U264 P2_R1170_U194 ; P2_R1170_U196
g18337 or P2_U3476 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U197
g18338 nand P2_R1170_U197 P2_R1170_U66 ; P2_R1170_U198
g18339 nand P2_R1170_U273 P2_R1170_U272 P2_R1170_U47 P2_R1170_U198 ; P2_R1170_U199
g18340 nand P2_R1170_U180 P2_R1170_U47 ; P2_R1170_U200
g18341 nand P2_U3479 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U201
g18342 nand P2_R1170_U201 P2_R1170_U9 P2_R1170_U200 ; P2_R1170_U202
g18343 or P2_U3476 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U203
g18344 nand P2_R1170_U168 P2_R1170_U88 ; P2_R1170_U204
g18345 not P2_R1170_U67 ; P2_R1170_U205
g18346 or P2_U3464 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U206
g18347 nand P2_R1170_U206 P2_R1170_U67 ; P2_R1170_U207
g18348 nand P2_R1170_U294 P2_R1170_U293 P2_R1170_U91 P2_R1170_U207 ; P2_R1170_U208
g18349 nand P2_R1170_U205 P2_R1170_U91 ; P2_R1170_U209
g18350 nand P2_U3467 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U210
g18351 nand P2_R1170_U210 P2_R1170_U8 P2_R1170_U209 ; P2_R1170_U211
g18352 or P2_U3464 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U212
g18353 or P2_U3455 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U213
g18354 nand P2_R1170_U213 P2_R1170_U38 ; P2_R1170_U214
g18355 nand P2_R1170_U306 P2_R1170_U305 P2_R1170_U90 P2_R1170_U214 ; P2_R1170_U215
g18356 nand P2_R1170_U122 P2_R1170_U90 ; P2_R1170_U216
g18357 nand P2_U3458 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U217
g18358 nand P2_R1170_U217 P2_R1170_U7 P2_R1170_U216 ; P2_R1170_U218
g18359 nand P2_R1170_U123 P2_R1170_U90 ; P2_R1170_U219
g18360 nand P2_R1170_U120 P2_R1170_U49 ; P2_R1170_U220
g18361 nand P2_R1170_U130 P2_R1170_U20 ; P2_R1170_U221
g18362 nand P2_R1170_U144 P2_R1170_U32 ; P2_R1170_U222
g18363 nand P2_R1170_U147 P2_R1170_U96 ; P2_R1170_U223
g18364 nand P2_R1170_U203 P2_R1170_U47 ; P2_R1170_U224
g18365 nand P2_R1170_U212 P2_R1170_U91 ; P2_R1170_U225
g18366 nand P2_R1170_U168 P2_R1170_U56 ; P2_R1170_U226
g18367 nand P2_U3455 P2_R1170_U37 ; P2_R1170_U227
g18368 nand P2_R1170_U36 P2_REG2_REG_9__SCAN_IN ; P2_R1170_U228
g18369 nand P2_R1170_U228 P2_R1170_U227 ; P2_R1170_U229
g18370 nand P2_R1170_U219 P2_R1170_U38 ; P2_R1170_U230
g18371 nand P2_R1170_U229 P2_R1170_U122 ; P2_R1170_U231
g18372 nand P2_U3452 P2_R1170_U34 ; P2_R1170_U232
g18373 nand P2_R1170_U35 P2_REG2_REG_8__SCAN_IN ; P2_R1170_U233
g18374 nand P2_R1170_U233 P2_R1170_U232 ; P2_R1170_U234
g18375 nand P2_R1170_U220 P2_R1170_U81 ; P2_R1170_U235
g18376 nand P2_R1170_U119 P2_R1170_U234 ; P2_R1170_U236
g18377 nand P2_U3449 P2_R1170_U21 ; P2_R1170_U237
g18378 nand P2_R1170_U19 P2_REG2_REG_7__SCAN_IN ; P2_R1170_U238
g18379 nand P2_U3446 P2_R1170_U17 ; P2_R1170_U239
g18380 nand P2_R1170_U18 P2_REG2_REG_6__SCAN_IN ; P2_R1170_U240
g18381 nand P2_R1170_U240 P2_R1170_U239 ; P2_R1170_U241
g18382 nand P2_R1170_U221 P2_R1170_U39 ; P2_R1170_U242
g18383 nand P2_R1170_U241 P2_R1170_U111 ; P2_R1170_U243
g18384 nand P2_U3443 P2_R1170_U33 ; P2_R1170_U244
g18385 nand P2_R1170_U24 P2_REG2_REG_5__SCAN_IN ; P2_R1170_U245
g18386 nand P2_U3440 P2_R1170_U22 ; P2_R1170_U246
g18387 nand P2_R1170_U23 P2_REG2_REG_4__SCAN_IN ; P2_R1170_U247
g18388 nand P2_R1170_U247 P2_R1170_U246 ; P2_R1170_U248
g18389 nand P2_R1170_U222 P2_R1170_U42 ; P2_R1170_U249
g18390 nand P2_R1170_U248 P2_R1170_U137 ; P2_R1170_U250
g18391 nand P2_U3437 P2_R1170_U30 ; P2_R1170_U251
g18392 nand P2_R1170_U31 P2_REG2_REG_3__SCAN_IN ; P2_R1170_U252
g18393 nand P2_R1170_U252 P2_R1170_U251 ; P2_R1170_U253
g18394 nand P2_R1170_U223 P2_R1170_U82 ; P2_R1170_U254
g18395 nand P2_R1170_U146 P2_R1170_U253 ; P2_R1170_U255
g18396 nand P2_U3434 P2_R1170_U25 ; P2_R1170_U256
g18397 nand P2_R1170_U26 P2_REG2_REG_2__SCAN_IN ; P2_R1170_U257
g18398 nand P2_R1170_U98 P2_R1170_U83 ; P2_R1170_U258
g18399 nand P2_R1170_U153 P2_R1170_U29 ; P2_R1170_U259
g18400 nand P2_U3424 P2_R1170_U85 ; P2_R1170_U260
g18401 nand P2_R1170_U84 P2_REG2_REG_19__SCAN_IN ; P2_R1170_U261
g18402 nand P2_U3424 P2_R1170_U85 ; P2_R1170_U262
g18403 nand P2_R1170_U84 P2_REG2_REG_19__SCAN_IN ; P2_R1170_U263
g18404 nand P2_R1170_U263 P2_R1170_U262 ; P2_R1170_U264
g18405 nand P2_U3482 P2_R1170_U63 ; P2_R1170_U265
g18406 nand P2_R1170_U64 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U266
g18407 nand P2_U3482 P2_R1170_U63 ; P2_R1170_U267
g18408 nand P2_R1170_U64 P2_REG2_REG_18__SCAN_IN ; P2_R1170_U268
g18409 nand P2_R1170_U268 P2_R1170_U267 ; P2_R1170_U269
g18410 nand P2_R1170_U266 P2_R1170_U265 P2_R1170_U65 ; P2_R1170_U270
g18411 nand P2_R1170_U269 P2_R1170_U188 ; P2_R1170_U271
g18412 nand P2_U3479 P2_R1170_U48 ; P2_R1170_U272
g18413 nand P2_R1170_U46 P2_REG2_REG_17__SCAN_IN ; P2_R1170_U273
g18414 nand P2_U3476 P2_R1170_U44 ; P2_R1170_U274
g18415 nand P2_R1170_U45 P2_REG2_REG_16__SCAN_IN ; P2_R1170_U275
g18416 nand P2_R1170_U275 P2_R1170_U274 ; P2_R1170_U276
g18417 nand P2_R1170_U224 P2_R1170_U66 ; P2_R1170_U277
g18418 nand P2_R1170_U276 P2_R1170_U180 ; P2_R1170_U278
g18419 nand P2_U3473 P2_R1170_U61 ; P2_R1170_U279
g18420 nand P2_R1170_U62 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U280
g18421 nand P2_U3473 P2_R1170_U61 ; P2_R1170_U281
g18422 nand P2_R1170_U62 P2_REG2_REG_15__SCAN_IN ; P2_R1170_U282
g18423 nand P2_R1170_U282 P2_R1170_U281 ; P2_R1170_U283
g18424 nand P2_R1170_U280 P2_R1170_U279 P2_R1170_U86 ; P2_R1170_U284
g18425 nand P2_R1170_U176 P2_R1170_U283 ; P2_R1170_U285
g18426 nand P2_U3470 P2_R1170_U59 ; P2_R1170_U286
g18427 nand P2_R1170_U60 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U287
g18428 nand P2_U3470 P2_R1170_U59 ; P2_R1170_U288
g18429 nand P2_R1170_U60 P2_REG2_REG_14__SCAN_IN ; P2_R1170_U289
g18430 nand P2_R1170_U289 P2_R1170_U288 ; P2_R1170_U290
g18431 nand P2_R1170_U287 P2_R1170_U286 P2_R1170_U87 ; P2_R1170_U291
g18432 nand P2_R1170_U172 P2_R1170_U290 ; P2_R1170_U292
g18433 nand P2_U3467 P2_R1170_U57 ; P2_R1170_U293
g18434 nand P2_R1170_U58 P2_REG2_REG_13__SCAN_IN ; P2_R1170_U294
g18435 nand P2_U3464 P2_R1170_U52 ; P2_R1170_U295
g18436 nand P2_R1170_U53 P2_REG2_REG_12__SCAN_IN ; P2_R1170_U296
g18437 nand P2_R1170_U296 P2_R1170_U295 ; P2_R1170_U297
g18438 nand P2_R1170_U225 P2_R1170_U67 ; P2_R1170_U298
g18439 nand P2_R1170_U297 P2_R1170_U205 ; P2_R1170_U299
g18440 nand P2_U3461 P2_R1170_U54 ; P2_R1170_U300
g18441 nand P2_R1170_U55 P2_REG2_REG_11__SCAN_IN ; P2_R1170_U301
g18442 nand P2_R1170_U301 P2_R1170_U300 ; P2_R1170_U302
g18443 nand P2_R1170_U226 P2_R1170_U88 ; P2_R1170_U303
g18444 nand P2_R1170_U162 P2_R1170_U302 ; P2_R1170_U304
g18445 nand P2_U3458 P2_R1170_U50 ; P2_R1170_U305
g18446 nand P2_R1170_U51 P2_REG2_REG_10__SCAN_IN ; P2_R1170_U306
g18447 nand P2_U3425 P2_R1170_U27 ; P2_R1170_U307
g18448 nand P2_R1170_U28 P2_REG2_REG_0__SCAN_IN ; P2_R1170_U308
g18449 and P2_R1275_U135 P2_R1275_U35 ; P2_R1275_U6
g18450 and P2_R1275_U133 P2_R1275_U36 ; P2_R1275_U7
g18451 and P2_R1275_U132 P2_R1275_U37 ; P2_R1275_U8
g18452 and P2_R1275_U131 P2_R1275_U38 ; P2_R1275_U9
g18453 and P2_R1275_U129 P2_R1275_U39 ; P2_R1275_U10
g18454 and P2_R1275_U128 P2_R1275_U40 ; P2_R1275_U11
g18455 and P2_R1275_U127 P2_R1275_U41 ; P2_R1275_U12
g18456 and P2_R1275_U125 P2_R1275_U42 ; P2_R1275_U13
g18457 and P2_R1275_U123 P2_R1275_U43 ; P2_R1275_U14
g18458 and P2_R1275_U121 P2_R1275_U44 ; P2_R1275_U15
g18459 and P2_R1275_U119 P2_R1275_U45 ; P2_R1275_U16
g18460 and P2_R1275_U117 P2_R1275_U46 ; P2_R1275_U17
g18461 and P2_R1275_U115 P2_R1275_U25 ; P2_R1275_U18
g18462 and P2_R1275_U113 P2_R1275_U67 ; P2_R1275_U19
g18463 and P2_R1275_U98 P2_R1275_U26 ; P2_R1275_U20
g18464 and P2_R1275_U97 P2_R1275_U27 ; P2_R1275_U21
g18465 and P2_R1275_U96 P2_R1275_U28 ; P2_R1275_U22
g18466 and P2_R1275_U94 P2_R1275_U29 ; P2_R1275_U23
g18467 and P2_R1275_U93 P2_R1275_U30 ; P2_R1275_U24
g18468 or P2_U3432 P2_U3427 P2_U3435 ; P2_R1275_U25
g18469 nand P2_R1275_U87 P2_R1275_U34 ; P2_R1275_U26
g18470 nand P2_R1275_U88 P2_R1275_U33 ; P2_R1275_U27
g18471 nand P2_R1275_U56 P2_R1275_U89 ; P2_R1275_U28
g18472 nand P2_R1275_U90 P2_R1275_U32 ; P2_R1275_U29
g18473 nand P2_R1275_U91 P2_R1275_U31 ; P2_R1275_U30
g18474 not P2_U3453 ; P2_R1275_U31
g18475 not P2_U3450 ; P2_R1275_U32
g18476 not P2_U3441 ; P2_R1275_U33
g18477 not P2_U3438 ; P2_R1275_U34
g18478 nand P2_R1275_U57 P2_R1275_U92 ; P2_R1275_U35
g18479 nand P2_R1275_U99 P2_R1275_U54 ; P2_R1275_U36
g18480 nand P2_R1275_U100 P2_R1275_U53 ; P2_R1275_U37
g18481 nand P2_R1275_U58 P2_R1275_U101 ; P2_R1275_U38
g18482 nand P2_R1275_U102 P2_R1275_U52 ; P2_R1275_U39
g18483 nand P2_R1275_U103 P2_R1275_U51 ; P2_R1275_U40
g18484 nand P2_R1275_U59 P2_R1275_U104 ; P2_R1275_U41
g18485 nand P2_R1275_U60 P2_R1275_U105 ; P2_R1275_U42
g18486 nand P2_R1275_U61 P2_R1275_U106 ; P2_R1275_U43
g18487 nand P2_R1275_U107 P2_R1275_U75 P2_R1275_U50 ; P2_R1275_U44
g18488 nand P2_R1275_U108 P2_R1275_U73 P2_R1275_U49 ; P2_R1275_U45
g18489 nand P2_R1275_U109 P2_R1275_U71 P2_R1275_U48 ; P2_R1275_U46
g18490 not P2_U3959 ; P2_R1275_U47
g18491 not P2_U3949 ; P2_R1275_U48
g18492 not P2_U3951 ; P2_R1275_U49
g18493 not P2_U3953 ; P2_R1275_U50
g18494 not P2_U3477 ; P2_R1275_U51
g18495 not P2_U3474 ; P2_R1275_U52
g18496 not P2_U3465 ; P2_R1275_U53
g18497 not P2_U3462 ; P2_R1275_U54
g18498 nand P2_R1275_U153 P2_R1275_U152 ; P2_R1275_U55
g18499 nor P2_U3444 P2_U3447 ; P2_R1275_U56
g18500 nor P2_U3459 P2_U3456 ; P2_R1275_U57
g18501 nor P2_U3468 P2_U3471 ; P2_R1275_U58
g18502 nor P2_U3480 P2_U3483 ; P2_R1275_U59
g18503 nor P2_U3485 P2_U3957 ; P2_R1275_U60
g18504 nor P2_U3956 P2_U3955 ; P2_R1275_U61
g18505 not P2_U3456 ; P2_R1275_U62
g18506 and P2_R1275_U137 P2_R1275_U136 ; P2_R1275_U63
g18507 not P2_U3444 ; P2_R1275_U64
g18508 and P2_R1275_U139 P2_R1275_U138 ; P2_R1275_U65
g18509 not P2_U3958 ; P2_R1275_U66
g18510 nand P2_R1275_U110 P2_R1275_U69 P2_R1275_U47 ; P2_R1275_U67
g18511 and P2_R1275_U141 P2_R1275_U140 ; P2_R1275_U68
g18512 not P2_U3960 ; P2_R1275_U69
g18513 and P2_R1275_U143 P2_R1275_U142 ; P2_R1275_U70
g18514 not P2_U3950 ; P2_R1275_U71
g18515 and P2_R1275_U145 P2_R1275_U144 ; P2_R1275_U72
g18516 not P2_U3952 ; P2_R1275_U73
g18517 and P2_R1275_U147 P2_R1275_U146 ; P2_R1275_U74
g18518 not P2_U3954 ; P2_R1275_U75
g18519 and P2_R1275_U149 P2_R1275_U148 ; P2_R1275_U76
g18520 not P2_U3956 ; P2_R1275_U77
g18521 and P2_R1275_U151 P2_R1275_U150 ; P2_R1275_U78
g18522 not P2_U3432 ; P2_R1275_U79
g18523 not P2_U3427 ; P2_R1275_U80
g18524 not P2_U3485 ; P2_R1275_U81
g18525 and P2_R1275_U155 P2_R1275_U154 ; P2_R1275_U82
g18526 not P2_U3480 ; P2_R1275_U83
g18527 and P2_R1275_U157 P2_R1275_U156 ; P2_R1275_U84
g18528 not P2_U3468 ; P2_R1275_U85
g18529 and P2_R1275_U159 P2_R1275_U158 ; P2_R1275_U86
g18530 not P2_R1275_U25 ; P2_R1275_U87
g18531 not P2_R1275_U26 ; P2_R1275_U88
g18532 not P2_R1275_U27 ; P2_R1275_U89
g18533 not P2_R1275_U28 ; P2_R1275_U90
g18534 not P2_R1275_U29 ; P2_R1275_U91
g18535 not P2_R1275_U30 ; P2_R1275_U92
g18536 nand P2_U3453 P2_R1275_U29 ; P2_R1275_U93
g18537 nand P2_U3450 P2_R1275_U28 ; P2_R1275_U94
g18538 nand P2_R1275_U89 P2_R1275_U64 ; P2_R1275_U95
g18539 nand P2_U3447 P2_R1275_U95 ; P2_R1275_U96
g18540 nand P2_U3441 P2_R1275_U26 ; P2_R1275_U97
g18541 nand P2_U3438 P2_R1275_U25 ; P2_R1275_U98
g18542 not P2_R1275_U35 ; P2_R1275_U99
g18543 not P2_R1275_U36 ; P2_R1275_U100
g18544 not P2_R1275_U37 ; P2_R1275_U101
g18545 not P2_R1275_U38 ; P2_R1275_U102
g18546 not P2_R1275_U39 ; P2_R1275_U103
g18547 not P2_R1275_U40 ; P2_R1275_U104
g18548 not P2_R1275_U41 ; P2_R1275_U105
g18549 not P2_R1275_U42 ; P2_R1275_U106
g18550 not P2_R1275_U43 ; P2_R1275_U107
g18551 not P2_R1275_U44 ; P2_R1275_U108
g18552 not P2_R1275_U45 ; P2_R1275_U109
g18553 not P2_R1275_U46 ; P2_R1275_U110
g18554 not P2_R1275_U67 ; P2_R1275_U111
g18555 nand P2_R1275_U110 P2_R1275_U69 ; P2_R1275_U112
g18556 nand P2_U3959 P2_R1275_U112 ; P2_R1275_U113
g18557 or P2_U3432 P2_U3427 ; P2_R1275_U114
g18558 nand P2_U3435 P2_R1275_U114 ; P2_R1275_U115
g18559 nand P2_R1275_U109 P2_R1275_U71 ; P2_R1275_U116
g18560 nand P2_U3949 P2_R1275_U116 ; P2_R1275_U117
g18561 nand P2_R1275_U108 P2_R1275_U73 ; P2_R1275_U118
g18562 nand P2_U3951 P2_R1275_U118 ; P2_R1275_U119
g18563 nand P2_R1275_U107 P2_R1275_U75 ; P2_R1275_U120
g18564 nand P2_U3953 P2_R1275_U120 ; P2_R1275_U121
g18565 nand P2_R1275_U106 P2_R1275_U77 ; P2_R1275_U122
g18566 nand P2_U3955 P2_R1275_U122 ; P2_R1275_U123
g18567 nand P2_R1275_U105 P2_R1275_U81 ; P2_R1275_U124
g18568 nand P2_U3957 P2_R1275_U124 ; P2_R1275_U125
g18569 nand P2_R1275_U104 P2_R1275_U83 ; P2_R1275_U126
g18570 nand P2_U3483 P2_R1275_U126 ; P2_R1275_U127
g18571 nand P2_U3477 P2_R1275_U39 ; P2_R1275_U128
g18572 nand P2_U3474 P2_R1275_U38 ; P2_R1275_U129
g18573 nand P2_R1275_U101 P2_R1275_U85 ; P2_R1275_U130
g18574 nand P2_U3471 P2_R1275_U130 ; P2_R1275_U131
g18575 nand P2_U3465 P2_R1275_U36 ; P2_R1275_U132
g18576 nand P2_U3462 P2_R1275_U35 ; P2_R1275_U133
g18577 nand P2_R1275_U92 P2_R1275_U62 ; P2_R1275_U134
g18578 nand P2_U3459 P2_R1275_U134 ; P2_R1275_U135
g18579 nand P2_U3456 P2_R1275_U30 ; P2_R1275_U136
g18580 nand P2_R1275_U92 P2_R1275_U62 ; P2_R1275_U137
g18581 nand P2_U3444 P2_R1275_U27 ; P2_R1275_U138
g18582 nand P2_R1275_U89 P2_R1275_U64 ; P2_R1275_U139
g18583 nand P2_U3958 P2_R1275_U67 ; P2_R1275_U140
g18584 nand P2_R1275_U111 P2_R1275_U66 ; P2_R1275_U141
g18585 nand P2_U3960 P2_R1275_U46 ; P2_R1275_U142
g18586 nand P2_R1275_U110 P2_R1275_U69 ; P2_R1275_U143
g18587 nand P2_U3950 P2_R1275_U45 ; P2_R1275_U144
g18588 nand P2_R1275_U109 P2_R1275_U71 ; P2_R1275_U145
g18589 nand P2_U3952 P2_R1275_U44 ; P2_R1275_U146
g18590 nand P2_R1275_U108 P2_R1275_U73 ; P2_R1275_U147
g18591 nand P2_U3954 P2_R1275_U43 ; P2_R1275_U148
g18592 nand P2_R1275_U107 P2_R1275_U75 ; P2_R1275_U149
g18593 nand P2_U3956 P2_R1275_U42 ; P2_R1275_U150
g18594 nand P2_R1275_U106 P2_R1275_U77 ; P2_R1275_U151
g18595 nand P2_U3432 P2_R1275_U80 ; P2_R1275_U152
g18596 nand P2_U3427 P2_R1275_U79 ; P2_R1275_U153
g18597 nand P2_U3485 P2_R1275_U41 ; P2_R1275_U154
g18598 nand P2_R1275_U105 P2_R1275_U81 ; P2_R1275_U155
g18599 nand P2_U3480 P2_R1275_U40 ; P2_R1275_U156
g18600 nand P2_R1275_U104 P2_R1275_U83 ; P2_R1275_U157
g18601 nand P2_U3468 P2_R1275_U37 ; P2_R1275_U158
g18602 nand P2_R1275_U101 P2_R1275_U85 ; P2_R1275_U159
g18603 and P2_R1179_U202 P2_R1179_U201 ; P2_R1179_U6
g18604 and P2_R1179_U241 P2_R1179_U240 ; P2_R1179_U7
g18605 and P2_R1179_U181 P2_R1179_U256 ; P2_R1179_U8
g18606 and P2_R1179_U258 P2_R1179_U257 ; P2_R1179_U9
g18607 and P2_R1179_U182 P2_R1179_U282 ; P2_R1179_U10
g18608 and P2_R1179_U284 P2_R1179_U283 ; P2_R1179_U11
g18609 nand P2_R1179_U344 P2_R1179_U347 ; P2_R1179_U12
g18610 nand P2_R1179_U333 P2_R1179_U336 ; P2_R1179_U13
g18611 nand P2_R1179_U322 P2_R1179_U325 ; P2_R1179_U14
g18612 nand P2_R1179_U314 P2_R1179_U316 ; P2_R1179_U15
g18613 nand P2_R1179_U352 P2_R1179_U312 ; P2_R1179_U16
g18614 nand P2_R1179_U235 P2_R1179_U237 ; P2_R1179_U17
g18615 nand P2_R1179_U227 P2_R1179_U230 ; P2_R1179_U18
g18616 nand P2_R1179_U219 P2_R1179_U221 ; P2_R1179_U19
g18617 nand P2_R1179_U166 P2_R1179_U350 ; P2_R1179_U20
g18618 not P2_U3450 ; P2_R1179_U21
g18619 not P2_U3444 ; P2_R1179_U22
g18620 not P2_U3435 ; P2_R1179_U23
g18621 not P2_U3427 ; P2_R1179_U24
g18622 not P2_U3080 ; P2_R1179_U25
g18623 not P2_U3438 ; P2_R1179_U26
g18624 not P2_U3070 ; P2_R1179_U27
g18625 nand P2_U3070 P2_R1179_U23 ; P2_R1179_U28
g18626 not P2_U3066 ; P2_R1179_U29
g18627 not P2_U3447 ; P2_R1179_U30
g18628 not P2_U3441 ; P2_R1179_U31
g18629 not P2_U3073 ; P2_R1179_U32
g18630 not P2_U3069 ; P2_R1179_U33
g18631 not P2_U3062 ; P2_R1179_U34
g18632 nand P2_U3062 P2_R1179_U31 ; P2_R1179_U35
g18633 not P2_U3453 ; P2_R1179_U36
g18634 not P2_U3072 ; P2_R1179_U37
g18635 nand P2_U3072 P2_R1179_U21 ; P2_R1179_U38
g18636 not P2_U3086 ; P2_R1179_U39
g18637 not P2_U3456 ; P2_R1179_U40
g18638 not P2_U3085 ; P2_R1179_U41
g18639 nand P2_R1179_U208 P2_R1179_U207 ; P2_R1179_U42
g18640 nand P2_R1179_U35 P2_R1179_U223 ; P2_R1179_U43
g18641 nand P2_R1179_U192 P2_R1179_U176 P2_R1179_U351 ; P2_R1179_U44
g18642 not P2_U3951 ; P2_R1179_U45
g18643 not P2_U3459 ; P2_R1179_U46
g18644 not P2_U3462 ; P2_R1179_U47
g18645 not P2_U3065 ; P2_R1179_U48
g18646 not P2_U3064 ; P2_R1179_U49
g18647 nand P2_U3085 P2_R1179_U40 ; P2_R1179_U50
g18648 not P2_U3465 ; P2_R1179_U51
g18649 not P2_U3074 ; P2_R1179_U52
g18650 not P2_U3468 ; P2_R1179_U53
g18651 not P2_U3082 ; P2_R1179_U54
g18652 not P2_U3477 ; P2_R1179_U55
g18653 not P2_U3474 ; P2_R1179_U56
g18654 not P2_U3471 ; P2_R1179_U57
g18655 not P2_U3075 ; P2_R1179_U58
g18656 not P2_U3076 ; P2_R1179_U59
g18657 not P2_U3081 ; P2_R1179_U60
g18658 nand P2_U3081 P2_R1179_U57 ; P2_R1179_U61
g18659 not P2_U3480 ; P2_R1179_U62
g18660 not P2_U3071 ; P2_R1179_U63
g18661 nand P2_R1179_U268 P2_R1179_U267 ; P2_R1179_U64
g18662 not P2_U3084 ; P2_R1179_U65
g18663 not P2_U3485 ; P2_R1179_U66
g18664 not P2_U3083 ; P2_R1179_U67
g18665 not P2_U3957 ; P2_R1179_U68
g18666 not P2_U3078 ; P2_R1179_U69
g18667 not P2_U3954 ; P2_R1179_U70
g18668 not P2_U3955 ; P2_R1179_U71
g18669 not P2_U3956 ; P2_R1179_U72
g18670 not P2_U3068 ; P2_R1179_U73
g18671 not P2_U3063 ; P2_R1179_U74
g18672 not P2_U3077 ; P2_R1179_U75
g18673 nand P2_U3077 P2_R1179_U72 ; P2_R1179_U76
g18674 not P2_U3953 ; P2_R1179_U77
g18675 not P2_U3067 ; P2_R1179_U78
g18676 not P2_U3952 ; P2_R1179_U79
g18677 not P2_U3060 ; P2_R1179_U80
g18678 not P2_U3950 ; P2_R1179_U81
g18679 not P2_U3059 ; P2_R1179_U82
g18680 nand P2_U3059 P2_R1179_U45 ; P2_R1179_U83
g18681 not P2_U3055 ; P2_R1179_U84
g18682 not P2_U3949 ; P2_R1179_U85
g18683 not P2_U3056 ; P2_R1179_U86
g18684 nand P2_R1179_U128 P2_R1179_U301 ; P2_R1179_U87
g18685 nand P2_R1179_U298 P2_R1179_U297 ; P2_R1179_U88
g18686 nand P2_R1179_U76 P2_R1179_U318 ; P2_R1179_U89
g18687 nand P2_R1179_U61 P2_R1179_U329 ; P2_R1179_U90
g18688 nand P2_R1179_U50 P2_R1179_U340 ; P2_R1179_U91
g18689 not P2_U3079 ; P2_R1179_U92
g18690 nand P2_R1179_U395 P2_R1179_U394 ; P2_R1179_U93
g18691 nand P2_R1179_U409 P2_R1179_U408 ; P2_R1179_U94
g18692 nand P2_R1179_U414 P2_R1179_U413 ; P2_R1179_U95
g18693 nand P2_R1179_U430 P2_R1179_U429 ; P2_R1179_U96
g18694 nand P2_R1179_U435 P2_R1179_U434 ; P2_R1179_U97
g18695 nand P2_R1179_U440 P2_R1179_U439 ; P2_R1179_U98
g18696 nand P2_R1179_U445 P2_R1179_U444 ; P2_R1179_U99
g18697 nand P2_R1179_U450 P2_R1179_U449 ; P2_R1179_U100
g18698 nand P2_R1179_U466 P2_R1179_U465 ; P2_R1179_U101
g18699 nand P2_R1179_U471 P2_R1179_U470 ; P2_R1179_U102
g18700 nand P2_R1179_U356 P2_R1179_U355 ; P2_R1179_U103
g18701 nand P2_R1179_U365 P2_R1179_U364 ; P2_R1179_U104
g18702 nand P2_R1179_U372 P2_R1179_U371 ; P2_R1179_U105
g18703 nand P2_R1179_U376 P2_R1179_U375 ; P2_R1179_U106
g18704 nand P2_R1179_U385 P2_R1179_U384 ; P2_R1179_U107
g18705 nand P2_R1179_U404 P2_R1179_U403 ; P2_R1179_U108
g18706 nand P2_R1179_U421 P2_R1179_U420 ; P2_R1179_U109
g18707 nand P2_R1179_U425 P2_R1179_U424 ; P2_R1179_U110
g18708 nand P2_R1179_U457 P2_R1179_U456 ; P2_R1179_U111
g18709 nand P2_R1179_U461 P2_R1179_U460 ; P2_R1179_U112
g18710 nand P2_R1179_U478 P2_R1179_U477 ; P2_R1179_U113
g18711 and P2_R1179_U194 P2_R1179_U184 ; P2_R1179_U114
g18712 and P2_R1179_U197 P2_R1179_U198 ; P2_R1179_U115
g18713 and P2_R1179_U205 P2_R1179_U200 P2_R1179_U185 ; P2_R1179_U116
g18714 and P2_R1179_U210 P2_R1179_U186 ; P2_R1179_U117
g18715 and P2_R1179_U213 P2_R1179_U214 ; P2_R1179_U118
g18716 and P2_R1179_U358 P2_R1179_U357 P2_R1179_U38 ; P2_R1179_U119
g18717 and P2_R1179_U361 P2_R1179_U186 ; P2_R1179_U120
g18718 and P2_R1179_U229 P2_R1179_U6 ; P2_R1179_U121
g18719 and P2_R1179_U368 P2_R1179_U185 ; P2_R1179_U122
g18720 and P2_R1179_U378 P2_R1179_U377 P2_R1179_U28 ; P2_R1179_U123
g18721 and P2_R1179_U381 P2_R1179_U184 ; P2_R1179_U124
g18722 and P2_R1179_U239 P2_R1179_U216 P2_R1179_U180 ; P2_R1179_U125
g18723 and P2_R1179_U261 P2_R1179_U8 ; P2_R1179_U126
g18724 and P2_R1179_U287 P2_R1179_U10 ; P2_R1179_U127
g18725 and P2_R1179_U303 P2_R1179_U304 ; P2_R1179_U128
g18726 and P2_R1179_U387 P2_R1179_U386 P2_R1179_U311 ; P2_R1179_U129
g18727 and P2_R1179_U308 P2_R1179_U390 ; P2_R1179_U130
g18728 nand P2_R1179_U392 P2_R1179_U391 ; P2_R1179_U131
g18729 and P2_R1179_U397 P2_R1179_U396 P2_R1179_U83 ; P2_R1179_U132
g18730 and P2_R1179_U400 P2_R1179_U183 ; P2_R1179_U133
g18731 nand P2_R1179_U406 P2_R1179_U405 ; P2_R1179_U134
g18732 nand P2_R1179_U411 P2_R1179_U410 ; P2_R1179_U135
g18733 and P2_R1179_U324 P2_R1179_U11 ; P2_R1179_U136
g18734 and P2_R1179_U417 P2_R1179_U182 ; P2_R1179_U137
g18735 nand P2_R1179_U427 P2_R1179_U426 ; P2_R1179_U138
g18736 nand P2_R1179_U432 P2_R1179_U431 ; P2_R1179_U139
g18737 nand P2_R1179_U437 P2_R1179_U436 ; P2_R1179_U140
g18738 nand P2_R1179_U442 P2_R1179_U441 ; P2_R1179_U141
g18739 nand P2_R1179_U447 P2_R1179_U446 ; P2_R1179_U142
g18740 and P2_R1179_U335 P2_R1179_U9 ; P2_R1179_U143
g18741 and P2_R1179_U453 P2_R1179_U181 ; P2_R1179_U144
g18742 nand P2_R1179_U463 P2_R1179_U462 ; P2_R1179_U145
g18743 nand P2_R1179_U468 P2_R1179_U467 ; P2_R1179_U146
g18744 and P2_R1179_U346 P2_R1179_U7 ; P2_R1179_U147
g18745 and P2_R1179_U474 P2_R1179_U180 ; P2_R1179_U148
g18746 and P2_R1179_U354 P2_R1179_U353 ; P2_R1179_U149
g18747 nand P2_R1179_U118 P2_R1179_U211 ; P2_R1179_U150
g18748 and P2_R1179_U363 P2_R1179_U362 ; P2_R1179_U151
g18749 and P2_R1179_U370 P2_R1179_U369 ; P2_R1179_U152
g18750 and P2_R1179_U374 P2_R1179_U373 ; P2_R1179_U153
g18751 nand P2_R1179_U115 P2_R1179_U195 ; P2_R1179_U154
g18752 and P2_R1179_U383 P2_R1179_U382 ; P2_R1179_U155
g18753 not P2_U3960 ; P2_R1179_U156
g18754 not P2_U3057 ; P2_R1179_U157
g18755 and P2_R1179_U402 P2_R1179_U401 ; P2_R1179_U158
g18756 nand P2_R1179_U294 P2_R1179_U293 ; P2_R1179_U159
g18757 nand P2_R1179_U290 P2_R1179_U289 ; P2_R1179_U160
g18758 and P2_R1179_U419 P2_R1179_U418 ; P2_R1179_U161
g18759 and P2_R1179_U423 P2_R1179_U422 ; P2_R1179_U162
g18760 nand P2_R1179_U280 P2_R1179_U279 ; P2_R1179_U163
g18761 nand P2_R1179_U276 P2_R1179_U275 ; P2_R1179_U164
g18762 not P2_U3432 ; P2_R1179_U165
g18763 nand P2_U3427 P2_R1179_U92 ; P2_R1179_U166
g18764 nand P2_R1179_U272 P2_R1179_U271 ; P2_R1179_U167
g18765 not P2_U3483 ; P2_R1179_U168
g18766 nand P2_R1179_U264 P2_R1179_U263 ; P2_R1179_U169
g18767 and P2_R1179_U455 P2_R1179_U454 ; P2_R1179_U170
g18768 and P2_R1179_U459 P2_R1179_U458 ; P2_R1179_U171
g18769 nand P2_R1179_U254 P2_R1179_U253 ; P2_R1179_U172
g18770 nand P2_R1179_U250 P2_R1179_U249 ; P2_R1179_U173
g18771 nand P2_R1179_U246 P2_R1179_U245 ; P2_R1179_U174
g18772 and P2_R1179_U476 P2_R1179_U475 ; P2_R1179_U175
g18773 nand P2_R1179_U166 P2_R1179_U165 ; P2_R1179_U176
g18774 not P2_R1179_U83 ; P2_R1179_U177
g18775 not P2_R1179_U28 ; P2_R1179_U178
g18776 not P2_R1179_U38 ; P2_R1179_U179
g18777 nand P2_U3459 P2_R1179_U49 ; P2_R1179_U180
g18778 nand P2_U3474 P2_R1179_U59 ; P2_R1179_U181
g18779 nand P2_U3955 P2_R1179_U74 ; P2_R1179_U182
g18780 nand P2_U3951 P2_R1179_U82 ; P2_R1179_U183
g18781 nand P2_U3435 P2_R1179_U27 ; P2_R1179_U184
g18782 nand P2_U3444 P2_R1179_U33 ; P2_R1179_U185
g18783 nand P2_U3450 P2_R1179_U37 ; P2_R1179_U186
g18784 not P2_R1179_U61 ; P2_R1179_U187
g18785 not P2_R1179_U76 ; P2_R1179_U188
g18786 not P2_R1179_U35 ; P2_R1179_U189
g18787 not P2_R1179_U50 ; P2_R1179_U190
g18788 not P2_R1179_U166 ; P2_R1179_U191
g18789 nand P2_U3080 P2_R1179_U166 ; P2_R1179_U192
g18790 not P2_R1179_U44 ; P2_R1179_U193
g18791 nand P2_U3438 P2_R1179_U29 ; P2_R1179_U194
g18792 nand P2_R1179_U114 P2_R1179_U44 ; P2_R1179_U195
g18793 nand P2_R1179_U29 P2_R1179_U28 ; P2_R1179_U196
g18794 nand P2_R1179_U196 P2_R1179_U26 ; P2_R1179_U197
g18795 nand P2_U3066 P2_R1179_U178 ; P2_R1179_U198
g18796 not P2_R1179_U154 ; P2_R1179_U199
g18797 nand P2_U3447 P2_R1179_U32 ; P2_R1179_U200
g18798 nand P2_U3073 P2_R1179_U30 ; P2_R1179_U201
g18799 nand P2_U3069 P2_R1179_U22 ; P2_R1179_U202
g18800 nand P2_R1179_U189 P2_R1179_U185 ; P2_R1179_U203
g18801 nand P2_R1179_U6 P2_R1179_U203 ; P2_R1179_U204
g18802 nand P2_U3441 P2_R1179_U34 ; P2_R1179_U205
g18803 nand P2_U3447 P2_R1179_U32 ; P2_R1179_U206
g18804 nand P2_R1179_U154 P2_R1179_U116 ; P2_R1179_U207
g18805 nand P2_R1179_U206 P2_R1179_U204 ; P2_R1179_U208
g18806 not P2_R1179_U42 ; P2_R1179_U209
g18807 nand P2_U3453 P2_R1179_U39 ; P2_R1179_U210
g18808 nand P2_R1179_U117 P2_R1179_U42 ; P2_R1179_U211
g18809 nand P2_R1179_U39 P2_R1179_U38 ; P2_R1179_U212
g18810 nand P2_R1179_U212 P2_R1179_U36 ; P2_R1179_U213
g18811 nand P2_U3086 P2_R1179_U179 ; P2_R1179_U214
g18812 not P2_R1179_U150 ; P2_R1179_U215
g18813 nand P2_U3456 P2_R1179_U41 ; P2_R1179_U216
g18814 nand P2_R1179_U216 P2_R1179_U50 ; P2_R1179_U217
g18815 nand P2_R1179_U209 P2_R1179_U38 ; P2_R1179_U218
g18816 nand P2_R1179_U120 P2_R1179_U218 ; P2_R1179_U219
g18817 nand P2_R1179_U42 P2_R1179_U186 ; P2_R1179_U220
g18818 nand P2_R1179_U119 P2_R1179_U220 ; P2_R1179_U221
g18819 nand P2_R1179_U38 P2_R1179_U186 ; P2_R1179_U222
g18820 nand P2_R1179_U205 P2_R1179_U154 ; P2_R1179_U223
g18821 not P2_R1179_U43 ; P2_R1179_U224
g18822 nand P2_U3069 P2_R1179_U22 ; P2_R1179_U225
g18823 nand P2_R1179_U224 P2_R1179_U225 ; P2_R1179_U226
g18824 nand P2_R1179_U122 P2_R1179_U226 ; P2_R1179_U227
g18825 nand P2_R1179_U43 P2_R1179_U185 ; P2_R1179_U228
g18826 nand P2_U3447 P2_R1179_U32 ; P2_R1179_U229
g18827 nand P2_R1179_U121 P2_R1179_U228 ; P2_R1179_U230
g18828 nand P2_U3069 P2_R1179_U22 ; P2_R1179_U231
g18829 nand P2_R1179_U185 P2_R1179_U231 ; P2_R1179_U232
g18830 nand P2_R1179_U205 P2_R1179_U35 ; P2_R1179_U233
g18831 nand P2_R1179_U193 P2_R1179_U28 ; P2_R1179_U234
g18832 nand P2_R1179_U124 P2_R1179_U234 ; P2_R1179_U235
g18833 nand P2_R1179_U44 P2_R1179_U184 ; P2_R1179_U236
g18834 nand P2_R1179_U123 P2_R1179_U236 ; P2_R1179_U237
g18835 nand P2_R1179_U28 P2_R1179_U184 ; P2_R1179_U238
g18836 nand P2_U3462 P2_R1179_U48 ; P2_R1179_U239
g18837 nand P2_U3065 P2_R1179_U47 ; P2_R1179_U240
g18838 nand P2_U3064 P2_R1179_U46 ; P2_R1179_U241
g18839 nand P2_R1179_U190 P2_R1179_U180 ; P2_R1179_U242
g18840 nand P2_R1179_U7 P2_R1179_U242 ; P2_R1179_U243
g18841 nand P2_U3462 P2_R1179_U48 ; P2_R1179_U244
g18842 nand P2_R1179_U150 P2_R1179_U125 ; P2_R1179_U245
g18843 nand P2_R1179_U244 P2_R1179_U243 ; P2_R1179_U246
g18844 not P2_R1179_U174 ; P2_R1179_U247
g18845 nand P2_U3465 P2_R1179_U52 ; P2_R1179_U248
g18846 nand P2_R1179_U248 P2_R1179_U174 ; P2_R1179_U249
g18847 nand P2_U3074 P2_R1179_U51 ; P2_R1179_U250
g18848 not P2_R1179_U173 ; P2_R1179_U251
g18849 nand P2_U3468 P2_R1179_U54 ; P2_R1179_U252
g18850 nand P2_R1179_U252 P2_R1179_U173 ; P2_R1179_U253
g18851 nand P2_U3082 P2_R1179_U53 ; P2_R1179_U254
g18852 not P2_R1179_U172 ; P2_R1179_U255
g18853 nand P2_U3477 P2_R1179_U58 ; P2_R1179_U256
g18854 nand P2_U3075 P2_R1179_U55 ; P2_R1179_U257
g18855 nand P2_U3076 P2_R1179_U56 ; P2_R1179_U258
g18856 nand P2_R1179_U187 P2_R1179_U8 ; P2_R1179_U259
g18857 nand P2_R1179_U9 P2_R1179_U259 ; P2_R1179_U260
g18858 nand P2_U3471 P2_R1179_U60 ; P2_R1179_U261
g18859 nand P2_U3477 P2_R1179_U58 ; P2_R1179_U262
g18860 nand P2_R1179_U126 P2_R1179_U172 ; P2_R1179_U263
g18861 nand P2_R1179_U262 P2_R1179_U260 ; P2_R1179_U264
g18862 not P2_R1179_U169 ; P2_R1179_U265
g18863 nand P2_U3480 P2_R1179_U63 ; P2_R1179_U266
g18864 nand P2_R1179_U266 P2_R1179_U169 ; P2_R1179_U267
g18865 nand P2_U3071 P2_R1179_U62 ; P2_R1179_U268
g18866 not P2_R1179_U64 ; P2_R1179_U269
g18867 nand P2_R1179_U269 P2_R1179_U65 ; P2_R1179_U270
g18868 nand P2_R1179_U270 P2_R1179_U168 ; P2_R1179_U271
g18869 nand P2_U3084 P2_R1179_U64 ; P2_R1179_U272
g18870 not P2_R1179_U167 ; P2_R1179_U273
g18871 nand P2_U3485 P2_R1179_U67 ; P2_R1179_U274
g18872 nand P2_R1179_U274 P2_R1179_U167 ; P2_R1179_U275
g18873 nand P2_U3083 P2_R1179_U66 ; P2_R1179_U276
g18874 not P2_R1179_U164 ; P2_R1179_U277
g18875 nand P2_U3957 P2_R1179_U69 ; P2_R1179_U278
g18876 nand P2_R1179_U278 P2_R1179_U164 ; P2_R1179_U279
g18877 nand P2_U3078 P2_R1179_U68 ; P2_R1179_U280
g18878 not P2_R1179_U163 ; P2_R1179_U281
g18879 nand P2_U3954 P2_R1179_U73 ; P2_R1179_U282
g18880 nand P2_U3068 P2_R1179_U70 ; P2_R1179_U283
g18881 nand P2_U3063 P2_R1179_U71 ; P2_R1179_U284
g18882 nand P2_R1179_U188 P2_R1179_U10 ; P2_R1179_U285
g18883 nand P2_R1179_U11 P2_R1179_U285 ; P2_R1179_U286
g18884 nand P2_U3956 P2_R1179_U75 ; P2_R1179_U287
g18885 nand P2_U3954 P2_R1179_U73 ; P2_R1179_U288
g18886 nand P2_R1179_U127 P2_R1179_U163 ; P2_R1179_U289
g18887 nand P2_R1179_U288 P2_R1179_U286 ; P2_R1179_U290
g18888 not P2_R1179_U160 ; P2_R1179_U291
g18889 nand P2_U3953 P2_R1179_U78 ; P2_R1179_U292
g18890 nand P2_R1179_U292 P2_R1179_U160 ; P2_R1179_U293
g18891 nand P2_U3067 P2_R1179_U77 ; P2_R1179_U294
g18892 not P2_R1179_U159 ; P2_R1179_U295
g18893 nand P2_U3952 P2_R1179_U80 ; P2_R1179_U296
g18894 nand P2_R1179_U296 P2_R1179_U159 ; P2_R1179_U297
g18895 nand P2_U3060 P2_R1179_U79 ; P2_R1179_U298
g18896 not P2_R1179_U88 ; P2_R1179_U299
g18897 nand P2_U3950 P2_R1179_U84 ; P2_R1179_U300
g18898 nand P2_R1179_U88 P2_R1179_U183 P2_R1179_U300 ; P2_R1179_U301
g18899 nand P2_R1179_U84 P2_R1179_U83 ; P2_R1179_U302
g18900 nand P2_R1179_U302 P2_R1179_U81 ; P2_R1179_U303
g18901 nand P2_U3055 P2_R1179_U177 ; P2_R1179_U304
g18902 not P2_R1179_U87 ; P2_R1179_U305
g18903 nand P2_U3056 P2_R1179_U85 ; P2_R1179_U306
g18904 nand P2_R1179_U305 P2_R1179_U306 ; P2_R1179_U307
g18905 nand P2_U3949 P2_R1179_U86 ; P2_R1179_U308
g18906 nand P2_U3949 P2_R1179_U86 ; P2_R1179_U309
g18907 nand P2_R1179_U309 P2_R1179_U87 ; P2_R1179_U310
g18908 nand P2_U3056 P2_R1179_U85 ; P2_R1179_U311
g18909 nand P2_R1179_U129 P2_R1179_U310 ; P2_R1179_U312
g18910 nand P2_R1179_U299 P2_R1179_U83 ; P2_R1179_U313
g18911 nand P2_R1179_U133 P2_R1179_U313 ; P2_R1179_U314
g18912 nand P2_R1179_U88 P2_R1179_U183 ; P2_R1179_U315
g18913 nand P2_R1179_U132 P2_R1179_U315 ; P2_R1179_U316
g18914 nand P2_R1179_U83 P2_R1179_U183 ; P2_R1179_U317
g18915 nand P2_R1179_U287 P2_R1179_U163 ; P2_R1179_U318
g18916 not P2_R1179_U89 ; P2_R1179_U319
g18917 nand P2_U3063 P2_R1179_U71 ; P2_R1179_U320
g18918 nand P2_R1179_U319 P2_R1179_U320 ; P2_R1179_U321
g18919 nand P2_R1179_U137 P2_R1179_U321 ; P2_R1179_U322
g18920 nand P2_R1179_U89 P2_R1179_U182 ; P2_R1179_U323
g18921 nand P2_U3954 P2_R1179_U73 ; P2_R1179_U324
g18922 nand P2_R1179_U136 P2_R1179_U323 ; P2_R1179_U325
g18923 nand P2_U3063 P2_R1179_U71 ; P2_R1179_U326
g18924 nand P2_R1179_U182 P2_R1179_U326 ; P2_R1179_U327
g18925 nand P2_R1179_U287 P2_R1179_U76 ; P2_R1179_U328
g18926 nand P2_R1179_U261 P2_R1179_U172 ; P2_R1179_U329
g18927 not P2_R1179_U90 ; P2_R1179_U330
g18928 nand P2_U3076 P2_R1179_U56 ; P2_R1179_U331
g18929 nand P2_R1179_U330 P2_R1179_U331 ; P2_R1179_U332
g18930 nand P2_R1179_U144 P2_R1179_U332 ; P2_R1179_U333
g18931 nand P2_R1179_U90 P2_R1179_U181 ; P2_R1179_U334
g18932 nand P2_U3477 P2_R1179_U58 ; P2_R1179_U335
g18933 nand P2_R1179_U143 P2_R1179_U334 ; P2_R1179_U336
g18934 nand P2_U3076 P2_R1179_U56 ; P2_R1179_U337
g18935 nand P2_R1179_U181 P2_R1179_U337 ; P2_R1179_U338
g18936 nand P2_R1179_U261 P2_R1179_U61 ; P2_R1179_U339
g18937 nand P2_R1179_U216 P2_R1179_U150 ; P2_R1179_U340
g18938 not P2_R1179_U91 ; P2_R1179_U341
g18939 nand P2_U3064 P2_R1179_U46 ; P2_R1179_U342
g18940 nand P2_R1179_U341 P2_R1179_U342 ; P2_R1179_U343
g18941 nand P2_R1179_U148 P2_R1179_U343 ; P2_R1179_U344
g18942 nand P2_R1179_U91 P2_R1179_U180 ; P2_R1179_U345
g18943 nand P2_U3462 P2_R1179_U48 ; P2_R1179_U346
g18944 nand P2_R1179_U147 P2_R1179_U345 ; P2_R1179_U347
g18945 nand P2_U3064 P2_R1179_U46 ; P2_R1179_U348
g18946 nand P2_R1179_U180 P2_R1179_U348 ; P2_R1179_U349
g18947 nand P2_U3079 P2_R1179_U24 ; P2_R1179_U350
g18948 nand P2_U3080 P2_R1179_U165 ; P2_R1179_U351
g18949 nand P2_R1179_U130 P2_R1179_U307 ; P2_R1179_U352
g18950 nand P2_U3456 P2_R1179_U41 ; P2_R1179_U353
g18951 nand P2_U3085 P2_R1179_U40 ; P2_R1179_U354
g18952 nand P2_R1179_U217 P2_R1179_U150 ; P2_R1179_U355
g18953 nand P2_R1179_U215 P2_R1179_U149 ; P2_R1179_U356
g18954 nand P2_U3453 P2_R1179_U39 ; P2_R1179_U357
g18955 nand P2_U3086 P2_R1179_U36 ; P2_R1179_U358
g18956 nand P2_U3453 P2_R1179_U39 ; P2_R1179_U359
g18957 nand P2_U3086 P2_R1179_U36 ; P2_R1179_U360
g18958 nand P2_R1179_U360 P2_R1179_U359 ; P2_R1179_U361
g18959 nand P2_U3450 P2_R1179_U37 ; P2_R1179_U362
g18960 nand P2_U3072 P2_R1179_U21 ; P2_R1179_U363
g18961 nand P2_R1179_U222 P2_R1179_U42 ; P2_R1179_U364
g18962 nand P2_R1179_U151 P2_R1179_U209 ; P2_R1179_U365
g18963 nand P2_U3447 P2_R1179_U32 ; P2_R1179_U366
g18964 nand P2_U3073 P2_R1179_U30 ; P2_R1179_U367
g18965 nand P2_R1179_U367 P2_R1179_U366 ; P2_R1179_U368
g18966 nand P2_U3444 P2_R1179_U33 ; P2_R1179_U369
g18967 nand P2_U3069 P2_R1179_U22 ; P2_R1179_U370
g18968 nand P2_R1179_U232 P2_R1179_U43 ; P2_R1179_U371
g18969 nand P2_R1179_U152 P2_R1179_U224 ; P2_R1179_U372
g18970 nand P2_U3441 P2_R1179_U34 ; P2_R1179_U373
g18971 nand P2_U3062 P2_R1179_U31 ; P2_R1179_U374
g18972 nand P2_R1179_U233 P2_R1179_U154 ; P2_R1179_U375
g18973 nand P2_R1179_U199 P2_R1179_U153 ; P2_R1179_U376
g18974 nand P2_U3438 P2_R1179_U29 ; P2_R1179_U377
g18975 nand P2_U3066 P2_R1179_U26 ; P2_R1179_U378
g18976 nand P2_U3438 P2_R1179_U29 ; P2_R1179_U379
g18977 nand P2_U3066 P2_R1179_U26 ; P2_R1179_U380
g18978 nand P2_R1179_U380 P2_R1179_U379 ; P2_R1179_U381
g18979 nand P2_U3435 P2_R1179_U27 ; P2_R1179_U382
g18980 nand P2_U3070 P2_R1179_U23 ; P2_R1179_U383
g18981 nand P2_R1179_U238 P2_R1179_U44 ; P2_R1179_U384
g18982 nand P2_R1179_U155 P2_R1179_U193 ; P2_R1179_U385
g18983 nand P2_U3960 P2_R1179_U157 ; P2_R1179_U386
g18984 nand P2_U3057 P2_R1179_U156 ; P2_R1179_U387
g18985 nand P2_U3960 P2_R1179_U157 ; P2_R1179_U388
g18986 nand P2_U3057 P2_R1179_U156 ; P2_R1179_U389
g18987 nand P2_R1179_U389 P2_R1179_U388 ; P2_R1179_U390
g18988 nand P2_U3949 P2_R1179_U86 ; P2_R1179_U391
g18989 nand P2_U3056 P2_R1179_U85 ; P2_R1179_U392
g18990 not P2_R1179_U131 ; P2_R1179_U393
g18991 nand P2_R1179_U393 P2_R1179_U305 ; P2_R1179_U394
g18992 nand P2_R1179_U131 P2_R1179_U87 ; P2_R1179_U395
g18993 nand P2_U3950 P2_R1179_U84 ; P2_R1179_U396
g18994 nand P2_U3055 P2_R1179_U81 ; P2_R1179_U397
g18995 nand P2_U3950 P2_R1179_U84 ; P2_R1179_U398
g18996 nand P2_U3055 P2_R1179_U81 ; P2_R1179_U399
g18997 nand P2_R1179_U399 P2_R1179_U398 ; P2_R1179_U400
g18998 nand P2_U3951 P2_R1179_U82 ; P2_R1179_U401
g18999 nand P2_U3059 P2_R1179_U45 ; P2_R1179_U402
g19000 nand P2_R1179_U317 P2_R1179_U88 ; P2_R1179_U403
g19001 nand P2_R1179_U158 P2_R1179_U299 ; P2_R1179_U404
g19002 nand P2_U3952 P2_R1179_U80 ; P2_R1179_U405
g19003 nand P2_U3060 P2_R1179_U79 ; P2_R1179_U406
g19004 not P2_R1179_U134 ; P2_R1179_U407
g19005 nand P2_R1179_U295 P2_R1179_U407 ; P2_R1179_U408
g19006 nand P2_R1179_U134 P2_R1179_U159 ; P2_R1179_U409
g19007 nand P2_U3953 P2_R1179_U78 ; P2_R1179_U410
g19008 nand P2_U3067 P2_R1179_U77 ; P2_R1179_U411
g19009 not P2_R1179_U135 ; P2_R1179_U412
g19010 nand P2_R1179_U291 P2_R1179_U412 ; P2_R1179_U413
g19011 nand P2_R1179_U135 P2_R1179_U160 ; P2_R1179_U414
g19012 nand P2_U3954 P2_R1179_U73 ; P2_R1179_U415
g19013 nand P2_U3068 P2_R1179_U70 ; P2_R1179_U416
g19014 nand P2_R1179_U416 P2_R1179_U415 ; P2_R1179_U417
g19015 nand P2_U3955 P2_R1179_U74 ; P2_R1179_U418
g19016 nand P2_U3063 P2_R1179_U71 ; P2_R1179_U419
g19017 nand P2_R1179_U327 P2_R1179_U89 ; P2_R1179_U420
g19018 nand P2_R1179_U161 P2_R1179_U319 ; P2_R1179_U421
g19019 nand P2_U3956 P2_R1179_U75 ; P2_R1179_U422
g19020 nand P2_U3077 P2_R1179_U72 ; P2_R1179_U423
g19021 nand P2_R1179_U328 P2_R1179_U163 ; P2_R1179_U424
g19022 nand P2_R1179_U281 P2_R1179_U162 ; P2_R1179_U425
g19023 nand P2_U3957 P2_R1179_U69 ; P2_R1179_U426
g19024 nand P2_U3078 P2_R1179_U68 ; P2_R1179_U427
g19025 not P2_R1179_U138 ; P2_R1179_U428
g19026 nand P2_R1179_U277 P2_R1179_U428 ; P2_R1179_U429
g19027 nand P2_R1179_U138 P2_R1179_U164 ; P2_R1179_U430
g19028 nand P2_U3432 P2_R1179_U25 ; P2_R1179_U431
g19029 nand P2_U3080 P2_R1179_U165 ; P2_R1179_U432
g19030 not P2_R1179_U139 ; P2_R1179_U433
g19031 nand P2_R1179_U191 P2_R1179_U433 ; P2_R1179_U434
g19032 nand P2_R1179_U139 P2_R1179_U166 ; P2_R1179_U435
g19033 nand P2_U3485 P2_R1179_U67 ; P2_R1179_U436
g19034 nand P2_U3083 P2_R1179_U66 ; P2_R1179_U437
g19035 not P2_R1179_U140 ; P2_R1179_U438
g19036 nand P2_R1179_U273 P2_R1179_U438 ; P2_R1179_U439
g19037 nand P2_R1179_U140 P2_R1179_U167 ; P2_R1179_U440
g19038 nand P2_U3483 P2_R1179_U65 ; P2_R1179_U441
g19039 nand P2_U3084 P2_R1179_U168 ; P2_R1179_U442
g19040 not P2_R1179_U141 ; P2_R1179_U443
g19041 nand P2_R1179_U443 P2_R1179_U269 ; P2_R1179_U444
g19042 nand P2_R1179_U141 P2_R1179_U64 ; P2_R1179_U445
g19043 nand P2_U3480 P2_R1179_U63 ; P2_R1179_U446
g19044 nand P2_U3071 P2_R1179_U62 ; P2_R1179_U447
g19045 not P2_R1179_U142 ; P2_R1179_U448
g19046 nand P2_R1179_U265 P2_R1179_U448 ; P2_R1179_U449
g19047 nand P2_R1179_U142 P2_R1179_U169 ; P2_R1179_U450
g19048 nand P2_U3477 P2_R1179_U58 ; P2_R1179_U451
g19049 nand P2_U3075 P2_R1179_U55 ; P2_R1179_U452
g19050 nand P2_R1179_U452 P2_R1179_U451 ; P2_R1179_U453
g19051 nand P2_U3474 P2_R1179_U59 ; P2_R1179_U454
g19052 nand P2_U3076 P2_R1179_U56 ; P2_R1179_U455
g19053 nand P2_R1179_U338 P2_R1179_U90 ; P2_R1179_U456
g19054 nand P2_R1179_U170 P2_R1179_U330 ; P2_R1179_U457
g19055 nand P2_U3471 P2_R1179_U60 ; P2_R1179_U458
g19056 nand P2_U3081 P2_R1179_U57 ; P2_R1179_U459
g19057 nand P2_R1179_U339 P2_R1179_U172 ; P2_R1179_U460
g19058 nand P2_R1179_U255 P2_R1179_U171 ; P2_R1179_U461
g19059 nand P2_U3468 P2_R1179_U54 ; P2_R1179_U462
g19060 nand P2_U3082 P2_R1179_U53 ; P2_R1179_U463
g19061 not P2_R1179_U145 ; P2_R1179_U464
g19062 nand P2_R1179_U251 P2_R1179_U464 ; P2_R1179_U465
g19063 nand P2_R1179_U145 P2_R1179_U173 ; P2_R1179_U466
g19064 nand P2_U3465 P2_R1179_U52 ; P2_R1179_U467
g19065 nand P2_U3074 P2_R1179_U51 ; P2_R1179_U468
g19066 not P2_R1179_U146 ; P2_R1179_U469
g19067 nand P2_R1179_U247 P2_R1179_U469 ; P2_R1179_U470
g19068 nand P2_R1179_U146 P2_R1179_U174 ; P2_R1179_U471
g19069 nand P2_U3462 P2_R1179_U48 ; P2_R1179_U472
g19070 nand P2_U3065 P2_R1179_U47 ; P2_R1179_U473
g19071 nand P2_R1179_U473 P2_R1179_U472 ; P2_R1179_U474
g19072 nand P2_U3459 P2_R1179_U49 ; P2_R1179_U475
g19073 nand P2_U3064 P2_R1179_U46 ; P2_R1179_U476
g19074 nand P2_R1179_U349 P2_R1179_U91 ; P2_R1179_U477
g19075 nand P2_R1179_U175 P2_R1179_U341 ; P2_R1179_U478
g19076 and P2_R1215_U179 P2_R1215_U178 ; P2_R1215_U4
g19077 and P2_R1215_U180 P2_R1215_U181 ; P2_R1215_U5
g19078 and P2_R1215_U197 P2_R1215_U196 ; P2_R1215_U6
g19079 and P2_R1215_U237 P2_R1215_U236 ; P2_R1215_U7
g19080 and P2_R1215_U246 P2_R1215_U245 ; P2_R1215_U8
g19081 and P2_R1215_U264 P2_R1215_U263 ; P2_R1215_U9
g19082 and P2_R1215_U272 P2_R1215_U271 ; P2_R1215_U10
g19083 and P2_R1215_U351 P2_R1215_U348 ; P2_R1215_U11
g19084 and P2_R1215_U344 P2_R1215_U341 ; P2_R1215_U12
g19085 and P2_R1215_U335 P2_R1215_U332 ; P2_R1215_U13
g19086 and P2_R1215_U326 P2_R1215_U323 ; P2_R1215_U14
g19087 and P2_R1215_U320 P2_R1215_U318 ; P2_R1215_U15
g19088 and P2_R1215_U313 P2_R1215_U310 ; P2_R1215_U16
g19089 and P2_R1215_U235 P2_R1215_U232 ; P2_R1215_U17
g19090 and P2_R1215_U227 P2_R1215_U224 ; P2_R1215_U18
g19091 and P2_R1215_U213 P2_R1215_U210 ; P2_R1215_U19
g19092 not P2_U3447 ; P2_R1215_U20
g19093 not P2_U3073 ; P2_R1215_U21
g19094 not P2_U3072 ; P2_R1215_U22
g19095 nand P2_U3073 P2_U3447 ; P2_R1215_U23
g19096 not P2_U3450 ; P2_R1215_U24
g19097 not P2_U3441 ; P2_R1215_U25
g19098 not P2_U3062 ; P2_R1215_U26
g19099 not P2_U3069 ; P2_R1215_U27
g19100 not P2_U3435 ; P2_R1215_U28
g19101 not P2_U3070 ; P2_R1215_U29
g19102 not P2_U3427 ; P2_R1215_U30
g19103 not P2_U3079 ; P2_R1215_U31
g19104 nand P2_U3079 P2_U3427 ; P2_R1215_U32
g19105 not P2_U3438 ; P2_R1215_U33
g19106 not P2_U3066 ; P2_R1215_U34
g19107 nand P2_U3062 P2_U3441 ; P2_R1215_U35
g19108 not P2_U3444 ; P2_R1215_U36
g19109 not P2_U3453 ; P2_R1215_U37
g19110 not P2_U3086 ; P2_R1215_U38
g19111 not P2_U3085 ; P2_R1215_U39
g19112 not P2_U3456 ; P2_R1215_U40
g19113 nand P2_R1215_U62 P2_R1215_U205 ; P2_R1215_U41
g19114 nand P2_R1215_U118 P2_R1215_U193 ; P2_R1215_U42
g19115 nand P2_R1215_U182 P2_R1215_U183 ; P2_R1215_U43
g19116 nand P2_U3432 P2_U3080 ; P2_R1215_U44
g19117 nand P2_R1215_U122 P2_R1215_U219 ; P2_R1215_U45
g19118 nand P2_R1215_U216 P2_R1215_U215 ; P2_R1215_U46
g19119 not P2_U3950 ; P2_R1215_U47
g19120 not P2_U3055 ; P2_R1215_U48
g19121 not P2_U3059 ; P2_R1215_U49
g19122 not P2_U3951 ; P2_R1215_U50
g19123 not P2_U3952 ; P2_R1215_U51
g19124 not P2_U3060 ; P2_R1215_U52
g19125 not P2_U3953 ; P2_R1215_U53
g19126 not P2_U3067 ; P2_R1215_U54
g19127 not P2_U3956 ; P2_R1215_U55
g19128 not P2_U3077 ; P2_R1215_U56
g19129 not P2_U3477 ; P2_R1215_U57
g19130 not P2_U3075 ; P2_R1215_U58
g19131 not P2_U3071 ; P2_R1215_U59
g19132 nand P2_U3075 P2_U3477 ; P2_R1215_U60
g19133 not P2_U3480 ; P2_R1215_U61
g19134 nand P2_U3086 P2_U3453 ; P2_R1215_U62
g19135 not P2_U3459 ; P2_R1215_U63
g19136 not P2_U3064 ; P2_R1215_U64
g19137 not P2_U3465 ; P2_R1215_U65
g19138 not P2_U3074 ; P2_R1215_U66
g19139 not P2_U3462 ; P2_R1215_U67
g19140 not P2_U3065 ; P2_R1215_U68
g19141 nand P2_U3065 P2_U3462 ; P2_R1215_U69
g19142 not P2_U3468 ; P2_R1215_U70
g19143 not P2_U3082 ; P2_R1215_U71
g19144 not P2_U3471 ; P2_R1215_U72
g19145 not P2_U3081 ; P2_R1215_U73
g19146 not P2_U3474 ; P2_R1215_U74
g19147 not P2_U3076 ; P2_R1215_U75
g19148 not P2_U3483 ; P2_R1215_U76
g19149 not P2_U3084 ; P2_R1215_U77
g19150 nand P2_U3084 P2_U3483 ; P2_R1215_U78
g19151 not P2_U3485 ; P2_R1215_U79
g19152 not P2_U3083 ; P2_R1215_U80
g19153 nand P2_U3083 P2_U3485 ; P2_R1215_U81
g19154 not P2_U3957 ; P2_R1215_U82
g19155 not P2_U3955 ; P2_R1215_U83
g19156 not P2_U3063 ; P2_R1215_U84
g19157 not P2_U3954 ; P2_R1215_U85
g19158 not P2_U3068 ; P2_R1215_U86
g19159 nand P2_U3951 P2_U3059 ; P2_R1215_U87
g19160 not P2_U3056 ; P2_R1215_U88
g19161 not P2_U3949 ; P2_R1215_U89
g19162 nand P2_R1215_U306 P2_R1215_U176 ; P2_R1215_U90
g19163 not P2_U3078 ; P2_R1215_U91
g19164 nand P2_R1215_U78 P2_R1215_U315 ; P2_R1215_U92
g19165 nand P2_R1215_U261 P2_R1215_U260 ; P2_R1215_U93
g19166 nand P2_R1215_U69 P2_R1215_U337 ; P2_R1215_U94
g19167 nand P2_R1215_U457 P2_R1215_U456 ; P2_R1215_U95
g19168 nand P2_R1215_U504 P2_R1215_U503 ; P2_R1215_U96
g19169 nand P2_R1215_U375 P2_R1215_U374 ; P2_R1215_U97
g19170 nand P2_R1215_U380 P2_R1215_U379 ; P2_R1215_U98
g19171 nand P2_R1215_U387 P2_R1215_U386 ; P2_R1215_U99
g19172 nand P2_R1215_U394 P2_R1215_U393 ; P2_R1215_U100
g19173 nand P2_R1215_U399 P2_R1215_U398 ; P2_R1215_U101
g19174 nand P2_R1215_U408 P2_R1215_U407 ; P2_R1215_U102
g19175 nand P2_R1215_U415 P2_R1215_U414 ; P2_R1215_U103
g19176 nand P2_R1215_U422 P2_R1215_U421 ; P2_R1215_U104
g19177 nand P2_R1215_U429 P2_R1215_U428 ; P2_R1215_U105
g19178 nand P2_R1215_U434 P2_R1215_U433 ; P2_R1215_U106
g19179 nand P2_R1215_U441 P2_R1215_U440 ; P2_R1215_U107
g19180 nand P2_R1215_U448 P2_R1215_U447 ; P2_R1215_U108
g19181 nand P2_R1215_U462 P2_R1215_U461 ; P2_R1215_U109
g19182 nand P2_R1215_U467 P2_R1215_U466 ; P2_R1215_U110
g19183 nand P2_R1215_U474 P2_R1215_U473 ; P2_R1215_U111
g19184 nand P2_R1215_U481 P2_R1215_U480 ; P2_R1215_U112
g19185 nand P2_R1215_U488 P2_R1215_U487 ; P2_R1215_U113
g19186 nand P2_R1215_U495 P2_R1215_U494 ; P2_R1215_U114
g19187 nand P2_R1215_U500 P2_R1215_U499 ; P2_R1215_U115
g19188 and P2_U3435 P2_U3070 ; P2_R1215_U116
g19189 and P2_R1215_U189 P2_R1215_U187 ; P2_R1215_U117
g19190 and P2_R1215_U194 P2_R1215_U192 ; P2_R1215_U118
g19191 and P2_R1215_U201 P2_R1215_U200 ; P2_R1215_U119
g19192 and P2_R1215_U382 P2_R1215_U381 P2_R1215_U23 ; P2_R1215_U120
g19193 and P2_R1215_U212 P2_R1215_U6 ; P2_R1215_U121
g19194 and P2_R1215_U220 P2_R1215_U218 ; P2_R1215_U122
g19195 and P2_R1215_U389 P2_R1215_U388 P2_R1215_U35 ; P2_R1215_U123
g19196 and P2_R1215_U226 P2_R1215_U4 ; P2_R1215_U124
g19197 and P2_R1215_U234 P2_R1215_U181 ; P2_R1215_U125
g19198 and P2_R1215_U204 P2_R1215_U7 ; P2_R1215_U126
g19199 and P2_R1215_U239 P2_R1215_U171 ; P2_R1215_U127
g19200 and P2_R1215_U250 P2_R1215_U8 ; P2_R1215_U128
g19201 and P2_R1215_U248 P2_R1215_U172 ; P2_R1215_U129
g19202 and P2_R1215_U268 P2_R1215_U267 ; P2_R1215_U130
g19203 and P2_R1215_U10 P2_R1215_U282 ; P2_R1215_U131
g19204 and P2_R1215_U285 P2_R1215_U280 ; P2_R1215_U132
g19205 and P2_R1215_U301 P2_R1215_U298 ; P2_R1215_U133
g19206 and P2_R1215_U368 P2_R1215_U302 ; P2_R1215_U134
g19207 and P2_R1215_U160 P2_R1215_U278 ; P2_R1215_U135
g19208 and P2_R1215_U455 P2_R1215_U454 P2_R1215_U81 ; P2_R1215_U136
g19209 and P2_R1215_U325 P2_R1215_U10 ; P2_R1215_U137
g19210 and P2_R1215_U469 P2_R1215_U468 P2_R1215_U60 ; P2_R1215_U138
g19211 and P2_R1215_U334 P2_R1215_U9 ; P2_R1215_U139
g19212 and P2_R1215_U490 P2_R1215_U489 P2_R1215_U172 ; P2_R1215_U140
g19213 and P2_R1215_U343 P2_R1215_U8 ; P2_R1215_U141
g19214 and P2_R1215_U502 P2_R1215_U501 P2_R1215_U171 ; P2_R1215_U142
g19215 and P2_R1215_U350 P2_R1215_U7 ; P2_R1215_U143
g19216 nand P2_R1215_U119 P2_R1215_U202 ; P2_R1215_U144
g19217 nand P2_R1215_U217 P2_R1215_U229 ; P2_R1215_U145
g19218 not P2_U3057 ; P2_R1215_U146
g19219 not P2_U3960 ; P2_R1215_U147
g19220 and P2_R1215_U403 P2_R1215_U402 ; P2_R1215_U148
g19221 nand P2_R1215_U304 P2_R1215_U169 P2_R1215_U364 ; P2_R1215_U149
g19222 and P2_R1215_U410 P2_R1215_U409 ; P2_R1215_U150
g19223 nand P2_R1215_U370 P2_R1215_U369 P2_R1215_U134 ; P2_R1215_U151
g19224 and P2_R1215_U417 P2_R1215_U416 ; P2_R1215_U152
g19225 nand P2_R1215_U365 P2_R1215_U299 P2_R1215_U87 ; P2_R1215_U153
g19226 and P2_R1215_U424 P2_R1215_U423 ; P2_R1215_U154
g19227 nand P2_R1215_U293 P2_R1215_U292 ; P2_R1215_U155
g19228 and P2_R1215_U436 P2_R1215_U435 ; P2_R1215_U156
g19229 nand P2_R1215_U289 P2_R1215_U288 ; P2_R1215_U157
g19230 and P2_R1215_U443 P2_R1215_U442 ; P2_R1215_U158
g19231 nand P2_R1215_U132 P2_R1215_U284 ; P2_R1215_U159
g19232 and P2_R1215_U450 P2_R1215_U449 ; P2_R1215_U160
g19233 nand P2_R1215_U44 P2_R1215_U327 ; P2_R1215_U161
g19234 nand P2_R1215_U130 P2_R1215_U269 ; P2_R1215_U162
g19235 and P2_R1215_U476 P2_R1215_U475 ; P2_R1215_U163
g19236 nand P2_R1215_U257 P2_R1215_U256 ; P2_R1215_U164
g19237 and P2_R1215_U483 P2_R1215_U482 ; P2_R1215_U165
g19238 nand P2_R1215_U253 P2_R1215_U252 ; P2_R1215_U166
g19239 nand P2_R1215_U243 P2_R1215_U242 ; P2_R1215_U167
g19240 nand P2_R1215_U367 P2_R1215_U366 ; P2_R1215_U168
g19241 nand P2_U3056 P2_R1215_U151 ; P2_R1215_U169
g19242 not P2_R1215_U35 ; P2_R1215_U170
g19243 nand P2_U3456 P2_U3085 ; P2_R1215_U171
g19244 nand P2_U3074 P2_U3465 ; P2_R1215_U172
g19245 nand P2_U3060 P2_U3952 ; P2_R1215_U173
g19246 not P2_R1215_U69 ; P2_R1215_U174
g19247 not P2_R1215_U78 ; P2_R1215_U175
g19248 nand P2_U3067 P2_U3953 ; P2_R1215_U176
g19249 not P2_R1215_U62 ; P2_R1215_U177
g19250 or P2_U3069 P2_U3444 ; P2_R1215_U178
g19251 or P2_U3062 P2_U3441 ; P2_R1215_U179
g19252 or P2_U3438 P2_U3066 ; P2_R1215_U180
g19253 or P2_U3435 P2_U3070 ; P2_R1215_U181
g19254 not P2_R1215_U32 ; P2_R1215_U182
g19255 or P2_U3432 P2_U3080 ; P2_R1215_U183
g19256 not P2_R1215_U43 ; P2_R1215_U184
g19257 not P2_R1215_U44 ; P2_R1215_U185
g19258 nand P2_R1215_U43 P2_R1215_U44 ; P2_R1215_U186
g19259 nand P2_R1215_U116 P2_R1215_U180 ; P2_R1215_U187
g19260 nand P2_R1215_U5 P2_R1215_U186 ; P2_R1215_U188
g19261 nand P2_U3066 P2_U3438 ; P2_R1215_U189
g19262 nand P2_R1215_U117 P2_R1215_U188 ; P2_R1215_U190
g19263 nand P2_R1215_U36 P2_R1215_U35 ; P2_R1215_U191
g19264 nand P2_U3069 P2_R1215_U191 ; P2_R1215_U192
g19265 nand P2_R1215_U4 P2_R1215_U190 ; P2_R1215_U193
g19266 nand P2_U3444 P2_R1215_U170 ; P2_R1215_U194
g19267 not P2_R1215_U42 ; P2_R1215_U195
g19268 or P2_U3072 P2_U3450 ; P2_R1215_U196
g19269 or P2_U3073 P2_U3447 ; P2_R1215_U197
g19270 not P2_R1215_U23 ; P2_R1215_U198
g19271 nand P2_R1215_U24 P2_R1215_U23 ; P2_R1215_U199
g19272 nand P2_U3072 P2_R1215_U199 ; P2_R1215_U200
g19273 nand P2_U3450 P2_R1215_U198 ; P2_R1215_U201
g19274 nand P2_R1215_U6 P2_R1215_U42 ; P2_R1215_U202
g19275 not P2_R1215_U144 ; P2_R1215_U203
g19276 or P2_U3453 P2_U3086 ; P2_R1215_U204
g19277 nand P2_R1215_U204 P2_R1215_U144 ; P2_R1215_U205
g19278 not P2_R1215_U41 ; P2_R1215_U206
g19279 or P2_U3085 P2_U3456 ; P2_R1215_U207
g19280 or P2_U3447 P2_U3073 ; P2_R1215_U208
g19281 nand P2_R1215_U208 P2_R1215_U42 ; P2_R1215_U209
g19282 nand P2_R1215_U120 P2_R1215_U209 ; P2_R1215_U210
g19283 nand P2_R1215_U195 P2_R1215_U23 ; P2_R1215_U211
g19284 nand P2_U3450 P2_U3072 ; P2_R1215_U212
g19285 nand P2_R1215_U121 P2_R1215_U211 ; P2_R1215_U213
g19286 or P2_U3073 P2_U3447 ; P2_R1215_U214
g19287 nand P2_R1215_U185 P2_R1215_U181 ; P2_R1215_U215
g19288 nand P2_U3070 P2_U3435 ; P2_R1215_U216
g19289 not P2_R1215_U46 ; P2_R1215_U217
g19290 nand P2_R1215_U184 P2_R1215_U5 ; P2_R1215_U218
g19291 nand P2_R1215_U46 P2_R1215_U180 ; P2_R1215_U219
g19292 nand P2_U3066 P2_U3438 ; P2_R1215_U220
g19293 not P2_R1215_U45 ; P2_R1215_U221
g19294 or P2_U3441 P2_U3062 ; P2_R1215_U222
g19295 nand P2_R1215_U222 P2_R1215_U45 ; P2_R1215_U223
g19296 nand P2_R1215_U123 P2_R1215_U223 ; P2_R1215_U224
g19297 nand P2_R1215_U221 P2_R1215_U35 ; P2_R1215_U225
g19298 nand P2_U3444 P2_U3069 ; P2_R1215_U226
g19299 nand P2_R1215_U124 P2_R1215_U225 ; P2_R1215_U227
g19300 or P2_U3062 P2_U3441 ; P2_R1215_U228
g19301 nand P2_R1215_U184 P2_R1215_U181 ; P2_R1215_U229
g19302 not P2_R1215_U145 ; P2_R1215_U230
g19303 nand P2_U3066 P2_U3438 ; P2_R1215_U231
g19304 nand P2_R1215_U401 P2_R1215_U400 P2_R1215_U44 P2_R1215_U43 ; P2_R1215_U232
g19305 nand P2_R1215_U44 P2_R1215_U43 ; P2_R1215_U233
g19306 nand P2_U3070 P2_U3435 ; P2_R1215_U234
g19307 nand P2_R1215_U125 P2_R1215_U233 ; P2_R1215_U235
g19308 or P2_U3085 P2_U3456 ; P2_R1215_U236
g19309 or P2_U3064 P2_U3459 ; P2_R1215_U237
g19310 nand P2_R1215_U177 P2_R1215_U7 ; P2_R1215_U238
g19311 nand P2_U3064 P2_U3459 ; P2_R1215_U239
g19312 nand P2_R1215_U127 P2_R1215_U238 ; P2_R1215_U240
g19313 or P2_U3459 P2_U3064 ; P2_R1215_U241
g19314 nand P2_R1215_U126 P2_R1215_U144 ; P2_R1215_U242
g19315 nand P2_R1215_U241 P2_R1215_U240 ; P2_R1215_U243
g19316 not P2_R1215_U167 ; P2_R1215_U244
g19317 or P2_U3082 P2_U3468 ; P2_R1215_U245
g19318 or P2_U3074 P2_U3465 ; P2_R1215_U246
g19319 nand P2_R1215_U174 P2_R1215_U8 ; P2_R1215_U247
g19320 nand P2_U3082 P2_U3468 ; P2_R1215_U248
g19321 nand P2_R1215_U129 P2_R1215_U247 ; P2_R1215_U249
g19322 or P2_U3462 P2_U3065 ; P2_R1215_U250
g19323 or P2_U3468 P2_U3082 ; P2_R1215_U251
g19324 nand P2_R1215_U128 P2_R1215_U167 ; P2_R1215_U252
g19325 nand P2_R1215_U251 P2_R1215_U249 ; P2_R1215_U253
g19326 not P2_R1215_U166 ; P2_R1215_U254
g19327 or P2_U3471 P2_U3081 ; P2_R1215_U255
g19328 nand P2_R1215_U255 P2_R1215_U166 ; P2_R1215_U256
g19329 nand P2_U3081 P2_U3471 ; P2_R1215_U257
g19330 not P2_R1215_U164 ; P2_R1215_U258
g19331 or P2_U3474 P2_U3076 ; P2_R1215_U259
g19332 nand P2_R1215_U259 P2_R1215_U164 ; P2_R1215_U260
g19333 nand P2_U3076 P2_U3474 ; P2_R1215_U261
g19334 not P2_R1215_U93 ; P2_R1215_U262
g19335 or P2_U3071 P2_U3480 ; P2_R1215_U263
g19336 or P2_U3075 P2_U3477 ; P2_R1215_U264
g19337 not P2_R1215_U60 ; P2_R1215_U265
g19338 nand P2_R1215_U61 P2_R1215_U60 ; P2_R1215_U266
g19339 nand P2_U3071 P2_R1215_U266 ; P2_R1215_U267
g19340 nand P2_U3480 P2_R1215_U265 ; P2_R1215_U268
g19341 nand P2_R1215_U9 P2_R1215_U93 ; P2_R1215_U269
g19342 not P2_R1215_U162 ; P2_R1215_U270
g19343 or P2_U3078 P2_U3957 ; P2_R1215_U271
g19344 or P2_U3083 P2_U3485 ; P2_R1215_U272
g19345 or P2_U3077 P2_U3956 ; P2_R1215_U273
g19346 not P2_R1215_U81 ; P2_R1215_U274
g19347 nand P2_U3957 P2_R1215_U274 ; P2_R1215_U275
g19348 nand P2_R1215_U275 P2_R1215_U91 ; P2_R1215_U276
g19349 nand P2_R1215_U81 P2_R1215_U82 ; P2_R1215_U277
g19350 nand P2_R1215_U277 P2_R1215_U276 ; P2_R1215_U278
g19351 nand P2_R1215_U175 P2_R1215_U10 ; P2_R1215_U279
g19352 nand P2_U3077 P2_U3956 ; P2_R1215_U280
g19353 nand P2_R1215_U278 P2_R1215_U279 ; P2_R1215_U281
g19354 or P2_U3483 P2_U3084 ; P2_R1215_U282
g19355 or P2_U3956 P2_U3077 ; P2_R1215_U283
g19356 nand P2_R1215_U273 P2_R1215_U162 P2_R1215_U131 ; P2_R1215_U284
g19357 nand P2_R1215_U283 P2_R1215_U281 ; P2_R1215_U285
g19358 not P2_R1215_U159 ; P2_R1215_U286
g19359 or P2_U3955 P2_U3063 ; P2_R1215_U287
g19360 nand P2_R1215_U287 P2_R1215_U159 ; P2_R1215_U288
g19361 nand P2_U3063 P2_U3955 ; P2_R1215_U289
g19362 not P2_R1215_U157 ; P2_R1215_U290
g19363 or P2_U3954 P2_U3068 ; P2_R1215_U291
g19364 nand P2_R1215_U291 P2_R1215_U157 ; P2_R1215_U292
g19365 nand P2_U3068 P2_U3954 ; P2_R1215_U293
g19366 not P2_R1215_U155 ; P2_R1215_U294
g19367 or P2_U3060 P2_U3952 ; P2_R1215_U295
g19368 nand P2_R1215_U176 P2_R1215_U173 ; P2_R1215_U296
g19369 not P2_R1215_U87 ; P2_R1215_U297
g19370 or P2_U3953 P2_U3067 ; P2_R1215_U298
g19371 nand P2_R1215_U155 P2_R1215_U298 P2_R1215_U168 ; P2_R1215_U299
g19372 not P2_R1215_U153 ; P2_R1215_U300
g19373 or P2_U3950 P2_U3055 ; P2_R1215_U301
g19374 nand P2_U3055 P2_U3950 ; P2_R1215_U302
g19375 not P2_R1215_U151 ; P2_R1215_U303
g19376 nand P2_U3949 P2_R1215_U151 ; P2_R1215_U304
g19377 not P2_R1215_U149 ; P2_R1215_U305
g19378 nand P2_R1215_U298 P2_R1215_U155 ; P2_R1215_U306
g19379 not P2_R1215_U90 ; P2_R1215_U307
g19380 or P2_U3952 P2_U3060 ; P2_R1215_U308
g19381 nand P2_R1215_U308 P2_R1215_U90 ; P2_R1215_U309
g19382 nand P2_R1215_U309 P2_R1215_U173 P2_R1215_U154 ; P2_R1215_U310
g19383 nand P2_R1215_U307 P2_R1215_U173 ; P2_R1215_U311
g19384 nand P2_U3951 P2_U3059 ; P2_R1215_U312
g19385 nand P2_R1215_U311 P2_R1215_U312 P2_R1215_U168 ; P2_R1215_U313
g19386 or P2_U3060 P2_U3952 ; P2_R1215_U314
g19387 nand P2_R1215_U282 P2_R1215_U162 ; P2_R1215_U315
g19388 not P2_R1215_U92 ; P2_R1215_U316
g19389 nand P2_R1215_U10 P2_R1215_U92 ; P2_R1215_U317
g19390 nand P2_R1215_U135 P2_R1215_U317 ; P2_R1215_U318
g19391 nand P2_R1215_U317 P2_R1215_U278 ; P2_R1215_U319
g19392 nand P2_R1215_U453 P2_R1215_U319 ; P2_R1215_U320
g19393 or P2_U3485 P2_U3083 ; P2_R1215_U321
g19394 nand P2_R1215_U321 P2_R1215_U92 ; P2_R1215_U322
g19395 nand P2_R1215_U136 P2_R1215_U322 ; P2_R1215_U323
g19396 nand P2_R1215_U316 P2_R1215_U81 ; P2_R1215_U324
g19397 nand P2_U3078 P2_U3957 ; P2_R1215_U325
g19398 nand P2_R1215_U137 P2_R1215_U324 ; P2_R1215_U326
g19399 or P2_U3432 P2_U3080 ; P2_R1215_U327
g19400 not P2_R1215_U161 ; P2_R1215_U328
g19401 or P2_U3083 P2_U3485 ; P2_R1215_U329
g19402 or P2_U3477 P2_U3075 ; P2_R1215_U330
g19403 nand P2_R1215_U330 P2_R1215_U93 ; P2_R1215_U331
g19404 nand P2_R1215_U138 P2_R1215_U331 ; P2_R1215_U332
g19405 nand P2_R1215_U262 P2_R1215_U60 ; P2_R1215_U333
g19406 nand P2_U3480 P2_U3071 ; P2_R1215_U334
g19407 nand P2_R1215_U139 P2_R1215_U333 ; P2_R1215_U335
g19408 or P2_U3075 P2_U3477 ; P2_R1215_U336
g19409 nand P2_R1215_U250 P2_R1215_U167 ; P2_R1215_U337
g19410 not P2_R1215_U94 ; P2_R1215_U338
g19411 or P2_U3465 P2_U3074 ; P2_R1215_U339
g19412 nand P2_R1215_U339 P2_R1215_U94 ; P2_R1215_U340
g19413 nand P2_R1215_U140 P2_R1215_U340 ; P2_R1215_U341
g19414 nand P2_R1215_U338 P2_R1215_U172 ; P2_R1215_U342
g19415 nand P2_U3082 P2_U3468 ; P2_R1215_U343
g19416 nand P2_R1215_U141 P2_R1215_U342 ; P2_R1215_U344
g19417 or P2_U3074 P2_U3465 ; P2_R1215_U345
g19418 or P2_U3456 P2_U3085 ; P2_R1215_U346
g19419 nand P2_R1215_U346 P2_R1215_U41 ; P2_R1215_U347
g19420 nand P2_R1215_U142 P2_R1215_U347 ; P2_R1215_U348
g19421 nand P2_R1215_U206 P2_R1215_U171 ; P2_R1215_U349
g19422 nand P2_U3064 P2_U3459 ; P2_R1215_U350
g19423 nand P2_R1215_U143 P2_R1215_U349 ; P2_R1215_U351
g19424 nand P2_R1215_U207 P2_R1215_U171 ; P2_R1215_U352
g19425 nand P2_R1215_U204 P2_R1215_U62 ; P2_R1215_U353
g19426 nand P2_R1215_U214 P2_R1215_U23 ; P2_R1215_U354
g19427 nand P2_R1215_U228 P2_R1215_U35 ; P2_R1215_U355
g19428 nand P2_R1215_U231 P2_R1215_U180 ; P2_R1215_U356
g19429 nand P2_R1215_U314 P2_R1215_U173 ; P2_R1215_U357
g19430 nand P2_R1215_U298 P2_R1215_U176 ; P2_R1215_U358
g19431 nand P2_R1215_U329 P2_R1215_U81 ; P2_R1215_U359
g19432 nand P2_R1215_U282 P2_R1215_U78 ; P2_R1215_U360
g19433 nand P2_R1215_U336 P2_R1215_U60 ; P2_R1215_U361
g19434 nand P2_R1215_U345 P2_R1215_U172 ; P2_R1215_U362
g19435 nand P2_R1215_U250 P2_R1215_U69 ; P2_R1215_U363
g19436 nand P2_U3949 P2_U3056 ; P2_R1215_U364
g19437 nand P2_R1215_U296 P2_R1215_U168 ; P2_R1215_U365
g19438 nand P2_U3059 P2_R1215_U295 ; P2_R1215_U366
g19439 nand P2_U3951 P2_R1215_U295 ; P2_R1215_U367
g19440 nand P2_R1215_U296 P2_R1215_U168 P2_R1215_U301 ; P2_R1215_U368
g19441 nand P2_R1215_U155 P2_R1215_U168 P2_R1215_U133 ; P2_R1215_U369
g19442 nand P2_R1215_U297 P2_R1215_U301 ; P2_R1215_U370
g19443 nand P2_U3085 P2_R1215_U40 ; P2_R1215_U371
g19444 nand P2_U3456 P2_R1215_U39 ; P2_R1215_U372
g19445 nand P2_R1215_U372 P2_R1215_U371 ; P2_R1215_U373
g19446 nand P2_R1215_U352 P2_R1215_U41 ; P2_R1215_U374
g19447 nand P2_R1215_U373 P2_R1215_U206 ; P2_R1215_U375
g19448 nand P2_U3086 P2_R1215_U37 ; P2_R1215_U376
g19449 nand P2_U3453 P2_R1215_U38 ; P2_R1215_U377
g19450 nand P2_R1215_U377 P2_R1215_U376 ; P2_R1215_U378
g19451 nand P2_R1215_U353 P2_R1215_U144 ; P2_R1215_U379
g19452 nand P2_R1215_U203 P2_R1215_U378 ; P2_R1215_U380
g19453 nand P2_U3072 P2_R1215_U24 ; P2_R1215_U381
g19454 nand P2_U3450 P2_R1215_U22 ; P2_R1215_U382
g19455 nand P2_U3073 P2_R1215_U20 ; P2_R1215_U383
g19456 nand P2_U3447 P2_R1215_U21 ; P2_R1215_U384
g19457 nand P2_R1215_U384 P2_R1215_U383 ; P2_R1215_U385
g19458 nand P2_R1215_U354 P2_R1215_U42 ; P2_R1215_U386
g19459 nand P2_R1215_U385 P2_R1215_U195 ; P2_R1215_U387
g19460 nand P2_U3069 P2_R1215_U36 ; P2_R1215_U388
g19461 nand P2_U3444 P2_R1215_U27 ; P2_R1215_U389
g19462 nand P2_U3062 P2_R1215_U25 ; P2_R1215_U390
g19463 nand P2_U3441 P2_R1215_U26 ; P2_R1215_U391
g19464 nand P2_R1215_U391 P2_R1215_U390 ; P2_R1215_U392
g19465 nand P2_R1215_U355 P2_R1215_U45 ; P2_R1215_U393
g19466 nand P2_R1215_U392 P2_R1215_U221 ; P2_R1215_U394
g19467 nand P2_U3066 P2_R1215_U33 ; P2_R1215_U395
g19468 nand P2_U3438 P2_R1215_U34 ; P2_R1215_U396
g19469 nand P2_R1215_U396 P2_R1215_U395 ; P2_R1215_U397
g19470 nand P2_R1215_U356 P2_R1215_U145 ; P2_R1215_U398
g19471 nand P2_R1215_U230 P2_R1215_U397 ; P2_R1215_U399
g19472 nand P2_U3070 P2_R1215_U28 ; P2_R1215_U400
g19473 nand P2_U3435 P2_R1215_U29 ; P2_R1215_U401
g19474 nand P2_U3057 P2_R1215_U147 ; P2_R1215_U402
g19475 nand P2_U3960 P2_R1215_U146 ; P2_R1215_U403
g19476 nand P2_U3057 P2_R1215_U147 ; P2_R1215_U404
g19477 nand P2_U3960 P2_R1215_U146 ; P2_R1215_U405
g19478 nand P2_R1215_U405 P2_R1215_U404 ; P2_R1215_U406
g19479 nand P2_R1215_U148 P2_R1215_U149 ; P2_R1215_U407
g19480 nand P2_R1215_U305 P2_R1215_U406 ; P2_R1215_U408
g19481 nand P2_U3056 P2_R1215_U89 ; P2_R1215_U409
g19482 nand P2_U3949 P2_R1215_U88 ; P2_R1215_U410
g19483 nand P2_U3056 P2_R1215_U89 ; P2_R1215_U411
g19484 nand P2_U3949 P2_R1215_U88 ; P2_R1215_U412
g19485 nand P2_R1215_U412 P2_R1215_U411 ; P2_R1215_U413
g19486 nand P2_R1215_U150 P2_R1215_U151 ; P2_R1215_U414
g19487 nand P2_R1215_U303 P2_R1215_U413 ; P2_R1215_U415
g19488 nand P2_U3055 P2_R1215_U47 ; P2_R1215_U416
g19489 nand P2_U3950 P2_R1215_U48 ; P2_R1215_U417
g19490 nand P2_U3055 P2_R1215_U47 ; P2_R1215_U418
g19491 nand P2_U3950 P2_R1215_U48 ; P2_R1215_U419
g19492 nand P2_R1215_U419 P2_R1215_U418 ; P2_R1215_U420
g19493 nand P2_R1215_U152 P2_R1215_U153 ; P2_R1215_U421
g19494 nand P2_R1215_U300 P2_R1215_U420 ; P2_R1215_U422
g19495 nand P2_U3059 P2_R1215_U50 ; P2_R1215_U423
g19496 nand P2_U3951 P2_R1215_U49 ; P2_R1215_U424
g19497 nand P2_U3060 P2_R1215_U51 ; P2_R1215_U425
g19498 nand P2_U3952 P2_R1215_U52 ; P2_R1215_U426
g19499 nand P2_R1215_U426 P2_R1215_U425 ; P2_R1215_U427
g19500 nand P2_R1215_U357 P2_R1215_U90 ; P2_R1215_U428
g19501 nand P2_R1215_U427 P2_R1215_U307 ; P2_R1215_U429
g19502 nand P2_U3067 P2_R1215_U53 ; P2_R1215_U430
g19503 nand P2_U3953 P2_R1215_U54 ; P2_R1215_U431
g19504 nand P2_R1215_U431 P2_R1215_U430 ; P2_R1215_U432
g19505 nand P2_R1215_U358 P2_R1215_U155 ; P2_R1215_U433
g19506 nand P2_R1215_U294 P2_R1215_U432 ; P2_R1215_U434
g19507 nand P2_U3068 P2_R1215_U85 ; P2_R1215_U435
g19508 nand P2_U3954 P2_R1215_U86 ; P2_R1215_U436
g19509 nand P2_U3068 P2_R1215_U85 ; P2_R1215_U437
g19510 nand P2_U3954 P2_R1215_U86 ; P2_R1215_U438
g19511 nand P2_R1215_U438 P2_R1215_U437 ; P2_R1215_U439
g19512 nand P2_R1215_U156 P2_R1215_U157 ; P2_R1215_U440
g19513 nand P2_R1215_U290 P2_R1215_U439 ; P2_R1215_U441
g19514 nand P2_U3063 P2_R1215_U83 ; P2_R1215_U442
g19515 nand P2_U3955 P2_R1215_U84 ; P2_R1215_U443
g19516 nand P2_U3063 P2_R1215_U83 ; P2_R1215_U444
g19517 nand P2_U3955 P2_R1215_U84 ; P2_R1215_U445
g19518 nand P2_R1215_U445 P2_R1215_U444 ; P2_R1215_U446
g19519 nand P2_R1215_U158 P2_R1215_U159 ; P2_R1215_U447
g19520 nand P2_R1215_U286 P2_R1215_U446 ; P2_R1215_U448
g19521 nand P2_U3077 P2_R1215_U55 ; P2_R1215_U449
g19522 nand P2_U3956 P2_R1215_U56 ; P2_R1215_U450
g19523 nand P2_U3077 P2_R1215_U55 ; P2_R1215_U451
g19524 nand P2_U3956 P2_R1215_U56 ; P2_R1215_U452
g19525 nand P2_R1215_U452 P2_R1215_U451 ; P2_R1215_U453
g19526 nand P2_U3078 P2_R1215_U82 ; P2_R1215_U454
g19527 nand P2_U3957 P2_R1215_U91 ; P2_R1215_U455
g19528 nand P2_R1215_U182 P2_R1215_U161 ; P2_R1215_U456
g19529 nand P2_R1215_U328 P2_R1215_U32 ; P2_R1215_U457
g19530 nand P2_U3083 P2_R1215_U79 ; P2_R1215_U458
g19531 nand P2_U3485 P2_R1215_U80 ; P2_R1215_U459
g19532 nand P2_R1215_U459 P2_R1215_U458 ; P2_R1215_U460
g19533 nand P2_R1215_U359 P2_R1215_U92 ; P2_R1215_U461
g19534 nand P2_R1215_U460 P2_R1215_U316 ; P2_R1215_U462
g19535 nand P2_U3084 P2_R1215_U76 ; P2_R1215_U463
g19536 nand P2_U3483 P2_R1215_U77 ; P2_R1215_U464
g19537 nand P2_R1215_U464 P2_R1215_U463 ; P2_R1215_U465
g19538 nand P2_R1215_U360 P2_R1215_U162 ; P2_R1215_U466
g19539 nand P2_R1215_U270 P2_R1215_U465 ; P2_R1215_U467
g19540 nand P2_U3071 P2_R1215_U61 ; P2_R1215_U468
g19541 nand P2_U3480 P2_R1215_U59 ; P2_R1215_U469
g19542 nand P2_U3075 P2_R1215_U57 ; P2_R1215_U470
g19543 nand P2_U3477 P2_R1215_U58 ; P2_R1215_U471
g19544 nand P2_R1215_U471 P2_R1215_U470 ; P2_R1215_U472
g19545 nand P2_R1215_U361 P2_R1215_U93 ; P2_R1215_U473
g19546 nand P2_R1215_U472 P2_R1215_U262 ; P2_R1215_U474
g19547 nand P2_U3076 P2_R1215_U74 ; P2_R1215_U475
g19548 nand P2_U3474 P2_R1215_U75 ; P2_R1215_U476
g19549 nand P2_U3076 P2_R1215_U74 ; P2_R1215_U477
g19550 nand P2_U3474 P2_R1215_U75 ; P2_R1215_U478
g19551 nand P2_R1215_U478 P2_R1215_U477 ; P2_R1215_U479
g19552 nand P2_R1215_U163 P2_R1215_U164 ; P2_R1215_U480
g19553 nand P2_R1215_U258 P2_R1215_U479 ; P2_R1215_U481
g19554 nand P2_U3081 P2_R1215_U72 ; P2_R1215_U482
g19555 nand P2_U3471 P2_R1215_U73 ; P2_R1215_U483
g19556 nand P2_U3081 P2_R1215_U72 ; P2_R1215_U484
g19557 nand P2_U3471 P2_R1215_U73 ; P2_R1215_U485
g19558 nand P2_R1215_U485 P2_R1215_U484 ; P2_R1215_U486
g19559 nand P2_R1215_U165 P2_R1215_U166 ; P2_R1215_U487
g19560 nand P2_R1215_U254 P2_R1215_U486 ; P2_R1215_U488
g19561 nand P2_U3082 P2_R1215_U70 ; P2_R1215_U489
g19562 nand P2_U3468 P2_R1215_U71 ; P2_R1215_U490
g19563 nand P2_U3074 P2_R1215_U65 ; P2_R1215_U491
g19564 nand P2_U3465 P2_R1215_U66 ; P2_R1215_U492
g19565 nand P2_R1215_U492 P2_R1215_U491 ; P2_R1215_U493
g19566 nand P2_R1215_U362 P2_R1215_U94 ; P2_R1215_U494
g19567 nand P2_R1215_U493 P2_R1215_U338 ; P2_R1215_U495
g19568 nand P2_U3065 P2_R1215_U67 ; P2_R1215_U496
g19569 nand P2_U3462 P2_R1215_U68 ; P2_R1215_U497
g19570 nand P2_R1215_U497 P2_R1215_U496 ; P2_R1215_U498
g19571 nand P2_R1215_U363 P2_R1215_U167 ; P2_R1215_U499
g19572 nand P2_R1215_U244 P2_R1215_U498 ; P2_R1215_U500
g19573 nand P2_U3064 P2_R1215_U63 ; P2_R1215_U501
g19574 nand P2_U3459 P2_R1215_U64 ; P2_R1215_U502
g19575 nand P2_U3079 P2_R1215_U30 ; P2_R1215_U503
g19576 nand P2_U3427 P2_R1215_U31 ; P2_R1215_U504
g19577 and P2_R1164_U179 P2_R1164_U178 ; P2_R1164_U4
g19578 and P2_R1164_U197 P2_R1164_U196 ; P2_R1164_U5
g19579 and P2_R1164_U237 P2_R1164_U236 ; P2_R1164_U6
g19580 and P2_R1164_U246 P2_R1164_U245 ; P2_R1164_U7
g19581 and P2_R1164_U264 P2_R1164_U263 ; P2_R1164_U8
g19582 and P2_R1164_U272 P2_R1164_U271 ; P2_R1164_U9
g19583 and P2_R1164_U351 P2_R1164_U348 ; P2_R1164_U10
g19584 and P2_R1164_U344 P2_R1164_U341 ; P2_R1164_U11
g19585 and P2_R1164_U335 P2_R1164_U332 ; P2_R1164_U12
g19586 and P2_R1164_U326 P2_R1164_U323 ; P2_R1164_U13
g19587 and P2_R1164_U320 P2_R1164_U318 ; P2_R1164_U14
g19588 and P2_R1164_U313 P2_R1164_U310 ; P2_R1164_U15
g19589 and P2_R1164_U235 P2_R1164_U232 ; P2_R1164_U16
g19590 and P2_R1164_U227 P2_R1164_U224 ; P2_R1164_U17
g19591 and P2_R1164_U213 P2_R1164_U210 ; P2_R1164_U18
g19592 not P2_U3447 ; P2_R1164_U19
g19593 not P2_U3073 ; P2_R1164_U20
g19594 not P2_U3072 ; P2_R1164_U21
g19595 nand P2_U3073 P2_U3447 ; P2_R1164_U22
g19596 not P2_U3450 ; P2_R1164_U23
g19597 not P2_U3441 ; P2_R1164_U24
g19598 not P2_U3062 ; P2_R1164_U25
g19599 not P2_U3069 ; P2_R1164_U26
g19600 not P2_U3435 ; P2_R1164_U27
g19601 not P2_U3070 ; P2_R1164_U28
g19602 not P2_U3427 ; P2_R1164_U29
g19603 not P2_U3079 ; P2_R1164_U30
g19604 nand P2_U3079 P2_U3427 ; P2_R1164_U31
g19605 not P2_U3438 ; P2_R1164_U32
g19606 not P2_U3066 ; P2_R1164_U33
g19607 nand P2_U3062 P2_U3441 ; P2_R1164_U34
g19608 not P2_U3444 ; P2_R1164_U35
g19609 not P2_U3453 ; P2_R1164_U36
g19610 not P2_U3086 ; P2_R1164_U37
g19611 not P2_U3085 ; P2_R1164_U38
g19612 not P2_U3456 ; P2_R1164_U39
g19613 nand P2_R1164_U61 P2_R1164_U205 ; P2_R1164_U40
g19614 nand P2_R1164_U117 P2_R1164_U193 ; P2_R1164_U41
g19615 nand P2_R1164_U182 P2_R1164_U183 ; P2_R1164_U42
g19616 nand P2_U3432 P2_U3080 ; P2_R1164_U43
g19617 nand P2_R1164_U122 P2_R1164_U219 ; P2_R1164_U44
g19618 nand P2_R1164_U216 P2_R1164_U215 ; P2_R1164_U45
g19619 not P2_U3950 ; P2_R1164_U46
g19620 not P2_U3055 ; P2_R1164_U47
g19621 not P2_U3059 ; P2_R1164_U48
g19622 not P2_U3951 ; P2_R1164_U49
g19623 not P2_U3952 ; P2_R1164_U50
g19624 not P2_U3060 ; P2_R1164_U51
g19625 not P2_U3953 ; P2_R1164_U52
g19626 not P2_U3067 ; P2_R1164_U53
g19627 not P2_U3956 ; P2_R1164_U54
g19628 not P2_U3077 ; P2_R1164_U55
g19629 not P2_U3477 ; P2_R1164_U56
g19630 not P2_U3075 ; P2_R1164_U57
g19631 not P2_U3071 ; P2_R1164_U58
g19632 nand P2_U3075 P2_U3477 ; P2_R1164_U59
g19633 not P2_U3480 ; P2_R1164_U60
g19634 nand P2_U3086 P2_U3453 ; P2_R1164_U61
g19635 not P2_U3459 ; P2_R1164_U62
g19636 not P2_U3064 ; P2_R1164_U63
g19637 not P2_U3465 ; P2_R1164_U64
g19638 not P2_U3074 ; P2_R1164_U65
g19639 not P2_U3462 ; P2_R1164_U66
g19640 not P2_U3065 ; P2_R1164_U67
g19641 nand P2_U3065 P2_U3462 ; P2_R1164_U68
g19642 not P2_U3468 ; P2_R1164_U69
g19643 not P2_U3082 ; P2_R1164_U70
g19644 not P2_U3471 ; P2_R1164_U71
g19645 not P2_U3081 ; P2_R1164_U72
g19646 not P2_U3474 ; P2_R1164_U73
g19647 not P2_U3076 ; P2_R1164_U74
g19648 not P2_U3483 ; P2_R1164_U75
g19649 not P2_U3084 ; P2_R1164_U76
g19650 nand P2_U3084 P2_U3483 ; P2_R1164_U77
g19651 not P2_U3485 ; P2_R1164_U78
g19652 not P2_U3083 ; P2_R1164_U79
g19653 nand P2_U3083 P2_U3485 ; P2_R1164_U80
g19654 not P2_U3957 ; P2_R1164_U81
g19655 not P2_U3955 ; P2_R1164_U82
g19656 not P2_U3063 ; P2_R1164_U83
g19657 not P2_U3954 ; P2_R1164_U84
g19658 not P2_U3068 ; P2_R1164_U85
g19659 nand P2_U3951 P2_U3059 ; P2_R1164_U86
g19660 not P2_U3056 ; P2_R1164_U87
g19661 not P2_U3949 ; P2_R1164_U88
g19662 nand P2_R1164_U306 P2_R1164_U176 ; P2_R1164_U89
g19663 not P2_U3078 ; P2_R1164_U90
g19664 nand P2_R1164_U77 P2_R1164_U315 ; P2_R1164_U91
g19665 nand P2_R1164_U261 P2_R1164_U260 ; P2_R1164_U92
g19666 nand P2_R1164_U68 P2_R1164_U337 ; P2_R1164_U93
g19667 nand P2_R1164_U457 P2_R1164_U456 ; P2_R1164_U94
g19668 nand P2_R1164_U504 P2_R1164_U503 ; P2_R1164_U95
g19669 nand P2_R1164_U375 P2_R1164_U374 ; P2_R1164_U96
g19670 nand P2_R1164_U380 P2_R1164_U379 ; P2_R1164_U97
g19671 nand P2_R1164_U387 P2_R1164_U386 ; P2_R1164_U98
g19672 nand P2_R1164_U394 P2_R1164_U393 ; P2_R1164_U99
g19673 nand P2_R1164_U399 P2_R1164_U398 ; P2_R1164_U100
g19674 nand P2_R1164_U408 P2_R1164_U407 ; P2_R1164_U101
g19675 nand P2_R1164_U415 P2_R1164_U414 ; P2_R1164_U102
g19676 nand P2_R1164_U422 P2_R1164_U421 ; P2_R1164_U103
g19677 nand P2_R1164_U429 P2_R1164_U428 ; P2_R1164_U104
g19678 nand P2_R1164_U434 P2_R1164_U433 ; P2_R1164_U105
g19679 nand P2_R1164_U441 P2_R1164_U440 ; P2_R1164_U106
g19680 nand P2_R1164_U448 P2_R1164_U447 ; P2_R1164_U107
g19681 nand P2_R1164_U462 P2_R1164_U461 ; P2_R1164_U108
g19682 nand P2_R1164_U467 P2_R1164_U466 ; P2_R1164_U109
g19683 nand P2_R1164_U474 P2_R1164_U473 ; P2_R1164_U110
g19684 nand P2_R1164_U481 P2_R1164_U480 ; P2_R1164_U111
g19685 nand P2_R1164_U488 P2_R1164_U487 ; P2_R1164_U112
g19686 nand P2_R1164_U495 P2_R1164_U494 ; P2_R1164_U113
g19687 nand P2_R1164_U500 P2_R1164_U499 ; P2_R1164_U114
g19688 and P2_R1164_U189 P2_R1164_U187 ; P2_R1164_U115
g19689 and P2_R1164_U4 P2_R1164_U180 ; P2_R1164_U116
g19690 and P2_R1164_U194 P2_R1164_U192 ; P2_R1164_U117
g19691 and P2_R1164_U201 P2_R1164_U200 ; P2_R1164_U118
g19692 and P2_R1164_U382 P2_R1164_U381 P2_R1164_U22 ; P2_R1164_U119
g19693 and P2_R1164_U212 P2_R1164_U5 ; P2_R1164_U120
g19694 and P2_R1164_U181 P2_R1164_U180 ; P2_R1164_U121
g19695 and P2_R1164_U220 P2_R1164_U218 ; P2_R1164_U122
g19696 and P2_R1164_U389 P2_R1164_U388 P2_R1164_U34 ; P2_R1164_U123
g19697 and P2_R1164_U226 P2_R1164_U4 ; P2_R1164_U124
g19698 and P2_R1164_U234 P2_R1164_U181 ; P2_R1164_U125
g19699 and P2_R1164_U204 P2_R1164_U6 ; P2_R1164_U126
g19700 and P2_R1164_U239 P2_R1164_U171 ; P2_R1164_U127
g19701 and P2_R1164_U250 P2_R1164_U7 ; P2_R1164_U128
g19702 and P2_R1164_U248 P2_R1164_U172 ; P2_R1164_U129
g19703 and P2_R1164_U268 P2_R1164_U267 ; P2_R1164_U130
g19704 and P2_R1164_U9 P2_R1164_U282 ; P2_R1164_U131
g19705 and P2_R1164_U285 P2_R1164_U280 ; P2_R1164_U132
g19706 and P2_R1164_U301 P2_R1164_U298 ; P2_R1164_U133
g19707 and P2_R1164_U368 P2_R1164_U302 ; P2_R1164_U134
g19708 and P2_R1164_U160 P2_R1164_U278 ; P2_R1164_U135
g19709 and P2_R1164_U455 P2_R1164_U454 P2_R1164_U80 ; P2_R1164_U136
g19710 and P2_R1164_U325 P2_R1164_U9 ; P2_R1164_U137
g19711 and P2_R1164_U469 P2_R1164_U468 P2_R1164_U59 ; P2_R1164_U138
g19712 and P2_R1164_U334 P2_R1164_U8 ; P2_R1164_U139
g19713 and P2_R1164_U490 P2_R1164_U489 P2_R1164_U172 ; P2_R1164_U140
g19714 and P2_R1164_U343 P2_R1164_U7 ; P2_R1164_U141
g19715 and P2_R1164_U502 P2_R1164_U501 P2_R1164_U171 ; P2_R1164_U142
g19716 and P2_R1164_U350 P2_R1164_U6 ; P2_R1164_U143
g19717 nand P2_R1164_U118 P2_R1164_U202 ; P2_R1164_U144
g19718 nand P2_R1164_U217 P2_R1164_U229 ; P2_R1164_U145
g19719 not P2_U3057 ; P2_R1164_U146
g19720 not P2_U3960 ; P2_R1164_U147
g19721 and P2_R1164_U403 P2_R1164_U402 ; P2_R1164_U148
g19722 nand P2_R1164_U304 P2_R1164_U169 P2_R1164_U364 ; P2_R1164_U149
g19723 and P2_R1164_U410 P2_R1164_U409 ; P2_R1164_U150
g19724 nand P2_R1164_U370 P2_R1164_U369 P2_R1164_U134 ; P2_R1164_U151
g19725 and P2_R1164_U417 P2_R1164_U416 ; P2_R1164_U152
g19726 nand P2_R1164_U365 P2_R1164_U299 P2_R1164_U86 ; P2_R1164_U153
g19727 and P2_R1164_U424 P2_R1164_U423 ; P2_R1164_U154
g19728 nand P2_R1164_U293 P2_R1164_U292 ; P2_R1164_U155
g19729 and P2_R1164_U436 P2_R1164_U435 ; P2_R1164_U156
g19730 nand P2_R1164_U289 P2_R1164_U288 ; P2_R1164_U157
g19731 and P2_R1164_U443 P2_R1164_U442 ; P2_R1164_U158
g19732 nand P2_R1164_U132 P2_R1164_U284 ; P2_R1164_U159
g19733 and P2_R1164_U450 P2_R1164_U449 ; P2_R1164_U160
g19734 nand P2_R1164_U43 P2_R1164_U327 ; P2_R1164_U161
g19735 nand P2_R1164_U130 P2_R1164_U269 ; P2_R1164_U162
g19736 and P2_R1164_U476 P2_R1164_U475 ; P2_R1164_U163
g19737 nand P2_R1164_U257 P2_R1164_U256 ; P2_R1164_U164
g19738 and P2_R1164_U483 P2_R1164_U482 ; P2_R1164_U165
g19739 nand P2_R1164_U253 P2_R1164_U252 ; P2_R1164_U166
g19740 nand P2_R1164_U243 P2_R1164_U242 ; P2_R1164_U167
g19741 nand P2_R1164_U367 P2_R1164_U366 ; P2_R1164_U168
g19742 nand P2_U3056 P2_R1164_U151 ; P2_R1164_U169
g19743 not P2_R1164_U34 ; P2_R1164_U170
g19744 nand P2_U3456 P2_U3085 ; P2_R1164_U171
g19745 nand P2_U3074 P2_U3465 ; P2_R1164_U172
g19746 nand P2_U3060 P2_U3952 ; P2_R1164_U173
g19747 not P2_R1164_U68 ; P2_R1164_U174
g19748 not P2_R1164_U77 ; P2_R1164_U175
g19749 nand P2_U3067 P2_U3953 ; P2_R1164_U176
g19750 not P2_R1164_U61 ; P2_R1164_U177
g19751 or P2_U3069 P2_U3444 ; P2_R1164_U178
g19752 or P2_U3062 P2_U3441 ; P2_R1164_U179
g19753 or P2_U3438 P2_U3066 ; P2_R1164_U180
g19754 or P2_U3435 P2_U3070 ; P2_R1164_U181
g19755 not P2_R1164_U31 ; P2_R1164_U182
g19756 or P2_U3432 P2_U3080 ; P2_R1164_U183
g19757 not P2_R1164_U42 ; P2_R1164_U184
g19758 not P2_R1164_U43 ; P2_R1164_U185
g19759 nand P2_R1164_U42 P2_R1164_U43 ; P2_R1164_U186
g19760 nand P2_U3070 P2_U3435 ; P2_R1164_U187
g19761 nand P2_R1164_U186 P2_R1164_U181 ; P2_R1164_U188
g19762 nand P2_U3066 P2_U3438 ; P2_R1164_U189
g19763 nand P2_R1164_U115 P2_R1164_U188 ; P2_R1164_U190
g19764 nand P2_R1164_U35 P2_R1164_U34 ; P2_R1164_U191
g19765 nand P2_U3069 P2_R1164_U191 ; P2_R1164_U192
g19766 nand P2_R1164_U116 P2_R1164_U190 ; P2_R1164_U193
g19767 nand P2_U3444 P2_R1164_U170 ; P2_R1164_U194
g19768 not P2_R1164_U41 ; P2_R1164_U195
g19769 or P2_U3072 P2_U3450 ; P2_R1164_U196
g19770 or P2_U3073 P2_U3447 ; P2_R1164_U197
g19771 not P2_R1164_U22 ; P2_R1164_U198
g19772 nand P2_R1164_U23 P2_R1164_U22 ; P2_R1164_U199
g19773 nand P2_U3072 P2_R1164_U199 ; P2_R1164_U200
g19774 nand P2_U3450 P2_R1164_U198 ; P2_R1164_U201
g19775 nand P2_R1164_U5 P2_R1164_U41 ; P2_R1164_U202
g19776 not P2_R1164_U144 ; P2_R1164_U203
g19777 or P2_U3453 P2_U3086 ; P2_R1164_U204
g19778 nand P2_R1164_U204 P2_R1164_U144 ; P2_R1164_U205
g19779 not P2_R1164_U40 ; P2_R1164_U206
g19780 or P2_U3085 P2_U3456 ; P2_R1164_U207
g19781 or P2_U3447 P2_U3073 ; P2_R1164_U208
g19782 nand P2_R1164_U208 P2_R1164_U41 ; P2_R1164_U209
g19783 nand P2_R1164_U119 P2_R1164_U209 ; P2_R1164_U210
g19784 nand P2_R1164_U195 P2_R1164_U22 ; P2_R1164_U211
g19785 nand P2_U3450 P2_U3072 ; P2_R1164_U212
g19786 nand P2_R1164_U120 P2_R1164_U211 ; P2_R1164_U213
g19787 or P2_U3073 P2_U3447 ; P2_R1164_U214
g19788 nand P2_R1164_U185 P2_R1164_U181 ; P2_R1164_U215
g19789 nand P2_U3070 P2_U3435 ; P2_R1164_U216
g19790 not P2_R1164_U45 ; P2_R1164_U217
g19791 nand P2_R1164_U121 P2_R1164_U184 ; P2_R1164_U218
g19792 nand P2_R1164_U45 P2_R1164_U180 ; P2_R1164_U219
g19793 nand P2_U3066 P2_U3438 ; P2_R1164_U220
g19794 not P2_R1164_U44 ; P2_R1164_U221
g19795 or P2_U3441 P2_U3062 ; P2_R1164_U222
g19796 nand P2_R1164_U222 P2_R1164_U44 ; P2_R1164_U223
g19797 nand P2_R1164_U123 P2_R1164_U223 ; P2_R1164_U224
g19798 nand P2_R1164_U221 P2_R1164_U34 ; P2_R1164_U225
g19799 nand P2_U3444 P2_U3069 ; P2_R1164_U226
g19800 nand P2_R1164_U124 P2_R1164_U225 ; P2_R1164_U227
g19801 or P2_U3062 P2_U3441 ; P2_R1164_U228
g19802 nand P2_R1164_U184 P2_R1164_U181 ; P2_R1164_U229
g19803 not P2_R1164_U145 ; P2_R1164_U230
g19804 nand P2_U3066 P2_U3438 ; P2_R1164_U231
g19805 nand P2_R1164_U401 P2_R1164_U400 P2_R1164_U43 P2_R1164_U42 ; P2_R1164_U232
g19806 nand P2_R1164_U43 P2_R1164_U42 ; P2_R1164_U233
g19807 nand P2_U3070 P2_U3435 ; P2_R1164_U234
g19808 nand P2_R1164_U125 P2_R1164_U233 ; P2_R1164_U235
g19809 or P2_U3085 P2_U3456 ; P2_R1164_U236
g19810 or P2_U3064 P2_U3459 ; P2_R1164_U237
g19811 nand P2_R1164_U177 P2_R1164_U6 ; P2_R1164_U238
g19812 nand P2_U3064 P2_U3459 ; P2_R1164_U239
g19813 nand P2_R1164_U127 P2_R1164_U238 ; P2_R1164_U240
g19814 or P2_U3459 P2_U3064 ; P2_R1164_U241
g19815 nand P2_R1164_U126 P2_R1164_U144 ; P2_R1164_U242
g19816 nand P2_R1164_U241 P2_R1164_U240 ; P2_R1164_U243
g19817 not P2_R1164_U167 ; P2_R1164_U244
g19818 or P2_U3082 P2_U3468 ; P2_R1164_U245
g19819 or P2_U3074 P2_U3465 ; P2_R1164_U246
g19820 nand P2_R1164_U174 P2_R1164_U7 ; P2_R1164_U247
g19821 nand P2_U3082 P2_U3468 ; P2_R1164_U248
g19822 nand P2_R1164_U129 P2_R1164_U247 ; P2_R1164_U249
g19823 or P2_U3462 P2_U3065 ; P2_R1164_U250
g19824 or P2_U3468 P2_U3082 ; P2_R1164_U251
g19825 nand P2_R1164_U128 P2_R1164_U167 ; P2_R1164_U252
g19826 nand P2_R1164_U251 P2_R1164_U249 ; P2_R1164_U253
g19827 not P2_R1164_U166 ; P2_R1164_U254
g19828 or P2_U3471 P2_U3081 ; P2_R1164_U255
g19829 nand P2_R1164_U255 P2_R1164_U166 ; P2_R1164_U256
g19830 nand P2_U3081 P2_U3471 ; P2_R1164_U257
g19831 not P2_R1164_U164 ; P2_R1164_U258
g19832 or P2_U3474 P2_U3076 ; P2_R1164_U259
g19833 nand P2_R1164_U259 P2_R1164_U164 ; P2_R1164_U260
g19834 nand P2_U3076 P2_U3474 ; P2_R1164_U261
g19835 not P2_R1164_U92 ; P2_R1164_U262
g19836 or P2_U3071 P2_U3480 ; P2_R1164_U263
g19837 or P2_U3075 P2_U3477 ; P2_R1164_U264
g19838 not P2_R1164_U59 ; P2_R1164_U265
g19839 nand P2_R1164_U60 P2_R1164_U59 ; P2_R1164_U266
g19840 nand P2_U3071 P2_R1164_U266 ; P2_R1164_U267
g19841 nand P2_U3480 P2_R1164_U265 ; P2_R1164_U268
g19842 nand P2_R1164_U8 P2_R1164_U92 ; P2_R1164_U269
g19843 not P2_R1164_U162 ; P2_R1164_U270
g19844 or P2_U3078 P2_U3957 ; P2_R1164_U271
g19845 or P2_U3083 P2_U3485 ; P2_R1164_U272
g19846 or P2_U3077 P2_U3956 ; P2_R1164_U273
g19847 not P2_R1164_U80 ; P2_R1164_U274
g19848 nand P2_U3957 P2_R1164_U274 ; P2_R1164_U275
g19849 nand P2_R1164_U275 P2_R1164_U90 ; P2_R1164_U276
g19850 nand P2_R1164_U80 P2_R1164_U81 ; P2_R1164_U277
g19851 nand P2_R1164_U277 P2_R1164_U276 ; P2_R1164_U278
g19852 nand P2_R1164_U175 P2_R1164_U9 ; P2_R1164_U279
g19853 nand P2_U3077 P2_U3956 ; P2_R1164_U280
g19854 nand P2_R1164_U278 P2_R1164_U279 ; P2_R1164_U281
g19855 or P2_U3483 P2_U3084 ; P2_R1164_U282
g19856 or P2_U3956 P2_U3077 ; P2_R1164_U283
g19857 nand P2_R1164_U273 P2_R1164_U162 P2_R1164_U131 ; P2_R1164_U284
g19858 nand P2_R1164_U283 P2_R1164_U281 ; P2_R1164_U285
g19859 not P2_R1164_U159 ; P2_R1164_U286
g19860 or P2_U3955 P2_U3063 ; P2_R1164_U287
g19861 nand P2_R1164_U287 P2_R1164_U159 ; P2_R1164_U288
g19862 nand P2_U3063 P2_U3955 ; P2_R1164_U289
g19863 not P2_R1164_U157 ; P2_R1164_U290
g19864 or P2_U3954 P2_U3068 ; P2_R1164_U291
g19865 nand P2_R1164_U291 P2_R1164_U157 ; P2_R1164_U292
g19866 nand P2_U3068 P2_U3954 ; P2_R1164_U293
g19867 not P2_R1164_U155 ; P2_R1164_U294
g19868 or P2_U3060 P2_U3952 ; P2_R1164_U295
g19869 nand P2_R1164_U176 P2_R1164_U173 ; P2_R1164_U296
g19870 not P2_R1164_U86 ; P2_R1164_U297
g19871 or P2_U3953 P2_U3067 ; P2_R1164_U298
g19872 nand P2_R1164_U155 P2_R1164_U298 P2_R1164_U168 ; P2_R1164_U299
g19873 not P2_R1164_U153 ; P2_R1164_U300
g19874 or P2_U3950 P2_U3055 ; P2_R1164_U301
g19875 nand P2_U3055 P2_U3950 ; P2_R1164_U302
g19876 not P2_R1164_U151 ; P2_R1164_U303
g19877 nand P2_U3949 P2_R1164_U151 ; P2_R1164_U304
g19878 not P2_R1164_U149 ; P2_R1164_U305
g19879 nand P2_R1164_U298 P2_R1164_U155 ; P2_R1164_U306
g19880 not P2_R1164_U89 ; P2_R1164_U307
g19881 or P2_U3952 P2_U3060 ; P2_R1164_U308
g19882 nand P2_R1164_U308 P2_R1164_U89 ; P2_R1164_U309
g19883 nand P2_R1164_U309 P2_R1164_U173 P2_R1164_U154 ; P2_R1164_U310
g19884 nand P2_R1164_U307 P2_R1164_U173 ; P2_R1164_U311
g19885 nand P2_U3951 P2_U3059 ; P2_R1164_U312
g19886 nand P2_R1164_U311 P2_R1164_U312 P2_R1164_U168 ; P2_R1164_U313
g19887 or P2_U3060 P2_U3952 ; P2_R1164_U314
g19888 nand P2_R1164_U282 P2_R1164_U162 ; P2_R1164_U315
g19889 not P2_R1164_U91 ; P2_R1164_U316
g19890 nand P2_R1164_U9 P2_R1164_U91 ; P2_R1164_U317
g19891 nand P2_R1164_U135 P2_R1164_U317 ; P2_R1164_U318
g19892 nand P2_R1164_U317 P2_R1164_U278 ; P2_R1164_U319
g19893 nand P2_R1164_U453 P2_R1164_U319 ; P2_R1164_U320
g19894 or P2_U3485 P2_U3083 ; P2_R1164_U321
g19895 nand P2_R1164_U321 P2_R1164_U91 ; P2_R1164_U322
g19896 nand P2_R1164_U136 P2_R1164_U322 ; P2_R1164_U323
g19897 nand P2_R1164_U316 P2_R1164_U80 ; P2_R1164_U324
g19898 nand P2_U3078 P2_U3957 ; P2_R1164_U325
g19899 nand P2_R1164_U137 P2_R1164_U324 ; P2_R1164_U326
g19900 or P2_U3432 P2_U3080 ; P2_R1164_U327
g19901 not P2_R1164_U161 ; P2_R1164_U328
g19902 or P2_U3083 P2_U3485 ; P2_R1164_U329
g19903 or P2_U3477 P2_U3075 ; P2_R1164_U330
g19904 nand P2_R1164_U330 P2_R1164_U92 ; P2_R1164_U331
g19905 nand P2_R1164_U138 P2_R1164_U331 ; P2_R1164_U332
g19906 nand P2_R1164_U262 P2_R1164_U59 ; P2_R1164_U333
g19907 nand P2_U3480 P2_U3071 ; P2_R1164_U334
g19908 nand P2_R1164_U139 P2_R1164_U333 ; P2_R1164_U335
g19909 or P2_U3075 P2_U3477 ; P2_R1164_U336
g19910 nand P2_R1164_U250 P2_R1164_U167 ; P2_R1164_U337
g19911 not P2_R1164_U93 ; P2_R1164_U338
g19912 or P2_U3465 P2_U3074 ; P2_R1164_U339
g19913 nand P2_R1164_U339 P2_R1164_U93 ; P2_R1164_U340
g19914 nand P2_R1164_U140 P2_R1164_U340 ; P2_R1164_U341
g19915 nand P2_R1164_U338 P2_R1164_U172 ; P2_R1164_U342
g19916 nand P2_U3082 P2_U3468 ; P2_R1164_U343
g19917 nand P2_R1164_U141 P2_R1164_U342 ; P2_R1164_U344
g19918 or P2_U3074 P2_U3465 ; P2_R1164_U345
g19919 or P2_U3456 P2_U3085 ; P2_R1164_U346
g19920 nand P2_R1164_U346 P2_R1164_U40 ; P2_R1164_U347
g19921 nand P2_R1164_U142 P2_R1164_U347 ; P2_R1164_U348
g19922 nand P2_R1164_U206 P2_R1164_U171 ; P2_R1164_U349
g19923 nand P2_U3064 P2_U3459 ; P2_R1164_U350
g19924 nand P2_R1164_U143 P2_R1164_U349 ; P2_R1164_U351
g19925 nand P2_R1164_U207 P2_R1164_U171 ; P2_R1164_U352
g19926 nand P2_R1164_U204 P2_R1164_U61 ; P2_R1164_U353
g19927 nand P2_R1164_U214 P2_R1164_U22 ; P2_R1164_U354
g19928 nand P2_R1164_U228 P2_R1164_U34 ; P2_R1164_U355
g19929 nand P2_R1164_U231 P2_R1164_U180 ; P2_R1164_U356
g19930 nand P2_R1164_U314 P2_R1164_U173 ; P2_R1164_U357
g19931 nand P2_R1164_U298 P2_R1164_U176 ; P2_R1164_U358
g19932 nand P2_R1164_U329 P2_R1164_U80 ; P2_R1164_U359
g19933 nand P2_R1164_U282 P2_R1164_U77 ; P2_R1164_U360
g19934 nand P2_R1164_U336 P2_R1164_U59 ; P2_R1164_U361
g19935 nand P2_R1164_U345 P2_R1164_U172 ; P2_R1164_U362
g19936 nand P2_R1164_U250 P2_R1164_U68 ; P2_R1164_U363
g19937 nand P2_U3949 P2_U3056 ; P2_R1164_U364
g19938 nand P2_R1164_U296 P2_R1164_U168 ; P2_R1164_U365
g19939 nand P2_U3059 P2_R1164_U295 ; P2_R1164_U366
g19940 nand P2_U3951 P2_R1164_U295 ; P2_R1164_U367
g19941 nand P2_R1164_U296 P2_R1164_U168 P2_R1164_U301 ; P2_R1164_U368
g19942 nand P2_R1164_U155 P2_R1164_U168 P2_R1164_U133 ; P2_R1164_U369
g19943 nand P2_R1164_U297 P2_R1164_U301 ; P2_R1164_U370
g19944 nand P2_U3085 P2_R1164_U39 ; P2_R1164_U371
g19945 nand P2_U3456 P2_R1164_U38 ; P2_R1164_U372
g19946 nand P2_R1164_U372 P2_R1164_U371 ; P2_R1164_U373
g19947 nand P2_R1164_U352 P2_R1164_U40 ; P2_R1164_U374
g19948 nand P2_R1164_U373 P2_R1164_U206 ; P2_R1164_U375
g19949 nand P2_U3086 P2_R1164_U36 ; P2_R1164_U376
g19950 nand P2_U3453 P2_R1164_U37 ; P2_R1164_U377
g19951 nand P2_R1164_U377 P2_R1164_U376 ; P2_R1164_U378
g19952 nand P2_R1164_U353 P2_R1164_U144 ; P2_R1164_U379
g19953 nand P2_R1164_U203 P2_R1164_U378 ; P2_R1164_U380
g19954 nand P2_U3072 P2_R1164_U23 ; P2_R1164_U381
g19955 nand P2_U3450 P2_R1164_U21 ; P2_R1164_U382
g19956 nand P2_U3073 P2_R1164_U19 ; P2_R1164_U383
g19957 nand P2_U3447 P2_R1164_U20 ; P2_R1164_U384
g19958 nand P2_R1164_U384 P2_R1164_U383 ; P2_R1164_U385
g19959 nand P2_R1164_U354 P2_R1164_U41 ; P2_R1164_U386
g19960 nand P2_R1164_U385 P2_R1164_U195 ; P2_R1164_U387
g19961 nand P2_U3069 P2_R1164_U35 ; P2_R1164_U388
g19962 nand P2_U3444 P2_R1164_U26 ; P2_R1164_U389
g19963 nand P2_U3062 P2_R1164_U24 ; P2_R1164_U390
g19964 nand P2_U3441 P2_R1164_U25 ; P2_R1164_U391
g19965 nand P2_R1164_U391 P2_R1164_U390 ; P2_R1164_U392
g19966 nand P2_R1164_U355 P2_R1164_U44 ; P2_R1164_U393
g19967 nand P2_R1164_U392 P2_R1164_U221 ; P2_R1164_U394
g19968 nand P2_U3066 P2_R1164_U32 ; P2_R1164_U395
g19969 nand P2_U3438 P2_R1164_U33 ; P2_R1164_U396
g19970 nand P2_R1164_U396 P2_R1164_U395 ; P2_R1164_U397
g19971 nand P2_R1164_U356 P2_R1164_U145 ; P2_R1164_U398
g19972 nand P2_R1164_U230 P2_R1164_U397 ; P2_R1164_U399
g19973 nand P2_U3070 P2_R1164_U27 ; P2_R1164_U400
g19974 nand P2_U3435 P2_R1164_U28 ; P2_R1164_U401
g19975 nand P2_U3057 P2_R1164_U147 ; P2_R1164_U402
g19976 nand P2_U3960 P2_R1164_U146 ; P2_R1164_U403
g19977 nand P2_U3057 P2_R1164_U147 ; P2_R1164_U404
g19978 nand P2_U3960 P2_R1164_U146 ; P2_R1164_U405
g19979 nand P2_R1164_U405 P2_R1164_U404 ; P2_R1164_U406
g19980 nand P2_R1164_U148 P2_R1164_U149 ; P2_R1164_U407
g19981 nand P2_R1164_U305 P2_R1164_U406 ; P2_R1164_U408
g19982 nand P2_U3056 P2_R1164_U88 ; P2_R1164_U409
g19983 nand P2_U3949 P2_R1164_U87 ; P2_R1164_U410
g19984 nand P2_U3056 P2_R1164_U88 ; P2_R1164_U411
g19985 nand P2_U3949 P2_R1164_U87 ; P2_R1164_U412
g19986 nand P2_R1164_U412 P2_R1164_U411 ; P2_R1164_U413
g19987 nand P2_R1164_U150 P2_R1164_U151 ; P2_R1164_U414
g19988 nand P2_R1164_U303 P2_R1164_U413 ; P2_R1164_U415
g19989 nand P2_U3055 P2_R1164_U46 ; P2_R1164_U416
g19990 nand P2_U3950 P2_R1164_U47 ; P2_R1164_U417
g19991 nand P2_U3055 P2_R1164_U46 ; P2_R1164_U418
g19992 nand P2_U3950 P2_R1164_U47 ; P2_R1164_U419
g19993 nand P2_R1164_U419 P2_R1164_U418 ; P2_R1164_U420
g19994 nand P2_R1164_U152 P2_R1164_U153 ; P2_R1164_U421
g19995 nand P2_R1164_U300 P2_R1164_U420 ; P2_R1164_U422
g19996 nand P2_U3059 P2_R1164_U49 ; P2_R1164_U423
g19997 nand P2_U3951 P2_R1164_U48 ; P2_R1164_U424
g19998 nand P2_U3060 P2_R1164_U50 ; P2_R1164_U425
g19999 nand P2_U3952 P2_R1164_U51 ; P2_R1164_U426
g20000 nand P2_R1164_U426 P2_R1164_U425 ; P2_R1164_U427
g20001 nand P2_R1164_U357 P2_R1164_U89 ; P2_R1164_U428
g20002 nand P2_R1164_U427 P2_R1164_U307 ; P2_R1164_U429
g20003 nand P2_U3067 P2_R1164_U52 ; P2_R1164_U430
g20004 nand P2_U3953 P2_R1164_U53 ; P2_R1164_U431
g20005 nand P2_R1164_U431 P2_R1164_U430 ; P2_R1164_U432
g20006 nand P2_R1164_U358 P2_R1164_U155 ; P2_R1164_U433
g20007 nand P2_R1164_U294 P2_R1164_U432 ; P2_R1164_U434
g20008 nand P2_U3068 P2_R1164_U84 ; P2_R1164_U435
g20009 nand P2_U3954 P2_R1164_U85 ; P2_R1164_U436
g20010 nand P2_U3068 P2_R1164_U84 ; P2_R1164_U437
g20011 nand P2_U3954 P2_R1164_U85 ; P2_R1164_U438
g20012 nand P2_R1164_U438 P2_R1164_U437 ; P2_R1164_U439
g20013 nand P2_R1164_U156 P2_R1164_U157 ; P2_R1164_U440
g20014 nand P2_R1164_U290 P2_R1164_U439 ; P2_R1164_U441
g20015 nand P2_U3063 P2_R1164_U82 ; P2_R1164_U442
g20016 nand P2_U3955 P2_R1164_U83 ; P2_R1164_U443
g20017 nand P2_U3063 P2_R1164_U82 ; P2_R1164_U444
g20018 nand P2_U3955 P2_R1164_U83 ; P2_R1164_U445
g20019 nand P2_R1164_U445 P2_R1164_U444 ; P2_R1164_U446
g20020 nand P2_R1164_U158 P2_R1164_U159 ; P2_R1164_U447
g20021 nand P2_R1164_U286 P2_R1164_U446 ; P2_R1164_U448
g20022 nand P2_U3077 P2_R1164_U54 ; P2_R1164_U449
g20023 nand P2_U3956 P2_R1164_U55 ; P2_R1164_U450
g20024 nand P2_U3077 P2_R1164_U54 ; P2_R1164_U451
g20025 nand P2_U3956 P2_R1164_U55 ; P2_R1164_U452
g20026 nand P2_R1164_U452 P2_R1164_U451 ; P2_R1164_U453
g20027 nand P2_U3078 P2_R1164_U81 ; P2_R1164_U454
g20028 nand P2_U3957 P2_R1164_U90 ; P2_R1164_U455
g20029 nand P2_R1164_U182 P2_R1164_U161 ; P2_R1164_U456
g20030 nand P2_R1164_U328 P2_R1164_U31 ; P2_R1164_U457
g20031 nand P2_U3083 P2_R1164_U78 ; P2_R1164_U458
g20032 nand P2_U3485 P2_R1164_U79 ; P2_R1164_U459
g20033 nand P2_R1164_U459 P2_R1164_U458 ; P2_R1164_U460
g20034 nand P2_R1164_U359 P2_R1164_U91 ; P2_R1164_U461
g20035 nand P2_R1164_U460 P2_R1164_U316 ; P2_R1164_U462
g20036 nand P2_U3084 P2_R1164_U75 ; P2_R1164_U463
g20037 nand P2_U3483 P2_R1164_U76 ; P2_R1164_U464
g20038 nand P2_R1164_U464 P2_R1164_U463 ; P2_R1164_U465
g20039 nand P2_R1164_U360 P2_R1164_U162 ; P2_R1164_U466
g20040 nand P2_R1164_U270 P2_R1164_U465 ; P2_R1164_U467
g20041 nand P2_U3071 P2_R1164_U60 ; P2_R1164_U468
g20042 nand P2_U3480 P2_R1164_U58 ; P2_R1164_U469
g20043 nand P2_U3075 P2_R1164_U56 ; P2_R1164_U470
g20044 nand P2_U3477 P2_R1164_U57 ; P2_R1164_U471
g20045 nand P2_R1164_U471 P2_R1164_U470 ; P2_R1164_U472
g20046 nand P2_R1164_U361 P2_R1164_U92 ; P2_R1164_U473
g20047 nand P2_R1164_U472 P2_R1164_U262 ; P2_R1164_U474
g20048 nand P2_U3076 P2_R1164_U73 ; P2_R1164_U475
g20049 nand P2_U3474 P2_R1164_U74 ; P2_R1164_U476
g20050 nand P2_U3076 P2_R1164_U73 ; P2_R1164_U477
g20051 nand P2_U3474 P2_R1164_U74 ; P2_R1164_U478
g20052 nand P2_R1164_U478 P2_R1164_U477 ; P2_R1164_U479
g20053 nand P2_R1164_U163 P2_R1164_U164 ; P2_R1164_U480
g20054 nand P2_R1164_U258 P2_R1164_U479 ; P2_R1164_U481
g20055 nand P2_U3081 P2_R1164_U71 ; P2_R1164_U482
g20056 nand P2_U3471 P2_R1164_U72 ; P2_R1164_U483
g20057 nand P2_U3081 P2_R1164_U71 ; P2_R1164_U484
g20058 nand P2_U3471 P2_R1164_U72 ; P2_R1164_U485
g20059 nand P2_R1164_U485 P2_R1164_U484 ; P2_R1164_U486
g20060 nand P2_R1164_U165 P2_R1164_U166 ; P2_R1164_U487
g20061 nand P2_R1164_U254 P2_R1164_U486 ; P2_R1164_U488
g20062 nand P2_U3082 P2_R1164_U69 ; P2_R1164_U489
g20063 nand P2_U3468 P2_R1164_U70 ; P2_R1164_U490
g20064 nand P2_U3074 P2_R1164_U64 ; P2_R1164_U491
g20065 nand P2_U3465 P2_R1164_U65 ; P2_R1164_U492
g20066 nand P2_R1164_U492 P2_R1164_U491 ; P2_R1164_U493
g20067 nand P2_R1164_U362 P2_R1164_U93 ; P2_R1164_U494
g20068 nand P2_R1164_U493 P2_R1164_U338 ; P2_R1164_U495
g20069 nand P2_U3065 P2_R1164_U66 ; P2_R1164_U496
g20070 nand P2_U3462 P2_R1164_U67 ; P2_R1164_U497
g20071 nand P2_R1164_U497 P2_R1164_U496 ; P2_R1164_U498
g20072 nand P2_R1164_U363 P2_R1164_U167 ; P2_R1164_U499
g20073 nand P2_R1164_U244 P2_R1164_U498 ; P2_R1164_U500
g20074 nand P2_U3064 P2_R1164_U62 ; P2_R1164_U501
g20075 nand P2_U3459 P2_R1164_U63 ; P2_R1164_U502
g20076 nand P2_U3079 P2_R1164_U29 ; P2_R1164_U503
g20077 nand P2_U3427 P2_R1164_U30 ; P2_R1164_U504
g20078 and P2_R1233_U179 P2_R1233_U178 ; P2_R1233_U4
g20079 and P2_R1233_U197 P2_R1233_U196 ; P2_R1233_U5
g20080 and P2_R1233_U237 P2_R1233_U236 ; P2_R1233_U6
g20081 and P2_R1233_U246 P2_R1233_U245 ; P2_R1233_U7
g20082 and P2_R1233_U264 P2_R1233_U263 ; P2_R1233_U8
g20083 and P2_R1233_U272 P2_R1233_U271 ; P2_R1233_U9
g20084 and P2_R1233_U351 P2_R1233_U348 ; P2_R1233_U10
g20085 and P2_R1233_U344 P2_R1233_U341 ; P2_R1233_U11
g20086 and P2_R1233_U335 P2_R1233_U332 ; P2_R1233_U12
g20087 and P2_R1233_U326 P2_R1233_U323 ; P2_R1233_U13
g20088 and P2_R1233_U320 P2_R1233_U318 ; P2_R1233_U14
g20089 and P2_R1233_U313 P2_R1233_U310 ; P2_R1233_U15
g20090 and P2_R1233_U235 P2_R1233_U232 ; P2_R1233_U16
g20091 and P2_R1233_U227 P2_R1233_U224 ; P2_R1233_U17
g20092 and P2_R1233_U213 P2_R1233_U210 ; P2_R1233_U18
g20093 not P2_U3447 ; P2_R1233_U19
g20094 not P2_U3073 ; P2_R1233_U20
g20095 not P2_U3072 ; P2_R1233_U21
g20096 nand P2_U3073 P2_U3447 ; P2_R1233_U22
g20097 not P2_U3450 ; P2_R1233_U23
g20098 not P2_U3441 ; P2_R1233_U24
g20099 not P2_U3062 ; P2_R1233_U25
g20100 not P2_U3069 ; P2_R1233_U26
g20101 not P2_U3435 ; P2_R1233_U27
g20102 not P2_U3070 ; P2_R1233_U28
g20103 not P2_U3427 ; P2_R1233_U29
g20104 not P2_U3079 ; P2_R1233_U30
g20105 nand P2_U3079 P2_U3427 ; P2_R1233_U31
g20106 not P2_U3438 ; P2_R1233_U32
g20107 not P2_U3066 ; P2_R1233_U33
g20108 nand P2_U3062 P2_U3441 ; P2_R1233_U34
g20109 not P2_U3444 ; P2_R1233_U35
g20110 not P2_U3453 ; P2_R1233_U36
g20111 not P2_U3086 ; P2_R1233_U37
g20112 not P2_U3085 ; P2_R1233_U38
g20113 not P2_U3456 ; P2_R1233_U39
g20114 nand P2_R1233_U61 P2_R1233_U205 ; P2_R1233_U40
g20115 nand P2_R1233_U117 P2_R1233_U193 ; P2_R1233_U41
g20116 nand P2_R1233_U182 P2_R1233_U183 ; P2_R1233_U42
g20117 nand P2_U3432 P2_U3080 ; P2_R1233_U43
g20118 nand P2_R1233_U122 P2_R1233_U219 ; P2_R1233_U44
g20119 nand P2_R1233_U216 P2_R1233_U215 ; P2_R1233_U45
g20120 not P2_U3950 ; P2_R1233_U46
g20121 not P2_U3055 ; P2_R1233_U47
g20122 not P2_U3059 ; P2_R1233_U48
g20123 not P2_U3951 ; P2_R1233_U49
g20124 not P2_U3952 ; P2_R1233_U50
g20125 not P2_U3060 ; P2_R1233_U51
g20126 not P2_U3953 ; P2_R1233_U52
g20127 not P2_U3067 ; P2_R1233_U53
g20128 not P2_U3956 ; P2_R1233_U54
g20129 not P2_U3077 ; P2_R1233_U55
g20130 not P2_U3477 ; P2_R1233_U56
g20131 not P2_U3075 ; P2_R1233_U57
g20132 not P2_U3071 ; P2_R1233_U58
g20133 nand P2_U3075 P2_U3477 ; P2_R1233_U59
g20134 not P2_U3480 ; P2_R1233_U60
g20135 nand P2_U3086 P2_U3453 ; P2_R1233_U61
g20136 not P2_U3459 ; P2_R1233_U62
g20137 not P2_U3064 ; P2_R1233_U63
g20138 not P2_U3465 ; P2_R1233_U64
g20139 not P2_U3074 ; P2_R1233_U65
g20140 not P2_U3462 ; P2_R1233_U66
g20141 not P2_U3065 ; P2_R1233_U67
g20142 nand P2_U3065 P2_U3462 ; P2_R1233_U68
g20143 not P2_U3468 ; P2_R1233_U69
g20144 not P2_U3082 ; P2_R1233_U70
g20145 not P2_U3471 ; P2_R1233_U71
g20146 not P2_U3081 ; P2_R1233_U72
g20147 not P2_U3474 ; P2_R1233_U73
g20148 not P2_U3076 ; P2_R1233_U74
g20149 not P2_U3483 ; P2_R1233_U75
g20150 not P2_U3084 ; P2_R1233_U76
g20151 nand P2_U3084 P2_U3483 ; P2_R1233_U77
g20152 not P2_U3485 ; P2_R1233_U78
g20153 not P2_U3083 ; P2_R1233_U79
g20154 nand P2_U3083 P2_U3485 ; P2_R1233_U80
g20155 not P2_U3957 ; P2_R1233_U81
g20156 not P2_U3955 ; P2_R1233_U82
g20157 not P2_U3063 ; P2_R1233_U83
g20158 not P2_U3954 ; P2_R1233_U84
g20159 not P2_U3068 ; P2_R1233_U85
g20160 nand P2_U3951 P2_U3059 ; P2_R1233_U86
g20161 not P2_U3056 ; P2_R1233_U87
g20162 not P2_U3949 ; P2_R1233_U88
g20163 nand P2_R1233_U306 P2_R1233_U176 ; P2_R1233_U89
g20164 not P2_U3078 ; P2_R1233_U90
g20165 nand P2_R1233_U77 P2_R1233_U315 ; P2_R1233_U91
g20166 nand P2_R1233_U261 P2_R1233_U260 ; P2_R1233_U92
g20167 nand P2_R1233_U68 P2_R1233_U337 ; P2_R1233_U93
g20168 nand P2_R1233_U457 P2_R1233_U456 ; P2_R1233_U94
g20169 nand P2_R1233_U504 P2_R1233_U503 ; P2_R1233_U95
g20170 nand P2_R1233_U375 P2_R1233_U374 ; P2_R1233_U96
g20171 nand P2_R1233_U380 P2_R1233_U379 ; P2_R1233_U97
g20172 nand P2_R1233_U387 P2_R1233_U386 ; P2_R1233_U98
g20173 nand P2_R1233_U394 P2_R1233_U393 ; P2_R1233_U99
g20174 nand P2_R1233_U399 P2_R1233_U398 ; P2_R1233_U100
g20175 nand P2_R1233_U408 P2_R1233_U407 ; P2_R1233_U101
g20176 nand P2_R1233_U415 P2_R1233_U414 ; P2_R1233_U102
g20177 nand P2_R1233_U422 P2_R1233_U421 ; P2_R1233_U103
g20178 nand P2_R1233_U429 P2_R1233_U428 ; P2_R1233_U104
g20179 nand P2_R1233_U434 P2_R1233_U433 ; P2_R1233_U105
g20180 nand P2_R1233_U441 P2_R1233_U440 ; P2_R1233_U106
g20181 nand P2_R1233_U448 P2_R1233_U447 ; P2_R1233_U107
g20182 nand P2_R1233_U462 P2_R1233_U461 ; P2_R1233_U108
g20183 nand P2_R1233_U467 P2_R1233_U466 ; P2_R1233_U109
g20184 nand P2_R1233_U474 P2_R1233_U473 ; P2_R1233_U110
g20185 nand P2_R1233_U481 P2_R1233_U480 ; P2_R1233_U111
g20186 nand P2_R1233_U488 P2_R1233_U487 ; P2_R1233_U112
g20187 nand P2_R1233_U495 P2_R1233_U494 ; P2_R1233_U113
g20188 nand P2_R1233_U500 P2_R1233_U499 ; P2_R1233_U114
g20189 and P2_R1233_U189 P2_R1233_U187 ; P2_R1233_U115
g20190 and P2_R1233_U4 P2_R1233_U180 ; P2_R1233_U116
g20191 and P2_R1233_U194 P2_R1233_U192 ; P2_R1233_U117
g20192 and P2_R1233_U201 P2_R1233_U200 ; P2_R1233_U118
g20193 and P2_R1233_U382 P2_R1233_U381 P2_R1233_U22 ; P2_R1233_U119
g20194 and P2_R1233_U212 P2_R1233_U5 ; P2_R1233_U120
g20195 and P2_R1233_U181 P2_R1233_U180 ; P2_R1233_U121
g20196 and P2_R1233_U220 P2_R1233_U218 ; P2_R1233_U122
g20197 and P2_R1233_U389 P2_R1233_U388 P2_R1233_U34 ; P2_R1233_U123
g20198 and P2_R1233_U226 P2_R1233_U4 ; P2_R1233_U124
g20199 and P2_R1233_U234 P2_R1233_U181 ; P2_R1233_U125
g20200 and P2_R1233_U204 P2_R1233_U6 ; P2_R1233_U126
g20201 and P2_R1233_U239 P2_R1233_U171 ; P2_R1233_U127
g20202 and P2_R1233_U250 P2_R1233_U7 ; P2_R1233_U128
g20203 and P2_R1233_U248 P2_R1233_U172 ; P2_R1233_U129
g20204 and P2_R1233_U268 P2_R1233_U267 ; P2_R1233_U130
g20205 and P2_R1233_U9 P2_R1233_U282 ; P2_R1233_U131
g20206 and P2_R1233_U285 P2_R1233_U280 ; P2_R1233_U132
g20207 and P2_R1233_U301 P2_R1233_U298 ; P2_R1233_U133
g20208 and P2_R1233_U368 P2_R1233_U302 ; P2_R1233_U134
g20209 and P2_R1233_U160 P2_R1233_U278 ; P2_R1233_U135
g20210 and P2_R1233_U455 P2_R1233_U454 P2_R1233_U80 ; P2_R1233_U136
g20211 and P2_R1233_U325 P2_R1233_U9 ; P2_R1233_U137
g20212 and P2_R1233_U469 P2_R1233_U468 P2_R1233_U59 ; P2_R1233_U138
g20213 and P2_R1233_U334 P2_R1233_U8 ; P2_R1233_U139
g20214 and P2_R1233_U490 P2_R1233_U489 P2_R1233_U172 ; P2_R1233_U140
g20215 and P2_R1233_U343 P2_R1233_U7 ; P2_R1233_U141
g20216 and P2_R1233_U502 P2_R1233_U501 P2_R1233_U171 ; P2_R1233_U142
g20217 and P2_R1233_U350 P2_R1233_U6 ; P2_R1233_U143
g20218 nand P2_R1233_U118 P2_R1233_U202 ; P2_R1233_U144
g20219 nand P2_R1233_U217 P2_R1233_U229 ; P2_R1233_U145
g20220 not P2_U3057 ; P2_R1233_U146
g20221 not P2_U3960 ; P2_R1233_U147
g20222 and P2_R1233_U403 P2_R1233_U402 ; P2_R1233_U148
g20223 nand P2_R1233_U304 P2_R1233_U169 P2_R1233_U364 ; P2_R1233_U149
g20224 and P2_R1233_U410 P2_R1233_U409 ; P2_R1233_U150
g20225 nand P2_R1233_U370 P2_R1233_U369 P2_R1233_U134 ; P2_R1233_U151
g20226 and P2_R1233_U417 P2_R1233_U416 ; P2_R1233_U152
g20227 nand P2_R1233_U365 P2_R1233_U299 P2_R1233_U86 ; P2_R1233_U153
g20228 and P2_R1233_U424 P2_R1233_U423 ; P2_R1233_U154
g20229 nand P2_R1233_U293 P2_R1233_U292 ; P2_R1233_U155
g20230 and P2_R1233_U436 P2_R1233_U435 ; P2_R1233_U156
g20231 nand P2_R1233_U289 P2_R1233_U288 ; P2_R1233_U157
g20232 and P2_R1233_U443 P2_R1233_U442 ; P2_R1233_U158
g20233 nand P2_R1233_U132 P2_R1233_U284 ; P2_R1233_U159
g20234 and P2_R1233_U450 P2_R1233_U449 ; P2_R1233_U160
g20235 nand P2_R1233_U43 P2_R1233_U327 ; P2_R1233_U161
g20236 nand P2_R1233_U130 P2_R1233_U269 ; P2_R1233_U162
g20237 and P2_R1233_U476 P2_R1233_U475 ; P2_R1233_U163
g20238 nand P2_R1233_U257 P2_R1233_U256 ; P2_R1233_U164
g20239 and P2_R1233_U483 P2_R1233_U482 ; P2_R1233_U165
g20240 nand P2_R1233_U253 P2_R1233_U252 ; P2_R1233_U166
g20241 nand P2_R1233_U243 P2_R1233_U242 ; P2_R1233_U167
g20242 nand P2_R1233_U367 P2_R1233_U366 ; P2_R1233_U168
g20243 nand P2_U3056 P2_R1233_U151 ; P2_R1233_U169
g20244 not P2_R1233_U34 ; P2_R1233_U170
g20245 nand P2_U3456 P2_U3085 ; P2_R1233_U171
g20246 nand P2_U3074 P2_U3465 ; P2_R1233_U172
g20247 nand P2_U3060 P2_U3952 ; P2_R1233_U173
g20248 not P2_R1233_U68 ; P2_R1233_U174
g20249 not P2_R1233_U77 ; P2_R1233_U175
g20250 nand P2_U3067 P2_U3953 ; P2_R1233_U176
g20251 not P2_R1233_U61 ; P2_R1233_U177
g20252 or P2_U3069 P2_U3444 ; P2_R1233_U178
g20253 or P2_U3062 P2_U3441 ; P2_R1233_U179
g20254 or P2_U3438 P2_U3066 ; P2_R1233_U180
g20255 or P2_U3435 P2_U3070 ; P2_R1233_U181
g20256 not P2_R1233_U31 ; P2_R1233_U182
g20257 or P2_U3432 P2_U3080 ; P2_R1233_U183
g20258 not P2_R1233_U42 ; P2_R1233_U184
g20259 not P2_R1233_U43 ; P2_R1233_U185
g20260 nand P2_R1233_U42 P2_R1233_U43 ; P2_R1233_U186
g20261 nand P2_U3070 P2_U3435 ; P2_R1233_U187
g20262 nand P2_R1233_U186 P2_R1233_U181 ; P2_R1233_U188
g20263 nand P2_U3066 P2_U3438 ; P2_R1233_U189
g20264 nand P2_R1233_U115 P2_R1233_U188 ; P2_R1233_U190
g20265 nand P2_R1233_U35 P2_R1233_U34 ; P2_R1233_U191
g20266 nand P2_U3069 P2_R1233_U191 ; P2_R1233_U192
g20267 nand P2_R1233_U116 P2_R1233_U190 ; P2_R1233_U193
g20268 nand P2_U3444 P2_R1233_U170 ; P2_R1233_U194
g20269 not P2_R1233_U41 ; P2_R1233_U195
g20270 or P2_U3072 P2_U3450 ; P2_R1233_U196
g20271 or P2_U3073 P2_U3447 ; P2_R1233_U197
g20272 not P2_R1233_U22 ; P2_R1233_U198
g20273 nand P2_R1233_U23 P2_R1233_U22 ; P2_R1233_U199
g20274 nand P2_U3072 P2_R1233_U199 ; P2_R1233_U200
g20275 nand P2_U3450 P2_R1233_U198 ; P2_R1233_U201
g20276 nand P2_R1233_U5 P2_R1233_U41 ; P2_R1233_U202
g20277 not P2_R1233_U144 ; P2_R1233_U203
g20278 or P2_U3453 P2_U3086 ; P2_R1233_U204
g20279 nand P2_R1233_U204 P2_R1233_U144 ; P2_R1233_U205
g20280 not P2_R1233_U40 ; P2_R1233_U206
g20281 or P2_U3085 P2_U3456 ; P2_R1233_U207
g20282 or P2_U3447 P2_U3073 ; P2_R1233_U208
g20283 nand P2_R1233_U208 P2_R1233_U41 ; P2_R1233_U209
g20284 nand P2_R1233_U119 P2_R1233_U209 ; P2_R1233_U210
g20285 nand P2_R1233_U195 P2_R1233_U22 ; P2_R1233_U211
g20286 nand P2_U3450 P2_U3072 ; P2_R1233_U212
g20287 nand P2_R1233_U120 P2_R1233_U211 ; P2_R1233_U213
g20288 or P2_U3073 P2_U3447 ; P2_R1233_U214
g20289 nand P2_R1233_U185 P2_R1233_U181 ; P2_R1233_U215
g20290 nand P2_U3070 P2_U3435 ; P2_R1233_U216
g20291 not P2_R1233_U45 ; P2_R1233_U217
g20292 nand P2_R1233_U121 P2_R1233_U184 ; P2_R1233_U218
g20293 nand P2_R1233_U45 P2_R1233_U180 ; P2_R1233_U219
g20294 nand P2_U3066 P2_U3438 ; P2_R1233_U220
g20295 not P2_R1233_U44 ; P2_R1233_U221
g20296 or P2_U3441 P2_U3062 ; P2_R1233_U222
g20297 nand P2_R1233_U222 P2_R1233_U44 ; P2_R1233_U223
g20298 nand P2_R1233_U123 P2_R1233_U223 ; P2_R1233_U224
g20299 nand P2_R1233_U221 P2_R1233_U34 ; P2_R1233_U225
g20300 nand P2_U3444 P2_U3069 ; P2_R1233_U226
g20301 nand P2_R1233_U124 P2_R1233_U225 ; P2_R1233_U227
g20302 or P2_U3062 P2_U3441 ; P2_R1233_U228
g20303 nand P2_R1233_U184 P2_R1233_U181 ; P2_R1233_U229
g20304 not P2_R1233_U145 ; P2_R1233_U230
g20305 nand P2_U3066 P2_U3438 ; P2_R1233_U231
g20306 nand P2_R1233_U401 P2_R1233_U400 P2_R1233_U43 P2_R1233_U42 ; P2_R1233_U232
g20307 nand P2_R1233_U43 P2_R1233_U42 ; P2_R1233_U233
g20308 nand P2_U3070 P2_U3435 ; P2_R1233_U234
g20309 nand P2_R1233_U125 P2_R1233_U233 ; P2_R1233_U235
g20310 or P2_U3085 P2_U3456 ; P2_R1233_U236
g20311 or P2_U3064 P2_U3459 ; P2_R1233_U237
g20312 nand P2_R1233_U177 P2_R1233_U6 ; P2_R1233_U238
g20313 nand P2_U3064 P2_U3459 ; P2_R1233_U239
g20314 nand P2_R1233_U127 P2_R1233_U238 ; P2_R1233_U240
g20315 or P2_U3459 P2_U3064 ; P2_R1233_U241
g20316 nand P2_R1233_U126 P2_R1233_U144 ; P2_R1233_U242
g20317 nand P2_R1233_U241 P2_R1233_U240 ; P2_R1233_U243
g20318 not P2_R1233_U167 ; P2_R1233_U244
g20319 or P2_U3082 P2_U3468 ; P2_R1233_U245
g20320 or P2_U3074 P2_U3465 ; P2_R1233_U246
g20321 nand P2_R1233_U174 P2_R1233_U7 ; P2_R1233_U247
g20322 nand P2_U3082 P2_U3468 ; P2_R1233_U248
g20323 nand P2_R1233_U129 P2_R1233_U247 ; P2_R1233_U249
g20324 or P2_U3462 P2_U3065 ; P2_R1233_U250
g20325 or P2_U3468 P2_U3082 ; P2_R1233_U251
g20326 nand P2_R1233_U128 P2_R1233_U167 ; P2_R1233_U252
g20327 nand P2_R1233_U251 P2_R1233_U249 ; P2_R1233_U253
g20328 not P2_R1233_U166 ; P2_R1233_U254
g20329 or P2_U3471 P2_U3081 ; P2_R1233_U255
g20330 nand P2_R1233_U255 P2_R1233_U166 ; P2_R1233_U256
g20331 nand P2_U3081 P2_U3471 ; P2_R1233_U257
g20332 not P2_R1233_U164 ; P2_R1233_U258
g20333 or P2_U3474 P2_U3076 ; P2_R1233_U259
g20334 nand P2_R1233_U259 P2_R1233_U164 ; P2_R1233_U260
g20335 nand P2_U3076 P2_U3474 ; P2_R1233_U261
g20336 not P2_R1233_U92 ; P2_R1233_U262
g20337 or P2_U3071 P2_U3480 ; P2_R1233_U263
g20338 or P2_U3075 P2_U3477 ; P2_R1233_U264
g20339 not P2_R1233_U59 ; P2_R1233_U265
g20340 nand P2_R1233_U60 P2_R1233_U59 ; P2_R1233_U266
g20341 nand P2_U3071 P2_R1233_U266 ; P2_R1233_U267
g20342 nand P2_U3480 P2_R1233_U265 ; P2_R1233_U268
g20343 nand P2_R1233_U8 P2_R1233_U92 ; P2_R1233_U269
g20344 not P2_R1233_U162 ; P2_R1233_U270
g20345 or P2_U3078 P2_U3957 ; P2_R1233_U271
g20346 or P2_U3083 P2_U3485 ; P2_R1233_U272
g20347 or P2_U3077 P2_U3956 ; P2_R1233_U273
g20348 not P2_R1233_U80 ; P2_R1233_U274
g20349 nand P2_U3957 P2_R1233_U274 ; P2_R1233_U275
g20350 nand P2_R1233_U275 P2_R1233_U90 ; P2_R1233_U276
g20351 nand P2_R1233_U80 P2_R1233_U81 ; P2_R1233_U277
g20352 nand P2_R1233_U277 P2_R1233_U276 ; P2_R1233_U278
g20353 nand P2_R1233_U175 P2_R1233_U9 ; P2_R1233_U279
g20354 nand P2_U3077 P2_U3956 ; P2_R1233_U280
g20355 nand P2_R1233_U278 P2_R1233_U279 ; P2_R1233_U281
g20356 or P2_U3483 P2_U3084 ; P2_R1233_U282
g20357 or P2_U3956 P2_U3077 ; P2_R1233_U283
g20358 nand P2_R1233_U273 P2_R1233_U162 P2_R1233_U131 ; P2_R1233_U284
g20359 nand P2_R1233_U283 P2_R1233_U281 ; P2_R1233_U285
g20360 not P2_R1233_U159 ; P2_R1233_U286
g20361 or P2_U3955 P2_U3063 ; P2_R1233_U287
g20362 nand P2_R1233_U287 P2_R1233_U159 ; P2_R1233_U288
g20363 nand P2_U3063 P2_U3955 ; P2_R1233_U289
g20364 not P2_R1233_U157 ; P2_R1233_U290
g20365 or P2_U3954 P2_U3068 ; P2_R1233_U291
g20366 nand P2_R1233_U291 P2_R1233_U157 ; P2_R1233_U292
g20367 nand P2_U3068 P2_U3954 ; P2_R1233_U293
g20368 not P2_R1233_U155 ; P2_R1233_U294
g20369 or P2_U3060 P2_U3952 ; P2_R1233_U295
g20370 nand P2_R1233_U176 P2_R1233_U173 ; P2_R1233_U296
g20371 not P2_R1233_U86 ; P2_R1233_U297
g20372 or P2_U3953 P2_U3067 ; P2_R1233_U298
g20373 nand P2_R1233_U155 P2_R1233_U298 P2_R1233_U168 ; P2_R1233_U299
g20374 not P2_R1233_U153 ; P2_R1233_U300
g20375 or P2_U3950 P2_U3055 ; P2_R1233_U301
g20376 nand P2_U3055 P2_U3950 ; P2_R1233_U302
g20377 not P2_R1233_U151 ; P2_R1233_U303
g20378 nand P2_U3949 P2_R1233_U151 ; P2_R1233_U304
g20379 not P2_R1233_U149 ; P2_R1233_U305
g20380 nand P2_R1233_U298 P2_R1233_U155 ; P2_R1233_U306
g20381 not P2_R1233_U89 ; P2_R1233_U307
g20382 or P2_U3952 P2_U3060 ; P2_R1233_U308
g20383 nand P2_R1233_U308 P2_R1233_U89 ; P2_R1233_U309
g20384 nand P2_R1233_U309 P2_R1233_U173 P2_R1233_U154 ; P2_R1233_U310
g20385 nand P2_R1233_U307 P2_R1233_U173 ; P2_R1233_U311
g20386 nand P2_U3951 P2_U3059 ; P2_R1233_U312
g20387 nand P2_R1233_U311 P2_R1233_U312 P2_R1233_U168 ; P2_R1233_U313
g20388 or P2_U3060 P2_U3952 ; P2_R1233_U314
g20389 nand P2_R1233_U282 P2_R1233_U162 ; P2_R1233_U315
g20390 not P2_R1233_U91 ; P2_R1233_U316
g20391 nand P2_R1233_U9 P2_R1233_U91 ; P2_R1233_U317
g20392 nand P2_R1233_U135 P2_R1233_U317 ; P2_R1233_U318
g20393 nand P2_R1233_U317 P2_R1233_U278 ; P2_R1233_U319
g20394 nand P2_R1233_U453 P2_R1233_U319 ; P2_R1233_U320
g20395 or P2_U3485 P2_U3083 ; P2_R1233_U321
g20396 nand P2_R1233_U321 P2_R1233_U91 ; P2_R1233_U322
g20397 nand P2_R1233_U136 P2_R1233_U322 ; P2_R1233_U323
g20398 nand P2_R1233_U316 P2_R1233_U80 ; P2_R1233_U324
g20399 nand P2_U3078 P2_U3957 ; P2_R1233_U325
g20400 nand P2_R1233_U137 P2_R1233_U324 ; P2_R1233_U326
g20401 or P2_U3432 P2_U3080 ; P2_R1233_U327
g20402 not P2_R1233_U161 ; P2_R1233_U328
g20403 or P2_U3083 P2_U3485 ; P2_R1233_U329
g20404 or P2_U3477 P2_U3075 ; P2_R1233_U330
g20405 nand P2_R1233_U330 P2_R1233_U92 ; P2_R1233_U331
g20406 nand P2_R1233_U138 P2_R1233_U331 ; P2_R1233_U332
g20407 nand P2_R1233_U262 P2_R1233_U59 ; P2_R1233_U333
g20408 nand P2_U3480 P2_U3071 ; P2_R1233_U334
g20409 nand P2_R1233_U139 P2_R1233_U333 ; P2_R1233_U335
g20410 or P2_U3075 P2_U3477 ; P2_R1233_U336
g20411 nand P2_R1233_U250 P2_R1233_U167 ; P2_R1233_U337
g20412 not P2_R1233_U93 ; P2_R1233_U338
g20413 or P2_U3465 P2_U3074 ; P2_R1233_U339
g20414 nand P2_R1233_U339 P2_R1233_U93 ; P2_R1233_U340
g20415 nand P2_R1233_U140 P2_R1233_U340 ; P2_R1233_U341
g20416 nand P2_R1233_U338 P2_R1233_U172 ; P2_R1233_U342
g20417 nand P2_U3082 P2_U3468 ; P2_R1233_U343
g20418 nand P2_R1233_U141 P2_R1233_U342 ; P2_R1233_U344
g20419 or P2_U3074 P2_U3465 ; P2_R1233_U345
g20420 or P2_U3456 P2_U3085 ; P2_R1233_U346
g20421 nand P2_R1233_U346 P2_R1233_U40 ; P2_R1233_U347
g20422 nand P2_R1233_U142 P2_R1233_U347 ; P2_R1233_U348
g20423 nand P2_R1233_U206 P2_R1233_U171 ; P2_R1233_U349
g20424 nand P2_U3064 P2_U3459 ; P2_R1233_U350
g20425 nand P2_R1233_U143 P2_R1233_U349 ; P2_R1233_U351
g20426 nand P2_R1233_U207 P2_R1233_U171 ; P2_R1233_U352
g20427 nand P2_R1233_U204 P2_R1233_U61 ; P2_R1233_U353
g20428 nand P2_R1233_U214 P2_R1233_U22 ; P2_R1233_U354
g20429 nand P2_R1233_U228 P2_R1233_U34 ; P2_R1233_U355
g20430 nand P2_R1233_U231 P2_R1233_U180 ; P2_R1233_U356
g20431 nand P2_R1233_U314 P2_R1233_U173 ; P2_R1233_U357
g20432 nand P2_R1233_U298 P2_R1233_U176 ; P2_R1233_U358
g20433 nand P2_R1233_U329 P2_R1233_U80 ; P2_R1233_U359
g20434 nand P2_R1233_U282 P2_R1233_U77 ; P2_R1233_U360
g20435 nand P2_R1233_U336 P2_R1233_U59 ; P2_R1233_U361
g20436 nand P2_R1233_U345 P2_R1233_U172 ; P2_R1233_U362
g20437 nand P2_R1233_U250 P2_R1233_U68 ; P2_R1233_U363
g20438 nand P2_U3949 P2_U3056 ; P2_R1233_U364
g20439 nand P2_R1233_U296 P2_R1233_U168 ; P2_R1233_U365
g20440 nand P2_U3059 P2_R1233_U295 ; P2_R1233_U366
g20441 nand P2_U3951 P2_R1233_U295 ; P2_R1233_U367
g20442 nand P2_R1233_U296 P2_R1233_U168 P2_R1233_U301 ; P2_R1233_U368
g20443 nand P2_R1233_U155 P2_R1233_U168 P2_R1233_U133 ; P2_R1233_U369
g20444 nand P2_R1233_U297 P2_R1233_U301 ; P2_R1233_U370
g20445 nand P2_U3085 P2_R1233_U39 ; P2_R1233_U371
g20446 nand P2_U3456 P2_R1233_U38 ; P2_R1233_U372
g20447 nand P2_R1233_U372 P2_R1233_U371 ; P2_R1233_U373
g20448 nand P2_R1233_U352 P2_R1233_U40 ; P2_R1233_U374
g20449 nand P2_R1233_U373 P2_R1233_U206 ; P2_R1233_U375
g20450 nand P2_U3086 P2_R1233_U36 ; P2_R1233_U376
g20451 nand P2_U3453 P2_R1233_U37 ; P2_R1233_U377
g20452 nand P2_R1233_U377 P2_R1233_U376 ; P2_R1233_U378
g20453 nand P2_R1233_U353 P2_R1233_U144 ; P2_R1233_U379
g20454 nand P2_R1233_U203 P2_R1233_U378 ; P2_R1233_U380
g20455 nand P2_U3072 P2_R1233_U23 ; P2_R1233_U381
g20456 nand P2_U3450 P2_R1233_U21 ; P2_R1233_U382
g20457 nand P2_U3073 P2_R1233_U19 ; P2_R1233_U383
g20458 nand P2_U3447 P2_R1233_U20 ; P2_R1233_U384
g20459 nand P2_R1233_U384 P2_R1233_U383 ; P2_R1233_U385
g20460 nand P2_R1233_U354 P2_R1233_U41 ; P2_R1233_U386
g20461 nand P2_R1233_U385 P2_R1233_U195 ; P2_R1233_U387
g20462 nand P2_U3069 P2_R1233_U35 ; P2_R1233_U388
g20463 nand P2_U3444 P2_R1233_U26 ; P2_R1233_U389
g20464 nand P2_U3062 P2_R1233_U24 ; P2_R1233_U390
g20465 nand P2_U3441 P2_R1233_U25 ; P2_R1233_U391
g20466 nand P2_R1233_U391 P2_R1233_U390 ; P2_R1233_U392
g20467 nand P2_R1233_U355 P2_R1233_U44 ; P2_R1233_U393
g20468 nand P2_R1233_U392 P2_R1233_U221 ; P2_R1233_U394
g20469 nand P2_U3066 P2_R1233_U32 ; P2_R1233_U395
g20470 nand P2_U3438 P2_R1233_U33 ; P2_R1233_U396
g20471 nand P2_R1233_U396 P2_R1233_U395 ; P2_R1233_U397
g20472 nand P2_R1233_U356 P2_R1233_U145 ; P2_R1233_U398
g20473 nand P2_R1233_U230 P2_R1233_U397 ; P2_R1233_U399
g20474 nand P2_U3070 P2_R1233_U27 ; P2_R1233_U400
g20475 nand P2_U3435 P2_R1233_U28 ; P2_R1233_U401
g20476 nand P2_U3057 P2_R1233_U147 ; P2_R1233_U402
g20477 nand P2_U3960 P2_R1233_U146 ; P2_R1233_U403
g20478 nand P2_U3057 P2_R1233_U147 ; P2_R1233_U404
g20479 nand P2_U3960 P2_R1233_U146 ; P2_R1233_U405
g20480 nand P2_R1233_U405 P2_R1233_U404 ; P2_R1233_U406
g20481 nand P2_R1233_U148 P2_R1233_U149 ; P2_R1233_U407
g20482 nand P2_R1233_U305 P2_R1233_U406 ; P2_R1233_U408
g20483 nand P2_U3056 P2_R1233_U88 ; P2_R1233_U409
g20484 nand P2_U3949 P2_R1233_U87 ; P2_R1233_U410
g20485 nand P2_U3056 P2_R1233_U88 ; P2_R1233_U411
g20486 nand P2_U3949 P2_R1233_U87 ; P2_R1233_U412
g20487 nand P2_R1233_U412 P2_R1233_U411 ; P2_R1233_U413
g20488 nand P2_R1233_U150 P2_R1233_U151 ; P2_R1233_U414
g20489 nand P2_R1233_U303 P2_R1233_U413 ; P2_R1233_U415
g20490 nand P2_U3055 P2_R1233_U46 ; P2_R1233_U416
g20491 nand P2_U3950 P2_R1233_U47 ; P2_R1233_U417
g20492 nand P2_U3055 P2_R1233_U46 ; P2_R1233_U418
g20493 nand P2_U3950 P2_R1233_U47 ; P2_R1233_U419
g20494 nand P2_R1233_U419 P2_R1233_U418 ; P2_R1233_U420
g20495 nand P2_R1233_U152 P2_R1233_U153 ; P2_R1233_U421
g20496 nand P2_R1233_U300 P2_R1233_U420 ; P2_R1233_U422
g20497 nand P2_U3059 P2_R1233_U49 ; P2_R1233_U423
g20498 nand P2_U3951 P2_R1233_U48 ; P2_R1233_U424
g20499 nand P2_U3060 P2_R1233_U50 ; P2_R1233_U425
g20500 nand P2_U3952 P2_R1233_U51 ; P2_R1233_U426
g20501 nand P2_R1233_U426 P2_R1233_U425 ; P2_R1233_U427
g20502 nand P2_R1233_U357 P2_R1233_U89 ; P2_R1233_U428
g20503 nand P2_R1233_U427 P2_R1233_U307 ; P2_R1233_U429
g20504 nand P2_U3067 P2_R1233_U52 ; P2_R1233_U430
g20505 nand P2_U3953 P2_R1233_U53 ; P2_R1233_U431
g20506 nand P2_R1233_U431 P2_R1233_U430 ; P2_R1233_U432
g20507 nand P2_R1233_U358 P2_R1233_U155 ; P2_R1233_U433
g20508 nand P2_R1233_U294 P2_R1233_U432 ; P2_R1233_U434
g20509 nand P2_U3068 P2_R1233_U84 ; P2_R1233_U435
g20510 nand P2_U3954 P2_R1233_U85 ; P2_R1233_U436
g20511 nand P2_U3068 P2_R1233_U84 ; P2_R1233_U437
g20512 nand P2_U3954 P2_R1233_U85 ; P2_R1233_U438
g20513 nand P2_R1233_U438 P2_R1233_U437 ; P2_R1233_U439
g20514 nand P2_R1233_U156 P2_R1233_U157 ; P2_R1233_U440
g20515 nand P2_R1233_U290 P2_R1233_U439 ; P2_R1233_U441
g20516 nand P2_U3063 P2_R1233_U82 ; P2_R1233_U442
g20517 nand P2_U3955 P2_R1233_U83 ; P2_R1233_U443
g20518 nand P2_U3063 P2_R1233_U82 ; P2_R1233_U444
g20519 nand P2_U3955 P2_R1233_U83 ; P2_R1233_U445
g20520 nand P2_R1233_U445 P2_R1233_U444 ; P2_R1233_U446
g20521 nand P2_R1233_U158 P2_R1233_U159 ; P2_R1233_U447
g20522 nand P2_R1233_U286 P2_R1233_U446 ; P2_R1233_U448
g20523 nand P2_U3077 P2_R1233_U54 ; P2_R1233_U449
g20524 nand P2_U3956 P2_R1233_U55 ; P2_R1233_U450
g20525 nand P2_U3077 P2_R1233_U54 ; P2_R1233_U451
g20526 nand P2_U3956 P2_R1233_U55 ; P2_R1233_U452
g20527 nand P2_R1233_U452 P2_R1233_U451 ; P2_R1233_U453
g20528 nand P2_U3078 P2_R1233_U81 ; P2_R1233_U454
g20529 nand P2_U3957 P2_R1233_U90 ; P2_R1233_U455
g20530 nand P2_R1233_U182 P2_R1233_U161 ; P2_R1233_U456
g20531 nand P2_R1233_U328 P2_R1233_U31 ; P2_R1233_U457
g20532 nand P2_U3083 P2_R1233_U78 ; P2_R1233_U458
g20533 nand P2_U3485 P2_R1233_U79 ; P2_R1233_U459
g20534 nand P2_R1233_U459 P2_R1233_U458 ; P2_R1233_U460
g20535 nand P2_R1233_U359 P2_R1233_U91 ; P2_R1233_U461
g20536 nand P2_R1233_U460 P2_R1233_U316 ; P2_R1233_U462
g20537 nand P2_U3084 P2_R1233_U75 ; P2_R1233_U463
g20538 nand P2_U3483 P2_R1233_U76 ; P2_R1233_U464
g20539 nand P2_R1233_U464 P2_R1233_U463 ; P2_R1233_U465
g20540 nand P2_R1233_U360 P2_R1233_U162 ; P2_R1233_U466
g20541 nand P2_R1233_U270 P2_R1233_U465 ; P2_R1233_U467
g20542 nand P2_U3071 P2_R1233_U60 ; P2_R1233_U468
g20543 nand P2_U3480 P2_R1233_U58 ; P2_R1233_U469
g20544 nand P2_U3075 P2_R1233_U56 ; P2_R1233_U470
g20545 nand P2_U3477 P2_R1233_U57 ; P2_R1233_U471
g20546 nand P2_R1233_U471 P2_R1233_U470 ; P2_R1233_U472
g20547 nand P2_R1233_U361 P2_R1233_U92 ; P2_R1233_U473
g20548 nand P2_R1233_U472 P2_R1233_U262 ; P2_R1233_U474
g20549 nand P2_U3076 P2_R1233_U73 ; P2_R1233_U475
g20550 nand P2_U3474 P2_R1233_U74 ; P2_R1233_U476
g20551 nand P2_U3076 P2_R1233_U73 ; P2_R1233_U477
g20552 nand P2_U3474 P2_R1233_U74 ; P2_R1233_U478
g20553 nand P2_R1233_U478 P2_R1233_U477 ; P2_R1233_U479
g20554 nand P2_R1233_U163 P2_R1233_U164 ; P2_R1233_U480
g20555 nand P2_R1233_U258 P2_R1233_U479 ; P2_R1233_U481
g20556 nand P2_U3081 P2_R1233_U71 ; P2_R1233_U482
g20557 nand P2_U3471 P2_R1233_U72 ; P2_R1233_U483
g20558 nand P2_U3081 P2_R1233_U71 ; P2_R1233_U484
g20559 nand P2_U3471 P2_R1233_U72 ; P2_R1233_U485
g20560 nand P2_R1233_U485 P2_R1233_U484 ; P2_R1233_U486
g20561 nand P2_R1233_U165 P2_R1233_U166 ; P2_R1233_U487
g20562 nand P2_R1233_U254 P2_R1233_U486 ; P2_R1233_U488
g20563 nand P2_U3082 P2_R1233_U69 ; P2_R1233_U489
g20564 nand P2_U3468 P2_R1233_U70 ; P2_R1233_U490
g20565 nand P2_U3074 P2_R1233_U64 ; P2_R1233_U491
g20566 nand P2_U3465 P2_R1233_U65 ; P2_R1233_U492
g20567 nand P2_R1233_U492 P2_R1233_U491 ; P2_R1233_U493
g20568 nand P2_R1233_U362 P2_R1233_U93 ; P2_R1233_U494
g20569 nand P2_R1233_U493 P2_R1233_U338 ; P2_R1233_U495
g20570 nand P2_U3065 P2_R1233_U66 ; P2_R1233_U496
g20571 nand P2_U3462 P2_R1233_U67 ; P2_R1233_U497
g20572 nand P2_R1233_U497 P2_R1233_U496 ; P2_R1233_U498
g20573 nand P2_R1233_U363 P2_R1233_U167 ; P2_R1233_U499
g20574 nand P2_R1233_U244 P2_R1233_U498 ; P2_R1233_U500
g20575 nand P2_U3064 P2_R1233_U62 ; P2_R1233_U501
g20576 nand P2_U3459 P2_R1233_U63 ; P2_R1233_U502
g20577 nand P2_U3079 P2_R1233_U29 ; P2_R1233_U503
g20578 nand P2_U3427 P2_R1233_U30 ; P2_R1233_U504
g20579 and P2_R1176_U221 P2_R1176_U220 ; P2_R1176_U4
g20580 and P2_R1176_U234 P2_R1176_U233 ; P2_R1176_U5
g20581 and P2_R1176_U264 P2_R1176_U263 ; P2_R1176_U6
g20582 and P2_R1176_U280 P2_R1176_U279 ; P2_R1176_U7
g20583 and P2_R1176_U292 P2_R1176_U291 ; P2_R1176_U8
g20584 and P2_R1176_U6 P2_R1176_U268 ; P2_R1176_U9
g20585 and P2_R1176_U5 P2_R1176_U229 ; P2_R1176_U10
g20586 and P2_R1176_U9 P2_R1176_U259 ; P2_R1176_U11
g20587 and P2_R1176_U528 P2_R1176_U527 ; P2_R1176_U12
g20588 and P2_R1176_U351 P2_R1176_U348 ; P2_R1176_U13
g20589 and P2_R1176_U342 P2_R1176_U339 ; P2_R1176_U14
g20590 and P2_R1176_U335 P2_R1176_U332 ; P2_R1176_U15
g20591 and P2_R1176_U326 P2_R1176_U323 P2_R1176_U385 ; P2_R1176_U16
g20592 and P2_R1176_U255 P2_R1176_U252 ; P2_R1176_U17
g20593 and P2_R1176_U248 P2_R1176_U245 ; P2_R1176_U18
g20594 not P2_U3184 ; P2_R1176_U19
g20595 not P2_U3175 ; P2_R1176_U20
g20596 not P2_U3181 ; P2_R1176_U21
g20597 nand P2_U3181 P2_R1176_U66 ; P2_R1176_U22
g20598 not P2_U3180 ; P2_R1176_U23
g20599 not P2_U3182 ; P2_R1176_U24
g20600 not P2_U3183 ; P2_R1176_U25
g20601 nand P2_U3184 P2_R1176_U69 ; P2_R1176_U26
g20602 not P2_U3179 ; P2_R1176_U27
g20603 not P2_U3177 ; P2_R1176_U28
g20604 nand P2_U3177 P2_R1176_U73 ; P2_R1176_U29
g20605 not P2_U3176 ; P2_R1176_U30
g20606 not P2_U3178 ; P2_R1176_U31
g20607 nand P2_U3178 P2_R1176_U71 ; P2_R1176_U32
g20608 not P2_U3174 ; P2_R1176_U33
g20609 nand P2_R1176_U238 P2_R1176_U237 P2_R1176_U369 ; P2_R1176_U34
g20610 nand P2_R1176_U32 P2_R1176_U230 ; P2_R1176_U35
g20611 nand P2_R1176_U366 P2_R1176_U218 P2_R1176_U365 ; P2_R1176_U36
g20612 not P2_U3156 ; P2_R1176_U37
g20613 not P2_U3158 ; P2_R1176_U38
g20614 not P2_U3159 ; P2_R1176_U39
g20615 not P2_U3157 ; P2_R1176_U40
g20616 not P2_U3167 ; P2_R1176_U41
g20617 nand P2_U3167 P2_R1176_U78 ; P2_R1176_U42
g20618 not P2_U3166 ; P2_R1176_U43
g20619 not P2_U3169 ; P2_R1176_U44
g20620 not P2_U3171 ; P2_R1176_U45
g20621 not P2_U3172 ; P2_R1176_U46
g20622 nand P2_U3172 P2_R1176_U82 ; P2_R1176_U47
g20623 not P2_U3170 ; P2_R1176_U48
g20624 not P2_U3173 ; P2_R1176_U49
g20625 nand P2_U3173 P2_R1176_U81 ; P2_R1176_U50
g20626 not P2_U3168 ; P2_R1176_U51
g20627 not P2_U3165 ; P2_R1176_U52
g20628 not P2_U3163 ; P2_R1176_U53
g20629 not P2_U3164 ; P2_R1176_U54
g20630 nand P2_U3164 P2_R1176_U87 ; P2_R1176_U55
g20631 not P2_U3162 ; P2_R1176_U56
g20632 not P2_U3161 ; P2_R1176_U57
g20633 not P2_U3160 ; P2_R1176_U58
g20634 nand P2_R1176_U212 P2_R1176_U321 ; P2_R1176_U59
g20635 nand P2_R1176_U55 P2_R1176_U328 ; P2_R1176_U60
g20636 nand P2_R1176_U277 P2_R1176_U276 ; P2_R1176_U61
g20637 nand P2_R1176_U374 P2_R1176_U270 ; P2_R1176_U62
g20638 nand P2_R1176_U47 P2_R1176_U344 ; P2_R1176_U63
g20639 nand P2_R1176_U387 P2_R1176_U386 ; P2_R1176_U64
g20640 nand P2_R1176_U419 P2_R1176_U418 ; P2_R1176_U65
g20641 nand P2_R1176_U407 P2_R1176_U406 ; P2_R1176_U66
g20642 nand P2_R1176_U404 P2_R1176_U403 ; P2_R1176_U67
g20643 nand P2_R1176_U398 P2_R1176_U397 ; P2_R1176_U68
g20644 nand P2_R1176_U401 P2_R1176_U400 ; P2_R1176_U69
g20645 nand P2_R1176_U395 P2_R1176_U394 ; P2_R1176_U70
g20646 nand P2_R1176_U410 P2_R1176_U409 ; P2_R1176_U71
g20647 nand P2_R1176_U413 P2_R1176_U412 ; P2_R1176_U72
g20648 nand P2_R1176_U416 P2_R1176_U415 ; P2_R1176_U73
g20649 nand P2_R1176_U459 P2_R1176_U458 ; P2_R1176_U74
g20650 nand P2_R1176_U507 P2_R1176_U506 ; P2_R1176_U75
g20651 nand P2_R1176_U510 P2_R1176_U509 ; P2_R1176_U76
g20652 nand P2_R1176_U462 P2_R1176_U461 ; P2_R1176_U77
g20653 nand P2_R1176_U486 P2_R1176_U485 ; P2_R1176_U78
g20654 nand P2_R1176_U483 P2_R1176_U482 ; P2_R1176_U79
g20655 nand P2_R1176_U477 P2_R1176_U476 ; P2_R1176_U80
g20656 nand P2_R1176_U465 P2_R1176_U464 ; P2_R1176_U81
g20657 nand P2_R1176_U468 P2_R1176_U467 ; P2_R1176_U82
g20658 nand P2_R1176_U471 P2_R1176_U470 ; P2_R1176_U83
g20659 nand P2_R1176_U474 P2_R1176_U473 ; P2_R1176_U84
g20660 nand P2_R1176_U480 P2_R1176_U479 ; P2_R1176_U85
g20661 nand P2_R1176_U489 P2_R1176_U488 ; P2_R1176_U86
g20662 nand P2_R1176_U498 P2_R1176_U497 ; P2_R1176_U87
g20663 nand P2_R1176_U492 P2_R1176_U491 ; P2_R1176_U88
g20664 nand P2_R1176_U495 P2_R1176_U494 ; P2_R1176_U89
g20665 nand P2_R1176_U501 P2_R1176_U500 ; P2_R1176_U90
g20666 nand P2_R1176_U504 P2_R1176_U503 ; P2_R1176_U91
g20667 nand P2_R1176_U516 P2_R1176_U515 ; P2_R1176_U92
g20668 nand P2_R1176_U623 P2_R1176_U622 ; P2_R1176_U93
g20669 nand P2_R1176_U422 P2_R1176_U421 ; P2_R1176_U94
g20670 nand P2_R1176_U429 P2_R1176_U428 ; P2_R1176_U95
g20671 nand P2_R1176_U436 P2_R1176_U435 ; P2_R1176_U96
g20672 nand P2_R1176_U443 P2_R1176_U442 ; P2_R1176_U97
g20673 nand P2_R1176_U450 P2_R1176_U449 ; P2_R1176_U98
g20674 nand P2_R1176_U457 P2_R1176_U456 ; P2_R1176_U99
g20675 nand P2_R1176_U519 P2_R1176_U518 ; P2_R1176_U100
g20676 nand P2_R1176_U526 P2_R1176_U525 ; P2_R1176_U101
g20677 nand P2_R1176_U533 P2_R1176_U532 ; P2_R1176_U102
g20678 nand P2_R1176_U538 P2_R1176_U537 ; P2_R1176_U103
g20679 nand P2_R1176_U545 P2_R1176_U544 ; P2_R1176_U104
g20680 nand P2_R1176_U552 P2_R1176_U551 ; P2_R1176_U105
g20681 nand P2_R1176_U559 P2_R1176_U558 ; P2_R1176_U106
g20682 nand P2_R1176_U566 P2_R1176_U565 ; P2_R1176_U107
g20683 nand P2_R1176_U571 P2_R1176_U570 ; P2_R1176_U108
g20684 nand P2_R1176_U578 P2_R1176_U577 ; P2_R1176_U109
g20685 nand P2_R1176_U585 P2_R1176_U584 ; P2_R1176_U110
g20686 nand P2_R1176_U592 P2_R1176_U591 ; P2_R1176_U111
g20687 nand P2_R1176_U599 P2_R1176_U598 ; P2_R1176_U112
g20688 nand P2_R1176_U606 P2_R1176_U605 ; P2_R1176_U113
g20689 nand P2_R1176_U611 P2_R1176_U610 ; P2_R1176_U114
g20690 nand P2_R1176_U618 P2_R1176_U617 ; P2_R1176_U115
g20691 and P2_R1176_U224 P2_R1176_U223 ; P2_R1176_U116
g20692 and P2_R1176_U240 P2_R1176_U10 ; P2_R1176_U117
g20693 and P2_R1176_U372 P2_R1176_U241 ; P2_R1176_U118
g20694 and P2_R1176_U431 P2_R1176_U430 P2_R1176_U29 ; P2_R1176_U119
g20695 and P2_R1176_U247 P2_R1176_U5 ; P2_R1176_U120
g20696 and P2_R1176_U452 P2_R1176_U451 P2_R1176_U22 ; P2_R1176_U121
g20697 and P2_R1176_U254 P2_R1176_U4 ; P2_R1176_U122
g20698 and P2_R1176_U272 P2_R1176_U11 ; P2_R1176_U123
g20699 and P2_R1176_U266 P2_R1176_U207 ; P2_R1176_U124
g20700 and P2_R1176_U380 P2_R1176_U273 ; P2_R1176_U125
g20701 and P2_R1176_U284 P2_R1176_U283 ; P2_R1176_U126
g20702 and P2_R1176_U296 P2_R1176_U8 ; P2_R1176_U127
g20703 and P2_R1176_U294 P2_R1176_U208 ; P2_R1176_U128
g20704 and P2_R1176_U312 P2_R1176_U203 ; P2_R1176_U129
g20705 and P2_R1176_U383 P2_R1176_U318 ; P2_R1176_U130
g20706 and P2_R1176_U320 P2_R1176_U310 ; P2_R1176_U131
g20707 and P2_R1176_U320 P2_R1176_U312 ; P2_R1176_U132
g20708 and P2_R1176_U381 P2_R1176_U319 ; P2_R1176_U133
g20709 nand P2_R1176_U513 P2_R1176_U512 ; P2_R1176_U134
g20710 and P2_R1176_U508 P2_R1176_U38 ; P2_R1176_U135
g20711 and P2_R1176_U212 P2_R1176_U209 ; P2_R1176_U136
g20712 and P2_R1176_U325 P2_R1176_U203 ; P2_R1176_U137
g20713 and P2_R1176_U12 P2_R1176_U209 ; P2_R1176_U138
g20714 and P2_R1176_U554 P2_R1176_U553 P2_R1176_U208 ; P2_R1176_U139
g20715 and P2_R1176_U334 P2_R1176_U8 ; P2_R1176_U140
g20716 and P2_R1176_U580 P2_R1176_U579 P2_R1176_U42 ; P2_R1176_U141
g20717 and P2_R1176_U341 P2_R1176_U7 ; P2_R1176_U142
g20718 and P2_R1176_U601 P2_R1176_U600 P2_R1176_U207 ; P2_R1176_U143
g20719 and P2_R1176_U350 P2_R1176_U6 ; P2_R1176_U144
g20720 nand P2_R1176_U620 P2_R1176_U619 ; P2_R1176_U145
g20721 not P2_U3456 ; P2_R1176_U146
g20722 and P2_R1176_U390 P2_R1176_U389 ; P2_R1176_U147
g20723 not P2_U3441 ; P2_R1176_U148
g20724 not P2_U3432 ; P2_R1176_U149
g20725 not P2_U3427 ; P2_R1176_U150
g20726 not P2_U3438 ; P2_R1176_U151
g20727 not P2_U3435 ; P2_R1176_U152
g20728 not P2_U3444 ; P2_R1176_U153
g20729 not P2_U3450 ; P2_R1176_U154
g20730 not P2_U3447 ; P2_R1176_U155
g20731 not P2_U3453 ; P2_R1176_U156
g20732 nand P2_R1176_U118 P2_R1176_U371 ; P2_R1176_U157
g20733 and P2_R1176_U424 P2_R1176_U423 ; P2_R1176_U158
g20734 nand P2_R1176_U370 P2_R1176_U368 ; P2_R1176_U159
g20735 and P2_R1176_U438 P2_R1176_U437 ; P2_R1176_U160
g20736 nand P2_R1176_U227 P2_R1176_U205 P2_R1176_U362 ; P2_R1176_U161
g20737 and P2_R1176_U445 P2_R1176_U444 ; P2_R1176_U162
g20738 nand P2_R1176_U116 P2_R1176_U225 ; P2_R1176_U163
g20739 not P2_U3950 ; P2_R1176_U164
g20740 not P2_U3951 ; P2_R1176_U165
g20741 not P2_U3459 ; P2_R1176_U166
g20742 not P2_U3462 ; P2_R1176_U167
g20743 not P2_U3468 ; P2_R1176_U168
g20744 not P2_U3465 ; P2_R1176_U169
g20745 not P2_U3471 ; P2_R1176_U170
g20746 not P2_U3474 ; P2_R1176_U171
g20747 not P2_U3480 ; P2_R1176_U172
g20748 not P2_U3477 ; P2_R1176_U173
g20749 not P2_U3483 ; P2_R1176_U174
g20750 not P2_U3956 ; P2_R1176_U175
g20751 not P2_U3957 ; P2_R1176_U176
g20752 not P2_U3485 ; P2_R1176_U177
g20753 not P2_U3955 ; P2_R1176_U178
g20754 not P2_U3954 ; P2_R1176_U179
g20755 not P2_U3952 ; P2_R1176_U180
g20756 not P2_U3953 ; P2_R1176_U181
g20757 not P2_U3949 ; P2_R1176_U182
g20758 not P2_U3155 ; P2_R1176_U183
g20759 and P2_R1176_U521 P2_R1176_U520 ; P2_R1176_U184
g20760 nand P2_R1176_U315 P2_R1176_U314 ; P2_R1176_U185
g20761 nand P2_R1176_U307 P2_R1176_U306 ; P2_R1176_U186
g20762 and P2_R1176_U540 P2_R1176_U539 ; P2_R1176_U187
g20763 nand P2_R1176_U303 P2_R1176_U302 ; P2_R1176_U188
g20764 and P2_R1176_U547 P2_R1176_U546 ; P2_R1176_U189
g20765 nand P2_R1176_U299 P2_R1176_U298 ; P2_R1176_U190
g20766 and P2_R1176_U561 P2_R1176_U560 ; P2_R1176_U191
g20767 nand P2_R1176_U26 P2_R1176_U214 ; P2_R1176_U192
g20768 nand P2_R1176_U289 P2_R1176_U288 ; P2_R1176_U193
g20769 and P2_R1176_U573 P2_R1176_U572 ; P2_R1176_U194
g20770 nand P2_R1176_U126 P2_R1176_U285 ; P2_R1176_U195
g20771 and P2_R1176_U587 P2_R1176_U586 ; P2_R1176_U196
g20772 nand P2_R1176_U125 P2_R1176_U379 ; P2_R1176_U197
g20773 and P2_R1176_U594 P2_R1176_U593 ; P2_R1176_U198
g20774 nand P2_R1176_U378 P2_R1176_U373 ; P2_R1176_U199
g20775 nand P2_R1176_U50 P2_R1176_U260 ; P2_R1176_U200
g20776 and P2_R1176_U613 P2_R1176_U612 ; P2_R1176_U201
g20777 nand P2_R1176_U257 P2_R1176_U204 P2_R1176_U363 ; P2_R1176_U202
g20778 nand P2_R1176_U377 P2_R1176_U376 ; P2_R1176_U203
g20779 nand P2_R1176_U64 P2_R1176_U157 ; P2_R1176_U204
g20780 nand P2_R1176_U70 P2_R1176_U163 ; P2_R1176_U205
g20781 not P2_R1176_U22 ; P2_R1176_U206
g20782 nand P2_U3171 P2_R1176_U84 ; P2_R1176_U207
g20783 nand P2_U3163 P2_R1176_U89 ; P2_R1176_U208
g20784 nand P2_U3158 P2_R1176_U75 ; P2_R1176_U209
g20785 not P2_R1176_U47 ; P2_R1176_U210
g20786 not P2_R1176_U55 ; P2_R1176_U211
g20787 nand P2_U3159 P2_R1176_U76 ; P2_R1176_U212
g20788 nand P2_R1176_U402 P2_R1176_U19 ; P2_R1176_U213
g20789 nand P2_U3183 P2_R1176_U213 ; P2_R1176_U214
g20790 not P2_R1176_U26 ; P2_R1176_U215
g20791 not P2_R1176_U192 ; P2_R1176_U216
g20792 nand P2_R1176_U399 P2_R1176_U24 ; P2_R1176_U217
g20793 nand P2_U3182 P2_R1176_U68 ; P2_R1176_U218
g20794 not P2_R1176_U36 ; P2_R1176_U219
g20795 nand P2_R1176_U405 P2_R1176_U23 ; P2_R1176_U220
g20796 nand P2_R1176_U408 P2_R1176_U21 ; P2_R1176_U221
g20797 nand P2_R1176_U23 P2_R1176_U22 ; P2_R1176_U222
g20798 nand P2_R1176_U67 P2_R1176_U222 ; P2_R1176_U223
g20799 nand P2_U3180 P2_R1176_U206 ; P2_R1176_U224
g20800 nand P2_R1176_U4 P2_R1176_U36 ; P2_R1176_U225
g20801 not P2_R1176_U163 ; P2_R1176_U226
g20802 nand P2_U3179 P2_R1176_U163 ; P2_R1176_U227
g20803 not P2_R1176_U161 ; P2_R1176_U228
g20804 nand P2_R1176_U411 P2_R1176_U31 ; P2_R1176_U229
g20805 nand P2_R1176_U229 P2_R1176_U161 ; P2_R1176_U230
g20806 not P2_R1176_U32 ; P2_R1176_U231
g20807 not P2_R1176_U35 ; P2_R1176_U232
g20808 nand P2_R1176_U414 P2_R1176_U30 ; P2_R1176_U233
g20809 nand P2_R1176_U417 P2_R1176_U28 ; P2_R1176_U234
g20810 not P2_R1176_U29 ; P2_R1176_U235
g20811 nand P2_R1176_U30 P2_R1176_U29 ; P2_R1176_U236
g20812 nand P2_R1176_U72 P2_R1176_U236 ; P2_R1176_U237
g20813 nand P2_U3176 P2_R1176_U235 ; P2_R1176_U238
g20814 not P2_R1176_U159 ; P2_R1176_U239
g20815 nand P2_R1176_U420 P2_R1176_U20 ; P2_R1176_U240
g20816 nand P2_U3175 P2_R1176_U65 ; P2_R1176_U241
g20817 not P2_R1176_U157 ; P2_R1176_U242
g20818 nand P2_R1176_U417 P2_R1176_U28 ; P2_R1176_U243
g20819 nand P2_R1176_U243 P2_R1176_U35 ; P2_R1176_U244
g20820 nand P2_R1176_U119 P2_R1176_U244 ; P2_R1176_U245
g20821 nand P2_R1176_U232 P2_R1176_U29 ; P2_R1176_U246
g20822 nand P2_U3176 P2_R1176_U72 ; P2_R1176_U247
g20823 nand P2_R1176_U120 P2_R1176_U246 ; P2_R1176_U248
g20824 nand P2_R1176_U417 P2_R1176_U28 ; P2_R1176_U249
g20825 nand P2_R1176_U408 P2_R1176_U21 ; P2_R1176_U250
g20826 nand P2_R1176_U250 P2_R1176_U36 ; P2_R1176_U251
g20827 nand P2_R1176_U121 P2_R1176_U251 ; P2_R1176_U252
g20828 nand P2_R1176_U219 P2_R1176_U22 ; P2_R1176_U253
g20829 nand P2_U3180 P2_R1176_U67 ; P2_R1176_U254
g20830 nand P2_R1176_U122 P2_R1176_U253 ; P2_R1176_U255
g20831 nand P2_R1176_U408 P2_R1176_U21 ; P2_R1176_U256
g20832 nand P2_U3174 P2_R1176_U157 ; P2_R1176_U257
g20833 not P2_R1176_U202 ; P2_R1176_U258
g20834 nand P2_R1176_U466 P2_R1176_U49 ; P2_R1176_U259
g20835 nand P2_R1176_U259 P2_R1176_U202 ; P2_R1176_U260
g20836 not P2_R1176_U50 ; P2_R1176_U261
g20837 not P2_R1176_U200 ; P2_R1176_U262
g20838 nand P2_R1176_U472 P2_R1176_U48 ; P2_R1176_U263
g20839 nand P2_R1176_U475 P2_R1176_U45 ; P2_R1176_U264
g20840 nand P2_R1176_U210 P2_R1176_U6 ; P2_R1176_U265
g20841 nand P2_U3170 P2_R1176_U83 ; P2_R1176_U266
g20842 nand P2_R1176_U124 P2_R1176_U265 ; P2_R1176_U267
g20843 nand P2_R1176_U469 P2_R1176_U46 ; P2_R1176_U268
g20844 nand P2_R1176_U472 P2_R1176_U48 ; P2_R1176_U269
g20845 nand P2_R1176_U269 P2_R1176_U267 ; P2_R1176_U270
g20846 not P2_R1176_U199 ; P2_R1176_U271
g20847 nand P2_R1176_U478 P2_R1176_U44 ; P2_R1176_U272
g20848 nand P2_U3169 P2_R1176_U80 ; P2_R1176_U273
g20849 not P2_R1176_U197 ; P2_R1176_U274
g20850 nand P2_R1176_U481 P2_R1176_U51 ; P2_R1176_U275
g20851 nand P2_R1176_U275 P2_R1176_U197 ; P2_R1176_U276
g20852 nand P2_U3168 P2_R1176_U85 ; P2_R1176_U277
g20853 not P2_R1176_U61 ; P2_R1176_U278
g20854 nand P2_R1176_U484 P2_R1176_U43 ; P2_R1176_U279
g20855 nand P2_R1176_U487 P2_R1176_U41 ; P2_R1176_U280
g20856 not P2_R1176_U42 ; P2_R1176_U281
g20857 nand P2_R1176_U43 P2_R1176_U42 ; P2_R1176_U282
g20858 nand P2_R1176_U79 P2_R1176_U282 ; P2_R1176_U283
g20859 nand P2_U3166 P2_R1176_U281 ; P2_R1176_U284
g20860 nand P2_R1176_U7 P2_R1176_U61 ; P2_R1176_U285
g20861 not P2_R1176_U195 ; P2_R1176_U286
g20862 nand P2_R1176_U490 P2_R1176_U52 ; P2_R1176_U287
g20863 nand P2_R1176_U287 P2_R1176_U195 ; P2_R1176_U288
g20864 nand P2_U3165 P2_R1176_U86 ; P2_R1176_U289
g20865 not P2_R1176_U193 ; P2_R1176_U290
g20866 nand P2_R1176_U493 P2_R1176_U56 ; P2_R1176_U291
g20867 nand P2_R1176_U496 P2_R1176_U53 ; P2_R1176_U292
g20868 nand P2_R1176_U211 P2_R1176_U8 ; P2_R1176_U293
g20869 nand P2_U3162 P2_R1176_U88 ; P2_R1176_U294
g20870 nand P2_R1176_U128 P2_R1176_U293 ; P2_R1176_U295
g20871 nand P2_R1176_U499 P2_R1176_U54 ; P2_R1176_U296
g20872 nand P2_R1176_U493 P2_R1176_U56 ; P2_R1176_U297
g20873 nand P2_R1176_U127 P2_R1176_U193 ; P2_R1176_U298
g20874 nand P2_R1176_U297 P2_R1176_U295 ; P2_R1176_U299
g20875 not P2_R1176_U190 ; P2_R1176_U300
g20876 nand P2_R1176_U502 P2_R1176_U57 ; P2_R1176_U301
g20877 nand P2_R1176_U301 P2_R1176_U190 ; P2_R1176_U302
g20878 nand P2_U3161 P2_R1176_U90 ; P2_R1176_U303
g20879 not P2_R1176_U188 ; P2_R1176_U304
g20880 nand P2_R1176_U505 P2_R1176_U58 ; P2_R1176_U305
g20881 nand P2_R1176_U305 P2_R1176_U188 ; P2_R1176_U306
g20882 nand P2_U3160 P2_R1176_U91 ; P2_R1176_U307
g20883 not P2_R1176_U186 ; P2_R1176_U308
g20884 nand P2_R1176_U508 P2_R1176_U38 ; P2_R1176_U309
g20885 nand P2_R1176_U212 P2_R1176_U209 P2_R1176_U311 ; P2_R1176_U310
g20886 nand P2_U3157 P2_R1176_U77 ; P2_R1176_U311
g20887 nand P2_R1176_U511 P2_R1176_U39 ; P2_R1176_U312
g20888 nand P2_R1176_U463 P2_R1176_U40 ; P2_R1176_U313
g20889 nand P2_R1176_U129 P2_R1176_U186 ; P2_R1176_U314
g20890 nand P2_R1176_U375 P2_R1176_U310 ; P2_R1176_U315
g20891 not P2_R1176_U185 ; P2_R1176_U316
g20892 nand P2_R1176_U460 P2_R1176_U37 ; P2_R1176_U317
g20893 nand P2_U3156 P2_R1176_U74 ; P2_R1176_U318
g20894 nand P2_U3156 P2_R1176_U74 ; P2_R1176_U319
g20895 nand P2_R1176_U460 P2_R1176_U37 ; P2_R1176_U320
g20896 nand P2_R1176_U312 P2_R1176_U186 ; P2_R1176_U321
g20897 not P2_R1176_U59 ; P2_R1176_U322
g20898 nand P2_R1176_U135 P2_R1176_U12 ; P2_R1176_U323
g20899 nand P2_R1176_U136 P2_R1176_U321 ; P2_R1176_U324
g20900 nand P2_U3157 P2_R1176_U77 ; P2_R1176_U325
g20901 nand P2_R1176_U137 P2_R1176_U324 ; P2_R1176_U326
g20902 nand P2_R1176_U508 P2_R1176_U38 ; P2_R1176_U327
g20903 nand P2_R1176_U296 P2_R1176_U193 ; P2_R1176_U328
g20904 not P2_R1176_U60 ; P2_R1176_U329
g20905 nand P2_R1176_U496 P2_R1176_U53 ; P2_R1176_U330
g20906 nand P2_R1176_U330 P2_R1176_U60 ; P2_R1176_U331
g20907 nand P2_R1176_U139 P2_R1176_U331 ; P2_R1176_U332
g20908 nand P2_R1176_U329 P2_R1176_U208 ; P2_R1176_U333
g20909 nand P2_U3162 P2_R1176_U88 ; P2_R1176_U334
g20910 nand P2_R1176_U140 P2_R1176_U333 ; P2_R1176_U335
g20911 nand P2_R1176_U496 P2_R1176_U53 ; P2_R1176_U336
g20912 nand P2_R1176_U487 P2_R1176_U41 ; P2_R1176_U337
g20913 nand P2_R1176_U337 P2_R1176_U61 ; P2_R1176_U338
g20914 nand P2_R1176_U141 P2_R1176_U338 ; P2_R1176_U339
g20915 nand P2_R1176_U278 P2_R1176_U42 ; P2_R1176_U340
g20916 nand P2_U3166 P2_R1176_U79 ; P2_R1176_U341
g20917 nand P2_R1176_U142 P2_R1176_U340 ; P2_R1176_U342
g20918 nand P2_R1176_U487 P2_R1176_U41 ; P2_R1176_U343
g20919 nand P2_R1176_U268 P2_R1176_U200 ; P2_R1176_U344
g20920 not P2_R1176_U63 ; P2_R1176_U345
g20921 nand P2_R1176_U475 P2_R1176_U45 ; P2_R1176_U346
g20922 nand P2_R1176_U346 P2_R1176_U63 ; P2_R1176_U347
g20923 nand P2_R1176_U143 P2_R1176_U347 ; P2_R1176_U348
g20924 nand P2_R1176_U345 P2_R1176_U207 ; P2_R1176_U349
g20925 nand P2_U3170 P2_R1176_U83 ; P2_R1176_U350
g20926 nand P2_R1176_U144 P2_R1176_U349 ; P2_R1176_U351
g20927 nand P2_R1176_U475 P2_R1176_U45 ; P2_R1176_U352
g20928 nand P2_R1176_U249 P2_R1176_U29 ; P2_R1176_U353
g20929 nand P2_R1176_U256 P2_R1176_U22 ; P2_R1176_U354
g20930 nand P2_R1176_U327 P2_R1176_U209 ; P2_R1176_U355
g20931 nand P2_R1176_U312 P2_R1176_U212 ; P2_R1176_U356
g20932 nand P2_R1176_U336 P2_R1176_U208 ; P2_R1176_U357
g20933 nand P2_R1176_U296 P2_R1176_U55 ; P2_R1176_U358
g20934 nand P2_R1176_U343 P2_R1176_U42 ; P2_R1176_U359
g20935 nand P2_R1176_U352 P2_R1176_U207 ; P2_R1176_U360
g20936 nand P2_R1176_U268 P2_R1176_U47 ; P2_R1176_U361
g20937 nand P2_U3179 P2_R1176_U70 ; P2_R1176_U362
g20938 nand P2_U3174 P2_R1176_U64 ; P2_R1176_U363
g20939 nand P2_R1176_U314 P2_R1176_U311 P2_R1176_U130 ; P2_R1176_U364
g20940 nand P2_U3183 P2_R1176_U213 P2_R1176_U367 ; P2_R1176_U365
g20941 nand P2_R1176_U215 P2_R1176_U217 ; P2_R1176_U366
g20942 nand P2_R1176_U399 P2_R1176_U24 ; P2_R1176_U367
g20943 nand P2_R1176_U10 P2_R1176_U161 ; P2_R1176_U368
g20944 nand P2_R1176_U231 P2_R1176_U5 ; P2_R1176_U369
g20945 not P2_R1176_U34 ; P2_R1176_U370
g20946 nand P2_R1176_U117 P2_R1176_U161 ; P2_R1176_U371
g20947 nand P2_R1176_U34 P2_R1176_U240 ; P2_R1176_U372
g20948 nand P2_R1176_U11 P2_R1176_U202 ; P2_R1176_U373
g20949 nand P2_R1176_U261 P2_R1176_U9 ; P2_R1176_U374
g20950 nand P2_R1176_U376 P2_R1176_U311 P2_R1176_U377 ; P2_R1176_U375
g20951 nand P2_R1176_U77 P2_R1176_U309 ; P2_R1176_U376
g20952 nand P2_U3157 P2_R1176_U309 ; P2_R1176_U377
g20953 not P2_R1176_U62 ; P2_R1176_U378
g20954 nand P2_R1176_U123 P2_R1176_U202 ; P2_R1176_U379
g20955 nand P2_R1176_U62 P2_R1176_U272 ; P2_R1176_U380
g20956 nand P2_R1176_U131 P2_R1176_U375 ; P2_R1176_U381
g20957 nand P2_R1176_U186 P2_R1176_U203 P2_R1176_U132 ; P2_R1176_U382
g20958 nand P2_R1176_U384 P2_R1176_U309 P2_R1176_U313 ; P2_R1176_U383
g20959 nand P2_R1176_U212 P2_R1176_U209 ; P2_R1176_U384
g20960 nand P2_R1176_U138 P2_R1176_U322 ; P2_R1176_U385
g20961 nand P2_U3184 P2_R1176_U146 ; P2_R1176_U386
g20962 nand P2_U3456 P2_R1176_U19 ; P2_R1176_U387
g20963 not P2_R1176_U64 ; P2_R1176_U388
g20964 nand P2_R1176_U388 P2_U3174 ; P2_R1176_U389
g20965 nand P2_R1176_U64 P2_R1176_U33 ; P2_R1176_U390
g20966 nand P2_R1176_U388 P2_U3174 ; P2_R1176_U391
g20967 nand P2_R1176_U64 P2_R1176_U33 ; P2_R1176_U392
g20968 nand P2_R1176_U392 P2_R1176_U391 ; P2_R1176_U393
g20969 nand P2_U3184 P2_R1176_U148 ; P2_R1176_U394
g20970 nand P2_U3441 P2_R1176_U19 ; P2_R1176_U395
g20971 not P2_R1176_U70 ; P2_R1176_U396
g20972 nand P2_U3184 P2_R1176_U149 ; P2_R1176_U397
g20973 nand P2_U3432 P2_R1176_U19 ; P2_R1176_U398
g20974 not P2_R1176_U68 ; P2_R1176_U399
g20975 nand P2_U3184 P2_R1176_U150 ; P2_R1176_U400
g20976 nand P2_U3427 P2_R1176_U19 ; P2_R1176_U401
g20977 not P2_R1176_U69 ; P2_R1176_U402
g20978 nand P2_U3184 P2_R1176_U151 ; P2_R1176_U403
g20979 nand P2_U3438 P2_R1176_U19 ; P2_R1176_U404
g20980 not P2_R1176_U67 ; P2_R1176_U405
g20981 nand P2_U3184 P2_R1176_U152 ; P2_R1176_U406
g20982 nand P2_U3435 P2_R1176_U19 ; P2_R1176_U407
g20983 not P2_R1176_U66 ; P2_R1176_U408
g20984 nand P2_U3184 P2_R1176_U153 ; P2_R1176_U409
g20985 nand P2_U3444 P2_R1176_U19 ; P2_R1176_U410
g20986 not P2_R1176_U71 ; P2_R1176_U411
g20987 nand P2_U3184 P2_R1176_U154 ; P2_R1176_U412
g20988 nand P2_U3450 P2_R1176_U19 ; P2_R1176_U413
g20989 not P2_R1176_U72 ; P2_R1176_U414
g20990 nand P2_U3184 P2_R1176_U155 ; P2_R1176_U415
g20991 nand P2_U3447 P2_R1176_U19 ; P2_R1176_U416
g20992 not P2_R1176_U73 ; P2_R1176_U417
g20993 nand P2_U3184 P2_R1176_U156 ; P2_R1176_U418
g20994 nand P2_U3453 P2_R1176_U19 ; P2_R1176_U419
g20995 not P2_R1176_U65 ; P2_R1176_U420
g20996 nand P2_R1176_U147 P2_R1176_U157 ; P2_R1176_U421
g20997 nand P2_R1176_U242 P2_R1176_U393 ; P2_R1176_U422
g20998 nand P2_R1176_U420 P2_U3175 ; P2_R1176_U423
g20999 nand P2_R1176_U65 P2_R1176_U20 ; P2_R1176_U424
g21000 nand P2_R1176_U420 P2_U3175 ; P2_R1176_U425
g21001 nand P2_R1176_U65 P2_R1176_U20 ; P2_R1176_U426
g21002 nand P2_R1176_U426 P2_R1176_U425 ; P2_R1176_U427
g21003 nand P2_R1176_U158 P2_R1176_U159 ; P2_R1176_U428
g21004 nand P2_R1176_U239 P2_R1176_U427 ; P2_R1176_U429
g21005 nand P2_R1176_U414 P2_U3176 ; P2_R1176_U430
g21006 nand P2_R1176_U72 P2_R1176_U30 ; P2_R1176_U431
g21007 nand P2_R1176_U417 P2_U3177 ; P2_R1176_U432
g21008 nand P2_R1176_U73 P2_R1176_U28 ; P2_R1176_U433
g21009 nand P2_R1176_U433 P2_R1176_U432 ; P2_R1176_U434
g21010 nand P2_R1176_U353 P2_R1176_U35 ; P2_R1176_U435
g21011 nand P2_R1176_U434 P2_R1176_U232 ; P2_R1176_U436
g21012 nand P2_R1176_U411 P2_U3178 ; P2_R1176_U437
g21013 nand P2_R1176_U71 P2_R1176_U31 ; P2_R1176_U438
g21014 nand P2_R1176_U411 P2_U3178 ; P2_R1176_U439
g21015 nand P2_R1176_U71 P2_R1176_U31 ; P2_R1176_U440
g21016 nand P2_R1176_U440 P2_R1176_U439 ; P2_R1176_U441
g21017 nand P2_R1176_U160 P2_R1176_U161 ; P2_R1176_U442
g21018 nand P2_R1176_U228 P2_R1176_U441 ; P2_R1176_U443
g21019 nand P2_R1176_U396 P2_U3179 ; P2_R1176_U444
g21020 nand P2_R1176_U70 P2_R1176_U27 ; P2_R1176_U445
g21021 nand P2_R1176_U396 P2_U3179 ; P2_R1176_U446
g21022 nand P2_R1176_U70 P2_R1176_U27 ; P2_R1176_U447
g21023 nand P2_R1176_U447 P2_R1176_U446 ; P2_R1176_U448
g21024 nand P2_R1176_U162 P2_R1176_U163 ; P2_R1176_U449
g21025 nand P2_R1176_U226 P2_R1176_U448 ; P2_R1176_U450
g21026 nand P2_R1176_U405 P2_U3180 ; P2_R1176_U451
g21027 nand P2_R1176_U67 P2_R1176_U23 ; P2_R1176_U452
g21028 nand P2_R1176_U408 P2_U3181 ; P2_R1176_U453
g21029 nand P2_R1176_U66 P2_R1176_U21 ; P2_R1176_U454
g21030 nand P2_R1176_U454 P2_R1176_U453 ; P2_R1176_U455
g21031 nand P2_R1176_U354 P2_R1176_U36 ; P2_R1176_U456
g21032 nand P2_R1176_U455 P2_R1176_U219 ; P2_R1176_U457
g21033 nand P2_U3184 P2_R1176_U164 ; P2_R1176_U458
g21034 nand P2_U3950 P2_R1176_U19 ; P2_R1176_U459
g21035 not P2_R1176_U74 ; P2_R1176_U460
g21036 nand P2_U3184 P2_R1176_U165 ; P2_R1176_U461
g21037 nand P2_U3951 P2_R1176_U19 ; P2_R1176_U462
g21038 not P2_R1176_U77 ; P2_R1176_U463
g21039 nand P2_U3184 P2_R1176_U166 ; P2_R1176_U464
g21040 nand P2_U3459 P2_R1176_U19 ; P2_R1176_U465
g21041 not P2_R1176_U81 ; P2_R1176_U466
g21042 nand P2_U3184 P2_R1176_U167 ; P2_R1176_U467
g21043 nand P2_U3462 P2_R1176_U19 ; P2_R1176_U468
g21044 not P2_R1176_U82 ; P2_R1176_U469
g21045 nand P2_U3184 P2_R1176_U168 ; P2_R1176_U470
g21046 nand P2_U3468 P2_R1176_U19 ; P2_R1176_U471
g21047 not P2_R1176_U83 ; P2_R1176_U472
g21048 nand P2_U3184 P2_R1176_U169 ; P2_R1176_U473
g21049 nand P2_U3465 P2_R1176_U19 ; P2_R1176_U474
g21050 not P2_R1176_U84 ; P2_R1176_U475
g21051 nand P2_U3184 P2_R1176_U170 ; P2_R1176_U476
g21052 nand P2_U3471 P2_R1176_U19 ; P2_R1176_U477
g21053 not P2_R1176_U80 ; P2_R1176_U478
g21054 nand P2_U3184 P2_R1176_U171 ; P2_R1176_U479
g21055 nand P2_U3474 P2_R1176_U19 ; P2_R1176_U480
g21056 not P2_R1176_U85 ; P2_R1176_U481
g21057 nand P2_U3184 P2_R1176_U172 ; P2_R1176_U482
g21058 nand P2_U3480 P2_R1176_U19 ; P2_R1176_U483
g21059 not P2_R1176_U79 ; P2_R1176_U484
g21060 nand P2_U3184 P2_R1176_U173 ; P2_R1176_U485
g21061 nand P2_U3477 P2_R1176_U19 ; P2_R1176_U486
g21062 not P2_R1176_U78 ; P2_R1176_U487
g21063 nand P2_U3184 P2_R1176_U174 ; P2_R1176_U488
g21064 nand P2_U3483 P2_R1176_U19 ; P2_R1176_U489
g21065 not P2_R1176_U86 ; P2_R1176_U490
g21066 nand P2_U3184 P2_R1176_U175 ; P2_R1176_U491
g21067 nand P2_U3956 P2_R1176_U19 ; P2_R1176_U492
g21068 not P2_R1176_U88 ; P2_R1176_U493
g21069 nand P2_U3184 P2_R1176_U176 ; P2_R1176_U494
g21070 nand P2_U3957 P2_R1176_U19 ; P2_R1176_U495
g21071 not P2_R1176_U89 ; P2_R1176_U496
g21072 nand P2_U3184 P2_R1176_U177 ; P2_R1176_U497
g21073 nand P2_U3485 P2_R1176_U19 ; P2_R1176_U498
g21074 not P2_R1176_U87 ; P2_R1176_U499
g21075 nand P2_U3184 P2_R1176_U178 ; P2_R1176_U500
g21076 nand P2_U3955 P2_R1176_U19 ; P2_R1176_U501
g21077 not P2_R1176_U90 ; P2_R1176_U502
g21078 nand P2_U3184 P2_R1176_U179 ; P2_R1176_U503
g21079 nand P2_U3954 P2_R1176_U19 ; P2_R1176_U504
g21080 not P2_R1176_U91 ; P2_R1176_U505
g21081 nand P2_U3184 P2_R1176_U180 ; P2_R1176_U506
g21082 nand P2_U3952 P2_R1176_U19 ; P2_R1176_U507
g21083 not P2_R1176_U75 ; P2_R1176_U508
g21084 nand P2_U3184 P2_R1176_U181 ; P2_R1176_U509
g21085 nand P2_U3953 P2_R1176_U19 ; P2_R1176_U510
g21086 not P2_R1176_U76 ; P2_R1176_U511
g21087 nand P2_U3184 P2_R1176_U182 ; P2_R1176_U512
g21088 nand P2_U3949 P2_R1176_U19 ; P2_R1176_U513
g21089 not P2_R1176_U134 ; P2_R1176_U514
g21090 nand P2_U3155 P2_R1176_U514 ; P2_R1176_U515
g21091 nand P2_R1176_U134 P2_R1176_U183 ; P2_R1176_U516
g21092 not P2_R1176_U92 ; P2_R1176_U517
g21093 nand P2_R1176_U364 P2_R1176_U317 P2_R1176_U517 ; P2_R1176_U518
g21094 nand P2_R1176_U133 P2_R1176_U382 P2_R1176_U92 ; P2_R1176_U519
g21095 nand P2_R1176_U460 P2_U3156 ; P2_R1176_U520
g21096 nand P2_R1176_U74 P2_R1176_U37 ; P2_R1176_U521
g21097 nand P2_R1176_U460 P2_U3156 ; P2_R1176_U522
g21098 nand P2_R1176_U74 P2_R1176_U37 ; P2_R1176_U523
g21099 nand P2_R1176_U523 P2_R1176_U522 ; P2_R1176_U524
g21100 nand P2_R1176_U184 P2_R1176_U185 ; P2_R1176_U525
g21101 nand P2_R1176_U316 P2_R1176_U524 ; P2_R1176_U526
g21102 nand P2_R1176_U463 P2_U3157 ; P2_R1176_U527
g21103 nand P2_R1176_U77 P2_R1176_U40 ; P2_R1176_U528
g21104 nand P2_R1176_U508 P2_U3158 ; P2_R1176_U529
g21105 nand P2_R1176_U75 P2_R1176_U38 ; P2_R1176_U530
g21106 nand P2_R1176_U530 P2_R1176_U529 ; P2_R1176_U531
g21107 nand P2_R1176_U355 P2_R1176_U59 ; P2_R1176_U532
g21108 nand P2_R1176_U531 P2_R1176_U322 ; P2_R1176_U533
g21109 nand P2_R1176_U511 P2_U3159 ; P2_R1176_U534
g21110 nand P2_R1176_U76 P2_R1176_U39 ; P2_R1176_U535
g21111 nand P2_R1176_U535 P2_R1176_U534 ; P2_R1176_U536
g21112 nand P2_R1176_U356 P2_R1176_U186 ; P2_R1176_U537
g21113 nand P2_R1176_U308 P2_R1176_U536 ; P2_R1176_U538
g21114 nand P2_R1176_U505 P2_U3160 ; P2_R1176_U539
g21115 nand P2_R1176_U91 P2_R1176_U58 ; P2_R1176_U540
g21116 nand P2_R1176_U505 P2_U3160 ; P2_R1176_U541
g21117 nand P2_R1176_U91 P2_R1176_U58 ; P2_R1176_U542
g21118 nand P2_R1176_U542 P2_R1176_U541 ; P2_R1176_U543
g21119 nand P2_R1176_U187 P2_R1176_U188 ; P2_R1176_U544
g21120 nand P2_R1176_U304 P2_R1176_U543 ; P2_R1176_U545
g21121 nand P2_R1176_U502 P2_U3161 ; P2_R1176_U546
g21122 nand P2_R1176_U90 P2_R1176_U57 ; P2_R1176_U547
g21123 nand P2_R1176_U502 P2_U3161 ; P2_R1176_U548
g21124 nand P2_R1176_U90 P2_R1176_U57 ; P2_R1176_U549
g21125 nand P2_R1176_U549 P2_R1176_U548 ; P2_R1176_U550
g21126 nand P2_R1176_U189 P2_R1176_U190 ; P2_R1176_U551
g21127 nand P2_R1176_U300 P2_R1176_U550 ; P2_R1176_U552
g21128 nand P2_R1176_U493 P2_U3162 ; P2_R1176_U553
g21129 nand P2_R1176_U88 P2_R1176_U56 ; P2_R1176_U554
g21130 nand P2_R1176_U496 P2_U3163 ; P2_R1176_U555
g21131 nand P2_R1176_U89 P2_R1176_U53 ; P2_R1176_U556
g21132 nand P2_R1176_U556 P2_R1176_U555 ; P2_R1176_U557
g21133 nand P2_R1176_U357 P2_R1176_U60 ; P2_R1176_U558
g21134 nand P2_R1176_U557 P2_R1176_U329 ; P2_R1176_U559
g21135 nand P2_R1176_U399 P2_U3182 ; P2_R1176_U560
g21136 nand P2_R1176_U68 P2_R1176_U24 ; P2_R1176_U561
g21137 nand P2_R1176_U399 P2_U3182 ; P2_R1176_U562
g21138 nand P2_R1176_U68 P2_R1176_U24 ; P2_R1176_U563
g21139 nand P2_R1176_U563 P2_R1176_U562 ; P2_R1176_U564
g21140 nand P2_R1176_U191 P2_R1176_U192 ; P2_R1176_U565
g21141 nand P2_R1176_U216 P2_R1176_U564 ; P2_R1176_U566
g21142 nand P2_R1176_U499 P2_U3164 ; P2_R1176_U567
g21143 nand P2_R1176_U87 P2_R1176_U54 ; P2_R1176_U568
g21144 nand P2_R1176_U568 P2_R1176_U567 ; P2_R1176_U569
g21145 nand P2_R1176_U358 P2_R1176_U193 ; P2_R1176_U570
g21146 nand P2_R1176_U290 P2_R1176_U569 ; P2_R1176_U571
g21147 nand P2_R1176_U490 P2_U3165 ; P2_R1176_U572
g21148 nand P2_R1176_U86 P2_R1176_U52 ; P2_R1176_U573
g21149 nand P2_R1176_U490 P2_U3165 ; P2_R1176_U574
g21150 nand P2_R1176_U86 P2_R1176_U52 ; P2_R1176_U575
g21151 nand P2_R1176_U575 P2_R1176_U574 ; P2_R1176_U576
g21152 nand P2_R1176_U194 P2_R1176_U195 ; P2_R1176_U577
g21153 nand P2_R1176_U286 P2_R1176_U576 ; P2_R1176_U578
g21154 nand P2_R1176_U484 P2_U3166 ; P2_R1176_U579
g21155 nand P2_R1176_U79 P2_R1176_U43 ; P2_R1176_U580
g21156 nand P2_R1176_U487 P2_U3167 ; P2_R1176_U581
g21157 nand P2_R1176_U78 P2_R1176_U41 ; P2_R1176_U582
g21158 nand P2_R1176_U582 P2_R1176_U581 ; P2_R1176_U583
g21159 nand P2_R1176_U359 P2_R1176_U61 ; P2_R1176_U584
g21160 nand P2_R1176_U583 P2_R1176_U278 ; P2_R1176_U585
g21161 nand P2_R1176_U481 P2_U3168 ; P2_R1176_U586
g21162 nand P2_R1176_U85 P2_R1176_U51 ; P2_R1176_U587
g21163 nand P2_R1176_U481 P2_U3168 ; P2_R1176_U588
g21164 nand P2_R1176_U85 P2_R1176_U51 ; P2_R1176_U589
g21165 nand P2_R1176_U589 P2_R1176_U588 ; P2_R1176_U590
g21166 nand P2_R1176_U196 P2_R1176_U197 ; P2_R1176_U591
g21167 nand P2_R1176_U274 P2_R1176_U590 ; P2_R1176_U592
g21168 nand P2_R1176_U478 P2_U3169 ; P2_R1176_U593
g21169 nand P2_R1176_U80 P2_R1176_U44 ; P2_R1176_U594
g21170 nand P2_R1176_U478 P2_U3169 ; P2_R1176_U595
g21171 nand P2_R1176_U80 P2_R1176_U44 ; P2_R1176_U596
g21172 nand P2_R1176_U596 P2_R1176_U595 ; P2_R1176_U597
g21173 nand P2_R1176_U198 P2_R1176_U199 ; P2_R1176_U598
g21174 nand P2_R1176_U271 P2_R1176_U597 ; P2_R1176_U599
g21175 nand P2_R1176_U472 P2_U3170 ; P2_R1176_U600
g21176 nand P2_R1176_U83 P2_R1176_U48 ; P2_R1176_U601
g21177 nand P2_R1176_U475 P2_U3171 ; P2_R1176_U602
g21178 nand P2_R1176_U84 P2_R1176_U45 ; P2_R1176_U603
g21179 nand P2_R1176_U603 P2_R1176_U602 ; P2_R1176_U604
g21180 nand P2_R1176_U360 P2_R1176_U63 ; P2_R1176_U605
g21181 nand P2_R1176_U604 P2_R1176_U345 ; P2_R1176_U606
g21182 nand P2_R1176_U469 P2_U3172 ; P2_R1176_U607
g21183 nand P2_R1176_U82 P2_R1176_U46 ; P2_R1176_U608
g21184 nand P2_R1176_U608 P2_R1176_U607 ; P2_R1176_U609
g21185 nand P2_R1176_U361 P2_R1176_U200 ; P2_R1176_U610
g21186 nand P2_R1176_U262 P2_R1176_U609 ; P2_R1176_U611
g21187 nand P2_R1176_U466 P2_U3173 ; P2_R1176_U612
g21188 nand P2_R1176_U81 P2_R1176_U49 ; P2_R1176_U613
g21189 nand P2_R1176_U466 P2_U3173 ; P2_R1176_U614
g21190 nand P2_R1176_U81 P2_R1176_U49 ; P2_R1176_U615
g21191 nand P2_R1176_U615 P2_R1176_U614 ; P2_R1176_U616
g21192 nand P2_R1176_U201 P2_R1176_U202 ; P2_R1176_U617
g21193 nand P2_R1176_U258 P2_R1176_U616 ; P2_R1176_U618
g21194 nand P2_R1176_U69 P2_R1176_U19 ; P2_R1176_U619
g21195 nand P2_R1176_U402 P2_U3184 ; P2_R1176_U620
g21196 not P2_R1176_U145 ; P2_R1176_U621
g21197 nand P2_R1176_U621 P2_U3183 ; P2_R1176_U622
g21198 nand P2_R1176_U145 P2_R1176_U25 ; P2_R1176_U623
g21199 and P2_R1131_U179 P2_R1131_U178 ; P2_R1131_U4
g21200 and P2_R1131_U197 P2_R1131_U196 ; P2_R1131_U5
g21201 and P2_R1131_U237 P2_R1131_U236 ; P2_R1131_U6
g21202 and P2_R1131_U246 P2_R1131_U245 ; P2_R1131_U7
g21203 and P2_R1131_U264 P2_R1131_U263 ; P2_R1131_U8
g21204 and P2_R1131_U272 P2_R1131_U271 ; P2_R1131_U9
g21205 and P2_R1131_U351 P2_R1131_U348 ; P2_R1131_U10
g21206 and P2_R1131_U344 P2_R1131_U341 ; P2_R1131_U11
g21207 and P2_R1131_U335 P2_R1131_U332 ; P2_R1131_U12
g21208 and P2_R1131_U326 P2_R1131_U323 ; P2_R1131_U13
g21209 and P2_R1131_U320 P2_R1131_U318 ; P2_R1131_U14
g21210 and P2_R1131_U313 P2_R1131_U310 ; P2_R1131_U15
g21211 and P2_R1131_U235 P2_R1131_U232 ; P2_R1131_U16
g21212 and P2_R1131_U227 P2_R1131_U224 ; P2_R1131_U17
g21213 and P2_R1131_U213 P2_R1131_U210 ; P2_R1131_U18
g21214 not P2_U3447 ; P2_R1131_U19
g21215 not P2_U3073 ; P2_R1131_U20
g21216 not P2_U3072 ; P2_R1131_U21
g21217 nand P2_U3073 P2_U3447 ; P2_R1131_U22
g21218 not P2_U3450 ; P2_R1131_U23
g21219 not P2_U3441 ; P2_R1131_U24
g21220 not P2_U3062 ; P2_R1131_U25
g21221 not P2_U3069 ; P2_R1131_U26
g21222 not P2_U3435 ; P2_R1131_U27
g21223 not P2_U3070 ; P2_R1131_U28
g21224 not P2_U3427 ; P2_R1131_U29
g21225 not P2_U3079 ; P2_R1131_U30
g21226 nand P2_U3079 P2_U3427 ; P2_R1131_U31
g21227 not P2_U3438 ; P2_R1131_U32
g21228 not P2_U3066 ; P2_R1131_U33
g21229 nand P2_U3062 P2_U3441 ; P2_R1131_U34
g21230 not P2_U3444 ; P2_R1131_U35
g21231 not P2_U3453 ; P2_R1131_U36
g21232 not P2_U3086 ; P2_R1131_U37
g21233 not P2_U3085 ; P2_R1131_U38
g21234 not P2_U3456 ; P2_R1131_U39
g21235 nand P2_R1131_U61 P2_R1131_U205 ; P2_R1131_U40
g21236 nand P2_R1131_U117 P2_R1131_U193 ; P2_R1131_U41
g21237 nand P2_R1131_U182 P2_R1131_U183 ; P2_R1131_U42
g21238 nand P2_U3432 P2_U3080 ; P2_R1131_U43
g21239 nand P2_R1131_U122 P2_R1131_U219 ; P2_R1131_U44
g21240 nand P2_R1131_U216 P2_R1131_U215 ; P2_R1131_U45
g21241 not P2_U3950 ; P2_R1131_U46
g21242 not P2_U3055 ; P2_R1131_U47
g21243 not P2_U3059 ; P2_R1131_U48
g21244 not P2_U3951 ; P2_R1131_U49
g21245 not P2_U3952 ; P2_R1131_U50
g21246 not P2_U3060 ; P2_R1131_U51
g21247 not P2_U3953 ; P2_R1131_U52
g21248 not P2_U3067 ; P2_R1131_U53
g21249 not P2_U3956 ; P2_R1131_U54
g21250 not P2_U3077 ; P2_R1131_U55
g21251 not P2_U3477 ; P2_R1131_U56
g21252 not P2_U3075 ; P2_R1131_U57
g21253 not P2_U3071 ; P2_R1131_U58
g21254 nand P2_U3075 P2_U3477 ; P2_R1131_U59
g21255 not P2_U3480 ; P2_R1131_U60
g21256 nand P2_U3086 P2_U3453 ; P2_R1131_U61
g21257 not P2_U3459 ; P2_R1131_U62
g21258 not P2_U3064 ; P2_R1131_U63
g21259 not P2_U3465 ; P2_R1131_U64
g21260 not P2_U3074 ; P2_R1131_U65
g21261 not P2_U3462 ; P2_R1131_U66
g21262 not P2_U3065 ; P2_R1131_U67
g21263 nand P2_U3065 P2_U3462 ; P2_R1131_U68
g21264 not P2_U3468 ; P2_R1131_U69
g21265 not P2_U3082 ; P2_R1131_U70
g21266 not P2_U3471 ; P2_R1131_U71
g21267 not P2_U3081 ; P2_R1131_U72
g21268 not P2_U3474 ; P2_R1131_U73
g21269 not P2_U3076 ; P2_R1131_U74
g21270 not P2_U3483 ; P2_R1131_U75
g21271 not P2_U3084 ; P2_R1131_U76
g21272 nand P2_U3084 P2_U3483 ; P2_R1131_U77
g21273 not P2_U3485 ; P2_R1131_U78
g21274 not P2_U3083 ; P2_R1131_U79
g21275 nand P2_U3083 P2_U3485 ; P2_R1131_U80
g21276 not P2_U3957 ; P2_R1131_U81
g21277 not P2_U3955 ; P2_R1131_U82
g21278 not P2_U3063 ; P2_R1131_U83
g21279 not P2_U3954 ; P2_R1131_U84
g21280 not P2_U3068 ; P2_R1131_U85
g21281 nand P2_U3951 P2_U3059 ; P2_R1131_U86
g21282 not P2_U3056 ; P2_R1131_U87
g21283 not P2_U3949 ; P2_R1131_U88
g21284 nand P2_R1131_U306 P2_R1131_U176 ; P2_R1131_U89
g21285 not P2_U3078 ; P2_R1131_U90
g21286 nand P2_R1131_U77 P2_R1131_U315 ; P2_R1131_U91
g21287 nand P2_R1131_U261 P2_R1131_U260 ; P2_R1131_U92
g21288 nand P2_R1131_U68 P2_R1131_U337 ; P2_R1131_U93
g21289 nand P2_R1131_U457 P2_R1131_U456 ; P2_R1131_U94
g21290 nand P2_R1131_U504 P2_R1131_U503 ; P2_R1131_U95
g21291 nand P2_R1131_U375 P2_R1131_U374 ; P2_R1131_U96
g21292 nand P2_R1131_U380 P2_R1131_U379 ; P2_R1131_U97
g21293 nand P2_R1131_U387 P2_R1131_U386 ; P2_R1131_U98
g21294 nand P2_R1131_U394 P2_R1131_U393 ; P2_R1131_U99
g21295 nand P2_R1131_U399 P2_R1131_U398 ; P2_R1131_U100
g21296 nand P2_R1131_U408 P2_R1131_U407 ; P2_R1131_U101
g21297 nand P2_R1131_U415 P2_R1131_U414 ; P2_R1131_U102
g21298 nand P2_R1131_U422 P2_R1131_U421 ; P2_R1131_U103
g21299 nand P2_R1131_U429 P2_R1131_U428 ; P2_R1131_U104
g21300 nand P2_R1131_U434 P2_R1131_U433 ; P2_R1131_U105
g21301 nand P2_R1131_U441 P2_R1131_U440 ; P2_R1131_U106
g21302 nand P2_R1131_U448 P2_R1131_U447 ; P2_R1131_U107
g21303 nand P2_R1131_U462 P2_R1131_U461 ; P2_R1131_U108
g21304 nand P2_R1131_U467 P2_R1131_U466 ; P2_R1131_U109
g21305 nand P2_R1131_U474 P2_R1131_U473 ; P2_R1131_U110
g21306 nand P2_R1131_U481 P2_R1131_U480 ; P2_R1131_U111
g21307 nand P2_R1131_U488 P2_R1131_U487 ; P2_R1131_U112
g21308 nand P2_R1131_U495 P2_R1131_U494 ; P2_R1131_U113
g21309 nand P2_R1131_U500 P2_R1131_U499 ; P2_R1131_U114
g21310 and P2_R1131_U189 P2_R1131_U187 ; P2_R1131_U115
g21311 and P2_R1131_U4 P2_R1131_U180 ; P2_R1131_U116
g21312 and P2_R1131_U194 P2_R1131_U192 ; P2_R1131_U117
g21313 and P2_R1131_U201 P2_R1131_U200 ; P2_R1131_U118
g21314 and P2_R1131_U382 P2_R1131_U381 P2_R1131_U22 ; P2_R1131_U119
g21315 and P2_R1131_U212 P2_R1131_U5 ; P2_R1131_U120
g21316 and P2_R1131_U181 P2_R1131_U180 ; P2_R1131_U121
g21317 and P2_R1131_U220 P2_R1131_U218 ; P2_R1131_U122
g21318 and P2_R1131_U389 P2_R1131_U388 P2_R1131_U34 ; P2_R1131_U123
g21319 and P2_R1131_U226 P2_R1131_U4 ; P2_R1131_U124
g21320 and P2_R1131_U234 P2_R1131_U181 ; P2_R1131_U125
g21321 and P2_R1131_U204 P2_R1131_U6 ; P2_R1131_U126
g21322 and P2_R1131_U239 P2_R1131_U171 ; P2_R1131_U127
g21323 and P2_R1131_U250 P2_R1131_U7 ; P2_R1131_U128
g21324 and P2_R1131_U248 P2_R1131_U172 ; P2_R1131_U129
g21325 and P2_R1131_U268 P2_R1131_U267 ; P2_R1131_U130
g21326 and P2_R1131_U9 P2_R1131_U282 ; P2_R1131_U131
g21327 and P2_R1131_U285 P2_R1131_U280 ; P2_R1131_U132
g21328 and P2_R1131_U301 P2_R1131_U298 ; P2_R1131_U133
g21329 and P2_R1131_U368 P2_R1131_U302 ; P2_R1131_U134
g21330 and P2_R1131_U160 P2_R1131_U278 ; P2_R1131_U135
g21331 and P2_R1131_U455 P2_R1131_U454 P2_R1131_U80 ; P2_R1131_U136
g21332 and P2_R1131_U325 P2_R1131_U9 ; P2_R1131_U137
g21333 and P2_R1131_U469 P2_R1131_U468 P2_R1131_U59 ; P2_R1131_U138
g21334 and P2_R1131_U334 P2_R1131_U8 ; P2_R1131_U139
g21335 and P2_R1131_U490 P2_R1131_U489 P2_R1131_U172 ; P2_R1131_U140
g21336 and P2_R1131_U343 P2_R1131_U7 ; P2_R1131_U141
g21337 and P2_R1131_U502 P2_R1131_U501 P2_R1131_U171 ; P2_R1131_U142
g21338 and P2_R1131_U350 P2_R1131_U6 ; P2_R1131_U143
g21339 nand P2_R1131_U118 P2_R1131_U202 ; P2_R1131_U144
g21340 nand P2_R1131_U217 P2_R1131_U229 ; P2_R1131_U145
g21341 not P2_U3057 ; P2_R1131_U146
g21342 not P2_U3960 ; P2_R1131_U147
g21343 and P2_R1131_U403 P2_R1131_U402 ; P2_R1131_U148
g21344 nand P2_R1131_U304 P2_R1131_U169 P2_R1131_U364 ; P2_R1131_U149
g21345 and P2_R1131_U410 P2_R1131_U409 ; P2_R1131_U150
g21346 nand P2_R1131_U370 P2_R1131_U369 P2_R1131_U134 ; P2_R1131_U151
g21347 and P2_R1131_U417 P2_R1131_U416 ; P2_R1131_U152
g21348 nand P2_R1131_U365 P2_R1131_U299 P2_R1131_U86 ; P2_R1131_U153
g21349 and P2_R1131_U424 P2_R1131_U423 ; P2_R1131_U154
g21350 nand P2_R1131_U293 P2_R1131_U292 ; P2_R1131_U155
g21351 and P2_R1131_U436 P2_R1131_U435 ; P2_R1131_U156
g21352 nand P2_R1131_U289 P2_R1131_U288 ; P2_R1131_U157
g21353 and P2_R1131_U443 P2_R1131_U442 ; P2_R1131_U158
g21354 nand P2_R1131_U132 P2_R1131_U284 ; P2_R1131_U159
g21355 and P2_R1131_U450 P2_R1131_U449 ; P2_R1131_U160
g21356 nand P2_R1131_U43 P2_R1131_U327 ; P2_R1131_U161
g21357 nand P2_R1131_U130 P2_R1131_U269 ; P2_R1131_U162
g21358 and P2_R1131_U476 P2_R1131_U475 ; P2_R1131_U163
g21359 nand P2_R1131_U257 P2_R1131_U256 ; P2_R1131_U164
g21360 and P2_R1131_U483 P2_R1131_U482 ; P2_R1131_U165
g21361 nand P2_R1131_U253 P2_R1131_U252 ; P2_R1131_U166
g21362 nand P2_R1131_U243 P2_R1131_U242 ; P2_R1131_U167
g21363 nand P2_R1131_U367 P2_R1131_U366 ; P2_R1131_U168
g21364 nand P2_U3056 P2_R1131_U151 ; P2_R1131_U169
g21365 not P2_R1131_U34 ; P2_R1131_U170
g21366 nand P2_U3456 P2_U3085 ; P2_R1131_U171
g21367 nand P2_U3074 P2_U3465 ; P2_R1131_U172
g21368 nand P2_U3060 P2_U3952 ; P2_R1131_U173
g21369 not P2_R1131_U68 ; P2_R1131_U174
g21370 not P2_R1131_U77 ; P2_R1131_U175
g21371 nand P2_U3067 P2_U3953 ; P2_R1131_U176
g21372 not P2_R1131_U61 ; P2_R1131_U177
g21373 or P2_U3069 P2_U3444 ; P2_R1131_U178
g21374 or P2_U3062 P2_U3441 ; P2_R1131_U179
g21375 or P2_U3438 P2_U3066 ; P2_R1131_U180
g21376 or P2_U3435 P2_U3070 ; P2_R1131_U181
g21377 not P2_R1131_U31 ; P2_R1131_U182
g21378 or P2_U3432 P2_U3080 ; P2_R1131_U183
g21379 not P2_R1131_U42 ; P2_R1131_U184
g21380 not P2_R1131_U43 ; P2_R1131_U185
g21381 nand P2_R1131_U42 P2_R1131_U43 ; P2_R1131_U186
g21382 nand P2_U3070 P2_U3435 ; P2_R1131_U187
g21383 nand P2_R1131_U186 P2_R1131_U181 ; P2_R1131_U188
g21384 nand P2_U3066 P2_U3438 ; P2_R1131_U189
g21385 nand P2_R1131_U115 P2_R1131_U188 ; P2_R1131_U190
g21386 nand P2_R1131_U35 P2_R1131_U34 ; P2_R1131_U191
g21387 nand P2_U3069 P2_R1131_U191 ; P2_R1131_U192
g21388 nand P2_R1131_U116 P2_R1131_U190 ; P2_R1131_U193
g21389 nand P2_U3444 P2_R1131_U170 ; P2_R1131_U194
g21390 not P2_R1131_U41 ; P2_R1131_U195
g21391 or P2_U3072 P2_U3450 ; P2_R1131_U196
g21392 or P2_U3073 P2_U3447 ; P2_R1131_U197
g21393 not P2_R1131_U22 ; P2_R1131_U198
g21394 nand P2_R1131_U23 P2_R1131_U22 ; P2_R1131_U199
g21395 nand P2_U3072 P2_R1131_U199 ; P2_R1131_U200
g21396 nand P2_U3450 P2_R1131_U198 ; P2_R1131_U201
g21397 nand P2_R1131_U5 P2_R1131_U41 ; P2_R1131_U202
g21398 not P2_R1131_U144 ; P2_R1131_U203
g21399 or P2_U3453 P2_U3086 ; P2_R1131_U204
g21400 nand P2_R1131_U204 P2_R1131_U144 ; P2_R1131_U205
g21401 not P2_R1131_U40 ; P2_R1131_U206
g21402 or P2_U3085 P2_U3456 ; P2_R1131_U207
g21403 or P2_U3447 P2_U3073 ; P2_R1131_U208
g21404 nand P2_R1131_U208 P2_R1131_U41 ; P2_R1131_U209
g21405 nand P2_R1131_U119 P2_R1131_U209 ; P2_R1131_U210
g21406 nand P2_R1131_U195 P2_R1131_U22 ; P2_R1131_U211
g21407 nand P2_U3450 P2_U3072 ; P2_R1131_U212
g21408 nand P2_R1131_U120 P2_R1131_U211 ; P2_R1131_U213
g21409 or P2_U3073 P2_U3447 ; P2_R1131_U214
g21410 nand P2_R1131_U185 P2_R1131_U181 ; P2_R1131_U215
g21411 nand P2_U3070 P2_U3435 ; P2_R1131_U216
g21412 not P2_R1131_U45 ; P2_R1131_U217
g21413 nand P2_R1131_U121 P2_R1131_U184 ; P2_R1131_U218
g21414 nand P2_R1131_U45 P2_R1131_U180 ; P2_R1131_U219
g21415 nand P2_U3066 P2_U3438 ; P2_R1131_U220
g21416 not P2_R1131_U44 ; P2_R1131_U221
g21417 or P2_U3441 P2_U3062 ; P2_R1131_U222
g21418 nand P2_R1131_U222 P2_R1131_U44 ; P2_R1131_U223
g21419 nand P2_R1131_U123 P2_R1131_U223 ; P2_R1131_U224
g21420 nand P2_R1131_U221 P2_R1131_U34 ; P2_R1131_U225
g21421 nand P2_U3444 P2_U3069 ; P2_R1131_U226
g21422 nand P2_R1131_U124 P2_R1131_U225 ; P2_R1131_U227
g21423 or P2_U3062 P2_U3441 ; P2_R1131_U228
g21424 nand P2_R1131_U184 P2_R1131_U181 ; P2_R1131_U229
g21425 not P2_R1131_U145 ; P2_R1131_U230
g21426 nand P2_U3066 P2_U3438 ; P2_R1131_U231
g21427 nand P2_R1131_U401 P2_R1131_U400 P2_R1131_U43 P2_R1131_U42 ; P2_R1131_U232
g21428 nand P2_R1131_U43 P2_R1131_U42 ; P2_R1131_U233
g21429 nand P2_U3070 P2_U3435 ; P2_R1131_U234
g21430 nand P2_R1131_U125 P2_R1131_U233 ; P2_R1131_U235
g21431 or P2_U3085 P2_U3456 ; P2_R1131_U236
g21432 or P2_U3064 P2_U3459 ; P2_R1131_U237
g21433 nand P2_R1131_U177 P2_R1131_U6 ; P2_R1131_U238
g21434 nand P2_U3064 P2_U3459 ; P2_R1131_U239
g21435 nand P2_R1131_U127 P2_R1131_U238 ; P2_R1131_U240
g21436 or P2_U3459 P2_U3064 ; P2_R1131_U241
g21437 nand P2_R1131_U126 P2_R1131_U144 ; P2_R1131_U242
g21438 nand P2_R1131_U241 P2_R1131_U240 ; P2_R1131_U243
g21439 not P2_R1131_U167 ; P2_R1131_U244
g21440 or P2_U3082 P2_U3468 ; P2_R1131_U245
g21441 or P2_U3074 P2_U3465 ; P2_R1131_U246
g21442 nand P2_R1131_U174 P2_R1131_U7 ; P2_R1131_U247
g21443 nand P2_U3082 P2_U3468 ; P2_R1131_U248
g21444 nand P2_R1131_U129 P2_R1131_U247 ; P2_R1131_U249
g21445 or P2_U3462 P2_U3065 ; P2_R1131_U250
g21446 or P2_U3468 P2_U3082 ; P2_R1131_U251
g21447 nand P2_R1131_U128 P2_R1131_U167 ; P2_R1131_U252
g21448 nand P2_R1131_U251 P2_R1131_U249 ; P2_R1131_U253
g21449 not P2_R1131_U166 ; P2_R1131_U254
g21450 or P2_U3471 P2_U3081 ; P2_R1131_U255
g21451 nand P2_R1131_U255 P2_R1131_U166 ; P2_R1131_U256
g21452 nand P2_U3081 P2_U3471 ; P2_R1131_U257
g21453 not P2_R1131_U164 ; P2_R1131_U258
g21454 or P2_U3474 P2_U3076 ; P2_R1131_U259
g21455 nand P2_R1131_U259 P2_R1131_U164 ; P2_R1131_U260
g21456 nand P2_U3076 P2_U3474 ; P2_R1131_U261
g21457 not P2_R1131_U92 ; P2_R1131_U262
g21458 or P2_U3071 P2_U3480 ; P2_R1131_U263
g21459 or P2_U3075 P2_U3477 ; P2_R1131_U264
g21460 not P2_R1131_U59 ; P2_R1131_U265
g21461 nand P2_R1131_U60 P2_R1131_U59 ; P2_R1131_U266
g21462 nand P2_U3071 P2_R1131_U266 ; P2_R1131_U267
g21463 nand P2_U3480 P2_R1131_U265 ; P2_R1131_U268
g21464 nand P2_R1131_U8 P2_R1131_U92 ; P2_R1131_U269
g21465 not P2_R1131_U162 ; P2_R1131_U270
g21466 or P2_U3078 P2_U3957 ; P2_R1131_U271
g21467 or P2_U3083 P2_U3485 ; P2_R1131_U272
g21468 or P2_U3077 P2_U3956 ; P2_R1131_U273
g21469 not P2_R1131_U80 ; P2_R1131_U274
g21470 nand P2_U3957 P2_R1131_U274 ; P2_R1131_U275
g21471 nand P2_R1131_U275 P2_R1131_U90 ; P2_R1131_U276
g21472 nand P2_R1131_U80 P2_R1131_U81 ; P2_R1131_U277
g21473 nand P2_R1131_U277 P2_R1131_U276 ; P2_R1131_U278
g21474 nand P2_R1131_U175 P2_R1131_U9 ; P2_R1131_U279
g21475 nand P2_U3077 P2_U3956 ; P2_R1131_U280
g21476 nand P2_R1131_U278 P2_R1131_U279 ; P2_R1131_U281
g21477 or P2_U3483 P2_U3084 ; P2_R1131_U282
g21478 or P2_U3956 P2_U3077 ; P2_R1131_U283
g21479 nand P2_R1131_U273 P2_R1131_U162 P2_R1131_U131 ; P2_R1131_U284
g21480 nand P2_R1131_U283 P2_R1131_U281 ; P2_R1131_U285
g21481 not P2_R1131_U159 ; P2_R1131_U286
g21482 or P2_U3955 P2_U3063 ; P2_R1131_U287
g21483 nand P2_R1131_U287 P2_R1131_U159 ; P2_R1131_U288
g21484 nand P2_U3063 P2_U3955 ; P2_R1131_U289
g21485 not P2_R1131_U157 ; P2_R1131_U290
g21486 or P2_U3954 P2_U3068 ; P2_R1131_U291
g21487 nand P2_R1131_U291 P2_R1131_U157 ; P2_R1131_U292
g21488 nand P2_U3068 P2_U3954 ; P2_R1131_U293
g21489 not P2_R1131_U155 ; P2_R1131_U294
g21490 or P2_U3060 P2_U3952 ; P2_R1131_U295
g21491 nand P2_R1131_U176 P2_R1131_U173 ; P2_R1131_U296
g21492 not P2_R1131_U86 ; P2_R1131_U297
g21493 or P2_U3953 P2_U3067 ; P2_R1131_U298
g21494 nand P2_R1131_U155 P2_R1131_U298 P2_R1131_U168 ; P2_R1131_U299
g21495 not P2_R1131_U153 ; P2_R1131_U300
g21496 or P2_U3950 P2_U3055 ; P2_R1131_U301
g21497 nand P2_U3055 P2_U3950 ; P2_R1131_U302
g21498 not P2_R1131_U151 ; P2_R1131_U303
g21499 nand P2_U3949 P2_R1131_U151 ; P2_R1131_U304
g21500 not P2_R1131_U149 ; P2_R1131_U305
g21501 nand P2_R1131_U298 P2_R1131_U155 ; P2_R1131_U306
g21502 not P2_R1131_U89 ; P2_R1131_U307
g21503 or P2_U3952 P2_U3060 ; P2_R1131_U308
g21504 nand P2_R1131_U308 P2_R1131_U89 ; P2_R1131_U309
g21505 nand P2_R1131_U309 P2_R1131_U173 P2_R1131_U154 ; P2_R1131_U310
g21506 nand P2_R1131_U307 P2_R1131_U173 ; P2_R1131_U311
g21507 nand P2_U3951 P2_U3059 ; P2_R1131_U312
g21508 nand P2_R1131_U311 P2_R1131_U312 P2_R1131_U168 ; P2_R1131_U313
g21509 or P2_U3060 P2_U3952 ; P2_R1131_U314
g21510 nand P2_R1131_U282 P2_R1131_U162 ; P2_R1131_U315
g21511 not P2_R1131_U91 ; P2_R1131_U316
g21512 nand P2_R1131_U9 P2_R1131_U91 ; P2_R1131_U317
g21513 nand P2_R1131_U135 P2_R1131_U317 ; P2_R1131_U318
g21514 nand P2_R1131_U317 P2_R1131_U278 ; P2_R1131_U319
g21515 nand P2_R1131_U453 P2_R1131_U319 ; P2_R1131_U320
g21516 or P2_U3485 P2_U3083 ; P2_R1131_U321
g21517 nand P2_R1131_U321 P2_R1131_U91 ; P2_R1131_U322
g21518 nand P2_R1131_U136 P2_R1131_U322 ; P2_R1131_U323
g21519 nand P2_R1131_U316 P2_R1131_U80 ; P2_R1131_U324
g21520 nand P2_U3078 P2_U3957 ; P2_R1131_U325
g21521 nand P2_R1131_U137 P2_R1131_U324 ; P2_R1131_U326
g21522 or P2_U3432 P2_U3080 ; P2_R1131_U327
g21523 not P2_R1131_U161 ; P2_R1131_U328
g21524 or P2_U3083 P2_U3485 ; P2_R1131_U329
g21525 or P2_U3477 P2_U3075 ; P2_R1131_U330
g21526 nand P2_R1131_U330 P2_R1131_U92 ; P2_R1131_U331
g21527 nand P2_R1131_U138 P2_R1131_U331 ; P2_R1131_U332
g21528 nand P2_R1131_U262 P2_R1131_U59 ; P2_R1131_U333
g21529 nand P2_U3480 P2_U3071 ; P2_R1131_U334
g21530 nand P2_R1131_U139 P2_R1131_U333 ; P2_R1131_U335
g21531 or P2_U3075 P2_U3477 ; P2_R1131_U336
g21532 nand P2_R1131_U250 P2_R1131_U167 ; P2_R1131_U337
g21533 not P2_R1131_U93 ; P2_R1131_U338
g21534 or P2_U3465 P2_U3074 ; P2_R1131_U339
g21535 nand P2_R1131_U339 P2_R1131_U93 ; P2_R1131_U340
g21536 nand P2_R1131_U140 P2_R1131_U340 ; P2_R1131_U341
g21537 nand P2_R1131_U338 P2_R1131_U172 ; P2_R1131_U342
g21538 nand P2_U3082 P2_U3468 ; P2_R1131_U343
g21539 nand P2_R1131_U141 P2_R1131_U342 ; P2_R1131_U344
g21540 or P2_U3074 P2_U3465 ; P2_R1131_U345
g21541 or P2_U3456 P2_U3085 ; P2_R1131_U346
g21542 nand P2_R1131_U346 P2_R1131_U40 ; P2_R1131_U347
g21543 nand P2_R1131_U142 P2_R1131_U347 ; P2_R1131_U348
g21544 nand P2_R1131_U206 P2_R1131_U171 ; P2_R1131_U349
g21545 nand P2_U3064 P2_U3459 ; P2_R1131_U350
g21546 nand P2_R1131_U143 P2_R1131_U349 ; P2_R1131_U351
g21547 nand P2_R1131_U207 P2_R1131_U171 ; P2_R1131_U352
g21548 nand P2_R1131_U204 P2_R1131_U61 ; P2_R1131_U353
g21549 nand P2_R1131_U214 P2_R1131_U22 ; P2_R1131_U354
g21550 nand P2_R1131_U228 P2_R1131_U34 ; P2_R1131_U355
g21551 nand P2_R1131_U231 P2_R1131_U180 ; P2_R1131_U356
g21552 nand P2_R1131_U314 P2_R1131_U173 ; P2_R1131_U357
g21553 nand P2_R1131_U298 P2_R1131_U176 ; P2_R1131_U358
g21554 nand P2_R1131_U329 P2_R1131_U80 ; P2_R1131_U359
g21555 nand P2_R1131_U282 P2_R1131_U77 ; P2_R1131_U360
g21556 nand P2_R1131_U336 P2_R1131_U59 ; P2_R1131_U361
g21557 nand P2_R1131_U345 P2_R1131_U172 ; P2_R1131_U362
g21558 nand P2_R1131_U250 P2_R1131_U68 ; P2_R1131_U363
g21559 nand P2_U3949 P2_U3056 ; P2_R1131_U364
g21560 nand P2_R1131_U296 P2_R1131_U168 ; P2_R1131_U365
g21561 nand P2_U3059 P2_R1131_U295 ; P2_R1131_U366
g21562 nand P2_U3951 P2_R1131_U295 ; P2_R1131_U367
g21563 nand P2_R1131_U296 P2_R1131_U168 P2_R1131_U301 ; P2_R1131_U368
g21564 nand P2_R1131_U155 P2_R1131_U168 P2_R1131_U133 ; P2_R1131_U369
g21565 nand P2_R1131_U297 P2_R1131_U301 ; P2_R1131_U370
g21566 nand P2_U3085 P2_R1131_U39 ; P2_R1131_U371
g21567 nand P2_U3456 P2_R1131_U38 ; P2_R1131_U372
g21568 nand P2_R1131_U372 P2_R1131_U371 ; P2_R1131_U373
g21569 nand P2_R1131_U352 P2_R1131_U40 ; P2_R1131_U374
g21570 nand P2_R1131_U373 P2_R1131_U206 ; P2_R1131_U375
g21571 nand P2_U3086 P2_R1131_U36 ; P2_R1131_U376
g21572 nand P2_U3453 P2_R1131_U37 ; P2_R1131_U377
g21573 nand P2_R1131_U377 P2_R1131_U376 ; P2_R1131_U378
g21574 nand P2_R1131_U353 P2_R1131_U144 ; P2_R1131_U379
g21575 nand P2_R1131_U203 P2_R1131_U378 ; P2_R1131_U380
g21576 nand P2_U3072 P2_R1131_U23 ; P2_R1131_U381
g21577 nand P2_U3450 P2_R1131_U21 ; P2_R1131_U382
g21578 nand P2_U3073 P2_R1131_U19 ; P2_R1131_U383
g21579 nand P2_U3447 P2_R1131_U20 ; P2_R1131_U384
g21580 nand P2_R1131_U384 P2_R1131_U383 ; P2_R1131_U385
g21581 nand P2_R1131_U354 P2_R1131_U41 ; P2_R1131_U386
g21582 nand P2_R1131_U385 P2_R1131_U195 ; P2_R1131_U387
g21583 nand P2_U3069 P2_R1131_U35 ; P2_R1131_U388
g21584 nand P2_U3444 P2_R1131_U26 ; P2_R1131_U389
g21585 nand P2_U3062 P2_R1131_U24 ; P2_R1131_U390
g21586 nand P2_U3441 P2_R1131_U25 ; P2_R1131_U391
g21587 nand P2_R1131_U391 P2_R1131_U390 ; P2_R1131_U392
g21588 nand P2_R1131_U355 P2_R1131_U44 ; P2_R1131_U393
g21589 nand P2_R1131_U392 P2_R1131_U221 ; P2_R1131_U394
g21590 nand P2_U3066 P2_R1131_U32 ; P2_R1131_U395
g21591 nand P2_U3438 P2_R1131_U33 ; P2_R1131_U396
g21592 nand P2_R1131_U396 P2_R1131_U395 ; P2_R1131_U397
g21593 nand P2_R1131_U356 P2_R1131_U145 ; P2_R1131_U398
g21594 nand P2_R1131_U230 P2_R1131_U397 ; P2_R1131_U399
g21595 nand P2_U3070 P2_R1131_U27 ; P2_R1131_U400
g21596 nand P2_U3435 P2_R1131_U28 ; P2_R1131_U401
g21597 nand P2_U3057 P2_R1131_U147 ; P2_R1131_U402
g21598 nand P2_U3960 P2_R1131_U146 ; P2_R1131_U403
g21599 nand P2_U3057 P2_R1131_U147 ; P2_R1131_U404
g21600 nand P2_U3960 P2_R1131_U146 ; P2_R1131_U405
g21601 nand P2_R1131_U405 P2_R1131_U404 ; P2_R1131_U406
g21602 nand P2_R1131_U148 P2_R1131_U149 ; P2_R1131_U407
g21603 nand P2_R1131_U305 P2_R1131_U406 ; P2_R1131_U408
g21604 nand P2_U3056 P2_R1131_U88 ; P2_R1131_U409
g21605 nand P2_U3949 P2_R1131_U87 ; P2_R1131_U410
g21606 nand P2_U3056 P2_R1131_U88 ; P2_R1131_U411
g21607 nand P2_U3949 P2_R1131_U87 ; P2_R1131_U412
g21608 nand P2_R1131_U412 P2_R1131_U411 ; P2_R1131_U413
g21609 nand P2_R1131_U150 P2_R1131_U151 ; P2_R1131_U414
g21610 nand P2_R1131_U303 P2_R1131_U413 ; P2_R1131_U415
g21611 nand P2_U3055 P2_R1131_U46 ; P2_R1131_U416
g21612 nand P2_U3950 P2_R1131_U47 ; P2_R1131_U417
g21613 nand P2_U3055 P2_R1131_U46 ; P2_R1131_U418
g21614 nand P2_U3950 P2_R1131_U47 ; P2_R1131_U419
g21615 nand P2_R1131_U419 P2_R1131_U418 ; P2_R1131_U420
g21616 nand P2_R1131_U152 P2_R1131_U153 ; P2_R1131_U421
g21617 nand P2_R1131_U300 P2_R1131_U420 ; P2_R1131_U422
g21618 nand P2_U3059 P2_R1131_U49 ; P2_R1131_U423
g21619 nand P2_U3951 P2_R1131_U48 ; P2_R1131_U424
g21620 nand P2_U3060 P2_R1131_U50 ; P2_R1131_U425
g21621 nand P2_U3952 P2_R1131_U51 ; P2_R1131_U426
g21622 nand P2_R1131_U426 P2_R1131_U425 ; P2_R1131_U427
g21623 nand P2_R1131_U357 P2_R1131_U89 ; P2_R1131_U428
g21624 nand P2_R1131_U427 P2_R1131_U307 ; P2_R1131_U429
g21625 nand P2_U3067 P2_R1131_U52 ; P2_R1131_U430
g21626 nand P2_U3953 P2_R1131_U53 ; P2_R1131_U431
g21627 nand P2_R1131_U431 P2_R1131_U430 ; P2_R1131_U432
g21628 nand P2_R1131_U358 P2_R1131_U155 ; P2_R1131_U433
g21629 nand P2_R1131_U294 P2_R1131_U432 ; P2_R1131_U434
g21630 nand P2_U3068 P2_R1131_U84 ; P2_R1131_U435
g21631 nand P2_U3954 P2_R1131_U85 ; P2_R1131_U436
g21632 nand P2_U3068 P2_R1131_U84 ; P2_R1131_U437
g21633 nand P2_U3954 P2_R1131_U85 ; P2_R1131_U438
g21634 nand P2_R1131_U438 P2_R1131_U437 ; P2_R1131_U439
g21635 nand P2_R1131_U156 P2_R1131_U157 ; P2_R1131_U440
g21636 nand P2_R1131_U290 P2_R1131_U439 ; P2_R1131_U441
g21637 nand P2_U3063 P2_R1131_U82 ; P2_R1131_U442
g21638 nand P2_U3955 P2_R1131_U83 ; P2_R1131_U443
g21639 nand P2_U3063 P2_R1131_U82 ; P2_R1131_U444
g21640 nand P2_U3955 P2_R1131_U83 ; P2_R1131_U445
g21641 nand P2_R1131_U445 P2_R1131_U444 ; P2_R1131_U446
g21642 nand P2_R1131_U158 P2_R1131_U159 ; P2_R1131_U447
g21643 nand P2_R1131_U286 P2_R1131_U446 ; P2_R1131_U448
g21644 nand P2_U3077 P2_R1131_U54 ; P2_R1131_U449
g21645 nand P2_U3956 P2_R1131_U55 ; P2_R1131_U450
g21646 nand P2_U3077 P2_R1131_U54 ; P2_R1131_U451
g21647 nand P2_U3956 P2_R1131_U55 ; P2_R1131_U452
g21648 nand P2_R1131_U452 P2_R1131_U451 ; P2_R1131_U453
g21649 nand P2_U3078 P2_R1131_U81 ; P2_R1131_U454
g21650 nand P2_U3957 P2_R1131_U90 ; P2_R1131_U455
g21651 nand P2_R1131_U182 P2_R1131_U161 ; P2_R1131_U456
g21652 nand P2_R1131_U328 P2_R1131_U31 ; P2_R1131_U457
g21653 nand P2_U3083 P2_R1131_U78 ; P2_R1131_U458
g21654 nand P2_U3485 P2_R1131_U79 ; P2_R1131_U459
g21655 nand P2_R1131_U459 P2_R1131_U458 ; P2_R1131_U460
g21656 nand P2_R1131_U359 P2_R1131_U91 ; P2_R1131_U461
g21657 nand P2_R1131_U460 P2_R1131_U316 ; P2_R1131_U462
g21658 nand P2_U3084 P2_R1131_U75 ; P2_R1131_U463
g21659 nand P2_U3483 P2_R1131_U76 ; P2_R1131_U464
g21660 nand P2_R1131_U464 P2_R1131_U463 ; P2_R1131_U465
g21661 nand P2_R1131_U360 P2_R1131_U162 ; P2_R1131_U466
g21662 nand P2_R1131_U270 P2_R1131_U465 ; P2_R1131_U467
g21663 nand P2_U3071 P2_R1131_U60 ; P2_R1131_U468
g21664 nand P2_U3480 P2_R1131_U58 ; P2_R1131_U469
g21665 nand P2_U3075 P2_R1131_U56 ; P2_R1131_U470
g21666 nand P2_U3477 P2_R1131_U57 ; P2_R1131_U471
g21667 nand P2_R1131_U471 P2_R1131_U470 ; P2_R1131_U472
g21668 nand P2_R1131_U361 P2_R1131_U92 ; P2_R1131_U473
g21669 nand P2_R1131_U472 P2_R1131_U262 ; P2_R1131_U474
g21670 nand P2_U3076 P2_R1131_U73 ; P2_R1131_U475
g21671 nand P2_U3474 P2_R1131_U74 ; P2_R1131_U476
g21672 nand P2_U3076 P2_R1131_U73 ; P2_R1131_U477
g21673 nand P2_U3474 P2_R1131_U74 ; P2_R1131_U478
g21674 nand P2_R1131_U478 P2_R1131_U477 ; P2_R1131_U479
g21675 nand P2_R1131_U163 P2_R1131_U164 ; P2_R1131_U480
g21676 nand P2_R1131_U258 P2_R1131_U479 ; P2_R1131_U481
g21677 nand P2_U3081 P2_R1131_U71 ; P2_R1131_U482
g21678 nand P2_U3471 P2_R1131_U72 ; P2_R1131_U483
g21679 nand P2_U3081 P2_R1131_U71 ; P2_R1131_U484
g21680 nand P2_U3471 P2_R1131_U72 ; P2_R1131_U485
g21681 nand P2_R1131_U485 P2_R1131_U484 ; P2_R1131_U486
g21682 nand P2_R1131_U165 P2_R1131_U166 ; P2_R1131_U487
g21683 nand P2_R1131_U254 P2_R1131_U486 ; P2_R1131_U488
g21684 nand P2_U3082 P2_R1131_U69 ; P2_R1131_U489
g21685 nand P2_U3468 P2_R1131_U70 ; P2_R1131_U490
g21686 nand P2_U3074 P2_R1131_U64 ; P2_R1131_U491
g21687 nand P2_U3465 P2_R1131_U65 ; P2_R1131_U492
g21688 nand P2_R1131_U492 P2_R1131_U491 ; P2_R1131_U493
g21689 nand P2_R1131_U362 P2_R1131_U93 ; P2_R1131_U494
g21690 nand P2_R1131_U493 P2_R1131_U338 ; P2_R1131_U495
g21691 nand P2_U3065 P2_R1131_U66 ; P2_R1131_U496
g21692 nand P2_U3462 P2_R1131_U67 ; P2_R1131_U497
g21693 nand P2_R1131_U497 P2_R1131_U496 ; P2_R1131_U498
g21694 nand P2_R1131_U363 P2_R1131_U167 ; P2_R1131_U499
g21695 nand P2_R1131_U244 P2_R1131_U498 ; P2_R1131_U500
g21696 nand P2_U3064 P2_R1131_U62 ; P2_R1131_U501
g21697 nand P2_U3459 P2_R1131_U63 ; P2_R1131_U502
g21698 nand P2_U3079 P2_R1131_U29 ; P2_R1131_U503
g21699 nand P2_U3427 P2_R1131_U30 ; P2_R1131_U504
g21700 and P2_R1146_U202 P2_R1146_U201 ; P2_R1146_U6
g21701 and P2_R1146_U241 P2_R1146_U240 ; P2_R1146_U7
g21702 and P2_R1146_U181 P2_R1146_U256 ; P2_R1146_U8
g21703 and P2_R1146_U258 P2_R1146_U257 ; P2_R1146_U9
g21704 and P2_R1146_U182 P2_R1146_U282 ; P2_R1146_U10
g21705 and P2_R1146_U284 P2_R1146_U283 ; P2_R1146_U11
g21706 nand P2_R1146_U344 P2_R1146_U347 ; P2_R1146_U12
g21707 nand P2_R1146_U333 P2_R1146_U336 ; P2_R1146_U13
g21708 nand P2_R1146_U322 P2_R1146_U325 ; P2_R1146_U14
g21709 nand P2_R1146_U314 P2_R1146_U316 ; P2_R1146_U15
g21710 nand P2_R1146_U352 P2_R1146_U312 ; P2_R1146_U16
g21711 nand P2_R1146_U235 P2_R1146_U237 ; P2_R1146_U17
g21712 nand P2_R1146_U227 P2_R1146_U230 ; P2_R1146_U18
g21713 nand P2_R1146_U219 P2_R1146_U221 ; P2_R1146_U19
g21714 nand P2_R1146_U166 P2_R1146_U350 ; P2_R1146_U20
g21715 not P2_U3450 ; P2_R1146_U21
g21716 not P2_U3444 ; P2_R1146_U22
g21717 not P2_U3435 ; P2_R1146_U23
g21718 not P2_U3427 ; P2_R1146_U24
g21719 not P2_U3080 ; P2_R1146_U25
g21720 not P2_U3438 ; P2_R1146_U26
g21721 not P2_U3070 ; P2_R1146_U27
g21722 nand P2_U3070 P2_R1146_U23 ; P2_R1146_U28
g21723 not P2_U3066 ; P2_R1146_U29
g21724 not P2_U3447 ; P2_R1146_U30
g21725 not P2_U3441 ; P2_R1146_U31
g21726 not P2_U3073 ; P2_R1146_U32
g21727 not P2_U3069 ; P2_R1146_U33
g21728 not P2_U3062 ; P2_R1146_U34
g21729 nand P2_U3062 P2_R1146_U31 ; P2_R1146_U35
g21730 not P2_U3453 ; P2_R1146_U36
g21731 not P2_U3072 ; P2_R1146_U37
g21732 nand P2_U3072 P2_R1146_U21 ; P2_R1146_U38
g21733 not P2_U3086 ; P2_R1146_U39
g21734 not P2_U3456 ; P2_R1146_U40
g21735 not P2_U3085 ; P2_R1146_U41
g21736 nand P2_R1146_U208 P2_R1146_U207 ; P2_R1146_U42
g21737 nand P2_R1146_U35 P2_R1146_U223 ; P2_R1146_U43
g21738 nand P2_R1146_U192 P2_R1146_U176 P2_R1146_U351 ; P2_R1146_U44
g21739 not P2_U3951 ; P2_R1146_U45
g21740 not P2_U3459 ; P2_R1146_U46
g21741 not P2_U3462 ; P2_R1146_U47
g21742 not P2_U3065 ; P2_R1146_U48
g21743 not P2_U3064 ; P2_R1146_U49
g21744 nand P2_U3085 P2_R1146_U40 ; P2_R1146_U50
g21745 not P2_U3465 ; P2_R1146_U51
g21746 not P2_U3074 ; P2_R1146_U52
g21747 not P2_U3468 ; P2_R1146_U53
g21748 not P2_U3082 ; P2_R1146_U54
g21749 not P2_U3477 ; P2_R1146_U55
g21750 not P2_U3474 ; P2_R1146_U56
g21751 not P2_U3471 ; P2_R1146_U57
g21752 not P2_U3075 ; P2_R1146_U58
g21753 not P2_U3076 ; P2_R1146_U59
g21754 not P2_U3081 ; P2_R1146_U60
g21755 nand P2_U3081 P2_R1146_U57 ; P2_R1146_U61
g21756 not P2_U3480 ; P2_R1146_U62
g21757 not P2_U3071 ; P2_R1146_U63
g21758 nand P2_R1146_U268 P2_R1146_U267 ; P2_R1146_U64
g21759 not P2_U3084 ; P2_R1146_U65
g21760 not P2_U3485 ; P2_R1146_U66
g21761 not P2_U3083 ; P2_R1146_U67
g21762 not P2_U3957 ; P2_R1146_U68
g21763 not P2_U3078 ; P2_R1146_U69
g21764 not P2_U3954 ; P2_R1146_U70
g21765 not P2_U3955 ; P2_R1146_U71
g21766 not P2_U3956 ; P2_R1146_U72
g21767 not P2_U3068 ; P2_R1146_U73
g21768 not P2_U3063 ; P2_R1146_U74
g21769 not P2_U3077 ; P2_R1146_U75
g21770 nand P2_U3077 P2_R1146_U72 ; P2_R1146_U76
g21771 not P2_U3953 ; P2_R1146_U77
g21772 not P2_U3067 ; P2_R1146_U78
g21773 not P2_U3952 ; P2_R1146_U79
g21774 not P2_U3060 ; P2_R1146_U80
g21775 not P2_U3950 ; P2_R1146_U81
g21776 not P2_U3059 ; P2_R1146_U82
g21777 nand P2_U3059 P2_R1146_U45 ; P2_R1146_U83
g21778 not P2_U3055 ; P2_R1146_U84
g21779 not P2_U3949 ; P2_R1146_U85
g21780 not P2_U3056 ; P2_R1146_U86
g21781 nand P2_R1146_U128 P2_R1146_U301 ; P2_R1146_U87
g21782 nand P2_R1146_U298 P2_R1146_U297 ; P2_R1146_U88
g21783 nand P2_R1146_U76 P2_R1146_U318 ; P2_R1146_U89
g21784 nand P2_R1146_U61 P2_R1146_U329 ; P2_R1146_U90
g21785 nand P2_R1146_U50 P2_R1146_U340 ; P2_R1146_U91
g21786 not P2_U3079 ; P2_R1146_U92
g21787 nand P2_R1146_U395 P2_R1146_U394 ; P2_R1146_U93
g21788 nand P2_R1146_U409 P2_R1146_U408 ; P2_R1146_U94
g21789 nand P2_R1146_U414 P2_R1146_U413 ; P2_R1146_U95
g21790 nand P2_R1146_U430 P2_R1146_U429 ; P2_R1146_U96
g21791 nand P2_R1146_U435 P2_R1146_U434 ; P2_R1146_U97
g21792 nand P2_R1146_U440 P2_R1146_U439 ; P2_R1146_U98
g21793 nand P2_R1146_U445 P2_R1146_U444 ; P2_R1146_U99
g21794 nand P2_R1146_U450 P2_R1146_U449 ; P2_R1146_U100
g21795 nand P2_R1146_U466 P2_R1146_U465 ; P2_R1146_U101
g21796 nand P2_R1146_U471 P2_R1146_U470 ; P2_R1146_U102
g21797 nand P2_R1146_U356 P2_R1146_U355 ; P2_R1146_U103
g21798 nand P2_R1146_U365 P2_R1146_U364 ; P2_R1146_U104
g21799 nand P2_R1146_U372 P2_R1146_U371 ; P2_R1146_U105
g21800 nand P2_R1146_U376 P2_R1146_U375 ; P2_R1146_U106
g21801 nand P2_R1146_U385 P2_R1146_U384 ; P2_R1146_U107
g21802 nand P2_R1146_U404 P2_R1146_U403 ; P2_R1146_U108
g21803 nand P2_R1146_U421 P2_R1146_U420 ; P2_R1146_U109
g21804 nand P2_R1146_U425 P2_R1146_U424 ; P2_R1146_U110
g21805 nand P2_R1146_U457 P2_R1146_U456 ; P2_R1146_U111
g21806 nand P2_R1146_U461 P2_R1146_U460 ; P2_R1146_U112
g21807 nand P2_R1146_U478 P2_R1146_U477 ; P2_R1146_U113
g21808 and P2_R1146_U194 P2_R1146_U184 ; P2_R1146_U114
g21809 and P2_R1146_U197 P2_R1146_U198 ; P2_R1146_U115
g21810 and P2_R1146_U205 P2_R1146_U200 P2_R1146_U185 ; P2_R1146_U116
g21811 and P2_R1146_U210 P2_R1146_U186 ; P2_R1146_U117
g21812 and P2_R1146_U213 P2_R1146_U214 ; P2_R1146_U118
g21813 and P2_R1146_U358 P2_R1146_U357 P2_R1146_U38 ; P2_R1146_U119
g21814 and P2_R1146_U361 P2_R1146_U186 ; P2_R1146_U120
g21815 and P2_R1146_U229 P2_R1146_U6 ; P2_R1146_U121
g21816 and P2_R1146_U368 P2_R1146_U185 ; P2_R1146_U122
g21817 and P2_R1146_U378 P2_R1146_U377 P2_R1146_U28 ; P2_R1146_U123
g21818 and P2_R1146_U381 P2_R1146_U184 ; P2_R1146_U124
g21819 and P2_R1146_U239 P2_R1146_U216 P2_R1146_U180 ; P2_R1146_U125
g21820 and P2_R1146_U261 P2_R1146_U8 ; P2_R1146_U126
g21821 and P2_R1146_U287 P2_R1146_U10 ; P2_R1146_U127
g21822 and P2_R1146_U303 P2_R1146_U304 ; P2_R1146_U128
g21823 and P2_R1146_U387 P2_R1146_U386 P2_R1146_U311 ; P2_R1146_U129
g21824 and P2_R1146_U308 P2_R1146_U390 ; P2_R1146_U130
g21825 nand P2_R1146_U392 P2_R1146_U391 ; P2_R1146_U131
g21826 and P2_R1146_U397 P2_R1146_U396 P2_R1146_U83 ; P2_R1146_U132
g21827 and P2_R1146_U400 P2_R1146_U183 ; P2_R1146_U133
g21828 nand P2_R1146_U406 P2_R1146_U405 ; P2_R1146_U134
g21829 nand P2_R1146_U411 P2_R1146_U410 ; P2_R1146_U135
g21830 and P2_R1146_U324 P2_R1146_U11 ; P2_R1146_U136
g21831 and P2_R1146_U417 P2_R1146_U182 ; P2_R1146_U137
g21832 nand P2_R1146_U427 P2_R1146_U426 ; P2_R1146_U138
g21833 nand P2_R1146_U432 P2_R1146_U431 ; P2_R1146_U139
g21834 nand P2_R1146_U437 P2_R1146_U436 ; P2_R1146_U140
g21835 nand P2_R1146_U442 P2_R1146_U441 ; P2_R1146_U141
g21836 nand P2_R1146_U447 P2_R1146_U446 ; P2_R1146_U142
g21837 and P2_R1146_U335 P2_R1146_U9 ; P2_R1146_U143
g21838 and P2_R1146_U453 P2_R1146_U181 ; P2_R1146_U144
g21839 nand P2_R1146_U463 P2_R1146_U462 ; P2_R1146_U145
g21840 nand P2_R1146_U468 P2_R1146_U467 ; P2_R1146_U146
g21841 and P2_R1146_U346 P2_R1146_U7 ; P2_R1146_U147
g21842 and P2_R1146_U474 P2_R1146_U180 ; P2_R1146_U148
g21843 and P2_R1146_U354 P2_R1146_U353 ; P2_R1146_U149
g21844 nand P2_R1146_U118 P2_R1146_U211 ; P2_R1146_U150
g21845 and P2_R1146_U363 P2_R1146_U362 ; P2_R1146_U151
g21846 and P2_R1146_U370 P2_R1146_U369 ; P2_R1146_U152
g21847 and P2_R1146_U374 P2_R1146_U373 ; P2_R1146_U153
g21848 nand P2_R1146_U115 P2_R1146_U195 ; P2_R1146_U154
g21849 and P2_R1146_U383 P2_R1146_U382 ; P2_R1146_U155
g21850 not P2_U3960 ; P2_R1146_U156
g21851 not P2_U3057 ; P2_R1146_U157
g21852 and P2_R1146_U402 P2_R1146_U401 ; P2_R1146_U158
g21853 nand P2_R1146_U294 P2_R1146_U293 ; P2_R1146_U159
g21854 nand P2_R1146_U290 P2_R1146_U289 ; P2_R1146_U160
g21855 and P2_R1146_U419 P2_R1146_U418 ; P2_R1146_U161
g21856 and P2_R1146_U423 P2_R1146_U422 ; P2_R1146_U162
g21857 nand P2_R1146_U280 P2_R1146_U279 ; P2_R1146_U163
g21858 nand P2_R1146_U276 P2_R1146_U275 ; P2_R1146_U164
g21859 not P2_U3432 ; P2_R1146_U165
g21860 nand P2_U3427 P2_R1146_U92 ; P2_R1146_U166
g21861 nand P2_R1146_U272 P2_R1146_U271 ; P2_R1146_U167
g21862 not P2_U3483 ; P2_R1146_U168
g21863 nand P2_R1146_U264 P2_R1146_U263 ; P2_R1146_U169
g21864 and P2_R1146_U455 P2_R1146_U454 ; P2_R1146_U170
g21865 and P2_R1146_U459 P2_R1146_U458 ; P2_R1146_U171
g21866 nand P2_R1146_U254 P2_R1146_U253 ; P2_R1146_U172
g21867 nand P2_R1146_U250 P2_R1146_U249 ; P2_R1146_U173
g21868 nand P2_R1146_U246 P2_R1146_U245 ; P2_R1146_U174
g21869 and P2_R1146_U476 P2_R1146_U475 ; P2_R1146_U175
g21870 nand P2_R1146_U166 P2_R1146_U165 ; P2_R1146_U176
g21871 not P2_R1146_U83 ; P2_R1146_U177
g21872 not P2_R1146_U28 ; P2_R1146_U178
g21873 not P2_R1146_U38 ; P2_R1146_U179
g21874 nand P2_U3459 P2_R1146_U49 ; P2_R1146_U180
g21875 nand P2_U3474 P2_R1146_U59 ; P2_R1146_U181
g21876 nand P2_U3955 P2_R1146_U74 ; P2_R1146_U182
g21877 nand P2_U3951 P2_R1146_U82 ; P2_R1146_U183
g21878 nand P2_U3435 P2_R1146_U27 ; P2_R1146_U184
g21879 nand P2_U3444 P2_R1146_U33 ; P2_R1146_U185
g21880 nand P2_U3450 P2_R1146_U37 ; P2_R1146_U186
g21881 not P2_R1146_U61 ; P2_R1146_U187
g21882 not P2_R1146_U76 ; P2_R1146_U188
g21883 not P2_R1146_U35 ; P2_R1146_U189
g21884 not P2_R1146_U50 ; P2_R1146_U190
g21885 not P2_R1146_U166 ; P2_R1146_U191
g21886 nand P2_U3080 P2_R1146_U166 ; P2_R1146_U192
g21887 not P2_R1146_U44 ; P2_R1146_U193
g21888 nand P2_U3438 P2_R1146_U29 ; P2_R1146_U194
g21889 nand P2_R1146_U114 P2_R1146_U44 ; P2_R1146_U195
g21890 nand P2_R1146_U29 P2_R1146_U28 ; P2_R1146_U196
g21891 nand P2_R1146_U196 P2_R1146_U26 ; P2_R1146_U197
g21892 nand P2_U3066 P2_R1146_U178 ; P2_R1146_U198
g21893 not P2_R1146_U154 ; P2_R1146_U199
g21894 nand P2_U3447 P2_R1146_U32 ; P2_R1146_U200
g21895 nand P2_U3073 P2_R1146_U30 ; P2_R1146_U201
g21896 nand P2_U3069 P2_R1146_U22 ; P2_R1146_U202
g21897 nand P2_R1146_U189 P2_R1146_U185 ; P2_R1146_U203
g21898 nand P2_R1146_U6 P2_R1146_U203 ; P2_R1146_U204
g21899 nand P2_U3441 P2_R1146_U34 ; P2_R1146_U205
g21900 nand P2_U3447 P2_R1146_U32 ; P2_R1146_U206
g21901 nand P2_R1146_U154 P2_R1146_U116 ; P2_R1146_U207
g21902 nand P2_R1146_U206 P2_R1146_U204 ; P2_R1146_U208
g21903 not P2_R1146_U42 ; P2_R1146_U209
g21904 nand P2_U3453 P2_R1146_U39 ; P2_R1146_U210
g21905 nand P2_R1146_U117 P2_R1146_U42 ; P2_R1146_U211
g21906 nand P2_R1146_U39 P2_R1146_U38 ; P2_R1146_U212
g21907 nand P2_R1146_U212 P2_R1146_U36 ; P2_R1146_U213
g21908 nand P2_U3086 P2_R1146_U179 ; P2_R1146_U214
g21909 not P2_R1146_U150 ; P2_R1146_U215
g21910 nand P2_U3456 P2_R1146_U41 ; P2_R1146_U216
g21911 nand P2_R1146_U216 P2_R1146_U50 ; P2_R1146_U217
g21912 nand P2_R1146_U209 P2_R1146_U38 ; P2_R1146_U218
g21913 nand P2_R1146_U120 P2_R1146_U218 ; P2_R1146_U219
g21914 nand P2_R1146_U42 P2_R1146_U186 ; P2_R1146_U220
g21915 nand P2_R1146_U119 P2_R1146_U220 ; P2_R1146_U221
g21916 nand P2_R1146_U38 P2_R1146_U186 ; P2_R1146_U222
g21917 nand P2_R1146_U205 P2_R1146_U154 ; P2_R1146_U223
g21918 not P2_R1146_U43 ; P2_R1146_U224
g21919 nand P2_U3069 P2_R1146_U22 ; P2_R1146_U225
g21920 nand P2_R1146_U224 P2_R1146_U225 ; P2_R1146_U226
g21921 nand P2_R1146_U122 P2_R1146_U226 ; P2_R1146_U227
g21922 nand P2_R1146_U43 P2_R1146_U185 ; P2_R1146_U228
g21923 nand P2_U3447 P2_R1146_U32 ; P2_R1146_U229
g21924 nand P2_R1146_U121 P2_R1146_U228 ; P2_R1146_U230
g21925 nand P2_U3069 P2_R1146_U22 ; P2_R1146_U231
g21926 nand P2_R1146_U185 P2_R1146_U231 ; P2_R1146_U232
g21927 nand P2_R1146_U205 P2_R1146_U35 ; P2_R1146_U233
g21928 nand P2_R1146_U193 P2_R1146_U28 ; P2_R1146_U234
g21929 nand P2_R1146_U124 P2_R1146_U234 ; P2_R1146_U235
g21930 nand P2_R1146_U44 P2_R1146_U184 ; P2_R1146_U236
g21931 nand P2_R1146_U123 P2_R1146_U236 ; P2_R1146_U237
g21932 nand P2_R1146_U28 P2_R1146_U184 ; P2_R1146_U238
g21933 nand P2_U3462 P2_R1146_U48 ; P2_R1146_U239
g21934 nand P2_U3065 P2_R1146_U47 ; P2_R1146_U240
g21935 nand P2_U3064 P2_R1146_U46 ; P2_R1146_U241
g21936 nand P2_R1146_U190 P2_R1146_U180 ; P2_R1146_U242
g21937 nand P2_R1146_U7 P2_R1146_U242 ; P2_R1146_U243
g21938 nand P2_U3462 P2_R1146_U48 ; P2_R1146_U244
g21939 nand P2_R1146_U150 P2_R1146_U125 ; P2_R1146_U245
g21940 nand P2_R1146_U244 P2_R1146_U243 ; P2_R1146_U246
g21941 not P2_R1146_U174 ; P2_R1146_U247
g21942 nand P2_U3465 P2_R1146_U52 ; P2_R1146_U248
g21943 nand P2_R1146_U248 P2_R1146_U174 ; P2_R1146_U249
g21944 nand P2_U3074 P2_R1146_U51 ; P2_R1146_U250
g21945 not P2_R1146_U173 ; P2_R1146_U251
g21946 nand P2_U3468 P2_R1146_U54 ; P2_R1146_U252
g21947 nand P2_R1146_U252 P2_R1146_U173 ; P2_R1146_U253
g21948 nand P2_U3082 P2_R1146_U53 ; P2_R1146_U254
g21949 not P2_R1146_U172 ; P2_R1146_U255
g21950 nand P2_U3477 P2_R1146_U58 ; P2_R1146_U256
g21951 nand P2_U3075 P2_R1146_U55 ; P2_R1146_U257
g21952 nand P2_U3076 P2_R1146_U56 ; P2_R1146_U258
g21953 nand P2_R1146_U187 P2_R1146_U8 ; P2_R1146_U259
g21954 nand P2_R1146_U9 P2_R1146_U259 ; P2_R1146_U260
g21955 nand P2_U3471 P2_R1146_U60 ; P2_R1146_U261
g21956 nand P2_U3477 P2_R1146_U58 ; P2_R1146_U262
g21957 nand P2_R1146_U126 P2_R1146_U172 ; P2_R1146_U263
g21958 nand P2_R1146_U262 P2_R1146_U260 ; P2_R1146_U264
g21959 not P2_R1146_U169 ; P2_R1146_U265
g21960 nand P2_U3480 P2_R1146_U63 ; P2_R1146_U266
g21961 nand P2_R1146_U266 P2_R1146_U169 ; P2_R1146_U267
g21962 nand P2_U3071 P2_R1146_U62 ; P2_R1146_U268
g21963 not P2_R1146_U64 ; P2_R1146_U269
g21964 nand P2_R1146_U269 P2_R1146_U65 ; P2_R1146_U270
g21965 nand P2_R1146_U270 P2_R1146_U168 ; P2_R1146_U271
g21966 nand P2_U3084 P2_R1146_U64 ; P2_R1146_U272
g21967 not P2_R1146_U167 ; P2_R1146_U273
g21968 nand P2_U3485 P2_R1146_U67 ; P2_R1146_U274
g21969 nand P2_R1146_U274 P2_R1146_U167 ; P2_R1146_U275
g21970 nand P2_U3083 P2_R1146_U66 ; P2_R1146_U276
g21971 not P2_R1146_U164 ; P2_R1146_U277
g21972 nand P2_U3957 P2_R1146_U69 ; P2_R1146_U278
g21973 nand P2_R1146_U278 P2_R1146_U164 ; P2_R1146_U279
g21974 nand P2_U3078 P2_R1146_U68 ; P2_R1146_U280
g21975 not P2_R1146_U163 ; P2_R1146_U281
g21976 nand P2_U3954 P2_R1146_U73 ; P2_R1146_U282
g21977 nand P2_U3068 P2_R1146_U70 ; P2_R1146_U283
g21978 nand P2_U3063 P2_R1146_U71 ; P2_R1146_U284
g21979 nand P2_R1146_U188 P2_R1146_U10 ; P2_R1146_U285
g21980 nand P2_R1146_U11 P2_R1146_U285 ; P2_R1146_U286
g21981 nand P2_U3956 P2_R1146_U75 ; P2_R1146_U287
g21982 nand P2_U3954 P2_R1146_U73 ; P2_R1146_U288
g21983 nand P2_R1146_U127 P2_R1146_U163 ; P2_R1146_U289
g21984 nand P2_R1146_U288 P2_R1146_U286 ; P2_R1146_U290
g21985 not P2_R1146_U160 ; P2_R1146_U291
g21986 nand P2_U3953 P2_R1146_U78 ; P2_R1146_U292
g21987 nand P2_R1146_U292 P2_R1146_U160 ; P2_R1146_U293
g21988 nand P2_U3067 P2_R1146_U77 ; P2_R1146_U294
g21989 not P2_R1146_U159 ; P2_R1146_U295
g21990 nand P2_U3952 P2_R1146_U80 ; P2_R1146_U296
g21991 nand P2_R1146_U296 P2_R1146_U159 ; P2_R1146_U297
g21992 nand P2_U3060 P2_R1146_U79 ; P2_R1146_U298
g21993 not P2_R1146_U88 ; P2_R1146_U299
g21994 nand P2_U3950 P2_R1146_U84 ; P2_R1146_U300
g21995 nand P2_R1146_U88 P2_R1146_U183 P2_R1146_U300 ; P2_R1146_U301
g21996 nand P2_R1146_U84 P2_R1146_U83 ; P2_R1146_U302
g21997 nand P2_R1146_U302 P2_R1146_U81 ; P2_R1146_U303
g21998 nand P2_U3055 P2_R1146_U177 ; P2_R1146_U304
g21999 not P2_R1146_U87 ; P2_R1146_U305
g22000 nand P2_U3056 P2_R1146_U85 ; P2_R1146_U306
g22001 nand P2_R1146_U305 P2_R1146_U306 ; P2_R1146_U307
g22002 nand P2_U3949 P2_R1146_U86 ; P2_R1146_U308
g22003 nand P2_U3949 P2_R1146_U86 ; P2_R1146_U309
g22004 nand P2_R1146_U309 P2_R1146_U87 ; P2_R1146_U310
g22005 nand P2_U3056 P2_R1146_U85 ; P2_R1146_U311
g22006 nand P2_R1146_U129 P2_R1146_U310 ; P2_R1146_U312
g22007 nand P2_R1146_U299 P2_R1146_U83 ; P2_R1146_U313
g22008 nand P2_R1146_U133 P2_R1146_U313 ; P2_R1146_U314
g22009 nand P2_R1146_U88 P2_R1146_U183 ; P2_R1146_U315
g22010 nand P2_R1146_U132 P2_R1146_U315 ; P2_R1146_U316
g22011 nand P2_R1146_U83 P2_R1146_U183 ; P2_R1146_U317
g22012 nand P2_R1146_U287 P2_R1146_U163 ; P2_R1146_U318
g22013 not P2_R1146_U89 ; P2_R1146_U319
g22014 nand P2_U3063 P2_R1146_U71 ; P2_R1146_U320
g22015 nand P2_R1146_U319 P2_R1146_U320 ; P2_R1146_U321
g22016 nand P2_R1146_U137 P2_R1146_U321 ; P2_R1146_U322
g22017 nand P2_R1146_U89 P2_R1146_U182 ; P2_R1146_U323
g22018 nand P2_U3954 P2_R1146_U73 ; P2_R1146_U324
g22019 nand P2_R1146_U136 P2_R1146_U323 ; P2_R1146_U325
g22020 nand P2_U3063 P2_R1146_U71 ; P2_R1146_U326
g22021 nand P2_R1146_U182 P2_R1146_U326 ; P2_R1146_U327
g22022 nand P2_R1146_U287 P2_R1146_U76 ; P2_R1146_U328
g22023 nand P2_R1146_U261 P2_R1146_U172 ; P2_R1146_U329
g22024 not P2_R1146_U90 ; P2_R1146_U330
g22025 nand P2_U3076 P2_R1146_U56 ; P2_R1146_U331
g22026 nand P2_R1146_U330 P2_R1146_U331 ; P2_R1146_U332
g22027 nand P2_R1146_U144 P2_R1146_U332 ; P2_R1146_U333
g22028 nand P2_R1146_U90 P2_R1146_U181 ; P2_R1146_U334
g22029 nand P2_U3477 P2_R1146_U58 ; P2_R1146_U335
g22030 nand P2_R1146_U143 P2_R1146_U334 ; P2_R1146_U336
g22031 nand P2_U3076 P2_R1146_U56 ; P2_R1146_U337
g22032 nand P2_R1146_U181 P2_R1146_U337 ; P2_R1146_U338
g22033 nand P2_R1146_U261 P2_R1146_U61 ; P2_R1146_U339
g22034 nand P2_R1146_U216 P2_R1146_U150 ; P2_R1146_U340
g22035 not P2_R1146_U91 ; P2_R1146_U341
g22036 nand P2_U3064 P2_R1146_U46 ; P2_R1146_U342
g22037 nand P2_R1146_U341 P2_R1146_U342 ; P2_R1146_U343
g22038 nand P2_R1146_U148 P2_R1146_U343 ; P2_R1146_U344
g22039 nand P2_R1146_U91 P2_R1146_U180 ; P2_R1146_U345
g22040 nand P2_U3462 P2_R1146_U48 ; P2_R1146_U346
g22041 nand P2_R1146_U147 P2_R1146_U345 ; P2_R1146_U347
g22042 nand P2_U3064 P2_R1146_U46 ; P2_R1146_U348
g22043 nand P2_R1146_U180 P2_R1146_U348 ; P2_R1146_U349
g22044 nand P2_U3079 P2_R1146_U24 ; P2_R1146_U350
g22045 nand P2_U3080 P2_R1146_U165 ; P2_R1146_U351
g22046 nand P2_R1146_U130 P2_R1146_U307 ; P2_R1146_U352
g22047 nand P2_U3456 P2_R1146_U41 ; P2_R1146_U353
g22048 nand P2_U3085 P2_R1146_U40 ; P2_R1146_U354
g22049 nand P2_R1146_U217 P2_R1146_U150 ; P2_R1146_U355
g22050 nand P2_R1146_U215 P2_R1146_U149 ; P2_R1146_U356
g22051 nand P2_U3453 P2_R1146_U39 ; P2_R1146_U357
g22052 nand P2_U3086 P2_R1146_U36 ; P2_R1146_U358
g22053 nand P2_U3453 P2_R1146_U39 ; P2_R1146_U359
g22054 nand P2_U3086 P2_R1146_U36 ; P2_R1146_U360
g22055 nand P2_R1146_U360 P2_R1146_U359 ; P2_R1146_U361
g22056 nand P2_U3450 P2_R1146_U37 ; P2_R1146_U362
g22057 nand P2_U3072 P2_R1146_U21 ; P2_R1146_U363
g22058 nand P2_R1146_U222 P2_R1146_U42 ; P2_R1146_U364
g22059 nand P2_R1146_U151 P2_R1146_U209 ; P2_R1146_U365
g22060 nand P2_U3447 P2_R1146_U32 ; P2_R1146_U366
g22061 nand P2_U3073 P2_R1146_U30 ; P2_R1146_U367
g22062 nand P2_R1146_U367 P2_R1146_U366 ; P2_R1146_U368
g22063 nand P2_U3444 P2_R1146_U33 ; P2_R1146_U369
g22064 nand P2_U3069 P2_R1146_U22 ; P2_R1146_U370
g22065 nand P2_R1146_U232 P2_R1146_U43 ; P2_R1146_U371
g22066 nand P2_R1146_U152 P2_R1146_U224 ; P2_R1146_U372
g22067 nand P2_U3441 P2_R1146_U34 ; P2_R1146_U373
g22068 nand P2_U3062 P2_R1146_U31 ; P2_R1146_U374
g22069 nand P2_R1146_U233 P2_R1146_U154 ; P2_R1146_U375
g22070 nand P2_R1146_U199 P2_R1146_U153 ; P2_R1146_U376
g22071 nand P2_U3438 P2_R1146_U29 ; P2_R1146_U377
g22072 nand P2_U3066 P2_R1146_U26 ; P2_R1146_U378
g22073 nand P2_U3438 P2_R1146_U29 ; P2_R1146_U379
g22074 nand P2_U3066 P2_R1146_U26 ; P2_R1146_U380
g22075 nand P2_R1146_U380 P2_R1146_U379 ; P2_R1146_U381
g22076 nand P2_U3435 P2_R1146_U27 ; P2_R1146_U382
g22077 nand P2_U3070 P2_R1146_U23 ; P2_R1146_U383
g22078 nand P2_R1146_U238 P2_R1146_U44 ; P2_R1146_U384
g22079 nand P2_R1146_U155 P2_R1146_U193 ; P2_R1146_U385
g22080 nand P2_U3960 P2_R1146_U157 ; P2_R1146_U386
g22081 nand P2_U3057 P2_R1146_U156 ; P2_R1146_U387
g22082 nand P2_U3960 P2_R1146_U157 ; P2_R1146_U388
g22083 nand P2_U3057 P2_R1146_U156 ; P2_R1146_U389
g22084 nand P2_R1146_U389 P2_R1146_U388 ; P2_R1146_U390
g22085 nand P2_U3949 P2_R1146_U86 ; P2_R1146_U391
g22086 nand P2_U3056 P2_R1146_U85 ; P2_R1146_U392
g22087 not P2_R1146_U131 ; P2_R1146_U393
g22088 nand P2_R1146_U393 P2_R1146_U305 ; P2_R1146_U394
g22089 nand P2_R1146_U131 P2_R1146_U87 ; P2_R1146_U395
g22090 nand P2_U3950 P2_R1146_U84 ; P2_R1146_U396
g22091 nand P2_U3055 P2_R1146_U81 ; P2_R1146_U397
g22092 nand P2_U3950 P2_R1146_U84 ; P2_R1146_U398
g22093 nand P2_U3055 P2_R1146_U81 ; P2_R1146_U399
g22094 nand P2_R1146_U399 P2_R1146_U398 ; P2_R1146_U400
g22095 nand P2_U3951 P2_R1146_U82 ; P2_R1146_U401
g22096 nand P2_U3059 P2_R1146_U45 ; P2_R1146_U402
g22097 nand P2_R1146_U317 P2_R1146_U88 ; P2_R1146_U403
g22098 nand P2_R1146_U158 P2_R1146_U299 ; P2_R1146_U404
g22099 nand P2_U3952 P2_R1146_U80 ; P2_R1146_U405
g22100 nand P2_U3060 P2_R1146_U79 ; P2_R1146_U406
g22101 not P2_R1146_U134 ; P2_R1146_U407
g22102 nand P2_R1146_U295 P2_R1146_U407 ; P2_R1146_U408
g22103 nand P2_R1146_U134 P2_R1146_U159 ; P2_R1146_U409
g22104 nand P2_U3953 P2_R1146_U78 ; P2_R1146_U410
g22105 nand P2_U3067 P2_R1146_U77 ; P2_R1146_U411
g22106 not P2_R1146_U135 ; P2_R1146_U412
g22107 nand P2_R1146_U291 P2_R1146_U412 ; P2_R1146_U413
g22108 nand P2_R1146_U135 P2_R1146_U160 ; P2_R1146_U414
g22109 nand P2_U3954 P2_R1146_U73 ; P2_R1146_U415
g22110 nand P2_U3068 P2_R1146_U70 ; P2_R1146_U416
g22111 nand P2_R1146_U416 P2_R1146_U415 ; P2_R1146_U417
g22112 nand P2_U3955 P2_R1146_U74 ; P2_R1146_U418
g22113 nand P2_U3063 P2_R1146_U71 ; P2_R1146_U419
g22114 nand P2_R1146_U327 P2_R1146_U89 ; P2_R1146_U420
g22115 nand P2_R1146_U161 P2_R1146_U319 ; P2_R1146_U421
g22116 nand P2_U3956 P2_R1146_U75 ; P2_R1146_U422
g22117 nand P2_U3077 P2_R1146_U72 ; P2_R1146_U423
g22118 nand P2_R1146_U328 P2_R1146_U163 ; P2_R1146_U424
g22119 nand P2_R1146_U281 P2_R1146_U162 ; P2_R1146_U425
g22120 nand P2_U3957 P2_R1146_U69 ; P2_R1146_U426
g22121 nand P2_U3078 P2_R1146_U68 ; P2_R1146_U427
g22122 not P2_R1146_U138 ; P2_R1146_U428
g22123 nand P2_R1146_U277 P2_R1146_U428 ; P2_R1146_U429
g22124 nand P2_R1146_U138 P2_R1146_U164 ; P2_R1146_U430
g22125 nand P2_U3432 P2_R1146_U25 ; P2_R1146_U431
g22126 nand P2_U3080 P2_R1146_U165 ; P2_R1146_U432
g22127 not P2_R1146_U139 ; P2_R1146_U433
g22128 nand P2_R1146_U191 P2_R1146_U433 ; P2_R1146_U434
g22129 nand P2_R1146_U139 P2_R1146_U166 ; P2_R1146_U435
g22130 nand P2_U3485 P2_R1146_U67 ; P2_R1146_U436
g22131 nand P2_U3083 P2_R1146_U66 ; P2_R1146_U437
g22132 not P2_R1146_U140 ; P2_R1146_U438
g22133 nand P2_R1146_U273 P2_R1146_U438 ; P2_R1146_U439
g22134 nand P2_R1146_U140 P2_R1146_U167 ; P2_R1146_U440
g22135 nand P2_U3483 P2_R1146_U65 ; P2_R1146_U441
g22136 nand P2_U3084 P2_R1146_U168 ; P2_R1146_U442
g22137 not P2_R1146_U141 ; P2_R1146_U443
g22138 nand P2_R1146_U443 P2_R1146_U269 ; P2_R1146_U444
g22139 nand P2_R1146_U141 P2_R1146_U64 ; P2_R1146_U445
g22140 nand P2_U3480 P2_R1146_U63 ; P2_R1146_U446
g22141 nand P2_U3071 P2_R1146_U62 ; P2_R1146_U447
g22142 not P2_R1146_U142 ; P2_R1146_U448
g22143 nand P2_R1146_U265 P2_R1146_U448 ; P2_R1146_U449
g22144 nand P2_R1146_U142 P2_R1146_U169 ; P2_R1146_U450
g22145 nand P2_U3477 P2_R1146_U58 ; P2_R1146_U451
g22146 nand P2_U3075 P2_R1146_U55 ; P2_R1146_U452
g22147 nand P2_R1146_U452 P2_R1146_U451 ; P2_R1146_U453
g22148 nand P2_U3474 P2_R1146_U59 ; P2_R1146_U454
g22149 nand P2_U3076 P2_R1146_U56 ; P2_R1146_U455
g22150 nand P2_R1146_U338 P2_R1146_U90 ; P2_R1146_U456
g22151 nand P2_R1146_U170 P2_R1146_U330 ; P2_R1146_U457
g22152 nand P2_U3471 P2_R1146_U60 ; P2_R1146_U458
g22153 nand P2_U3081 P2_R1146_U57 ; P2_R1146_U459
g22154 nand P2_R1146_U339 P2_R1146_U172 ; P2_R1146_U460
g22155 nand P2_R1146_U255 P2_R1146_U171 ; P2_R1146_U461
g22156 nand P2_U3468 P2_R1146_U54 ; P2_R1146_U462
g22157 nand P2_U3082 P2_R1146_U53 ; P2_R1146_U463
g22158 not P2_R1146_U145 ; P2_R1146_U464
g22159 nand P2_R1146_U251 P2_R1146_U464 ; P2_R1146_U465
g22160 nand P2_R1146_U145 P2_R1146_U173 ; P2_R1146_U466
g22161 nand P2_U3465 P2_R1146_U52 ; P2_R1146_U467
g22162 nand P2_U3074 P2_R1146_U51 ; P2_R1146_U468
g22163 not P2_R1146_U146 ; P2_R1146_U469
g22164 nand P2_R1146_U247 P2_R1146_U469 ; P2_R1146_U470
g22165 nand P2_R1146_U146 P2_R1146_U174 ; P2_R1146_U471
g22166 nand P2_U3462 P2_R1146_U48 ; P2_R1146_U472
g22167 nand P2_U3065 P2_R1146_U47 ; P2_R1146_U473
g22168 nand P2_R1146_U473 P2_R1146_U472 ; P2_R1146_U474
g22169 nand P2_U3459 P2_R1146_U49 ; P2_R1146_U475
g22170 nand P2_U3064 P2_R1146_U46 ; P2_R1146_U476
g22171 nand P2_R1146_U349 P2_R1146_U91 ; P2_R1146_U477
g22172 nand P2_R1146_U175 P2_R1146_U341 ; P2_R1146_U478
g22173 and P2_R1203_U202 P2_R1203_U201 ; P2_R1203_U6
g22174 and P2_R1203_U241 P2_R1203_U240 ; P2_R1203_U7
g22175 and P2_R1203_U181 P2_R1203_U256 ; P2_R1203_U8
g22176 and P2_R1203_U258 P2_R1203_U257 ; P2_R1203_U9
g22177 and P2_R1203_U182 P2_R1203_U282 ; P2_R1203_U10
g22178 and P2_R1203_U284 P2_R1203_U283 ; P2_R1203_U11
g22179 nand P2_R1203_U344 P2_R1203_U347 ; P2_R1203_U12
g22180 nand P2_R1203_U333 P2_R1203_U336 ; P2_R1203_U13
g22181 nand P2_R1203_U322 P2_R1203_U325 ; P2_R1203_U14
g22182 nand P2_R1203_U314 P2_R1203_U316 ; P2_R1203_U15
g22183 nand P2_R1203_U352 P2_R1203_U312 ; P2_R1203_U16
g22184 nand P2_R1203_U235 P2_R1203_U237 ; P2_R1203_U17
g22185 nand P2_R1203_U227 P2_R1203_U230 ; P2_R1203_U18
g22186 nand P2_R1203_U219 P2_R1203_U221 ; P2_R1203_U19
g22187 nand P2_R1203_U166 P2_R1203_U350 ; P2_R1203_U20
g22188 not P2_U3450 ; P2_R1203_U21
g22189 not P2_U3444 ; P2_R1203_U22
g22190 not P2_U3435 ; P2_R1203_U23
g22191 not P2_U3427 ; P2_R1203_U24
g22192 not P2_U3080 ; P2_R1203_U25
g22193 not P2_U3438 ; P2_R1203_U26
g22194 not P2_U3070 ; P2_R1203_U27
g22195 nand P2_U3070 P2_R1203_U23 ; P2_R1203_U28
g22196 not P2_U3066 ; P2_R1203_U29
g22197 not P2_U3447 ; P2_R1203_U30
g22198 not P2_U3441 ; P2_R1203_U31
g22199 not P2_U3073 ; P2_R1203_U32
g22200 not P2_U3069 ; P2_R1203_U33
g22201 not P2_U3062 ; P2_R1203_U34
g22202 nand P2_U3062 P2_R1203_U31 ; P2_R1203_U35
g22203 not P2_U3453 ; P2_R1203_U36
g22204 not P2_U3072 ; P2_R1203_U37
g22205 nand P2_U3072 P2_R1203_U21 ; P2_R1203_U38
g22206 not P2_U3086 ; P2_R1203_U39
g22207 not P2_U3456 ; P2_R1203_U40
g22208 not P2_U3085 ; P2_R1203_U41
g22209 nand P2_R1203_U208 P2_R1203_U207 ; P2_R1203_U42
g22210 nand P2_R1203_U35 P2_R1203_U223 ; P2_R1203_U43
g22211 nand P2_R1203_U192 P2_R1203_U176 P2_R1203_U351 ; P2_R1203_U44
g22212 not P2_U3951 ; P2_R1203_U45
g22213 not P2_U3459 ; P2_R1203_U46
g22214 not P2_U3462 ; P2_R1203_U47
g22215 not P2_U3065 ; P2_R1203_U48
g22216 not P2_U3064 ; P2_R1203_U49
g22217 nand P2_U3085 P2_R1203_U40 ; P2_R1203_U50
g22218 not P2_U3465 ; P2_R1203_U51
g22219 not P2_U3074 ; P2_R1203_U52
g22220 not P2_U3468 ; P2_R1203_U53
g22221 not P2_U3082 ; P2_R1203_U54
g22222 not P2_U3477 ; P2_R1203_U55
g22223 not P2_U3474 ; P2_R1203_U56
g22224 not P2_U3471 ; P2_R1203_U57
g22225 not P2_U3075 ; P2_R1203_U58
g22226 not P2_U3076 ; P2_R1203_U59
g22227 not P2_U3081 ; P2_R1203_U60
g22228 nand P2_U3081 P2_R1203_U57 ; P2_R1203_U61
g22229 not P2_U3480 ; P2_R1203_U62
g22230 not P2_U3071 ; P2_R1203_U63
g22231 nand P2_R1203_U268 P2_R1203_U267 ; P2_R1203_U64
g22232 not P2_U3084 ; P2_R1203_U65
g22233 not P2_U3485 ; P2_R1203_U66
g22234 not P2_U3083 ; P2_R1203_U67
g22235 not P2_U3957 ; P2_R1203_U68
g22236 not P2_U3078 ; P2_R1203_U69
g22237 not P2_U3954 ; P2_R1203_U70
g22238 not P2_U3955 ; P2_R1203_U71
g22239 not P2_U3956 ; P2_R1203_U72
g22240 not P2_U3068 ; P2_R1203_U73
g22241 not P2_U3063 ; P2_R1203_U74
g22242 not P2_U3077 ; P2_R1203_U75
g22243 nand P2_U3077 P2_R1203_U72 ; P2_R1203_U76
g22244 not P2_U3953 ; P2_R1203_U77
g22245 not P2_U3067 ; P2_R1203_U78
g22246 not P2_U3952 ; P2_R1203_U79
g22247 not P2_U3060 ; P2_R1203_U80
g22248 not P2_U3950 ; P2_R1203_U81
g22249 not P2_U3059 ; P2_R1203_U82
g22250 nand P2_U3059 P2_R1203_U45 ; P2_R1203_U83
g22251 not P2_U3055 ; P2_R1203_U84
g22252 not P2_U3949 ; P2_R1203_U85
g22253 not P2_U3056 ; P2_R1203_U86
g22254 nand P2_R1203_U128 P2_R1203_U301 ; P2_R1203_U87
g22255 nand P2_R1203_U298 P2_R1203_U297 ; P2_R1203_U88
g22256 nand P2_R1203_U76 P2_R1203_U318 ; P2_R1203_U89
g22257 nand P2_R1203_U61 P2_R1203_U329 ; P2_R1203_U90
g22258 nand P2_R1203_U50 P2_R1203_U340 ; P2_R1203_U91
g22259 not P2_U3079 ; P2_R1203_U92
g22260 nand P2_R1203_U395 P2_R1203_U394 ; P2_R1203_U93
g22261 nand P2_R1203_U409 P2_R1203_U408 ; P2_R1203_U94
g22262 nand P2_R1203_U414 P2_R1203_U413 ; P2_R1203_U95
g22263 nand P2_R1203_U430 P2_R1203_U429 ; P2_R1203_U96
g22264 nand P2_R1203_U435 P2_R1203_U434 ; P2_R1203_U97
g22265 nand P2_R1203_U440 P2_R1203_U439 ; P2_R1203_U98
g22266 nand P2_R1203_U445 P2_R1203_U444 ; P2_R1203_U99
g22267 nand P2_R1203_U450 P2_R1203_U449 ; P2_R1203_U100
g22268 nand P2_R1203_U466 P2_R1203_U465 ; P2_R1203_U101
g22269 nand P2_R1203_U471 P2_R1203_U470 ; P2_R1203_U102
g22270 nand P2_R1203_U356 P2_R1203_U355 ; P2_R1203_U103
g22271 nand P2_R1203_U365 P2_R1203_U364 ; P2_R1203_U104
g22272 nand P2_R1203_U372 P2_R1203_U371 ; P2_R1203_U105
g22273 nand P2_R1203_U376 P2_R1203_U375 ; P2_R1203_U106
g22274 nand P2_R1203_U385 P2_R1203_U384 ; P2_R1203_U107
g22275 nand P2_R1203_U404 P2_R1203_U403 ; P2_R1203_U108
g22276 nand P2_R1203_U421 P2_R1203_U420 ; P2_R1203_U109
g22277 nand P2_R1203_U425 P2_R1203_U424 ; P2_R1203_U110
g22278 nand P2_R1203_U457 P2_R1203_U456 ; P2_R1203_U111
g22279 nand P2_R1203_U461 P2_R1203_U460 ; P2_R1203_U112
g22280 nand P2_R1203_U478 P2_R1203_U477 ; P2_R1203_U113
g22281 and P2_R1203_U194 P2_R1203_U184 ; P2_R1203_U114
g22282 and P2_R1203_U197 P2_R1203_U198 ; P2_R1203_U115
g22283 and P2_R1203_U205 P2_R1203_U200 P2_R1203_U185 ; P2_R1203_U116
g22284 and P2_R1203_U210 P2_R1203_U186 ; P2_R1203_U117
g22285 and P2_R1203_U213 P2_R1203_U214 ; P2_R1203_U118
g22286 and P2_R1203_U358 P2_R1203_U357 P2_R1203_U38 ; P2_R1203_U119
g22287 and P2_R1203_U361 P2_R1203_U186 ; P2_R1203_U120
g22288 and P2_R1203_U229 P2_R1203_U6 ; P2_R1203_U121
g22289 and P2_R1203_U368 P2_R1203_U185 ; P2_R1203_U122
g22290 and P2_R1203_U378 P2_R1203_U377 P2_R1203_U28 ; P2_R1203_U123
g22291 and P2_R1203_U381 P2_R1203_U184 ; P2_R1203_U124
g22292 and P2_R1203_U239 P2_R1203_U216 P2_R1203_U180 ; P2_R1203_U125
g22293 and P2_R1203_U261 P2_R1203_U8 ; P2_R1203_U126
g22294 and P2_R1203_U287 P2_R1203_U10 ; P2_R1203_U127
g22295 and P2_R1203_U303 P2_R1203_U304 ; P2_R1203_U128
g22296 and P2_R1203_U387 P2_R1203_U386 P2_R1203_U311 ; P2_R1203_U129
g22297 and P2_R1203_U308 P2_R1203_U390 ; P2_R1203_U130
g22298 nand P2_R1203_U392 P2_R1203_U391 ; P2_R1203_U131
g22299 and P2_R1203_U397 P2_R1203_U396 P2_R1203_U83 ; P2_R1203_U132
g22300 and P2_R1203_U400 P2_R1203_U183 ; P2_R1203_U133
g22301 nand P2_R1203_U406 P2_R1203_U405 ; P2_R1203_U134
g22302 nand P2_R1203_U411 P2_R1203_U410 ; P2_R1203_U135
g22303 and P2_R1203_U324 P2_R1203_U11 ; P2_R1203_U136
g22304 and P2_R1203_U417 P2_R1203_U182 ; P2_R1203_U137
g22305 nand P2_R1203_U427 P2_R1203_U426 ; P2_R1203_U138
g22306 nand P2_R1203_U432 P2_R1203_U431 ; P2_R1203_U139
g22307 nand P2_R1203_U437 P2_R1203_U436 ; P2_R1203_U140
g22308 nand P2_R1203_U442 P2_R1203_U441 ; P2_R1203_U141
g22309 nand P2_R1203_U447 P2_R1203_U446 ; P2_R1203_U142
g22310 and P2_R1203_U335 P2_R1203_U9 ; P2_R1203_U143
g22311 and P2_R1203_U453 P2_R1203_U181 ; P2_R1203_U144
g22312 nand P2_R1203_U463 P2_R1203_U462 ; P2_R1203_U145
g22313 nand P2_R1203_U468 P2_R1203_U467 ; P2_R1203_U146
g22314 and P2_R1203_U346 P2_R1203_U7 ; P2_R1203_U147
g22315 and P2_R1203_U474 P2_R1203_U180 ; P2_R1203_U148
g22316 and P2_R1203_U354 P2_R1203_U353 ; P2_R1203_U149
g22317 nand P2_R1203_U118 P2_R1203_U211 ; P2_R1203_U150
g22318 and P2_R1203_U363 P2_R1203_U362 ; P2_R1203_U151
g22319 and P2_R1203_U370 P2_R1203_U369 ; P2_R1203_U152
g22320 and P2_R1203_U374 P2_R1203_U373 ; P2_R1203_U153
g22321 nand P2_R1203_U115 P2_R1203_U195 ; P2_R1203_U154
g22322 and P2_R1203_U383 P2_R1203_U382 ; P2_R1203_U155
g22323 not P2_U3960 ; P2_R1203_U156
g22324 not P2_U3057 ; P2_R1203_U157
g22325 and P2_R1203_U402 P2_R1203_U401 ; P2_R1203_U158
g22326 nand P2_R1203_U294 P2_R1203_U293 ; P2_R1203_U159
g22327 nand P2_R1203_U290 P2_R1203_U289 ; P2_R1203_U160
g22328 and P2_R1203_U419 P2_R1203_U418 ; P2_R1203_U161
g22329 and P2_R1203_U423 P2_R1203_U422 ; P2_R1203_U162
g22330 nand P2_R1203_U280 P2_R1203_U279 ; P2_R1203_U163
g22331 nand P2_R1203_U276 P2_R1203_U275 ; P2_R1203_U164
g22332 not P2_U3432 ; P2_R1203_U165
g22333 nand P2_U3427 P2_R1203_U92 ; P2_R1203_U166
g22334 nand P2_R1203_U272 P2_R1203_U271 ; P2_R1203_U167
g22335 not P2_U3483 ; P2_R1203_U168
g22336 nand P2_R1203_U264 P2_R1203_U263 ; P2_R1203_U169
g22337 and P2_R1203_U455 P2_R1203_U454 ; P2_R1203_U170
g22338 and P2_R1203_U459 P2_R1203_U458 ; P2_R1203_U171
g22339 nand P2_R1203_U254 P2_R1203_U253 ; P2_R1203_U172
g22340 nand P2_R1203_U250 P2_R1203_U249 ; P2_R1203_U173
g22341 nand P2_R1203_U246 P2_R1203_U245 ; P2_R1203_U174
g22342 and P2_R1203_U476 P2_R1203_U475 ; P2_R1203_U175
g22343 nand P2_R1203_U166 P2_R1203_U165 ; P2_R1203_U176
g22344 not P2_R1203_U83 ; P2_R1203_U177
g22345 not P2_R1203_U28 ; P2_R1203_U178
g22346 not P2_R1203_U38 ; P2_R1203_U179
g22347 nand P2_U3459 P2_R1203_U49 ; P2_R1203_U180
g22348 nand P2_U3474 P2_R1203_U59 ; P2_R1203_U181
g22349 nand P2_U3955 P2_R1203_U74 ; P2_R1203_U182
g22350 nand P2_U3951 P2_R1203_U82 ; P2_R1203_U183
g22351 nand P2_U3435 P2_R1203_U27 ; P2_R1203_U184
g22352 nand P2_U3444 P2_R1203_U33 ; P2_R1203_U185
g22353 nand P2_U3450 P2_R1203_U37 ; P2_R1203_U186
g22354 not P2_R1203_U61 ; P2_R1203_U187
g22355 not P2_R1203_U76 ; P2_R1203_U188
g22356 not P2_R1203_U35 ; P2_R1203_U189
g22357 not P2_R1203_U50 ; P2_R1203_U190
g22358 not P2_R1203_U166 ; P2_R1203_U191
g22359 nand P2_U3080 P2_R1203_U166 ; P2_R1203_U192
g22360 not P2_R1203_U44 ; P2_R1203_U193
g22361 nand P2_U3438 P2_R1203_U29 ; P2_R1203_U194
g22362 nand P2_R1203_U114 P2_R1203_U44 ; P2_R1203_U195
g22363 nand P2_R1203_U29 P2_R1203_U28 ; P2_R1203_U196
g22364 nand P2_R1203_U196 P2_R1203_U26 ; P2_R1203_U197
g22365 nand P2_U3066 P2_R1203_U178 ; P2_R1203_U198
g22366 not P2_R1203_U154 ; P2_R1203_U199
g22367 nand P2_U3447 P2_R1203_U32 ; P2_R1203_U200
g22368 nand P2_U3073 P2_R1203_U30 ; P2_R1203_U201
g22369 nand P2_U3069 P2_R1203_U22 ; P2_R1203_U202
g22370 nand P2_R1203_U189 P2_R1203_U185 ; P2_R1203_U203
g22371 nand P2_R1203_U6 P2_R1203_U203 ; P2_R1203_U204
g22372 nand P2_U3441 P2_R1203_U34 ; P2_R1203_U205
g22373 nand P2_U3447 P2_R1203_U32 ; P2_R1203_U206
g22374 nand P2_R1203_U154 P2_R1203_U116 ; P2_R1203_U207
g22375 nand P2_R1203_U206 P2_R1203_U204 ; P2_R1203_U208
g22376 not P2_R1203_U42 ; P2_R1203_U209
g22377 nand P2_U3453 P2_R1203_U39 ; P2_R1203_U210
g22378 nand P2_R1203_U117 P2_R1203_U42 ; P2_R1203_U211
g22379 nand P2_R1203_U39 P2_R1203_U38 ; P2_R1203_U212
g22380 nand P2_R1203_U212 P2_R1203_U36 ; P2_R1203_U213
g22381 nand P2_U3086 P2_R1203_U179 ; P2_R1203_U214
g22382 not P2_R1203_U150 ; P2_R1203_U215
g22383 nand P2_U3456 P2_R1203_U41 ; P2_R1203_U216
g22384 nand P2_R1203_U216 P2_R1203_U50 ; P2_R1203_U217
g22385 nand P2_R1203_U209 P2_R1203_U38 ; P2_R1203_U218
g22386 nand P2_R1203_U120 P2_R1203_U218 ; P2_R1203_U219
g22387 nand P2_R1203_U42 P2_R1203_U186 ; P2_R1203_U220
g22388 nand P2_R1203_U119 P2_R1203_U220 ; P2_R1203_U221
g22389 nand P2_R1203_U38 P2_R1203_U186 ; P2_R1203_U222
g22390 nand P2_R1203_U205 P2_R1203_U154 ; P2_R1203_U223
g22391 not P2_R1203_U43 ; P2_R1203_U224
g22392 nand P2_U3069 P2_R1203_U22 ; P2_R1203_U225
g22393 nand P2_R1203_U224 P2_R1203_U225 ; P2_R1203_U226
g22394 nand P2_R1203_U122 P2_R1203_U226 ; P2_R1203_U227
g22395 nand P2_R1203_U43 P2_R1203_U185 ; P2_R1203_U228
g22396 nand P2_U3447 P2_R1203_U32 ; P2_R1203_U229
g22397 nand P2_R1203_U121 P2_R1203_U228 ; P2_R1203_U230
g22398 nand P2_U3069 P2_R1203_U22 ; P2_R1203_U231
g22399 nand P2_R1203_U185 P2_R1203_U231 ; P2_R1203_U232
g22400 nand P2_R1203_U205 P2_R1203_U35 ; P2_R1203_U233
g22401 nand P2_R1203_U193 P2_R1203_U28 ; P2_R1203_U234
g22402 nand P2_R1203_U124 P2_R1203_U234 ; P2_R1203_U235
g22403 nand P2_R1203_U44 P2_R1203_U184 ; P2_R1203_U236
g22404 nand P2_R1203_U123 P2_R1203_U236 ; P2_R1203_U237
g22405 nand P2_R1203_U28 P2_R1203_U184 ; P2_R1203_U238
g22406 nand P2_U3462 P2_R1203_U48 ; P2_R1203_U239
g22407 nand P2_U3065 P2_R1203_U47 ; P2_R1203_U240
g22408 nand P2_U3064 P2_R1203_U46 ; P2_R1203_U241
g22409 nand P2_R1203_U190 P2_R1203_U180 ; P2_R1203_U242
g22410 nand P2_R1203_U7 P2_R1203_U242 ; P2_R1203_U243
g22411 nand P2_U3462 P2_R1203_U48 ; P2_R1203_U244
g22412 nand P2_R1203_U150 P2_R1203_U125 ; P2_R1203_U245
g22413 nand P2_R1203_U244 P2_R1203_U243 ; P2_R1203_U246
g22414 not P2_R1203_U174 ; P2_R1203_U247
g22415 nand P2_U3465 P2_R1203_U52 ; P2_R1203_U248
g22416 nand P2_R1203_U248 P2_R1203_U174 ; P2_R1203_U249
g22417 nand P2_U3074 P2_R1203_U51 ; P2_R1203_U250
g22418 not P2_R1203_U173 ; P2_R1203_U251
g22419 nand P2_U3468 P2_R1203_U54 ; P2_R1203_U252
g22420 nand P2_R1203_U252 P2_R1203_U173 ; P2_R1203_U253
g22421 nand P2_U3082 P2_R1203_U53 ; P2_R1203_U254
g22422 not P2_R1203_U172 ; P2_R1203_U255
g22423 nand P2_U3477 P2_R1203_U58 ; P2_R1203_U256
g22424 nand P2_U3075 P2_R1203_U55 ; P2_R1203_U257
g22425 nand P2_U3076 P2_R1203_U56 ; P2_R1203_U258
g22426 nand P2_R1203_U187 P2_R1203_U8 ; P2_R1203_U259
g22427 nand P2_R1203_U9 P2_R1203_U259 ; P2_R1203_U260
g22428 nand P2_U3471 P2_R1203_U60 ; P2_R1203_U261
g22429 nand P2_U3477 P2_R1203_U58 ; P2_R1203_U262
g22430 nand P2_R1203_U126 P2_R1203_U172 ; P2_R1203_U263
g22431 nand P2_R1203_U262 P2_R1203_U260 ; P2_R1203_U264
g22432 not P2_R1203_U169 ; P2_R1203_U265
g22433 nand P2_U3480 P2_R1203_U63 ; P2_R1203_U266
g22434 nand P2_R1203_U266 P2_R1203_U169 ; P2_R1203_U267
g22435 nand P2_U3071 P2_R1203_U62 ; P2_R1203_U268
g22436 not P2_R1203_U64 ; P2_R1203_U269
g22437 nand P2_R1203_U269 P2_R1203_U65 ; P2_R1203_U270
g22438 nand P2_R1203_U270 P2_R1203_U168 ; P2_R1203_U271
g22439 nand P2_U3084 P2_R1203_U64 ; P2_R1203_U272
g22440 not P2_R1203_U167 ; P2_R1203_U273
g22441 nand P2_U3485 P2_R1203_U67 ; P2_R1203_U274
g22442 nand P2_R1203_U274 P2_R1203_U167 ; P2_R1203_U275
g22443 nand P2_U3083 P2_R1203_U66 ; P2_R1203_U276
g22444 not P2_R1203_U164 ; P2_R1203_U277
g22445 nand P2_U3957 P2_R1203_U69 ; P2_R1203_U278
g22446 nand P2_R1203_U278 P2_R1203_U164 ; P2_R1203_U279
g22447 nand P2_U3078 P2_R1203_U68 ; P2_R1203_U280
g22448 not P2_R1203_U163 ; P2_R1203_U281
g22449 nand P2_U3954 P2_R1203_U73 ; P2_R1203_U282
g22450 nand P2_U3068 P2_R1203_U70 ; P2_R1203_U283
g22451 nand P2_U3063 P2_R1203_U71 ; P2_R1203_U284
g22452 nand P2_R1203_U188 P2_R1203_U10 ; P2_R1203_U285
g22453 nand P2_R1203_U11 P2_R1203_U285 ; P2_R1203_U286
g22454 nand P2_U3956 P2_R1203_U75 ; P2_R1203_U287
g22455 nand P2_U3954 P2_R1203_U73 ; P2_R1203_U288
g22456 nand P2_R1203_U127 P2_R1203_U163 ; P2_R1203_U289
g22457 nand P2_R1203_U288 P2_R1203_U286 ; P2_R1203_U290
g22458 not P2_R1203_U160 ; P2_R1203_U291
g22459 nand P2_U3953 P2_R1203_U78 ; P2_R1203_U292
g22460 nand P2_R1203_U292 P2_R1203_U160 ; P2_R1203_U293
g22461 nand P2_U3067 P2_R1203_U77 ; P2_R1203_U294
g22462 not P2_R1203_U159 ; P2_R1203_U295
g22463 nand P2_U3952 P2_R1203_U80 ; P2_R1203_U296
g22464 nand P2_R1203_U296 P2_R1203_U159 ; P2_R1203_U297
g22465 nand P2_U3060 P2_R1203_U79 ; P2_R1203_U298
g22466 not P2_R1203_U88 ; P2_R1203_U299
g22467 nand P2_U3950 P2_R1203_U84 ; P2_R1203_U300
g22468 nand P2_R1203_U88 P2_R1203_U183 P2_R1203_U300 ; P2_R1203_U301
g22469 nand P2_R1203_U84 P2_R1203_U83 ; P2_R1203_U302
g22470 nand P2_R1203_U302 P2_R1203_U81 ; P2_R1203_U303
g22471 nand P2_U3055 P2_R1203_U177 ; P2_R1203_U304
g22472 not P2_R1203_U87 ; P2_R1203_U305
g22473 nand P2_U3056 P2_R1203_U85 ; P2_R1203_U306
g22474 nand P2_R1203_U305 P2_R1203_U306 ; P2_R1203_U307
g22475 nand P2_U3949 P2_R1203_U86 ; P2_R1203_U308
g22476 nand P2_U3949 P2_R1203_U86 ; P2_R1203_U309
g22477 nand P2_R1203_U309 P2_R1203_U87 ; P2_R1203_U310
g22478 nand P2_U3056 P2_R1203_U85 ; P2_R1203_U311
g22479 nand P2_R1203_U129 P2_R1203_U310 ; P2_R1203_U312
g22480 nand P2_R1203_U299 P2_R1203_U83 ; P2_R1203_U313
g22481 nand P2_R1203_U133 P2_R1203_U313 ; P2_R1203_U314
g22482 nand P2_R1203_U88 P2_R1203_U183 ; P2_R1203_U315
g22483 nand P2_R1203_U132 P2_R1203_U315 ; P2_R1203_U316
g22484 nand P2_R1203_U83 P2_R1203_U183 ; P2_R1203_U317
g22485 nand P2_R1203_U287 P2_R1203_U163 ; P2_R1203_U318
g22486 not P2_R1203_U89 ; P2_R1203_U319
g22487 nand P2_U3063 P2_R1203_U71 ; P2_R1203_U320
g22488 nand P2_R1203_U319 P2_R1203_U320 ; P2_R1203_U321
g22489 nand P2_R1203_U137 P2_R1203_U321 ; P2_R1203_U322
g22490 nand P2_R1203_U89 P2_R1203_U182 ; P2_R1203_U323
g22491 nand P2_U3954 P2_R1203_U73 ; P2_R1203_U324
g22492 nand P2_R1203_U136 P2_R1203_U323 ; P2_R1203_U325
g22493 nand P2_U3063 P2_R1203_U71 ; P2_R1203_U326
g22494 nand P2_R1203_U182 P2_R1203_U326 ; P2_R1203_U327
g22495 nand P2_R1203_U287 P2_R1203_U76 ; P2_R1203_U328
g22496 nand P2_R1203_U261 P2_R1203_U172 ; P2_R1203_U329
g22497 not P2_R1203_U90 ; P2_R1203_U330
g22498 nand P2_U3076 P2_R1203_U56 ; P2_R1203_U331
g22499 nand P2_R1203_U330 P2_R1203_U331 ; P2_R1203_U332
g22500 nand P2_R1203_U144 P2_R1203_U332 ; P2_R1203_U333
g22501 nand P2_R1203_U90 P2_R1203_U181 ; P2_R1203_U334
g22502 nand P2_U3477 P2_R1203_U58 ; P2_R1203_U335
g22503 nand P2_R1203_U143 P2_R1203_U334 ; P2_R1203_U336
g22504 nand P2_U3076 P2_R1203_U56 ; P2_R1203_U337
g22505 nand P2_R1203_U181 P2_R1203_U337 ; P2_R1203_U338
g22506 nand P2_R1203_U261 P2_R1203_U61 ; P2_R1203_U339
g22507 nand P2_R1203_U216 P2_R1203_U150 ; P2_R1203_U340
g22508 not P2_R1203_U91 ; P2_R1203_U341
g22509 nand P2_U3064 P2_R1203_U46 ; P2_R1203_U342
g22510 nand P2_R1203_U341 P2_R1203_U342 ; P2_R1203_U343
g22511 nand P2_R1203_U148 P2_R1203_U343 ; P2_R1203_U344
g22512 nand P2_R1203_U91 P2_R1203_U180 ; P2_R1203_U345
g22513 nand P2_U3462 P2_R1203_U48 ; P2_R1203_U346
g22514 nand P2_R1203_U147 P2_R1203_U345 ; P2_R1203_U347
g22515 nand P2_U3064 P2_R1203_U46 ; P2_R1203_U348
g22516 nand P2_R1203_U180 P2_R1203_U348 ; P2_R1203_U349
g22517 nand P2_U3079 P2_R1203_U24 ; P2_R1203_U350
g22518 nand P2_U3080 P2_R1203_U165 ; P2_R1203_U351
g22519 nand P2_R1203_U130 P2_R1203_U307 ; P2_R1203_U352
g22520 nand P2_U3456 P2_R1203_U41 ; P2_R1203_U353
g22521 nand P2_U3085 P2_R1203_U40 ; P2_R1203_U354
g22522 nand P2_R1203_U217 P2_R1203_U150 ; P2_R1203_U355
g22523 nand P2_R1203_U215 P2_R1203_U149 ; P2_R1203_U356
g22524 nand P2_U3453 P2_R1203_U39 ; P2_R1203_U357
g22525 nand P2_U3086 P2_R1203_U36 ; P2_R1203_U358
g22526 nand P2_U3453 P2_R1203_U39 ; P2_R1203_U359
g22527 nand P2_U3086 P2_R1203_U36 ; P2_R1203_U360
g22528 nand P2_R1203_U360 P2_R1203_U359 ; P2_R1203_U361
g22529 nand P2_U3450 P2_R1203_U37 ; P2_R1203_U362
g22530 nand P2_U3072 P2_R1203_U21 ; P2_R1203_U363
g22531 nand P2_R1203_U222 P2_R1203_U42 ; P2_R1203_U364
g22532 nand P2_R1203_U151 P2_R1203_U209 ; P2_R1203_U365
g22533 nand P2_U3447 P2_R1203_U32 ; P2_R1203_U366
g22534 nand P2_U3073 P2_R1203_U30 ; P2_R1203_U367
g22535 nand P2_R1203_U367 P2_R1203_U366 ; P2_R1203_U368
g22536 nand P2_U3444 P2_R1203_U33 ; P2_R1203_U369
g22537 nand P2_U3069 P2_R1203_U22 ; P2_R1203_U370
g22538 nand P2_R1203_U232 P2_R1203_U43 ; P2_R1203_U371
g22539 nand P2_R1203_U152 P2_R1203_U224 ; P2_R1203_U372
g22540 nand P2_U3441 P2_R1203_U34 ; P2_R1203_U373
g22541 nand P2_U3062 P2_R1203_U31 ; P2_R1203_U374
g22542 nand P2_R1203_U233 P2_R1203_U154 ; P2_R1203_U375
g22543 nand P2_R1203_U199 P2_R1203_U153 ; P2_R1203_U376
g22544 nand P2_U3438 P2_R1203_U29 ; P2_R1203_U377
g22545 nand P2_U3066 P2_R1203_U26 ; P2_R1203_U378
g22546 nand P2_U3438 P2_R1203_U29 ; P2_R1203_U379
g22547 nand P2_U3066 P2_R1203_U26 ; P2_R1203_U380
g22548 nand P2_R1203_U380 P2_R1203_U379 ; P2_R1203_U381
g22549 nand P2_U3435 P2_R1203_U27 ; P2_R1203_U382
g22550 nand P2_U3070 P2_R1203_U23 ; P2_R1203_U383
g22551 nand P2_R1203_U238 P2_R1203_U44 ; P2_R1203_U384
g22552 nand P2_R1203_U155 P2_R1203_U193 ; P2_R1203_U385
g22553 nand P2_U3960 P2_R1203_U157 ; P2_R1203_U386
g22554 nand P2_U3057 P2_R1203_U156 ; P2_R1203_U387
g22555 nand P2_U3960 P2_R1203_U157 ; P2_R1203_U388
g22556 nand P2_U3057 P2_R1203_U156 ; P2_R1203_U389
g22557 nand P2_R1203_U389 P2_R1203_U388 ; P2_R1203_U390
g22558 nand P2_U3949 P2_R1203_U86 ; P2_R1203_U391
g22559 nand P2_U3056 P2_R1203_U85 ; P2_R1203_U392
g22560 not P2_R1203_U131 ; P2_R1203_U393
g22561 nand P2_R1203_U393 P2_R1203_U305 ; P2_R1203_U394
g22562 nand P2_R1203_U131 P2_R1203_U87 ; P2_R1203_U395
g22563 nand P2_U3950 P2_R1203_U84 ; P2_R1203_U396
g22564 nand P2_U3055 P2_R1203_U81 ; P2_R1203_U397
g22565 nand P2_U3950 P2_R1203_U84 ; P2_R1203_U398
g22566 nand P2_U3055 P2_R1203_U81 ; P2_R1203_U399
g22567 nand P2_R1203_U399 P2_R1203_U398 ; P2_R1203_U400
g22568 nand P2_U3951 P2_R1203_U82 ; P2_R1203_U401
g22569 nand P2_U3059 P2_R1203_U45 ; P2_R1203_U402
g22570 nand P2_R1203_U317 P2_R1203_U88 ; P2_R1203_U403
g22571 nand P2_R1203_U158 P2_R1203_U299 ; P2_R1203_U404
g22572 nand P2_U3952 P2_R1203_U80 ; P2_R1203_U405
g22573 nand P2_U3060 P2_R1203_U79 ; P2_R1203_U406
g22574 not P2_R1203_U134 ; P2_R1203_U407
g22575 nand P2_R1203_U295 P2_R1203_U407 ; P2_R1203_U408
g22576 nand P2_R1203_U134 P2_R1203_U159 ; P2_R1203_U409
g22577 nand P2_U3953 P2_R1203_U78 ; P2_R1203_U410
g22578 nand P2_U3067 P2_R1203_U77 ; P2_R1203_U411
g22579 not P2_R1203_U135 ; P2_R1203_U412
g22580 nand P2_R1203_U291 P2_R1203_U412 ; P2_R1203_U413
g22581 nand P2_R1203_U135 P2_R1203_U160 ; P2_R1203_U414
g22582 nand P2_U3954 P2_R1203_U73 ; P2_R1203_U415
g22583 nand P2_U3068 P2_R1203_U70 ; P2_R1203_U416
g22584 nand P2_R1203_U416 P2_R1203_U415 ; P2_R1203_U417
g22585 nand P2_U3955 P2_R1203_U74 ; P2_R1203_U418
g22586 nand P2_U3063 P2_R1203_U71 ; P2_R1203_U419
g22587 nand P2_R1203_U327 P2_R1203_U89 ; P2_R1203_U420
g22588 nand P2_R1203_U161 P2_R1203_U319 ; P2_R1203_U421
g22589 nand P2_U3956 P2_R1203_U75 ; P2_R1203_U422
g22590 nand P2_U3077 P2_R1203_U72 ; P2_R1203_U423
g22591 nand P2_R1203_U328 P2_R1203_U163 ; P2_R1203_U424
g22592 nand P2_R1203_U281 P2_R1203_U162 ; P2_R1203_U425
g22593 nand P2_U3957 P2_R1203_U69 ; P2_R1203_U426
g22594 nand P2_U3078 P2_R1203_U68 ; P2_R1203_U427
g22595 not P2_R1203_U138 ; P2_R1203_U428
g22596 nand P2_R1203_U277 P2_R1203_U428 ; P2_R1203_U429
g22597 nand P2_R1203_U138 P2_R1203_U164 ; P2_R1203_U430
g22598 nand P2_U3432 P2_R1203_U25 ; P2_R1203_U431
g22599 nand P2_U3080 P2_R1203_U165 ; P2_R1203_U432
g22600 not P2_R1203_U139 ; P2_R1203_U433
g22601 nand P2_R1203_U191 P2_R1203_U433 ; P2_R1203_U434
g22602 nand P2_R1203_U139 P2_R1203_U166 ; P2_R1203_U435
g22603 nand P2_U3485 P2_R1203_U67 ; P2_R1203_U436
g22604 nand P2_U3083 P2_R1203_U66 ; P2_R1203_U437
g22605 not P2_R1203_U140 ; P2_R1203_U438
g22606 nand P2_R1203_U273 P2_R1203_U438 ; P2_R1203_U439
g22607 nand P2_R1203_U140 P2_R1203_U167 ; P2_R1203_U440
g22608 nand P2_U3483 P2_R1203_U65 ; P2_R1203_U441
g22609 nand P2_U3084 P2_R1203_U168 ; P2_R1203_U442
g22610 not P2_R1203_U141 ; P2_R1203_U443
g22611 nand P2_R1203_U443 P2_R1203_U269 ; P2_R1203_U444
g22612 nand P2_R1203_U141 P2_R1203_U64 ; P2_R1203_U445
g22613 nand P2_U3480 P2_R1203_U63 ; P2_R1203_U446
g22614 nand P2_U3071 P2_R1203_U62 ; P2_R1203_U447
g22615 not P2_R1203_U142 ; P2_R1203_U448
g22616 nand P2_R1203_U265 P2_R1203_U448 ; P2_R1203_U449
g22617 nand P2_R1203_U142 P2_R1203_U169 ; P2_R1203_U450
g22618 nand P2_U3477 P2_R1203_U58 ; P2_R1203_U451
g22619 nand P2_U3075 P2_R1203_U55 ; P2_R1203_U452
g22620 nand P2_R1203_U452 P2_R1203_U451 ; P2_R1203_U453
g22621 nand P2_U3474 P2_R1203_U59 ; P2_R1203_U454
g22622 nand P2_U3076 P2_R1203_U56 ; P2_R1203_U455
g22623 nand P2_R1203_U338 P2_R1203_U90 ; P2_R1203_U456
g22624 nand P2_R1203_U170 P2_R1203_U330 ; P2_R1203_U457
g22625 nand P2_U3471 P2_R1203_U60 ; P2_R1203_U458
g22626 nand P2_U3081 P2_R1203_U57 ; P2_R1203_U459
g22627 nand P2_R1203_U339 P2_R1203_U172 ; P2_R1203_U460
g22628 nand P2_R1203_U255 P2_R1203_U171 ; P2_R1203_U461
g22629 nand P2_U3468 P2_R1203_U54 ; P2_R1203_U462
g22630 nand P2_U3082 P2_R1203_U53 ; P2_R1203_U463
g22631 not P2_R1203_U145 ; P2_R1203_U464
g22632 nand P2_R1203_U251 P2_R1203_U464 ; P2_R1203_U465
g22633 nand P2_R1203_U145 P2_R1203_U173 ; P2_R1203_U466
g22634 nand P2_U3465 P2_R1203_U52 ; P2_R1203_U467
g22635 nand P2_U3074 P2_R1203_U51 ; P2_R1203_U468
g22636 not P2_R1203_U146 ; P2_R1203_U469
g22637 nand P2_R1203_U247 P2_R1203_U469 ; P2_R1203_U470
g22638 nand P2_R1203_U146 P2_R1203_U174 ; P2_R1203_U471
g22639 nand P2_U3462 P2_R1203_U48 ; P2_R1203_U472
g22640 nand P2_U3065 P2_R1203_U47 ; P2_R1203_U473
g22641 nand P2_R1203_U473 P2_R1203_U472 ; P2_R1203_U474
g22642 nand P2_U3459 P2_R1203_U49 ; P2_R1203_U475
g22643 nand P2_U3064 P2_R1203_U46 ; P2_R1203_U476
g22644 nand P2_R1203_U349 P2_R1203_U91 ; P2_R1203_U477
g22645 nand P2_R1203_U175 P2_R1203_U341 ; P2_R1203_U478
g22646 and P2_R1113_U202 P2_R1113_U201 ; P2_R1113_U6
g22647 and P2_R1113_U241 P2_R1113_U240 ; P2_R1113_U7
g22648 and P2_R1113_U181 P2_R1113_U256 ; P2_R1113_U8
g22649 and P2_R1113_U258 P2_R1113_U257 ; P2_R1113_U9
g22650 and P2_R1113_U182 P2_R1113_U282 ; P2_R1113_U10
g22651 and P2_R1113_U284 P2_R1113_U283 ; P2_R1113_U11
g22652 nand P2_R1113_U344 P2_R1113_U347 ; P2_R1113_U12
g22653 nand P2_R1113_U333 P2_R1113_U336 ; P2_R1113_U13
g22654 nand P2_R1113_U322 P2_R1113_U325 ; P2_R1113_U14
g22655 nand P2_R1113_U314 P2_R1113_U316 ; P2_R1113_U15
g22656 nand P2_R1113_U352 P2_R1113_U312 ; P2_R1113_U16
g22657 nand P2_R1113_U235 P2_R1113_U237 ; P2_R1113_U17
g22658 nand P2_R1113_U227 P2_R1113_U230 ; P2_R1113_U18
g22659 nand P2_R1113_U219 P2_R1113_U221 ; P2_R1113_U19
g22660 nand P2_R1113_U166 P2_R1113_U350 ; P2_R1113_U20
g22661 not P2_U3450 ; P2_R1113_U21
g22662 not P2_U3444 ; P2_R1113_U22
g22663 not P2_U3435 ; P2_R1113_U23
g22664 not P2_U3427 ; P2_R1113_U24
g22665 not P2_U3080 ; P2_R1113_U25
g22666 not P2_U3438 ; P2_R1113_U26
g22667 not P2_U3070 ; P2_R1113_U27
g22668 nand P2_U3070 P2_R1113_U23 ; P2_R1113_U28
g22669 not P2_U3066 ; P2_R1113_U29
g22670 not P2_U3447 ; P2_R1113_U30
g22671 not P2_U3441 ; P2_R1113_U31
g22672 not P2_U3073 ; P2_R1113_U32
g22673 not P2_U3069 ; P2_R1113_U33
g22674 not P2_U3062 ; P2_R1113_U34
g22675 nand P2_U3062 P2_R1113_U31 ; P2_R1113_U35
g22676 not P2_U3453 ; P2_R1113_U36
g22677 not P2_U3072 ; P2_R1113_U37
g22678 nand P2_U3072 P2_R1113_U21 ; P2_R1113_U38
g22679 not P2_U3086 ; P2_R1113_U39
g22680 not P2_U3456 ; P2_R1113_U40
g22681 not P2_U3085 ; P2_R1113_U41
g22682 nand P2_R1113_U208 P2_R1113_U207 ; P2_R1113_U42
g22683 nand P2_R1113_U35 P2_R1113_U223 ; P2_R1113_U43
g22684 nand P2_R1113_U192 P2_R1113_U176 P2_R1113_U351 ; P2_R1113_U44
g22685 not P2_U3951 ; P2_R1113_U45
g22686 not P2_U3459 ; P2_R1113_U46
g22687 not P2_U3462 ; P2_R1113_U47
g22688 not P2_U3065 ; P2_R1113_U48
g22689 not P2_U3064 ; P2_R1113_U49
g22690 nand P2_U3085 P2_R1113_U40 ; P2_R1113_U50
g22691 not P2_U3465 ; P2_R1113_U51
g22692 not P2_U3074 ; P2_R1113_U52
g22693 not P2_U3468 ; P2_R1113_U53
g22694 not P2_U3082 ; P2_R1113_U54
g22695 not P2_U3477 ; P2_R1113_U55
g22696 not P2_U3474 ; P2_R1113_U56
g22697 not P2_U3471 ; P2_R1113_U57
g22698 not P2_U3075 ; P2_R1113_U58
g22699 not P2_U3076 ; P2_R1113_U59
g22700 not P2_U3081 ; P2_R1113_U60
g22701 nand P2_U3081 P2_R1113_U57 ; P2_R1113_U61
g22702 not P2_U3480 ; P2_R1113_U62
g22703 not P2_U3071 ; P2_R1113_U63
g22704 nand P2_R1113_U268 P2_R1113_U267 ; P2_R1113_U64
g22705 not P2_U3084 ; P2_R1113_U65
g22706 not P2_U3485 ; P2_R1113_U66
g22707 not P2_U3083 ; P2_R1113_U67
g22708 not P2_U3957 ; P2_R1113_U68
g22709 not P2_U3078 ; P2_R1113_U69
g22710 not P2_U3954 ; P2_R1113_U70
g22711 not P2_U3955 ; P2_R1113_U71
g22712 not P2_U3956 ; P2_R1113_U72
g22713 not P2_U3068 ; P2_R1113_U73
g22714 not P2_U3063 ; P2_R1113_U74
g22715 not P2_U3077 ; P2_R1113_U75
g22716 nand P2_U3077 P2_R1113_U72 ; P2_R1113_U76
g22717 not P2_U3953 ; P2_R1113_U77
g22718 not P2_U3067 ; P2_R1113_U78
g22719 not P2_U3952 ; P2_R1113_U79
g22720 not P2_U3060 ; P2_R1113_U80
g22721 not P2_U3950 ; P2_R1113_U81
g22722 not P2_U3059 ; P2_R1113_U82
g22723 nand P2_U3059 P2_R1113_U45 ; P2_R1113_U83
g22724 not P2_U3055 ; P2_R1113_U84
g22725 not P2_U3949 ; P2_R1113_U85
g22726 not P2_U3056 ; P2_R1113_U86
g22727 nand P2_R1113_U128 P2_R1113_U301 ; P2_R1113_U87
g22728 nand P2_R1113_U298 P2_R1113_U297 ; P2_R1113_U88
g22729 nand P2_R1113_U76 P2_R1113_U318 ; P2_R1113_U89
g22730 nand P2_R1113_U61 P2_R1113_U329 ; P2_R1113_U90
g22731 nand P2_R1113_U50 P2_R1113_U340 ; P2_R1113_U91
g22732 not P2_U3079 ; P2_R1113_U92
g22733 nand P2_R1113_U395 P2_R1113_U394 ; P2_R1113_U93
g22734 nand P2_R1113_U409 P2_R1113_U408 ; P2_R1113_U94
g22735 nand P2_R1113_U414 P2_R1113_U413 ; P2_R1113_U95
g22736 nand P2_R1113_U430 P2_R1113_U429 ; P2_R1113_U96
g22737 nand P2_R1113_U435 P2_R1113_U434 ; P2_R1113_U97
g22738 nand P2_R1113_U440 P2_R1113_U439 ; P2_R1113_U98
g22739 nand P2_R1113_U445 P2_R1113_U444 ; P2_R1113_U99
g22740 nand P2_R1113_U450 P2_R1113_U449 ; P2_R1113_U100
g22741 nand P2_R1113_U466 P2_R1113_U465 ; P2_R1113_U101
g22742 nand P2_R1113_U471 P2_R1113_U470 ; P2_R1113_U102
g22743 nand P2_R1113_U356 P2_R1113_U355 ; P2_R1113_U103
g22744 nand P2_R1113_U365 P2_R1113_U364 ; P2_R1113_U104
g22745 nand P2_R1113_U372 P2_R1113_U371 ; P2_R1113_U105
g22746 nand P2_R1113_U376 P2_R1113_U375 ; P2_R1113_U106
g22747 nand P2_R1113_U385 P2_R1113_U384 ; P2_R1113_U107
g22748 nand P2_R1113_U404 P2_R1113_U403 ; P2_R1113_U108
g22749 nand P2_R1113_U421 P2_R1113_U420 ; P2_R1113_U109
g22750 nand P2_R1113_U425 P2_R1113_U424 ; P2_R1113_U110
g22751 nand P2_R1113_U457 P2_R1113_U456 ; P2_R1113_U111
g22752 nand P2_R1113_U461 P2_R1113_U460 ; P2_R1113_U112
g22753 nand P2_R1113_U478 P2_R1113_U477 ; P2_R1113_U113
g22754 and P2_R1113_U194 P2_R1113_U184 ; P2_R1113_U114
g22755 and P2_R1113_U197 P2_R1113_U198 ; P2_R1113_U115
g22756 and P2_R1113_U205 P2_R1113_U200 P2_R1113_U185 ; P2_R1113_U116
g22757 and P2_R1113_U210 P2_R1113_U186 ; P2_R1113_U117
g22758 and P2_R1113_U213 P2_R1113_U214 ; P2_R1113_U118
g22759 and P2_R1113_U358 P2_R1113_U357 P2_R1113_U38 ; P2_R1113_U119
g22760 and P2_R1113_U361 P2_R1113_U186 ; P2_R1113_U120
g22761 and P2_R1113_U229 P2_R1113_U6 ; P2_R1113_U121
g22762 and P2_R1113_U368 P2_R1113_U185 ; P2_R1113_U122
g22763 and P2_R1113_U378 P2_R1113_U377 P2_R1113_U28 ; P2_R1113_U123
g22764 and P2_R1113_U381 P2_R1113_U184 ; P2_R1113_U124
g22765 and P2_R1113_U239 P2_R1113_U216 P2_R1113_U180 ; P2_R1113_U125
g22766 and P2_R1113_U261 P2_R1113_U8 ; P2_R1113_U126
g22767 and P2_R1113_U287 P2_R1113_U10 ; P2_R1113_U127
g22768 and P2_R1113_U303 P2_R1113_U304 ; P2_R1113_U128
g22769 and P2_R1113_U387 P2_R1113_U386 P2_R1113_U311 ; P2_R1113_U129
g22770 and P2_R1113_U308 P2_R1113_U390 ; P2_R1113_U130
g22771 nand P2_R1113_U392 P2_R1113_U391 ; P2_R1113_U131
g22772 and P2_R1113_U397 P2_R1113_U396 P2_R1113_U83 ; P2_R1113_U132
g22773 and P2_R1113_U400 P2_R1113_U183 ; P2_R1113_U133
g22774 nand P2_R1113_U406 P2_R1113_U405 ; P2_R1113_U134
g22775 nand P2_R1113_U411 P2_R1113_U410 ; P2_R1113_U135
g22776 and P2_R1113_U324 P2_R1113_U11 ; P2_R1113_U136
g22777 and P2_R1113_U417 P2_R1113_U182 ; P2_R1113_U137
g22778 nand P2_R1113_U427 P2_R1113_U426 ; P2_R1113_U138
g22779 nand P2_R1113_U432 P2_R1113_U431 ; P2_R1113_U139
g22780 nand P2_R1113_U437 P2_R1113_U436 ; P2_R1113_U140
g22781 nand P2_R1113_U442 P2_R1113_U441 ; P2_R1113_U141
g22782 nand P2_R1113_U447 P2_R1113_U446 ; P2_R1113_U142
g22783 and P2_R1113_U335 P2_R1113_U9 ; P2_R1113_U143
g22784 and P2_R1113_U453 P2_R1113_U181 ; P2_R1113_U144
g22785 nand P2_R1113_U463 P2_R1113_U462 ; P2_R1113_U145
g22786 nand P2_R1113_U468 P2_R1113_U467 ; P2_R1113_U146
g22787 and P2_R1113_U346 P2_R1113_U7 ; P2_R1113_U147
g22788 and P2_R1113_U474 P2_R1113_U180 ; P2_R1113_U148
g22789 and P2_R1113_U354 P2_R1113_U353 ; P2_R1113_U149
g22790 nand P2_R1113_U118 P2_R1113_U211 ; P2_R1113_U150
g22791 and P2_R1113_U363 P2_R1113_U362 ; P2_R1113_U151
g22792 and P2_R1113_U370 P2_R1113_U369 ; P2_R1113_U152
g22793 and P2_R1113_U374 P2_R1113_U373 ; P2_R1113_U153
g22794 nand P2_R1113_U115 P2_R1113_U195 ; P2_R1113_U154
g22795 and P2_R1113_U383 P2_R1113_U382 ; P2_R1113_U155
g22796 not P2_U3960 ; P2_R1113_U156
g22797 not P2_U3057 ; P2_R1113_U157
g22798 and P2_R1113_U402 P2_R1113_U401 ; P2_R1113_U158
g22799 nand P2_R1113_U294 P2_R1113_U293 ; P2_R1113_U159
g22800 nand P2_R1113_U290 P2_R1113_U289 ; P2_R1113_U160
g22801 and P2_R1113_U419 P2_R1113_U418 ; P2_R1113_U161
g22802 and P2_R1113_U423 P2_R1113_U422 ; P2_R1113_U162
g22803 nand P2_R1113_U280 P2_R1113_U279 ; P2_R1113_U163
g22804 nand P2_R1113_U276 P2_R1113_U275 ; P2_R1113_U164
g22805 not P2_U3432 ; P2_R1113_U165
g22806 nand P2_U3427 P2_R1113_U92 ; P2_R1113_U166
g22807 nand P2_R1113_U272 P2_R1113_U271 ; P2_R1113_U167
g22808 not P2_U3483 ; P2_R1113_U168
g22809 nand P2_R1113_U264 P2_R1113_U263 ; P2_R1113_U169
g22810 and P2_R1113_U455 P2_R1113_U454 ; P2_R1113_U170
g22811 and P2_R1113_U459 P2_R1113_U458 ; P2_R1113_U171
g22812 nand P2_R1113_U254 P2_R1113_U253 ; P2_R1113_U172
g22813 nand P2_R1113_U250 P2_R1113_U249 ; P2_R1113_U173
g22814 nand P2_R1113_U246 P2_R1113_U245 ; P2_R1113_U174
g22815 and P2_R1113_U476 P2_R1113_U475 ; P2_R1113_U175
g22816 nand P2_R1113_U166 P2_R1113_U165 ; P2_R1113_U176
g22817 not P2_R1113_U83 ; P2_R1113_U177
g22818 not P2_R1113_U28 ; P2_R1113_U178
g22819 not P2_R1113_U38 ; P2_R1113_U179
g22820 nand P2_U3459 P2_R1113_U49 ; P2_R1113_U180
g22821 nand P2_U3474 P2_R1113_U59 ; P2_R1113_U181
g22822 nand P2_U3955 P2_R1113_U74 ; P2_R1113_U182
g22823 nand P2_U3951 P2_R1113_U82 ; P2_R1113_U183
g22824 nand P2_U3435 P2_R1113_U27 ; P2_R1113_U184
g22825 nand P2_U3444 P2_R1113_U33 ; P2_R1113_U185
g22826 nand P2_U3450 P2_R1113_U37 ; P2_R1113_U186
g22827 not P2_R1113_U61 ; P2_R1113_U187
g22828 not P2_R1113_U76 ; P2_R1113_U188
g22829 not P2_R1113_U35 ; P2_R1113_U189
g22830 not P2_R1113_U50 ; P2_R1113_U190
g22831 not P2_R1113_U166 ; P2_R1113_U191
g22832 nand P2_U3080 P2_R1113_U166 ; P2_R1113_U192
g22833 not P2_R1113_U44 ; P2_R1113_U193
g22834 nand P2_U3438 P2_R1113_U29 ; P2_R1113_U194
g22835 nand P2_R1113_U114 P2_R1113_U44 ; P2_R1113_U195
g22836 nand P2_R1113_U29 P2_R1113_U28 ; P2_R1113_U196
g22837 nand P2_R1113_U196 P2_R1113_U26 ; P2_R1113_U197
g22838 nand P2_U3066 P2_R1113_U178 ; P2_R1113_U198
g22839 not P2_R1113_U154 ; P2_R1113_U199
g22840 nand P2_U3447 P2_R1113_U32 ; P2_R1113_U200
g22841 nand P2_U3073 P2_R1113_U30 ; P2_R1113_U201
g22842 nand P2_U3069 P2_R1113_U22 ; P2_R1113_U202
g22843 nand P2_R1113_U189 P2_R1113_U185 ; P2_R1113_U203
g22844 nand P2_R1113_U6 P2_R1113_U203 ; P2_R1113_U204
g22845 nand P2_U3441 P2_R1113_U34 ; P2_R1113_U205
g22846 nand P2_U3447 P2_R1113_U32 ; P2_R1113_U206
g22847 nand P2_R1113_U154 P2_R1113_U116 ; P2_R1113_U207
g22848 nand P2_R1113_U206 P2_R1113_U204 ; P2_R1113_U208
g22849 not P2_R1113_U42 ; P2_R1113_U209
g22850 nand P2_U3453 P2_R1113_U39 ; P2_R1113_U210
g22851 nand P2_R1113_U117 P2_R1113_U42 ; P2_R1113_U211
g22852 nand P2_R1113_U39 P2_R1113_U38 ; P2_R1113_U212
g22853 nand P2_R1113_U212 P2_R1113_U36 ; P2_R1113_U213
g22854 nand P2_U3086 P2_R1113_U179 ; P2_R1113_U214
g22855 not P2_R1113_U150 ; P2_R1113_U215
g22856 nand P2_U3456 P2_R1113_U41 ; P2_R1113_U216
g22857 nand P2_R1113_U216 P2_R1113_U50 ; P2_R1113_U217
g22858 nand P2_R1113_U209 P2_R1113_U38 ; P2_R1113_U218
g22859 nand P2_R1113_U120 P2_R1113_U218 ; P2_R1113_U219
g22860 nand P2_R1113_U42 P2_R1113_U186 ; P2_R1113_U220
g22861 nand P2_R1113_U119 P2_R1113_U220 ; P2_R1113_U221
g22862 nand P2_R1113_U38 P2_R1113_U186 ; P2_R1113_U222
g22863 nand P2_R1113_U205 P2_R1113_U154 ; P2_R1113_U223
g22864 not P2_R1113_U43 ; P2_R1113_U224
g22865 nand P2_U3069 P2_R1113_U22 ; P2_R1113_U225
g22866 nand P2_R1113_U224 P2_R1113_U225 ; P2_R1113_U226
g22867 nand P2_R1113_U122 P2_R1113_U226 ; P2_R1113_U227
g22868 nand P2_R1113_U43 P2_R1113_U185 ; P2_R1113_U228
g22869 nand P2_U3447 P2_R1113_U32 ; P2_R1113_U229
g22870 nand P2_R1113_U121 P2_R1113_U228 ; P2_R1113_U230
g22871 nand P2_U3069 P2_R1113_U22 ; P2_R1113_U231
g22872 nand P2_R1113_U185 P2_R1113_U231 ; P2_R1113_U232
g22873 nand P2_R1113_U205 P2_R1113_U35 ; P2_R1113_U233
g22874 nand P2_R1113_U193 P2_R1113_U28 ; P2_R1113_U234
g22875 nand P2_R1113_U124 P2_R1113_U234 ; P2_R1113_U235
g22876 nand P2_R1113_U44 P2_R1113_U184 ; P2_R1113_U236
g22877 nand P2_R1113_U123 P2_R1113_U236 ; P2_R1113_U237
g22878 nand P2_R1113_U28 P2_R1113_U184 ; P2_R1113_U238
g22879 nand P2_U3462 P2_R1113_U48 ; P2_R1113_U239
g22880 nand P2_U3065 P2_R1113_U47 ; P2_R1113_U240
g22881 nand P2_U3064 P2_R1113_U46 ; P2_R1113_U241
g22882 nand P2_R1113_U190 P2_R1113_U180 ; P2_R1113_U242
g22883 nand P2_R1113_U7 P2_R1113_U242 ; P2_R1113_U243
g22884 nand P2_U3462 P2_R1113_U48 ; P2_R1113_U244
g22885 nand P2_R1113_U150 P2_R1113_U125 ; P2_R1113_U245
g22886 nand P2_R1113_U244 P2_R1113_U243 ; P2_R1113_U246
g22887 not P2_R1113_U174 ; P2_R1113_U247
g22888 nand P2_U3465 P2_R1113_U52 ; P2_R1113_U248
g22889 nand P2_R1113_U248 P2_R1113_U174 ; P2_R1113_U249
g22890 nand P2_U3074 P2_R1113_U51 ; P2_R1113_U250
g22891 not P2_R1113_U173 ; P2_R1113_U251
g22892 nand P2_U3468 P2_R1113_U54 ; P2_R1113_U252
g22893 nand P2_R1113_U252 P2_R1113_U173 ; P2_R1113_U253
g22894 nand P2_U3082 P2_R1113_U53 ; P2_R1113_U254
g22895 not P2_R1113_U172 ; P2_R1113_U255
g22896 nand P2_U3477 P2_R1113_U58 ; P2_R1113_U256
g22897 nand P2_U3075 P2_R1113_U55 ; P2_R1113_U257
g22898 nand P2_U3076 P2_R1113_U56 ; P2_R1113_U258
g22899 nand P2_R1113_U187 P2_R1113_U8 ; P2_R1113_U259
g22900 nand P2_R1113_U9 P2_R1113_U259 ; P2_R1113_U260
g22901 nand P2_U3471 P2_R1113_U60 ; P2_R1113_U261
g22902 nand P2_U3477 P2_R1113_U58 ; P2_R1113_U262
g22903 nand P2_R1113_U126 P2_R1113_U172 ; P2_R1113_U263
g22904 nand P2_R1113_U262 P2_R1113_U260 ; P2_R1113_U264
g22905 not P2_R1113_U169 ; P2_R1113_U265
g22906 nand P2_U3480 P2_R1113_U63 ; P2_R1113_U266
g22907 nand P2_R1113_U266 P2_R1113_U169 ; P2_R1113_U267
g22908 nand P2_U3071 P2_R1113_U62 ; P2_R1113_U268
g22909 not P2_R1113_U64 ; P2_R1113_U269
g22910 nand P2_R1113_U269 P2_R1113_U65 ; P2_R1113_U270
g22911 nand P2_R1113_U270 P2_R1113_U168 ; P2_R1113_U271
g22912 nand P2_U3084 P2_R1113_U64 ; P2_R1113_U272
g22913 not P2_R1113_U167 ; P2_R1113_U273
g22914 nand P2_U3485 P2_R1113_U67 ; P2_R1113_U274
g22915 nand P2_R1113_U274 P2_R1113_U167 ; P2_R1113_U275
g22916 nand P2_U3083 P2_R1113_U66 ; P2_R1113_U276
g22917 not P2_R1113_U164 ; P2_R1113_U277
g22918 nand P2_U3957 P2_R1113_U69 ; P2_R1113_U278
g22919 nand P2_R1113_U278 P2_R1113_U164 ; P2_R1113_U279
g22920 nand P2_U3078 P2_R1113_U68 ; P2_R1113_U280
g22921 not P2_R1113_U163 ; P2_R1113_U281
g22922 nand P2_U3954 P2_R1113_U73 ; P2_R1113_U282
g22923 nand P2_U3068 P2_R1113_U70 ; P2_R1113_U283
g22924 nand P2_U3063 P2_R1113_U71 ; P2_R1113_U284
g22925 nand P2_R1113_U188 P2_R1113_U10 ; P2_R1113_U285
g22926 nand P2_R1113_U11 P2_R1113_U285 ; P2_R1113_U286
g22927 nand P2_U3956 P2_R1113_U75 ; P2_R1113_U287
g22928 nand P2_U3954 P2_R1113_U73 ; P2_R1113_U288
g22929 nand P2_R1113_U127 P2_R1113_U163 ; P2_R1113_U289
g22930 nand P2_R1113_U288 P2_R1113_U286 ; P2_R1113_U290
g22931 not P2_R1113_U160 ; P2_R1113_U291
g22932 nand P2_U3953 P2_R1113_U78 ; P2_R1113_U292
g22933 nand P2_R1113_U292 P2_R1113_U160 ; P2_R1113_U293
g22934 nand P2_U3067 P2_R1113_U77 ; P2_R1113_U294
g22935 not P2_R1113_U159 ; P2_R1113_U295
g22936 nand P2_U3952 P2_R1113_U80 ; P2_R1113_U296
g22937 nand P2_R1113_U296 P2_R1113_U159 ; P2_R1113_U297
g22938 nand P2_U3060 P2_R1113_U79 ; P2_R1113_U298
g22939 not P2_R1113_U88 ; P2_R1113_U299
g22940 nand P2_U3950 P2_R1113_U84 ; P2_R1113_U300
g22941 nand P2_R1113_U88 P2_R1113_U183 P2_R1113_U300 ; P2_R1113_U301
g22942 nand P2_R1113_U84 P2_R1113_U83 ; P2_R1113_U302
g22943 nand P2_R1113_U302 P2_R1113_U81 ; P2_R1113_U303
g22944 nand P2_U3055 P2_R1113_U177 ; P2_R1113_U304
g22945 not P2_R1113_U87 ; P2_R1113_U305
g22946 nand P2_U3056 P2_R1113_U85 ; P2_R1113_U306
g22947 nand P2_R1113_U305 P2_R1113_U306 ; P2_R1113_U307
g22948 nand P2_U3949 P2_R1113_U86 ; P2_R1113_U308
g22949 nand P2_U3949 P2_R1113_U86 ; P2_R1113_U309
g22950 nand P2_R1113_U309 P2_R1113_U87 ; P2_R1113_U310
g22951 nand P2_U3056 P2_R1113_U85 ; P2_R1113_U311
g22952 nand P2_R1113_U129 P2_R1113_U310 ; P2_R1113_U312
g22953 nand P2_R1113_U299 P2_R1113_U83 ; P2_R1113_U313
g22954 nand P2_R1113_U133 P2_R1113_U313 ; P2_R1113_U314
g22955 nand P2_R1113_U88 P2_R1113_U183 ; P2_R1113_U315
g22956 nand P2_R1113_U132 P2_R1113_U315 ; P2_R1113_U316
g22957 nand P2_R1113_U83 P2_R1113_U183 ; P2_R1113_U317
g22958 nand P2_R1113_U287 P2_R1113_U163 ; P2_R1113_U318
g22959 not P2_R1113_U89 ; P2_R1113_U319
g22960 nand P2_U3063 P2_R1113_U71 ; P2_R1113_U320
g22961 nand P2_R1113_U319 P2_R1113_U320 ; P2_R1113_U321
g22962 nand P2_R1113_U137 P2_R1113_U321 ; P2_R1113_U322
g22963 nand P2_R1113_U89 P2_R1113_U182 ; P2_R1113_U323
g22964 nand P2_U3954 P2_R1113_U73 ; P2_R1113_U324
g22965 nand P2_R1113_U136 P2_R1113_U323 ; P2_R1113_U325
g22966 nand P2_U3063 P2_R1113_U71 ; P2_R1113_U326
g22967 nand P2_R1113_U182 P2_R1113_U326 ; P2_R1113_U327
g22968 nand P2_R1113_U287 P2_R1113_U76 ; P2_R1113_U328
g22969 nand P2_R1113_U261 P2_R1113_U172 ; P2_R1113_U329
g22970 not P2_R1113_U90 ; P2_R1113_U330
g22971 nand P2_U3076 P2_R1113_U56 ; P2_R1113_U331
g22972 nand P2_R1113_U330 P2_R1113_U331 ; P2_R1113_U332
g22973 nand P2_R1113_U144 P2_R1113_U332 ; P2_R1113_U333
g22974 nand P2_R1113_U90 P2_R1113_U181 ; P2_R1113_U334
g22975 nand P2_U3477 P2_R1113_U58 ; P2_R1113_U335
g22976 nand P2_R1113_U143 P2_R1113_U334 ; P2_R1113_U336
g22977 nand P2_U3076 P2_R1113_U56 ; P2_R1113_U337
g22978 nand P2_R1113_U181 P2_R1113_U337 ; P2_R1113_U338
g22979 nand P2_R1113_U261 P2_R1113_U61 ; P2_R1113_U339
g22980 nand P2_R1113_U216 P2_R1113_U150 ; P2_R1113_U340
g22981 not P2_R1113_U91 ; P2_R1113_U341
g22982 nand P2_U3064 P2_R1113_U46 ; P2_R1113_U342
g22983 nand P2_R1113_U341 P2_R1113_U342 ; P2_R1113_U343
g22984 nand P2_R1113_U148 P2_R1113_U343 ; P2_R1113_U344
g22985 nand P2_R1113_U91 P2_R1113_U180 ; P2_R1113_U345
g22986 nand P2_U3462 P2_R1113_U48 ; P2_R1113_U346
g22987 nand P2_R1113_U147 P2_R1113_U345 ; P2_R1113_U347
g22988 nand P2_U3064 P2_R1113_U46 ; P2_R1113_U348
g22989 nand P2_R1113_U180 P2_R1113_U348 ; P2_R1113_U349
g22990 nand P2_U3079 P2_R1113_U24 ; P2_R1113_U350
g22991 nand P2_U3080 P2_R1113_U165 ; P2_R1113_U351
g22992 nand P2_R1113_U130 P2_R1113_U307 ; P2_R1113_U352
g22993 nand P2_U3456 P2_R1113_U41 ; P2_R1113_U353
g22994 nand P2_U3085 P2_R1113_U40 ; P2_R1113_U354
g22995 nand P2_R1113_U217 P2_R1113_U150 ; P2_R1113_U355
g22996 nand P2_R1113_U215 P2_R1113_U149 ; P2_R1113_U356
g22997 nand P2_U3453 P2_R1113_U39 ; P2_R1113_U357
g22998 nand P2_U3086 P2_R1113_U36 ; P2_R1113_U358
g22999 nand P2_U3453 P2_R1113_U39 ; P2_R1113_U359
g23000 nand P2_U3086 P2_R1113_U36 ; P2_R1113_U360
g23001 nand P2_R1113_U360 P2_R1113_U359 ; P2_R1113_U361
g23002 nand P2_U3450 P2_R1113_U37 ; P2_R1113_U362
g23003 nand P2_U3072 P2_R1113_U21 ; P2_R1113_U363
g23004 nand P2_R1113_U222 P2_R1113_U42 ; P2_R1113_U364
g23005 nand P2_R1113_U151 P2_R1113_U209 ; P2_R1113_U365
g23006 nand P2_U3447 P2_R1113_U32 ; P2_R1113_U366
g23007 nand P2_U3073 P2_R1113_U30 ; P2_R1113_U367
g23008 nand P2_R1113_U367 P2_R1113_U366 ; P2_R1113_U368
g23009 nand P2_U3444 P2_R1113_U33 ; P2_R1113_U369
g23010 nand P2_U3069 P2_R1113_U22 ; P2_R1113_U370
g23011 nand P2_R1113_U232 P2_R1113_U43 ; P2_R1113_U371
g23012 nand P2_R1113_U152 P2_R1113_U224 ; P2_R1113_U372
g23013 nand P2_U3441 P2_R1113_U34 ; P2_R1113_U373
g23014 nand P2_U3062 P2_R1113_U31 ; P2_R1113_U374
g23015 nand P2_R1113_U233 P2_R1113_U154 ; P2_R1113_U375
g23016 nand P2_R1113_U199 P2_R1113_U153 ; P2_R1113_U376
g23017 nand P2_U3438 P2_R1113_U29 ; P2_R1113_U377
g23018 nand P2_U3066 P2_R1113_U26 ; P2_R1113_U378
g23019 nand P2_U3438 P2_R1113_U29 ; P2_R1113_U379
g23020 nand P2_U3066 P2_R1113_U26 ; P2_R1113_U380
g23021 nand P2_R1113_U380 P2_R1113_U379 ; P2_R1113_U381
g23022 nand P2_U3435 P2_R1113_U27 ; P2_R1113_U382
g23023 nand P2_U3070 P2_R1113_U23 ; P2_R1113_U383
g23024 nand P2_R1113_U238 P2_R1113_U44 ; P2_R1113_U384
g23025 nand P2_R1113_U155 P2_R1113_U193 ; P2_R1113_U385
g23026 nand P2_U3960 P2_R1113_U157 ; P2_R1113_U386
g23027 nand P2_U3057 P2_R1113_U156 ; P2_R1113_U387
g23028 nand P2_U3960 P2_R1113_U157 ; P2_R1113_U388
g23029 nand P2_U3057 P2_R1113_U156 ; P2_R1113_U389
g23030 nand P2_R1113_U389 P2_R1113_U388 ; P2_R1113_U390
g23031 nand P2_U3949 P2_R1113_U86 ; P2_R1113_U391
g23032 nand P2_U3056 P2_R1113_U85 ; P2_R1113_U392
g23033 not P2_R1113_U131 ; P2_R1113_U393
g23034 nand P2_R1113_U393 P2_R1113_U305 ; P2_R1113_U394
g23035 nand P2_R1113_U131 P2_R1113_U87 ; P2_R1113_U395
g23036 nand P2_U3950 P2_R1113_U84 ; P2_R1113_U396
g23037 nand P2_U3055 P2_R1113_U81 ; P2_R1113_U397
g23038 nand P2_U3950 P2_R1113_U84 ; P2_R1113_U398
g23039 nand P2_U3055 P2_R1113_U81 ; P2_R1113_U399
g23040 nand P2_R1113_U399 P2_R1113_U398 ; P2_R1113_U400
g23041 nand P2_U3951 P2_R1113_U82 ; P2_R1113_U401
g23042 nand P2_U3059 P2_R1113_U45 ; P2_R1113_U402
g23043 nand P2_R1113_U317 P2_R1113_U88 ; P2_R1113_U403
g23044 nand P2_R1113_U158 P2_R1113_U299 ; P2_R1113_U404
g23045 nand P2_U3952 P2_R1113_U80 ; P2_R1113_U405
g23046 nand P2_U3060 P2_R1113_U79 ; P2_R1113_U406
g23047 not P2_R1113_U134 ; P2_R1113_U407
g23048 nand P2_R1113_U295 P2_R1113_U407 ; P2_R1113_U408
g23049 nand P2_R1113_U134 P2_R1113_U159 ; P2_R1113_U409
g23050 nand P2_U3953 P2_R1113_U78 ; P2_R1113_U410
g23051 nand P2_U3067 P2_R1113_U77 ; P2_R1113_U411
g23052 not P2_R1113_U135 ; P2_R1113_U412
g23053 nand P2_R1113_U291 P2_R1113_U412 ; P2_R1113_U413
g23054 nand P2_R1113_U135 P2_R1113_U160 ; P2_R1113_U414
g23055 nand P2_U3954 P2_R1113_U73 ; P2_R1113_U415
g23056 nand P2_U3068 P2_R1113_U70 ; P2_R1113_U416
g23057 nand P2_R1113_U416 P2_R1113_U415 ; P2_R1113_U417
g23058 nand P2_U3955 P2_R1113_U74 ; P2_R1113_U418
g23059 nand P2_U3063 P2_R1113_U71 ; P2_R1113_U419
g23060 nand P2_R1113_U327 P2_R1113_U89 ; P2_R1113_U420
g23061 nand P2_R1113_U161 P2_R1113_U319 ; P2_R1113_U421
g23062 nand P2_U3956 P2_R1113_U75 ; P2_R1113_U422
g23063 nand P2_U3077 P2_R1113_U72 ; P2_R1113_U423
g23064 nand P2_R1113_U328 P2_R1113_U163 ; P2_R1113_U424
g23065 nand P2_R1113_U281 P2_R1113_U162 ; P2_R1113_U425
g23066 nand P2_U3957 P2_R1113_U69 ; P2_R1113_U426
g23067 nand P2_U3078 P2_R1113_U68 ; P2_R1113_U427
g23068 not P2_R1113_U138 ; P2_R1113_U428
g23069 nand P2_R1113_U277 P2_R1113_U428 ; P2_R1113_U429
g23070 nand P2_R1113_U138 P2_R1113_U164 ; P2_R1113_U430
g23071 nand P2_U3432 P2_R1113_U25 ; P2_R1113_U431
g23072 nand P2_U3080 P2_R1113_U165 ; P2_R1113_U432
g23073 not P2_R1113_U139 ; P2_R1113_U433
g23074 nand P2_R1113_U191 P2_R1113_U433 ; P2_R1113_U434
g23075 nand P2_R1113_U139 P2_R1113_U166 ; P2_R1113_U435
g23076 nand P2_U3485 P2_R1113_U67 ; P2_R1113_U436
g23077 nand P2_U3083 P2_R1113_U66 ; P2_R1113_U437
g23078 not P2_R1113_U140 ; P2_R1113_U438
g23079 nand P2_R1113_U273 P2_R1113_U438 ; P2_R1113_U439
g23080 nand P2_R1113_U140 P2_R1113_U167 ; P2_R1113_U440
g23081 nand P2_U3483 P2_R1113_U65 ; P2_R1113_U441
g23082 nand P2_U3084 P2_R1113_U168 ; P2_R1113_U442
g23083 not P2_R1113_U141 ; P2_R1113_U443
g23084 nand P2_R1113_U443 P2_R1113_U269 ; P2_R1113_U444
g23085 nand P2_R1113_U141 P2_R1113_U64 ; P2_R1113_U445
g23086 nand P2_U3480 P2_R1113_U63 ; P2_R1113_U446
g23087 nand P2_U3071 P2_R1113_U62 ; P2_R1113_U447
g23088 not P2_R1113_U142 ; P2_R1113_U448
g23089 nand P2_R1113_U265 P2_R1113_U448 ; P2_R1113_U449
g23090 nand P2_R1113_U142 P2_R1113_U169 ; P2_R1113_U450
g23091 nand P2_U3477 P2_R1113_U58 ; P2_R1113_U451
g23092 nand P2_U3075 P2_R1113_U55 ; P2_R1113_U452
g23093 nand P2_R1113_U452 P2_R1113_U451 ; P2_R1113_U453
g23094 nand P2_U3474 P2_R1113_U59 ; P2_R1113_U454
g23095 nand P2_U3076 P2_R1113_U56 ; P2_R1113_U455
g23096 nand P2_R1113_U338 P2_R1113_U90 ; P2_R1113_U456
g23097 nand P2_R1113_U170 P2_R1113_U330 ; P2_R1113_U457
g23098 nand P2_U3471 P2_R1113_U60 ; P2_R1113_U458
g23099 nand P2_U3081 P2_R1113_U57 ; P2_R1113_U459
g23100 nand P2_R1113_U339 P2_R1113_U172 ; P2_R1113_U460
g23101 nand P2_R1113_U255 P2_R1113_U171 ; P2_R1113_U461
g23102 nand P2_U3468 P2_R1113_U54 ; P2_R1113_U462
g23103 nand P2_U3082 P2_R1113_U53 ; P2_R1113_U463
g23104 not P2_R1113_U145 ; P2_R1113_U464
g23105 nand P2_R1113_U251 P2_R1113_U464 ; P2_R1113_U465
g23106 nand P2_R1113_U145 P2_R1113_U173 ; P2_R1113_U466
g23107 nand P2_U3465 P2_R1113_U52 ; P2_R1113_U467
g23108 nand P2_U3074 P2_R1113_U51 ; P2_R1113_U468
g23109 not P2_R1113_U146 ; P2_R1113_U469
g23110 nand P2_R1113_U247 P2_R1113_U469 ; P2_R1113_U470
g23111 nand P2_R1113_U146 P2_R1113_U174 ; P2_R1113_U471
g23112 nand P2_U3462 P2_R1113_U48 ; P2_R1113_U472
g23113 nand P2_U3065 P2_R1113_U47 ; P2_R1113_U473
g23114 nand P2_R1113_U473 P2_R1113_U472 ; P2_R1113_U474
g23115 nand P2_U3459 P2_R1113_U49 ; P2_R1113_U475
g23116 nand P2_U3064 P2_R1113_U46 ; P2_R1113_U476
g23117 nand P2_R1113_U349 P2_R1113_U91 ; P2_R1113_U477
g23118 nand P2_R1113_U175 P2_R1113_U341 ; P2_R1113_U478
g23119 nor P3_IR_REG_17__SCAN_IN P3_IR_REG_18__SCAN_IN P3_IR_REG_19__SCAN_IN P3_IR_REG_20__SCAN_IN ; P3_SUB_598_U6
g23120 and P3_SUB_598_U136 P3_SUB_598_U49 ; P3_SUB_598_U7
g23121 and P3_SUB_598_U134 P3_SUB_598_U102 ; P3_SUB_598_U8
g23122 and P3_SUB_598_U133 P3_SUB_598_U46 ; P3_SUB_598_U9
g23123 and P3_SUB_598_U132 P3_SUB_598_U47 ; P3_SUB_598_U10
g23124 and P3_SUB_598_U130 P3_SUB_598_U105 ; P3_SUB_598_U11
g23125 and P3_SUB_598_U129 P3_SUB_598_U34 ; P3_SUB_598_U12
g23126 and P3_SUB_598_U128 P3_SUB_598_U44 ; P3_SUB_598_U13
g23127 and P3_SUB_598_U126 P3_SUB_598_U108 ; P3_SUB_598_U14
g23128 and P3_SUB_598_U125 P3_SUB_598_U40 ; P3_SUB_598_U15
g23129 and P3_SUB_598_U124 P3_SUB_598_U41 ; P3_SUB_598_U16
g23130 and P3_SUB_598_U122 P3_SUB_598_U111 ; P3_SUB_598_U17
g23131 and P3_SUB_598_U121 P3_SUB_598_U35 ; P3_SUB_598_U18
g23132 and P3_SUB_598_U120 P3_SUB_598_U78 ; P3_SUB_598_U19
g23133 and P3_SUB_598_U65 P3_SUB_598_U139 ; P3_SUB_598_U20
g23134 and P3_SUB_598_U118 P3_SUB_598_U37 ; P3_SUB_598_U21
g23135 and P3_SUB_598_U117 P3_SUB_598_U28 ; P3_SUB_598_U22
g23136 and P3_SUB_598_U100 P3_SUB_598_U90 ; P3_SUB_598_U23
g23137 and P3_SUB_598_U99 P3_SUB_598_U30 ; P3_SUB_598_U24
g23138 and P3_SUB_598_U98 P3_SUB_598_U31 ; P3_SUB_598_U25
g23139 and P3_SUB_598_U96 P3_SUB_598_U93 ; P3_SUB_598_U26
g23140 and P3_SUB_598_U95 P3_SUB_598_U29 ; P3_SUB_598_U27
g23141 or P3_IR_REG_0__SCAN_IN P3_IR_REG_1__SCAN_IN P3_IR_REG_2__SCAN_IN ; P3_SUB_598_U28
g23142 nand P3_SUB_598_U54 P3_SUB_598_U140 P3_SUB_598_U53 ; P3_SUB_598_U29
g23143 nand P3_SUB_598_U55 P3_SUB_598_U140 ; P3_SUB_598_U30
g23144 nand P3_SUB_598_U56 P3_SUB_598_U91 ; P3_SUB_598_U31
g23145 not P3_IR_REG_7__SCAN_IN ; P3_SUB_598_U32
g23146 not P3_IR_REG_3__SCAN_IN ; P3_SUB_598_U33
g23147 nand P3_SUB_598_U60 P3_SUB_598_U59 P3_SUB_598_U58 P3_SUB_598_U57 ; P3_SUB_598_U34
g23148 nand P3_SUB_598_U62 P3_SUB_598_U106 ; P3_SUB_598_U35
g23149 nand P3_SUB_598_U63 P3_SUB_598_U112 ; P3_SUB_598_U36
g23150 nand P3_SUB_598_U114 P3_SUB_598_U38 ; P3_SUB_598_U37
g23151 not P3_IR_REG_29__SCAN_IN ; P3_SUB_598_U38
g23152 not P3_IR_REG_27__SCAN_IN ; P3_SUB_598_U39
g23153 nand P3_SUB_598_U106 P3_SUB_598_U6 ; P3_SUB_598_U40
g23154 nand P3_SUB_598_U66 P3_SUB_598_U109 ; P3_SUB_598_U41
g23155 not P3_IR_REG_24__SCAN_IN ; P3_SUB_598_U42
g23156 not P3_IR_REG_23__SCAN_IN ; P3_SUB_598_U43
g23157 nand P3_SUB_598_U67 P3_SUB_598_U106 ; P3_SUB_598_U44
g23158 not P3_IR_REG_19__SCAN_IN ; P3_SUB_598_U45
g23159 nand P3_SUB_598_U68 P3_SUB_598_U94 ; P3_SUB_598_U46
g23160 nand P3_SUB_598_U69 P3_SUB_598_U103 ; P3_SUB_598_U47
g23161 not P3_IR_REG_15__SCAN_IN ; P3_SUB_598_U48
g23162 nand P3_SUB_598_U70 P3_SUB_598_U94 ; P3_SUB_598_U49
g23163 not P3_IR_REG_11__SCAN_IN ; P3_SUB_598_U50
g23164 nand P3_SUB_598_U156 P3_SUB_598_U155 ; P3_SUB_598_U51
g23165 nand P3_SUB_598_U146 P3_SUB_598_U145 ; P3_SUB_598_U52
g23166 nor P3_IR_REG_3__SCAN_IN P3_IR_REG_4__SCAN_IN P3_IR_REG_5__SCAN_IN P3_IR_REG_6__SCAN_IN ; P3_SUB_598_U53
g23167 nor P3_IR_REG_7__SCAN_IN P3_IR_REG_8__SCAN_IN ; P3_SUB_598_U54
g23168 nor P3_IR_REG_3__SCAN_IN P3_IR_REG_4__SCAN_IN ; P3_SUB_598_U55
g23169 nor P3_IR_REG_5__SCAN_IN P3_IR_REG_6__SCAN_IN ; P3_SUB_598_U56
g23170 nor P3_IR_REG_10__SCAN_IN P3_IR_REG_11__SCAN_IN P3_IR_REG_12__SCAN_IN P3_IR_REG_13__SCAN_IN P3_IR_REG_14__SCAN_IN ; P3_SUB_598_U57
g23171 nor P3_IR_REG_0__SCAN_IN P3_IR_REG_1__SCAN_IN P3_IR_REG_15__SCAN_IN P3_IR_REG_16__SCAN_IN ; P3_SUB_598_U58
g23172 nor P3_IR_REG_2__SCAN_IN P3_IR_REG_3__SCAN_IN P3_IR_REG_4__SCAN_IN P3_IR_REG_5__SCAN_IN ; P3_SUB_598_U59
g23173 nor P3_IR_REG_6__SCAN_IN P3_IR_REG_7__SCAN_IN P3_IR_REG_8__SCAN_IN P3_IR_REG_9__SCAN_IN ; P3_SUB_598_U60
g23174 nor P3_IR_REG_21__SCAN_IN P3_IR_REG_22__SCAN_IN P3_IR_REG_23__SCAN_IN ; P3_SUB_598_U61
g23175 and P3_SUB_598_U6 P3_SUB_598_U42 P3_SUB_598_U61 ; P3_SUB_598_U62
g23176 nor P3_IR_REG_25__SCAN_IN P3_IR_REG_26__SCAN_IN P3_IR_REG_27__SCAN_IN P3_IR_REG_28__SCAN_IN ; P3_SUB_598_U63
g23177 nor P3_IR_REG_25__SCAN_IN P3_IR_REG_26__SCAN_IN ; P3_SUB_598_U64
g23178 and P3_SUB_598_U138 P3_SUB_598_U36 ; P3_SUB_598_U65
g23179 nor P3_IR_REG_21__SCAN_IN P3_IR_REG_22__SCAN_IN ; P3_SUB_598_U66
g23180 nor P3_IR_REG_17__SCAN_IN P3_IR_REG_18__SCAN_IN ; P3_SUB_598_U67
g23181 nor P3_IR_REG_9__SCAN_IN P3_IR_REG_10__SCAN_IN P3_IR_REG_11__SCAN_IN P3_IR_REG_12__SCAN_IN ; P3_SUB_598_U68
g23182 nor P3_IR_REG_13__SCAN_IN P3_IR_REG_14__SCAN_IN ; P3_SUB_598_U69
g23183 nor P3_IR_REG_9__SCAN_IN P3_IR_REG_10__SCAN_IN ; P3_SUB_598_U70
g23184 not P3_IR_REG_9__SCAN_IN ; P3_SUB_598_U71
g23185 and P3_SUB_598_U142 P3_SUB_598_U141 ; P3_SUB_598_U72
g23186 not P3_IR_REG_5__SCAN_IN ; P3_SUB_598_U73
g23187 and P3_SUB_598_U144 P3_SUB_598_U143 ; P3_SUB_598_U74
g23188 not P3_IR_REG_31__SCAN_IN ; P3_SUB_598_U75
g23189 not P3_IR_REG_30__SCAN_IN ; P3_SUB_598_U76
g23190 and P3_SUB_598_U148 P3_SUB_598_U147 ; P3_SUB_598_U77
g23191 nand P3_SUB_598_U64 P3_SUB_598_U112 ; P3_SUB_598_U78
g23192 and P3_SUB_598_U150 P3_SUB_598_U149 ; P3_SUB_598_U79
g23193 not P3_IR_REG_25__SCAN_IN ; P3_SUB_598_U80
g23194 and P3_SUB_598_U152 P3_SUB_598_U151 ; P3_SUB_598_U81
g23195 not P3_IR_REG_21__SCAN_IN ; P3_SUB_598_U82
g23196 and P3_SUB_598_U154 P3_SUB_598_U153 ; P3_SUB_598_U83
g23197 not P3_IR_REG_1__SCAN_IN ; P3_SUB_598_U84
g23198 not P3_IR_REG_0__SCAN_IN ; P3_SUB_598_U85
g23199 not P3_IR_REG_17__SCAN_IN ; P3_SUB_598_U86
g23200 and P3_SUB_598_U158 P3_SUB_598_U157 ; P3_SUB_598_U87
g23201 not P3_IR_REG_13__SCAN_IN ; P3_SUB_598_U88
g23202 and P3_SUB_598_U160 P3_SUB_598_U159 ; P3_SUB_598_U89
g23203 nand P3_SUB_598_U140 P3_SUB_598_U33 ; P3_SUB_598_U90
g23204 not P3_SUB_598_U30 ; P3_SUB_598_U91
g23205 not P3_SUB_598_U31 ; P3_SUB_598_U92
g23206 nand P3_SUB_598_U92 P3_SUB_598_U32 ; P3_SUB_598_U93
g23207 not P3_SUB_598_U29 ; P3_SUB_598_U94
g23208 nand P3_SUB_598_U93 P3_IR_REG_8__SCAN_IN ; P3_SUB_598_U95
g23209 nand P3_SUB_598_U31 P3_IR_REG_7__SCAN_IN ; P3_SUB_598_U96
g23210 nand P3_SUB_598_U91 P3_SUB_598_U73 ; P3_SUB_598_U97
g23211 nand P3_SUB_598_U97 P3_IR_REG_6__SCAN_IN ; P3_SUB_598_U98
g23212 nand P3_SUB_598_U90 P3_IR_REG_4__SCAN_IN ; P3_SUB_598_U99
g23213 nand P3_SUB_598_U28 P3_IR_REG_3__SCAN_IN ; P3_SUB_598_U100
g23214 not P3_SUB_598_U49 ; P3_SUB_598_U101
g23215 nand P3_SUB_598_U101 P3_SUB_598_U50 ; P3_SUB_598_U102
g23216 not P3_SUB_598_U46 ; P3_SUB_598_U103
g23217 not P3_SUB_598_U47 ; P3_SUB_598_U104
g23218 nand P3_SUB_598_U104 P3_SUB_598_U48 ; P3_SUB_598_U105
g23219 not P3_SUB_598_U34 ; P3_SUB_598_U106
g23220 not P3_SUB_598_U44 ; P3_SUB_598_U107
g23221 nand P3_SUB_598_U107 P3_SUB_598_U45 ; P3_SUB_598_U108
g23222 not P3_SUB_598_U40 ; P3_SUB_598_U109
g23223 not P3_SUB_598_U41 ; P3_SUB_598_U110
g23224 nand P3_SUB_598_U110 P3_SUB_598_U43 ; P3_SUB_598_U111
g23225 not P3_SUB_598_U35 ; P3_SUB_598_U112
g23226 not P3_SUB_598_U78 ; P3_SUB_598_U113
g23227 not P3_SUB_598_U36 ; P3_SUB_598_U114
g23228 not P3_SUB_598_U37 ; P3_SUB_598_U115
g23229 or P3_IR_REG_0__SCAN_IN P3_IR_REG_1__SCAN_IN ; P3_SUB_598_U116
g23230 nand P3_SUB_598_U116 P3_IR_REG_2__SCAN_IN ; P3_SUB_598_U117
g23231 nand P3_SUB_598_U36 P3_IR_REG_29__SCAN_IN ; P3_SUB_598_U118
g23232 nand P3_SUB_598_U112 P3_SUB_598_U80 ; P3_SUB_598_U119
g23233 nand P3_SUB_598_U119 P3_IR_REG_26__SCAN_IN ; P3_SUB_598_U120
g23234 nand P3_SUB_598_U111 P3_IR_REG_24__SCAN_IN ; P3_SUB_598_U121
g23235 nand P3_SUB_598_U41 P3_IR_REG_23__SCAN_IN ; P3_SUB_598_U122
g23236 nand P3_SUB_598_U109 P3_SUB_598_U82 ; P3_SUB_598_U123
g23237 nand P3_SUB_598_U123 P3_IR_REG_22__SCAN_IN ; P3_SUB_598_U124
g23238 nand P3_SUB_598_U108 P3_IR_REG_20__SCAN_IN ; P3_SUB_598_U125
g23239 nand P3_SUB_598_U44 P3_IR_REG_19__SCAN_IN ; P3_SUB_598_U126
g23240 nand P3_SUB_598_U106 P3_SUB_598_U86 ; P3_SUB_598_U127
g23241 nand P3_SUB_598_U127 P3_IR_REG_18__SCAN_IN ; P3_SUB_598_U128
g23242 nand P3_SUB_598_U105 P3_IR_REG_16__SCAN_IN ; P3_SUB_598_U129
g23243 nand P3_SUB_598_U47 P3_IR_REG_15__SCAN_IN ; P3_SUB_598_U130
g23244 nand P3_SUB_598_U103 P3_SUB_598_U88 ; P3_SUB_598_U131
g23245 nand P3_SUB_598_U131 P3_IR_REG_14__SCAN_IN ; P3_SUB_598_U132
g23246 nand P3_SUB_598_U102 P3_IR_REG_12__SCAN_IN ; P3_SUB_598_U133
g23247 nand P3_SUB_598_U49 P3_IR_REG_11__SCAN_IN ; P3_SUB_598_U134
g23248 nand P3_SUB_598_U94 P3_SUB_598_U71 ; P3_SUB_598_U135
g23249 nand P3_SUB_598_U135 P3_IR_REG_10__SCAN_IN ; P3_SUB_598_U136
g23250 nand P3_SUB_598_U115 P3_SUB_598_U76 ; P3_SUB_598_U137
g23251 nand P3_IR_REG_27__SCAN_IN P3_IR_REG_28__SCAN_IN ; P3_SUB_598_U138
g23252 nand P3_SUB_598_U78 P3_IR_REG_28__SCAN_IN ; P3_SUB_598_U139
g23253 not P3_SUB_598_U28 ; P3_SUB_598_U140
g23254 nand P3_SUB_598_U29 P3_IR_REG_9__SCAN_IN ; P3_SUB_598_U141
g23255 nand P3_SUB_598_U94 P3_SUB_598_U71 ; P3_SUB_598_U142
g23256 nand P3_SUB_598_U30 P3_IR_REG_5__SCAN_IN ; P3_SUB_598_U143
g23257 nand P3_SUB_598_U91 P3_SUB_598_U73 ; P3_SUB_598_U144
g23258 nand P3_SUB_598_U137 P3_SUB_598_U75 ; P3_SUB_598_U145
g23259 nand P3_SUB_598_U115 P3_SUB_598_U76 P3_IR_REG_31__SCAN_IN ; P3_SUB_598_U146
g23260 nand P3_SUB_598_U37 P3_IR_REG_30__SCAN_IN ; P3_SUB_598_U147
g23261 nand P3_SUB_598_U115 P3_SUB_598_U76 ; P3_SUB_598_U148
g23262 nand P3_SUB_598_U78 P3_IR_REG_27__SCAN_IN ; P3_SUB_598_U149
g23263 nand P3_SUB_598_U113 P3_SUB_598_U39 ; P3_SUB_598_U150
g23264 nand P3_SUB_598_U35 P3_IR_REG_25__SCAN_IN ; P3_SUB_598_U151
g23265 nand P3_SUB_598_U112 P3_SUB_598_U80 ; P3_SUB_598_U152
g23266 nand P3_SUB_598_U40 P3_IR_REG_21__SCAN_IN ; P3_SUB_598_U153
g23267 nand P3_SUB_598_U109 P3_SUB_598_U82 ; P3_SUB_598_U154
g23268 nand P3_SUB_598_U85 P3_IR_REG_1__SCAN_IN ; P3_SUB_598_U155
g23269 nand P3_SUB_598_U84 P3_IR_REG_0__SCAN_IN ; P3_SUB_598_U156
g23270 nand P3_SUB_598_U34 P3_IR_REG_17__SCAN_IN ; P3_SUB_598_U157
g23271 nand P3_SUB_598_U106 P3_SUB_598_U86 ; P3_SUB_598_U158
g23272 nand P3_SUB_598_U46 P3_IR_REG_13__SCAN_IN ; P3_SUB_598_U159
g23273 nand P3_SUB_598_U103 P3_SUB_598_U88 ; P3_SUB_598_U160
g23274 and P3_R693_U113 P3_R693_U114 ; P3_R693_U6
g23275 and P3_R693_U115 P3_R693_U116 ; P3_R693_U7
g23276 and P3_R693_U80 P3_R693_U118 P3_R693_U120 P3_R693_U7 ; P3_R693_U8
g23277 and P3_R693_U126 P3_R693_U125 ; P3_R693_U9
g23278 and P3_R693_U130 P3_R693_U131 ; P3_R693_U10
g23279 and P3_R693_U84 P3_R693_U10 ; P3_R693_U11
g23280 and P3_R693_U142 P3_R693_U141 ; P3_R693_U12
g23281 and P3_R693_U178 P3_R693_U179 P3_R693_U177 ; P3_R693_U13
g23282 and P3_R693_U189 P3_R693_U188 P3_R693_U108 P3_R693_U109 ; P3_R693_U14
g23283 not P3_U3529 ; P3_R693_U15
g23284 not P3_U3537 ; P3_R693_U16
g23285 not P3_U3536 ; P3_R693_U17
g23286 not P3_U3905 ; P3_R693_U18
g23287 not P3_U3540 ; P3_R693_U19
g23288 not P3_U3906 ; P3_R693_U20
g23289 not P3_U3541 ; P3_R693_U21
g23290 not P3_U3543 ; P3_R693_U22
g23291 not P3_U3443 ; P3_R693_U23
g23292 not P3_U3544 ; P3_R693_U24
g23293 not P3_U3440 ; P3_R693_U25
g23294 not P3_U3445 ; P3_R693_U26
g23295 not P3_U3907 ; P3_R693_U27
g23296 not P3_U3545 ; P3_R693_U28
g23297 not P3_U3546 ; P3_R693_U29
g23298 not P3_U3437 ; P3_R693_U30
g23299 not P3_U3434 ; P3_R693_U31
g23300 not P3_U3526 ; P3_R693_U32
g23301 not P3_U3525 ; P3_R693_U33
g23302 not P3_U3404 ; P3_R693_U34
g23303 not P3_U3407 ; P3_R693_U35
g23304 not P3_U3416 ; P3_R693_U36
g23305 not P3_U3419 ; P3_R693_U37
g23306 not P3_U3410 ; P3_R693_U38
g23307 not P3_U3413 ; P3_R693_U39
g23308 not P3_U3398 ; P3_R693_U40
g23309 not P3_U3401 ; P3_R693_U41
g23310 not P3_U3553 ; P3_R693_U42
g23311 not P3_U3395 ; P3_R693_U43
g23312 not P3_U3392 ; P3_R693_U44
g23313 not P3_U3550 ; P3_R693_U45
g23314 not P3_U3549 ; P3_R693_U46
g23315 not P3_U3542 ; P3_R693_U47
g23316 not P3_U3531 ; P3_R693_U48
g23317 not P3_U3528 ; P3_R693_U49
g23318 not P3_U3527 ; P3_R693_U50
g23319 not P3_U3523 ; P3_R693_U51
g23320 not P3_U3524 ; P3_R693_U52
g23321 not P3_U3552 ; P3_R693_U53
g23322 not P3_U3551 ; P3_R693_U54
g23323 not P3_U3425 ; P3_R693_U55
g23324 not P3_U3422 ; P3_R693_U56
g23325 not P3_U3431 ; P3_R693_U57
g23326 not P3_U3428 ; P3_R693_U58
g23327 not P3_U3548 ; P3_R693_U59
g23328 not P3_U3547 ; P3_R693_U60
g23329 not P3_U3539 ; P3_R693_U61
g23330 not P3_U3538 ; P3_R693_U62
g23331 not P3_U3908 ; P3_R693_U63
g23332 not P3_U3900 ; P3_R693_U64
g23333 not P3_U3899 ; P3_R693_U65
g23334 not P3_U3904 ; P3_R693_U66
g23335 not P3_U3903 ; P3_R693_U67
g23336 not P3_U3902 ; P3_R693_U68
g23337 not P3_U3901 ; P3_R693_U69
g23338 not P3_U3533 ; P3_R693_U70
g23339 not P3_U3534 ; P3_R693_U71
g23340 not P3_U3872 ; P3_R693_U72
g23341 not P3_U3532 ; P3_R693_U73
g23342 not P3_U3535 ; P3_R693_U74
g23343 and P3_U3540 P3_R693_U20 ; P3_R693_U75
g23344 and P3_U3541 P3_R693_U27 ; P3_R693_U76
g23345 and P3_R693_U168 P3_R693_U167 ; P3_R693_U77
g23346 and P3_U3443 P3_R693_U24 ; P3_R693_U78
g23347 and P3_U3440 P3_R693_U28 ; P3_R693_U79
g23348 and P3_R693_U119 P3_R693_U117 ; P3_R693_U80
g23349 and P3_U3404 P3_R693_U50 ; P3_R693_U81
g23350 and P3_U3407 P3_R693_U32 ; P3_R693_U82
g23351 and P3_U3387 P3_R693_U111 ; P3_R693_U83
g23352 and P3_R693_U133 P3_R693_U132 ; P3_R693_U84
g23353 and P3_R693_U129 P3_R693_U86 ; P3_R693_U85
g23354 and P3_R693_U135 P3_R693_U134 ; P3_R693_U86
g23355 and P3_R693_U138 P3_R693_U137 ; P3_R693_U87
g23356 and P3_R693_U135 P3_R693_U134 ; P3_R693_U88
g23357 and P3_R693_U9 P3_R693_U148 ; P3_R693_U89
g23358 and P3_R693_U129 P3_R693_U127 P3_R693_U11 ; P3_R693_U90
g23359 and P3_U3523 P3_R693_U36 ; P3_R693_U91
g23360 and P3_U3524 P3_R693_U39 ; P3_R693_U92
g23361 and P3_R693_U152 P3_R693_U151 P3_R693_U95 ; P3_R693_U93
g23362 and P3_R693_U154 P3_R693_U153 ; P3_R693_U94
g23363 and P3_R693_U94 P3_R693_U12 ; P3_R693_U95
g23364 and P3_U3425 P3_R693_U45 ; P3_R693_U96
g23365 and P3_U3422 P3_R693_U54 ; P3_R693_U97
g23366 and P3_R693_U157 P3_R693_U100 ; P3_R693_U98
g23367 and P3_R693_U98 P3_R693_U158 ; P3_R693_U99
g23368 and P3_R693_U160 P3_R693_U159 ; P3_R693_U100
g23369 and P3_R693_U171 P3_R693_U170 P3_R693_U122 P3_R693_U123 ; P3_R693_U101
g23370 and P3_R693_U175 P3_R693_U174 ; P3_R693_U102
g23371 and P3_R693_U187 P3_R693_U186 ; P3_R693_U103
g23372 and P3_R693_U103 P3_R693_U13 ; P3_R693_U104
g23373 and P3_R693_U106 P3_R693_U190 ; P3_R693_U105
g23374 and P3_U3533 P3_R693_U65 ; P3_R693_U106
g23375 and P3_U3532 P3_R693_U63 ; P3_R693_U107
g23376 and P3_R693_U192 P3_R693_U191 ; P3_R693_U108
g23377 and P3_R693_U194 P3_R693_U193 P3_R693_U195 ; P3_R693_U109
g23378 not P3_U3873 ; P3_R693_U110
g23379 not P3_U3554 ; P3_R693_U111
g23380 nand P3_R693_U181 P3_R693_U196 ; P3_R693_U112
g23381 nand P3_U3543 P3_R693_U26 ; P3_R693_U113
g23382 nand P3_U3544 P3_R693_U23 ; P3_R693_U114
g23383 nand P3_U3905 P3_R693_U61 ; P3_R693_U115
g23384 nand P3_U3906 P3_R693_U19 ; P3_R693_U116
g23385 nand P3_R693_U78 P3_R693_U113 ; P3_R693_U117
g23386 nand P3_R693_U79 P3_R693_U6 ; P3_R693_U118
g23387 nand P3_U3445 P3_R693_U22 ; P3_R693_U119
g23388 nand P3_U3907 P3_R693_U21 ; P3_R693_U120
g23389 nand P3_U3437 P3_R693_U29 ; P3_R693_U121
g23390 nand P3_U3537 P3_R693_U67 ; P3_R693_U122
g23391 nand P3_U3536 P3_R693_U68 ; P3_R693_U123
g23392 nand P3_U3434 P3_R693_U60 ; P3_R693_U124
g23393 nand P3_U3526 P3_R693_U35 ; P3_R693_U125
g23394 nand P3_U3525 P3_R693_U38 ; P3_R693_U126
g23395 nand P3_R693_U81 P3_R693_U9 ; P3_R693_U127
g23396 nand P3_U3525 P3_R693_U38 ; P3_R693_U128
g23397 nand P3_R693_U82 P3_R693_U128 ; P3_R693_U129
g23398 nand P3_U3419 P3_R693_U53 ; P3_R693_U130
g23399 nand P3_U3416 P3_R693_U51 ; P3_R693_U131
g23400 nand P3_U3410 P3_R693_U33 ; P3_R693_U132
g23401 nand P3_U3413 P3_R693_U52 ; P3_R693_U133
g23402 nand P3_U3398 P3_R693_U48 ; P3_R693_U134
g23403 nand P3_U3401 P3_R693_U49 ; P3_R693_U135
g23404 nand P3_U3553 P3_R693_U44 ; P3_R693_U136
g23405 nand P3_R693_U83 P3_R693_U136 ; P3_R693_U137
g23406 nand P3_U3395 P3_R693_U47 ; P3_R693_U138
g23407 nand P3_U3392 P3_R693_U42 ; P3_R693_U139
g23408 nand P3_R693_U11 P3_R693_U139 P3_R693_U87 P3_R693_U127 P3_R693_U85 ; P3_R693_U140
g23409 nand P3_U3550 P3_R693_U55 ; P3_R693_U141
g23410 nand P3_U3549 P3_R693_U58 ; P3_R693_U142
g23411 nand P3_U3542 P3_R693_U43 ; P3_R693_U143
g23412 nand P3_U3531 P3_R693_U40 ; P3_R693_U144
g23413 nand P3_R693_U144 P3_R693_U143 ; P3_R693_U145
g23414 nand P3_R693_U88 P3_R693_U145 ; P3_R693_U146
g23415 nand P3_U3528 P3_R693_U41 ; P3_R693_U147
g23416 nand P3_U3527 P3_R693_U34 ; P3_R693_U148
g23417 nand P3_R693_U147 P3_R693_U146 P3_R693_U89 ; P3_R693_U149
g23418 nand P3_R693_U90 P3_R693_U149 ; P3_R693_U150
g23419 nand P3_R693_U91 P3_R693_U130 ; P3_R693_U151
g23420 nand P3_R693_U92 P3_R693_U10 ; P3_R693_U152
g23421 nand P3_U3552 P3_R693_U37 ; P3_R693_U153
g23422 nand P3_U3551 P3_R693_U56 ; P3_R693_U154
g23423 nand P3_R693_U150 P3_R693_U140 P3_R693_U93 ; P3_R693_U155
g23424 nand P3_U3549 P3_R693_U58 ; P3_R693_U156
g23425 nand P3_R693_U96 P3_R693_U156 ; P3_R693_U157
g23426 nand P3_R693_U97 P3_R693_U12 ; P3_R693_U158
g23427 nand P3_U3431 P3_R693_U59 ; P3_R693_U159
g23428 nand P3_U3428 P3_R693_U46 ; P3_R693_U160
g23429 nand P3_R693_U155 P3_R693_U99 ; P3_R693_U161
g23430 nand P3_U3548 P3_R693_U57 ; P3_R693_U162
g23431 nand P3_R693_U162 P3_R693_U161 ; P3_R693_U163
g23432 nand P3_R693_U163 P3_R693_U124 ; P3_R693_U164
g23433 nand P3_U3547 P3_R693_U31 ; P3_R693_U165
g23434 nand P3_R693_U165 P3_R693_U164 ; P3_R693_U166
g23435 nand P3_U3545 P3_R693_U25 ; P3_R693_U167
g23436 nand P3_U3546 P3_R693_U30 ; P3_R693_U168
g23437 nand P3_R693_U77 P3_R693_U6 ; P3_R693_U169
g23438 nand P3_R693_U75 P3_R693_U115 ; P3_R693_U170
g23439 nand P3_R693_U76 P3_R693_U7 ; P3_R693_U171
g23440 nand P3_R693_U8 P3_R693_U169 ; P3_R693_U172
g23441 nand P3_R693_U166 P3_R693_U121 P3_R693_U8 ; P3_R693_U173
g23442 nand P3_U3539 P3_R693_U18 ; P3_R693_U174
g23443 nand P3_U3538 P3_R693_U66 ; P3_R693_U175
g23444 nand P3_R693_U173 P3_R693_U172 P3_R693_U102 P3_R693_U101 ; P3_R693_U176
g23445 nand P3_U3908 P3_R693_U73 ; P3_R693_U177
g23446 nand P3_U3900 P3_R693_U71 ; P3_R693_U178
g23447 nand P3_U3899 P3_R693_U70 ; P3_R693_U179
g23448 nand P3_U3529 P3_R693_U72 ; P3_R693_U180
g23449 nand P3_R693_U180 P3_R693_U110 ; P3_R693_U181
g23450 nand P3_U3904 P3_R693_U62 ; P3_R693_U182
g23451 nand P3_U3903 P3_R693_U16 ; P3_R693_U183
g23452 nand P3_R693_U183 P3_R693_U182 ; P3_R693_U184
g23453 nand P3_R693_U184 P3_R693_U122 P3_R693_U123 ; P3_R693_U185
g23454 nand P3_U3902 P3_R693_U17 ; P3_R693_U186
g23455 nand P3_U3901 P3_R693_U74 ; P3_R693_U187
g23456 nand P3_R693_U176 P3_R693_U185 P3_R693_U112 P3_R693_U104 ; P3_R693_U188
g23457 nand P3_R693_U180 P3_U3530 P3_R693_U110 ; P3_R693_U189
g23458 nand P3_U3908 P3_R693_U73 ; P3_R693_U190
g23459 nand P3_R693_U112 P3_R693_U105 ; P3_R693_U191
g23460 nand P3_U3534 P3_R693_U13 P3_R693_U112 P3_R693_U64 ; P3_R693_U192
g23461 nand P3_U3872 P3_R693_U15 ; P3_R693_U193
g23462 nand P3_R693_U107 P3_R693_U112 ; P3_R693_U194
g23463 nand P3_U3535 P3_R693_U13 P3_R693_U112 P3_R693_U69 ; P3_R693_U195
g23464 nand P3_U3530 P3_R693_U180 ; P3_R693_U196
g23465 nand P3_SUB_609_U40 P3_SUB_609_U98 ; P3_SUB_609_U6
g23466 nand P3_SUB_609_U79 P3_SUB_609_U105 ; P3_SUB_609_U7
g23467 nand P3_SUB_609_U65 P3_SUB_609_U113 ; P3_SUB_609_U8
g23468 nand P3_SUB_609_U34 P3_SUB_609_U110 ; P3_SUB_609_U9
g23469 nand P3_SUB_609_U87 P3_SUB_609_U97 ; P3_SUB_609_U10
g23470 nand P3_SUB_609_U81 P3_SUB_609_U103 ; P3_SUB_609_U11
g23471 nand P3_SUB_609_U67 P3_SUB_609_U70 ; P3_SUB_609_U12
g23472 nand P3_SUB_609_U73 P3_SUB_609_U111 ; P3_SUB_609_U13
g23473 nand P3_SUB_609_U33 P3_SUB_609_U69 ; P3_SUB_609_U14
g23474 nand P3_SUB_609_U38 P3_SUB_609_U102 ; P3_SUB_609_U15
g23475 nand P3_SUB_609_U41 P3_SUB_609_U96 ; P3_SUB_609_U16
g23476 nand P3_SUB_609_U85 P3_SUB_609_U99 ; P3_SUB_609_U17
g23477 nand P3_SUB_609_U31 P3_SUB_609_U71 ; P3_SUB_609_U18
g23478 nand P3_SUB_609_U37 P3_SUB_609_U104 ; P3_SUB_609_U19
g23479 nand P3_SUB_609_U83 P3_SUB_609_U101 ; P3_SUB_609_U20
g23480 nand P3_SUB_609_U36 P3_SUB_609_U106 ; P3_SUB_609_U21
g23481 nand P3_SUB_609_U42 P3_SUB_609_U94 ; P3_SUB_609_U22
g23482 nand P3_SUB_609_U75 P3_SUB_609_U109 ; P3_SUB_609_U23
g23483 nand P3_SUB_609_U35 P3_SUB_609_U108 ; P3_SUB_609_U24
g23484 not P3_REG3_REG_3__SCAN_IN ; P3_SUB_609_U25
g23485 nand P3_SUB_609_U89 P3_SUB_609_U95 ; P3_SUB_609_U26
g23486 nand P3_SUB_609_U39 P3_SUB_609_U100 ; P3_SUB_609_U27
g23487 nand P3_SUB_609_U91 P3_SUB_609_U93 ; P3_SUB_609_U28
g23488 nand P3_SUB_609_U64 P3_SUB_609_U72 ; P3_SUB_609_U29
g23489 nand P3_SUB_609_U77 P3_SUB_609_U107 ; P3_SUB_609_U30
g23490 or P3_REG3_REG_6__SCAN_IN P3_REG3_REG_4__SCAN_IN P3_REG3_REG_5__SCAN_IN P3_REG3_REG_3__SCAN_IN P3_REG3_REG_7__SCAN_IN ; P3_SUB_609_U31
g23491 not P3_REG3_REG_8__SCAN_IN ; P3_SUB_609_U32
g23492 nand P3_SUB_609_U54 P3_SUB_609_U66 ; P3_SUB_609_U33
g23493 nand P3_SUB_609_U55 P3_SUB_609_U68 ; P3_SUB_609_U34
g23494 nand P3_SUB_609_U56 P3_SUB_609_U74 ; P3_SUB_609_U35
g23495 nand P3_SUB_609_U57 P3_SUB_609_U76 ; P3_SUB_609_U36
g23496 nand P3_SUB_609_U58 P3_SUB_609_U78 ; P3_SUB_609_U37
g23497 nand P3_SUB_609_U59 P3_SUB_609_U80 ; P3_SUB_609_U38
g23498 nand P3_SUB_609_U60 P3_SUB_609_U82 ; P3_SUB_609_U39
g23499 nand P3_SUB_609_U61 P3_SUB_609_U84 ; P3_SUB_609_U40
g23500 nand P3_SUB_609_U62 P3_SUB_609_U86 ; P3_SUB_609_U41
g23501 nand P3_SUB_609_U63 P3_SUB_609_U88 ; P3_SUB_609_U42
g23502 not P3_REG3_REG_28__SCAN_IN ; P3_SUB_609_U43
g23503 not P3_REG3_REG_26__SCAN_IN ; P3_SUB_609_U44
g23504 not P3_REG3_REG_24__SCAN_IN ; P3_SUB_609_U45
g23505 not P3_REG3_REG_22__SCAN_IN ; P3_SUB_609_U46
g23506 not P3_REG3_REG_20__SCAN_IN ; P3_SUB_609_U47
g23507 not P3_REG3_REG_18__SCAN_IN ; P3_SUB_609_U48
g23508 not P3_REG3_REG_16__SCAN_IN ; P3_SUB_609_U49
g23509 not P3_REG3_REG_14__SCAN_IN ; P3_SUB_609_U50
g23510 not P3_REG3_REG_12__SCAN_IN ; P3_SUB_609_U51
g23511 not P3_REG3_REG_10__SCAN_IN ; P3_SUB_609_U52
g23512 nand P3_SUB_609_U115 P3_SUB_609_U114 ; P3_SUB_609_U53
g23513 nor P3_REG3_REG_9__SCAN_IN P3_REG3_REG_8__SCAN_IN ; P3_SUB_609_U54
g23514 nor P3_REG3_REG_11__SCAN_IN P3_REG3_REG_10__SCAN_IN ; P3_SUB_609_U55
g23515 nor P3_REG3_REG_13__SCAN_IN P3_REG3_REG_12__SCAN_IN ; P3_SUB_609_U56
g23516 nor P3_REG3_REG_15__SCAN_IN P3_REG3_REG_14__SCAN_IN ; P3_SUB_609_U57
g23517 nor P3_REG3_REG_17__SCAN_IN P3_REG3_REG_16__SCAN_IN ; P3_SUB_609_U58
g23518 nor P3_REG3_REG_18__SCAN_IN P3_REG3_REG_19__SCAN_IN ; P3_SUB_609_U59
g23519 nor P3_REG3_REG_20__SCAN_IN P3_REG3_REG_21__SCAN_IN ; P3_SUB_609_U60
g23520 nor P3_REG3_REG_22__SCAN_IN P3_REG3_REG_23__SCAN_IN ; P3_SUB_609_U61
g23521 nor P3_REG3_REG_24__SCAN_IN P3_REG3_REG_25__SCAN_IN ; P3_SUB_609_U62
g23522 nor P3_REG3_REG_26__SCAN_IN P3_REG3_REG_27__SCAN_IN ; P3_SUB_609_U63
g23523 or P3_REG3_REG_4__SCAN_IN P3_REG3_REG_3__SCAN_IN ; P3_SUB_609_U64
g23524 or P3_REG3_REG_6__SCAN_IN P3_REG3_REG_4__SCAN_IN P3_REG3_REG_5__SCAN_IN P3_REG3_REG_3__SCAN_IN ; P3_SUB_609_U65
g23525 not P3_SUB_609_U31 ; P3_SUB_609_U66
g23526 nand P3_SUB_609_U66 P3_SUB_609_U32 ; P3_SUB_609_U67
g23527 not P3_SUB_609_U33 ; P3_SUB_609_U68
g23528 nand P3_SUB_609_U67 P3_REG3_REG_9__SCAN_IN ; P3_SUB_609_U69
g23529 nand P3_SUB_609_U31 P3_REG3_REG_8__SCAN_IN ; P3_SUB_609_U70
g23530 nand P3_SUB_609_U65 P3_REG3_REG_7__SCAN_IN ; P3_SUB_609_U71
g23531 nand P3_REG3_REG_4__SCAN_IN P3_REG3_REG_3__SCAN_IN ; P3_SUB_609_U72
g23532 nand P3_SUB_609_U68 P3_SUB_609_U52 ; P3_SUB_609_U73
g23533 not P3_SUB_609_U34 ; P3_SUB_609_U74
g23534 nand P3_SUB_609_U74 P3_SUB_609_U51 ; P3_SUB_609_U75
g23535 not P3_SUB_609_U35 ; P3_SUB_609_U76
g23536 nand P3_SUB_609_U76 P3_SUB_609_U50 ; P3_SUB_609_U77
g23537 not P3_SUB_609_U36 ; P3_SUB_609_U78
g23538 nand P3_SUB_609_U78 P3_SUB_609_U49 ; P3_SUB_609_U79
g23539 not P3_SUB_609_U37 ; P3_SUB_609_U80
g23540 nand P3_SUB_609_U80 P3_SUB_609_U48 ; P3_SUB_609_U81
g23541 not P3_SUB_609_U38 ; P3_SUB_609_U82
g23542 nand P3_SUB_609_U82 P3_SUB_609_U47 ; P3_SUB_609_U83
g23543 not P3_SUB_609_U39 ; P3_SUB_609_U84
g23544 nand P3_SUB_609_U84 P3_SUB_609_U46 ; P3_SUB_609_U85
g23545 not P3_SUB_609_U40 ; P3_SUB_609_U86
g23546 nand P3_SUB_609_U86 P3_SUB_609_U45 ; P3_SUB_609_U87
g23547 not P3_SUB_609_U41 ; P3_SUB_609_U88
g23548 nand P3_SUB_609_U88 P3_SUB_609_U44 ; P3_SUB_609_U89
g23549 not P3_SUB_609_U42 ; P3_SUB_609_U90
g23550 nand P3_SUB_609_U90 P3_SUB_609_U43 ; P3_SUB_609_U91
g23551 not P3_SUB_609_U91 ; P3_SUB_609_U92
g23552 nand P3_SUB_609_U42 P3_REG3_REG_28__SCAN_IN ; P3_SUB_609_U93
g23553 nand P3_SUB_609_U89 P3_REG3_REG_27__SCAN_IN ; P3_SUB_609_U94
g23554 nand P3_SUB_609_U41 P3_REG3_REG_26__SCAN_IN ; P3_SUB_609_U95
g23555 nand P3_SUB_609_U87 P3_REG3_REG_25__SCAN_IN ; P3_SUB_609_U96
g23556 nand P3_SUB_609_U40 P3_REG3_REG_24__SCAN_IN ; P3_SUB_609_U97
g23557 nand P3_SUB_609_U85 P3_REG3_REG_23__SCAN_IN ; P3_SUB_609_U98
g23558 nand P3_SUB_609_U39 P3_REG3_REG_22__SCAN_IN ; P3_SUB_609_U99
g23559 nand P3_SUB_609_U83 P3_REG3_REG_21__SCAN_IN ; P3_SUB_609_U100
g23560 nand P3_SUB_609_U38 P3_REG3_REG_20__SCAN_IN ; P3_SUB_609_U101
g23561 nand P3_SUB_609_U81 P3_REG3_REG_19__SCAN_IN ; P3_SUB_609_U102
g23562 nand P3_SUB_609_U37 P3_REG3_REG_18__SCAN_IN ; P3_SUB_609_U103
g23563 nand P3_SUB_609_U79 P3_REG3_REG_17__SCAN_IN ; P3_SUB_609_U104
g23564 nand P3_SUB_609_U36 P3_REG3_REG_16__SCAN_IN ; P3_SUB_609_U105
g23565 nand P3_SUB_609_U77 P3_REG3_REG_15__SCAN_IN ; P3_SUB_609_U106
g23566 nand P3_SUB_609_U35 P3_REG3_REG_14__SCAN_IN ; P3_SUB_609_U107
g23567 nand P3_SUB_609_U75 P3_REG3_REG_13__SCAN_IN ; P3_SUB_609_U108
g23568 nand P3_SUB_609_U34 P3_REG3_REG_12__SCAN_IN ; P3_SUB_609_U109
g23569 nand P3_SUB_609_U73 P3_REG3_REG_11__SCAN_IN ; P3_SUB_609_U110
g23570 nand P3_SUB_609_U33 P3_REG3_REG_10__SCAN_IN ; P3_SUB_609_U111
g23571 or P3_REG3_REG_4__SCAN_IN P3_REG3_REG_5__SCAN_IN P3_REG3_REG_3__SCAN_IN ; P3_SUB_609_U112
g23572 nand P3_SUB_609_U112 P3_REG3_REG_6__SCAN_IN ; P3_SUB_609_U113
g23573 nand P3_SUB_609_U64 P3_REG3_REG_5__SCAN_IN ; P3_SUB_609_U114
g23574 or P3_REG3_REG_4__SCAN_IN P3_REG3_REG_5__SCAN_IN P3_REG3_REG_3__SCAN_IN ; P3_SUB_609_U115
g23575 and P3_R1095_U210 P3_R1095_U209 ; P3_R1095_U6
g23576 and P3_R1095_U189 P3_R1095_U245 ; P3_R1095_U7
g23577 and P3_R1095_U247 P3_R1095_U246 ; P3_R1095_U8
g23578 and P3_R1095_U190 P3_R1095_U262 ; P3_R1095_U9
g23579 and P3_R1095_U264 P3_R1095_U263 ; P3_R1095_U10
g23580 and P3_R1095_U191 P3_R1095_U286 ; P3_R1095_U11
g23581 and P3_R1095_U288 P3_R1095_U287 ; P3_R1095_U12
g23582 and P3_R1095_U208 P3_R1095_U194 P3_R1095_U213 ; P3_R1095_U13
g23583 and P3_R1095_U218 P3_R1095_U195 ; P3_R1095_U14
g23584 and P3_R1095_U392 P3_R1095_U391 ; P3_R1095_U15
g23585 nand P3_R1095_U342 P3_R1095_U345 ; P3_R1095_U16
g23586 nand P3_R1095_U331 P3_R1095_U334 ; P3_R1095_U17
g23587 nand P3_R1095_U320 P3_R1095_U323 ; P3_R1095_U18
g23588 nand P3_R1095_U312 P3_R1095_U314 ; P3_R1095_U19
g23589 nand P3_R1095_U162 P3_R1095_U183 P3_R1095_U351 ; P3_R1095_U20
g23590 nand P3_R1095_U241 P3_R1095_U243 ; P3_R1095_U21
g23591 nand P3_R1095_U233 P3_R1095_U236 ; P3_R1095_U22
g23592 nand P3_R1095_U225 P3_R1095_U227 ; P3_R1095_U23
g23593 nand P3_R1095_U172 P3_R1095_U348 ; P3_R1095_U24
g23594 not P3_U3069 ; P3_R1095_U25
g23595 nand P3_U3069 P3_R1095_U39 ; P3_R1095_U26
g23596 not P3_U3083 ; P3_R1095_U27
g23597 not P3_U3413 ; P3_R1095_U28
g23598 not P3_U3395 ; P3_R1095_U29
g23599 not P3_U3387 ; P3_R1095_U30
g23600 not P3_U3077 ; P3_R1095_U31
g23601 not P3_U3398 ; P3_R1095_U32
g23602 not P3_U3067 ; P3_R1095_U33
g23603 nand P3_U3067 P3_R1095_U29 ; P3_R1095_U34
g23604 not P3_U3063 ; P3_R1095_U35
g23605 not P3_U3404 ; P3_R1095_U36
g23606 not P3_U3407 ; P3_R1095_U37
g23607 not P3_U3401 ; P3_R1095_U38
g23608 not P3_U3410 ; P3_R1095_U39
g23609 not P3_U3070 ; P3_R1095_U40
g23610 not P3_U3066 ; P3_R1095_U41
g23611 not P3_U3059 ; P3_R1095_U42
g23612 nand P3_U3059 P3_R1095_U38 ; P3_R1095_U43
g23613 nand P3_R1095_U214 P3_R1095_U212 ; P3_R1095_U44
g23614 not P3_U3416 ; P3_R1095_U45
g23615 not P3_U3082 ; P3_R1095_U46
g23616 nand P3_R1095_U44 P3_R1095_U215 ; P3_R1095_U47
g23617 nand P3_R1095_U43 P3_R1095_U229 ; P3_R1095_U48
g23618 nand P3_R1095_U201 P3_R1095_U185 P3_R1095_U349 ; P3_R1095_U49
g23619 not P3_U3901 ; P3_R1095_U50
g23620 not P3_U3422 ; P3_R1095_U51
g23621 not P3_U3419 ; P3_R1095_U52
g23622 not P3_U3062 ; P3_R1095_U53
g23623 not P3_U3061 ; P3_R1095_U54
g23624 nand P3_U3082 P3_R1095_U45 ; P3_R1095_U55
g23625 not P3_U3425 ; P3_R1095_U56
g23626 not P3_U3071 ; P3_R1095_U57
g23627 not P3_U3428 ; P3_R1095_U58
g23628 not P3_U3079 ; P3_R1095_U59
g23629 not P3_U3437 ; P3_R1095_U60
g23630 not P3_U3434 ; P3_R1095_U61
g23631 not P3_U3431 ; P3_R1095_U62
g23632 not P3_U3072 ; P3_R1095_U63
g23633 not P3_U3073 ; P3_R1095_U64
g23634 not P3_U3078 ; P3_R1095_U65
g23635 nand P3_U3078 P3_R1095_U62 ; P3_R1095_U66
g23636 not P3_U3440 ; P3_R1095_U67
g23637 not P3_U3068 ; P3_R1095_U68
g23638 not P3_U3081 ; P3_R1095_U69
g23639 not P3_U3445 ; P3_R1095_U70
g23640 not P3_U3080 ; P3_R1095_U71
g23641 not P3_U3907 ; P3_R1095_U72
g23642 not P3_U3075 ; P3_R1095_U73
g23643 not P3_U3904 ; P3_R1095_U74
g23644 not P3_U3905 ; P3_R1095_U75
g23645 not P3_U3906 ; P3_R1095_U76
g23646 not P3_U3065 ; P3_R1095_U77
g23647 not P3_U3060 ; P3_R1095_U78
g23648 not P3_U3074 ; P3_R1095_U79
g23649 nand P3_U3074 P3_R1095_U76 ; P3_R1095_U80
g23650 not P3_U3903 ; P3_R1095_U81
g23651 not P3_U3064 ; P3_R1095_U82
g23652 not P3_U3902 ; P3_R1095_U83
g23653 not P3_U3057 ; P3_R1095_U84
g23654 not P3_U3900 ; P3_R1095_U85
g23655 not P3_U3056 ; P3_R1095_U86
g23656 nand P3_U3056 P3_R1095_U50 ; P3_R1095_U87
g23657 not P3_U3052 ; P3_R1095_U88
g23658 not P3_U3899 ; P3_R1095_U89
g23659 not P3_U3053 ; P3_R1095_U90
g23660 nand P3_R1095_U302 P3_R1095_U301 ; P3_R1095_U91
g23661 nand P3_R1095_U80 P3_R1095_U316 ; P3_R1095_U92
g23662 nand P3_R1095_U66 P3_R1095_U327 ; P3_R1095_U93
g23663 nand P3_R1095_U55 P3_R1095_U338 ; P3_R1095_U94
g23664 not P3_U3076 ; P3_R1095_U95
g23665 nand P3_R1095_U402 P3_R1095_U401 ; P3_R1095_U96
g23666 nand P3_R1095_U416 P3_R1095_U415 ; P3_R1095_U97
g23667 nand P3_R1095_U421 P3_R1095_U420 ; P3_R1095_U98
g23668 nand P3_R1095_U437 P3_R1095_U436 ; P3_R1095_U99
g23669 nand P3_R1095_U442 P3_R1095_U441 ; P3_R1095_U100
g23670 nand P3_R1095_U447 P3_R1095_U446 ; P3_R1095_U101
g23671 nand P3_R1095_U452 P3_R1095_U451 ; P3_R1095_U102
g23672 nand P3_R1095_U457 P3_R1095_U456 ; P3_R1095_U103
g23673 nand P3_R1095_U473 P3_R1095_U472 ; P3_R1095_U104
g23674 nand P3_R1095_U478 P3_R1095_U477 ; P3_R1095_U105
g23675 nand P3_R1095_U361 P3_R1095_U360 ; P3_R1095_U106
g23676 nand P3_R1095_U370 P3_R1095_U369 ; P3_R1095_U107
g23677 nand P3_R1095_U377 P3_R1095_U376 ; P3_R1095_U108
g23678 nand P3_R1095_U381 P3_R1095_U380 ; P3_R1095_U109
g23679 nand P3_R1095_U390 P3_R1095_U389 ; P3_R1095_U110
g23680 nand P3_R1095_U411 P3_R1095_U410 ; P3_R1095_U111
g23681 nand P3_R1095_U428 P3_R1095_U427 ; P3_R1095_U112
g23682 nand P3_R1095_U432 P3_R1095_U431 ; P3_R1095_U113
g23683 nand P3_R1095_U464 P3_R1095_U463 ; P3_R1095_U114
g23684 nand P3_R1095_U468 P3_R1095_U467 ; P3_R1095_U115
g23685 nand P3_R1095_U485 P3_R1095_U484 ; P3_R1095_U116
g23686 and P3_R1095_U352 P3_R1095_U193 ; P3_R1095_U117
g23687 and P3_R1095_U205 P3_R1095_U206 ; P3_R1095_U118
g23688 and P3_R1095_U14 P3_R1095_U13 ; P3_R1095_U119
g23689 and P3_R1095_U357 P3_R1095_U354 ; P3_R1095_U120
g23690 and P3_R1095_U363 P3_R1095_U362 P3_R1095_U26 ; P3_R1095_U121
g23691 and P3_R1095_U366 P3_R1095_U195 ; P3_R1095_U122
g23692 and P3_R1095_U235 P3_R1095_U6 ; P3_R1095_U123
g23693 and P3_R1095_U373 P3_R1095_U194 ; P3_R1095_U124
g23694 and P3_R1095_U383 P3_R1095_U382 P3_R1095_U34 ; P3_R1095_U125
g23695 and P3_R1095_U386 P3_R1095_U193 ; P3_R1095_U126
g23696 and P3_R1095_U222 P3_R1095_U7 ; P3_R1095_U127
g23697 and P3_R1095_U267 P3_R1095_U9 ; P3_R1095_U128
g23698 and P3_R1095_U291 P3_R1095_U11 ; P3_R1095_U129
g23699 and P3_R1095_U355 P3_R1095_U192 ; P3_R1095_U130
g23700 and P3_R1095_U306 P3_R1095_U307 ; P3_R1095_U131
g23701 and P3_R1095_U309 P3_R1095_U395 ; P3_R1095_U132
g23702 and P3_R1095_U306 P3_R1095_U307 ; P3_R1095_U133
g23703 and P3_R1095_U15 P3_R1095_U310 ; P3_R1095_U134
g23704 nand P3_R1095_U399 P3_R1095_U398 ; P3_R1095_U135
g23705 and P3_R1095_U404 P3_R1095_U403 P3_R1095_U87 ; P3_R1095_U136
g23706 and P3_R1095_U407 P3_R1095_U192 ; P3_R1095_U137
g23707 nand P3_R1095_U413 P3_R1095_U412 ; P3_R1095_U138
g23708 nand P3_R1095_U418 P3_R1095_U417 ; P3_R1095_U139
g23709 and P3_R1095_U322 P3_R1095_U12 ; P3_R1095_U140
g23710 and P3_R1095_U424 P3_R1095_U191 ; P3_R1095_U141
g23711 nand P3_R1095_U434 P3_R1095_U433 ; P3_R1095_U142
g23712 nand P3_R1095_U439 P3_R1095_U438 ; P3_R1095_U143
g23713 nand P3_R1095_U444 P3_R1095_U443 ; P3_R1095_U144
g23714 nand P3_R1095_U449 P3_R1095_U448 ; P3_R1095_U145
g23715 nand P3_R1095_U454 P3_R1095_U453 ; P3_R1095_U146
g23716 and P3_R1095_U333 P3_R1095_U10 ; P3_R1095_U147
g23717 and P3_R1095_U460 P3_R1095_U190 ; P3_R1095_U148
g23718 nand P3_R1095_U470 P3_R1095_U469 ; P3_R1095_U149
g23719 nand P3_R1095_U475 P3_R1095_U474 ; P3_R1095_U150
g23720 and P3_R1095_U344 P3_R1095_U8 ; P3_R1095_U151
g23721 and P3_R1095_U481 P3_R1095_U189 ; P3_R1095_U152
g23722 and P3_R1095_U359 P3_R1095_U358 ; P3_R1095_U153
g23723 nand P3_R1095_U120 P3_R1095_U356 ; P3_R1095_U154
g23724 and P3_R1095_U368 P3_R1095_U367 ; P3_R1095_U155
g23725 and P3_R1095_U375 P3_R1095_U374 ; P3_R1095_U156
g23726 and P3_R1095_U379 P3_R1095_U378 ; P3_R1095_U157
g23727 nand P3_R1095_U118 P3_R1095_U203 ; P3_R1095_U158
g23728 and P3_R1095_U388 P3_R1095_U387 ; P3_R1095_U159
g23729 not P3_U3908 ; P3_R1095_U160
g23730 not P3_U3054 ; P3_R1095_U161
g23731 and P3_R1095_U397 P3_R1095_U396 ; P3_R1095_U162
g23732 nand P3_R1095_U131 P3_R1095_U304 ; P3_R1095_U163
g23733 and P3_R1095_U409 P3_R1095_U408 ; P3_R1095_U164
g23734 nand P3_R1095_U298 P3_R1095_U297 ; P3_R1095_U165
g23735 nand P3_R1095_U294 P3_R1095_U293 ; P3_R1095_U166
g23736 and P3_R1095_U426 P3_R1095_U425 ; P3_R1095_U167
g23737 and P3_R1095_U430 P3_R1095_U429 ; P3_R1095_U168
g23738 nand P3_R1095_U284 P3_R1095_U283 ; P3_R1095_U169
g23739 nand P3_R1095_U280 P3_R1095_U279 ; P3_R1095_U170
g23740 not P3_U3392 ; P3_R1095_U171
g23741 nand P3_U3387 P3_R1095_U95 ; P3_R1095_U172
g23742 nand P3_R1095_U276 P3_R1095_U184 P3_R1095_U350 ; P3_R1095_U173
g23743 not P3_U3443 ; P3_R1095_U174
g23744 nand P3_R1095_U274 P3_R1095_U273 ; P3_R1095_U175
g23745 nand P3_R1095_U270 P3_R1095_U269 ; P3_R1095_U176
g23746 and P3_R1095_U462 P3_R1095_U461 ; P3_R1095_U177
g23747 and P3_R1095_U466 P3_R1095_U465 ; P3_R1095_U178
g23748 nand P3_R1095_U260 P3_R1095_U259 ; P3_R1095_U179
g23749 nand P3_R1095_U256 P3_R1095_U255 ; P3_R1095_U180
g23750 nand P3_R1095_U252 P3_R1095_U251 ; P3_R1095_U181
g23751 and P3_R1095_U483 P3_R1095_U482 ; P3_R1095_U182
g23752 nand P3_R1095_U132 P3_R1095_U163 ; P3_R1095_U183
g23753 nand P3_R1095_U175 P3_R1095_U174 ; P3_R1095_U184
g23754 nand P3_R1095_U172 P3_R1095_U171 ; P3_R1095_U185
g23755 not P3_R1095_U87 ; P3_R1095_U186
g23756 not P3_R1095_U34 ; P3_R1095_U187
g23757 not P3_R1095_U26 ; P3_R1095_U188
g23758 nand P3_U3419 P3_R1095_U54 ; P3_R1095_U189
g23759 nand P3_U3434 P3_R1095_U64 ; P3_R1095_U190
g23760 nand P3_U3905 P3_R1095_U78 ; P3_R1095_U191
g23761 nand P3_U3901 P3_R1095_U86 ; P3_R1095_U192
g23762 nand P3_U3395 P3_R1095_U33 ; P3_R1095_U193
g23763 nand P3_U3404 P3_R1095_U41 ; P3_R1095_U194
g23764 nand P3_U3410 P3_R1095_U25 ; P3_R1095_U195
g23765 not P3_R1095_U66 ; P3_R1095_U196
g23766 not P3_R1095_U80 ; P3_R1095_U197
g23767 not P3_R1095_U43 ; P3_R1095_U198
g23768 not P3_R1095_U55 ; P3_R1095_U199
g23769 not P3_R1095_U172 ; P3_R1095_U200
g23770 nand P3_U3077 P3_R1095_U172 ; P3_R1095_U201
g23771 not P3_R1095_U49 ; P3_R1095_U202
g23772 nand P3_R1095_U117 P3_R1095_U49 ; P3_R1095_U203
g23773 nand P3_R1095_U35 P3_R1095_U34 ; P3_R1095_U204
g23774 nand P3_R1095_U204 P3_R1095_U32 ; P3_R1095_U205
g23775 nand P3_U3063 P3_R1095_U187 ; P3_R1095_U206
g23776 not P3_R1095_U158 ; P3_R1095_U207
g23777 nand P3_U3407 P3_R1095_U40 ; P3_R1095_U208
g23778 nand P3_U3070 P3_R1095_U37 ; P3_R1095_U209
g23779 nand P3_U3066 P3_R1095_U36 ; P3_R1095_U210
g23780 nand P3_R1095_U198 P3_R1095_U194 ; P3_R1095_U211
g23781 nand P3_R1095_U6 P3_R1095_U211 ; P3_R1095_U212
g23782 nand P3_U3401 P3_R1095_U42 ; P3_R1095_U213
g23783 nand P3_U3407 P3_R1095_U40 ; P3_R1095_U214
g23784 nand P3_R1095_U13 P3_R1095_U158 ; P3_R1095_U215
g23785 not P3_R1095_U44 ; P3_R1095_U216
g23786 not P3_R1095_U47 ; P3_R1095_U217
g23787 nand P3_U3413 P3_R1095_U27 ; P3_R1095_U218
g23788 nand P3_R1095_U27 P3_R1095_U26 ; P3_R1095_U219
g23789 nand P3_U3083 P3_R1095_U188 ; P3_R1095_U220
g23790 not P3_R1095_U154 ; P3_R1095_U221
g23791 nand P3_U3416 P3_R1095_U46 ; P3_R1095_U222
g23792 nand P3_R1095_U222 P3_R1095_U55 ; P3_R1095_U223
g23793 nand P3_R1095_U217 P3_R1095_U26 ; P3_R1095_U224
g23794 nand P3_R1095_U122 P3_R1095_U224 ; P3_R1095_U225
g23795 nand P3_R1095_U47 P3_R1095_U195 ; P3_R1095_U226
g23796 nand P3_R1095_U121 P3_R1095_U226 ; P3_R1095_U227
g23797 nand P3_R1095_U26 P3_R1095_U195 ; P3_R1095_U228
g23798 nand P3_R1095_U213 P3_R1095_U158 ; P3_R1095_U229
g23799 not P3_R1095_U48 ; P3_R1095_U230
g23800 nand P3_U3066 P3_R1095_U36 ; P3_R1095_U231
g23801 nand P3_R1095_U230 P3_R1095_U231 ; P3_R1095_U232
g23802 nand P3_R1095_U124 P3_R1095_U232 ; P3_R1095_U233
g23803 nand P3_R1095_U48 P3_R1095_U194 ; P3_R1095_U234
g23804 nand P3_U3407 P3_R1095_U40 ; P3_R1095_U235
g23805 nand P3_R1095_U123 P3_R1095_U234 ; P3_R1095_U236
g23806 nand P3_U3066 P3_R1095_U36 ; P3_R1095_U237
g23807 nand P3_R1095_U194 P3_R1095_U237 ; P3_R1095_U238
g23808 nand P3_R1095_U213 P3_R1095_U43 ; P3_R1095_U239
g23809 nand P3_R1095_U202 P3_R1095_U34 ; P3_R1095_U240
g23810 nand P3_R1095_U126 P3_R1095_U240 ; P3_R1095_U241
g23811 nand P3_R1095_U49 P3_R1095_U193 ; P3_R1095_U242
g23812 nand P3_R1095_U125 P3_R1095_U242 ; P3_R1095_U243
g23813 nand P3_R1095_U193 P3_R1095_U34 ; P3_R1095_U244
g23814 nand P3_U3422 P3_R1095_U53 ; P3_R1095_U245
g23815 nand P3_U3062 P3_R1095_U51 ; P3_R1095_U246
g23816 nand P3_U3061 P3_R1095_U52 ; P3_R1095_U247
g23817 nand P3_R1095_U199 P3_R1095_U7 ; P3_R1095_U248
g23818 nand P3_R1095_U8 P3_R1095_U248 ; P3_R1095_U249
g23819 nand P3_U3422 P3_R1095_U53 ; P3_R1095_U250
g23820 nand P3_R1095_U127 P3_R1095_U154 ; P3_R1095_U251
g23821 nand P3_R1095_U250 P3_R1095_U249 ; P3_R1095_U252
g23822 not P3_R1095_U181 ; P3_R1095_U253
g23823 nand P3_U3425 P3_R1095_U57 ; P3_R1095_U254
g23824 nand P3_R1095_U254 P3_R1095_U181 ; P3_R1095_U255
g23825 nand P3_U3071 P3_R1095_U56 ; P3_R1095_U256
g23826 not P3_R1095_U180 ; P3_R1095_U257
g23827 nand P3_U3428 P3_R1095_U59 ; P3_R1095_U258
g23828 nand P3_R1095_U258 P3_R1095_U180 ; P3_R1095_U259
g23829 nand P3_U3079 P3_R1095_U58 ; P3_R1095_U260
g23830 not P3_R1095_U179 ; P3_R1095_U261
g23831 nand P3_U3437 P3_R1095_U63 ; P3_R1095_U262
g23832 nand P3_U3072 P3_R1095_U60 ; P3_R1095_U263
g23833 nand P3_U3073 P3_R1095_U61 ; P3_R1095_U264
g23834 nand P3_R1095_U196 P3_R1095_U9 ; P3_R1095_U265
g23835 nand P3_R1095_U10 P3_R1095_U265 ; P3_R1095_U266
g23836 nand P3_U3431 P3_R1095_U65 ; P3_R1095_U267
g23837 nand P3_U3437 P3_R1095_U63 ; P3_R1095_U268
g23838 nand P3_R1095_U128 P3_R1095_U179 ; P3_R1095_U269
g23839 nand P3_R1095_U268 P3_R1095_U266 ; P3_R1095_U270
g23840 not P3_R1095_U176 ; P3_R1095_U271
g23841 nand P3_U3440 P3_R1095_U68 ; P3_R1095_U272
g23842 nand P3_R1095_U272 P3_R1095_U176 ; P3_R1095_U273
g23843 nand P3_U3068 P3_R1095_U67 ; P3_R1095_U274
g23844 not P3_R1095_U175 ; P3_R1095_U275
g23845 nand P3_U3081 P3_R1095_U175 ; P3_R1095_U276
g23846 not P3_R1095_U173 ; P3_R1095_U277
g23847 nand P3_U3445 P3_R1095_U71 ; P3_R1095_U278
g23848 nand P3_R1095_U278 P3_R1095_U173 ; P3_R1095_U279
g23849 nand P3_U3080 P3_R1095_U70 ; P3_R1095_U280
g23850 not P3_R1095_U170 ; P3_R1095_U281
g23851 nand P3_U3907 P3_R1095_U73 ; P3_R1095_U282
g23852 nand P3_R1095_U282 P3_R1095_U170 ; P3_R1095_U283
g23853 nand P3_U3075 P3_R1095_U72 ; P3_R1095_U284
g23854 not P3_R1095_U169 ; P3_R1095_U285
g23855 nand P3_U3904 P3_R1095_U77 ; P3_R1095_U286
g23856 nand P3_U3065 P3_R1095_U74 ; P3_R1095_U287
g23857 nand P3_U3060 P3_R1095_U75 ; P3_R1095_U288
g23858 nand P3_R1095_U197 P3_R1095_U11 ; P3_R1095_U289
g23859 nand P3_R1095_U12 P3_R1095_U289 ; P3_R1095_U290
g23860 nand P3_U3906 P3_R1095_U79 ; P3_R1095_U291
g23861 nand P3_U3904 P3_R1095_U77 ; P3_R1095_U292
g23862 nand P3_R1095_U129 P3_R1095_U169 ; P3_R1095_U293
g23863 nand P3_R1095_U292 P3_R1095_U290 ; P3_R1095_U294
g23864 not P3_R1095_U166 ; P3_R1095_U295
g23865 nand P3_U3903 P3_R1095_U82 ; P3_R1095_U296
g23866 nand P3_R1095_U296 P3_R1095_U166 ; P3_R1095_U297
g23867 nand P3_U3064 P3_R1095_U81 ; P3_R1095_U298
g23868 not P3_R1095_U165 ; P3_R1095_U299
g23869 nand P3_U3902 P3_R1095_U84 ; P3_R1095_U300
g23870 nand P3_R1095_U300 P3_R1095_U165 ; P3_R1095_U301
g23871 nand P3_U3057 P3_R1095_U83 ; P3_R1095_U302
g23872 not P3_R1095_U91 ; P3_R1095_U303
g23873 nand P3_R1095_U130 P3_R1095_U91 ; P3_R1095_U304
g23874 nand P3_R1095_U88 P3_R1095_U87 ; P3_R1095_U305
g23875 nand P3_R1095_U305 P3_R1095_U85 ; P3_R1095_U306
g23876 nand P3_U3052 P3_R1095_U186 ; P3_R1095_U307
g23877 not P3_R1095_U163 ; P3_R1095_U308
g23878 nand P3_U3899 P3_R1095_U90 ; P3_R1095_U309
g23879 nand P3_U3053 P3_R1095_U89 ; P3_R1095_U310
g23880 nand P3_R1095_U303 P3_R1095_U87 ; P3_R1095_U311
g23881 nand P3_R1095_U137 P3_R1095_U311 ; P3_R1095_U312
g23882 nand P3_R1095_U91 P3_R1095_U192 ; P3_R1095_U313
g23883 nand P3_R1095_U136 P3_R1095_U313 ; P3_R1095_U314
g23884 nand P3_R1095_U192 P3_R1095_U87 ; P3_R1095_U315
g23885 nand P3_R1095_U291 P3_R1095_U169 ; P3_R1095_U316
g23886 not P3_R1095_U92 ; P3_R1095_U317
g23887 nand P3_U3060 P3_R1095_U75 ; P3_R1095_U318
g23888 nand P3_R1095_U317 P3_R1095_U318 ; P3_R1095_U319
g23889 nand P3_R1095_U141 P3_R1095_U319 ; P3_R1095_U320
g23890 nand P3_R1095_U92 P3_R1095_U191 ; P3_R1095_U321
g23891 nand P3_U3904 P3_R1095_U77 ; P3_R1095_U322
g23892 nand P3_R1095_U140 P3_R1095_U321 ; P3_R1095_U323
g23893 nand P3_U3060 P3_R1095_U75 ; P3_R1095_U324
g23894 nand P3_R1095_U191 P3_R1095_U324 ; P3_R1095_U325
g23895 nand P3_R1095_U291 P3_R1095_U80 ; P3_R1095_U326
g23896 nand P3_R1095_U267 P3_R1095_U179 ; P3_R1095_U327
g23897 not P3_R1095_U93 ; P3_R1095_U328
g23898 nand P3_U3073 P3_R1095_U61 ; P3_R1095_U329
g23899 nand P3_R1095_U328 P3_R1095_U329 ; P3_R1095_U330
g23900 nand P3_R1095_U148 P3_R1095_U330 ; P3_R1095_U331
g23901 nand P3_R1095_U93 P3_R1095_U190 ; P3_R1095_U332
g23902 nand P3_U3437 P3_R1095_U63 ; P3_R1095_U333
g23903 nand P3_R1095_U147 P3_R1095_U332 ; P3_R1095_U334
g23904 nand P3_U3073 P3_R1095_U61 ; P3_R1095_U335
g23905 nand P3_R1095_U190 P3_R1095_U335 ; P3_R1095_U336
g23906 nand P3_R1095_U267 P3_R1095_U66 ; P3_R1095_U337
g23907 nand P3_R1095_U222 P3_R1095_U154 ; P3_R1095_U338
g23908 not P3_R1095_U94 ; P3_R1095_U339
g23909 nand P3_U3061 P3_R1095_U52 ; P3_R1095_U340
g23910 nand P3_R1095_U339 P3_R1095_U340 ; P3_R1095_U341
g23911 nand P3_R1095_U152 P3_R1095_U341 ; P3_R1095_U342
g23912 nand P3_R1095_U94 P3_R1095_U189 ; P3_R1095_U343
g23913 nand P3_U3422 P3_R1095_U53 ; P3_R1095_U344
g23914 nand P3_R1095_U151 P3_R1095_U343 ; P3_R1095_U345
g23915 nand P3_U3061 P3_R1095_U52 ; P3_R1095_U346
g23916 nand P3_R1095_U189 P3_R1095_U346 ; P3_R1095_U347
g23917 nand P3_U3076 P3_R1095_U30 ; P3_R1095_U348
g23918 nand P3_U3077 P3_R1095_U171 ; P3_R1095_U349
g23919 nand P3_U3081 P3_R1095_U174 ; P3_R1095_U350
g23920 nand P3_R1095_U133 P3_R1095_U304 P3_R1095_U134 ; P3_R1095_U351
g23921 nand P3_U3398 P3_R1095_U35 ; P3_R1095_U352
g23922 nand P3_U3413 P3_R1095_U220 ; P3_R1095_U353
g23923 nand P3_R1095_U353 P3_R1095_U219 ; P3_R1095_U354
g23924 nand P3_U3900 P3_R1095_U88 ; P3_R1095_U355
g23925 nand P3_R1095_U119 P3_R1095_U158 ; P3_R1095_U356
g23926 nand P3_R1095_U216 P3_R1095_U14 ; P3_R1095_U357
g23927 nand P3_U3416 P3_R1095_U46 ; P3_R1095_U358
g23928 nand P3_U3082 P3_R1095_U45 ; P3_R1095_U359
g23929 nand P3_R1095_U223 P3_R1095_U154 ; P3_R1095_U360
g23930 nand P3_R1095_U221 P3_R1095_U153 ; P3_R1095_U361
g23931 nand P3_U3413 P3_R1095_U27 ; P3_R1095_U362
g23932 nand P3_U3083 P3_R1095_U28 ; P3_R1095_U363
g23933 nand P3_U3413 P3_R1095_U27 ; P3_R1095_U364
g23934 nand P3_U3083 P3_R1095_U28 ; P3_R1095_U365
g23935 nand P3_R1095_U365 P3_R1095_U364 ; P3_R1095_U366
g23936 nand P3_U3410 P3_R1095_U25 ; P3_R1095_U367
g23937 nand P3_U3069 P3_R1095_U39 ; P3_R1095_U368
g23938 nand P3_R1095_U228 P3_R1095_U47 ; P3_R1095_U369
g23939 nand P3_R1095_U155 P3_R1095_U217 ; P3_R1095_U370
g23940 nand P3_U3407 P3_R1095_U40 ; P3_R1095_U371
g23941 nand P3_U3070 P3_R1095_U37 ; P3_R1095_U372
g23942 nand P3_R1095_U372 P3_R1095_U371 ; P3_R1095_U373
g23943 nand P3_U3404 P3_R1095_U41 ; P3_R1095_U374
g23944 nand P3_U3066 P3_R1095_U36 ; P3_R1095_U375
g23945 nand P3_R1095_U238 P3_R1095_U48 ; P3_R1095_U376
g23946 nand P3_R1095_U156 P3_R1095_U230 ; P3_R1095_U377
g23947 nand P3_U3401 P3_R1095_U42 ; P3_R1095_U378
g23948 nand P3_U3059 P3_R1095_U38 ; P3_R1095_U379
g23949 nand P3_R1095_U239 P3_R1095_U158 ; P3_R1095_U380
g23950 nand P3_R1095_U207 P3_R1095_U157 ; P3_R1095_U381
g23951 nand P3_U3398 P3_R1095_U35 ; P3_R1095_U382
g23952 nand P3_U3063 P3_R1095_U32 ; P3_R1095_U383
g23953 nand P3_U3398 P3_R1095_U35 ; P3_R1095_U384
g23954 nand P3_U3063 P3_R1095_U32 ; P3_R1095_U385
g23955 nand P3_R1095_U385 P3_R1095_U384 ; P3_R1095_U386
g23956 nand P3_U3395 P3_R1095_U33 ; P3_R1095_U387
g23957 nand P3_U3067 P3_R1095_U29 ; P3_R1095_U388
g23958 nand P3_R1095_U244 P3_R1095_U49 ; P3_R1095_U389
g23959 nand P3_R1095_U159 P3_R1095_U202 ; P3_R1095_U390
g23960 nand P3_U3908 P3_R1095_U161 ; P3_R1095_U391
g23961 nand P3_U3054 P3_R1095_U160 ; P3_R1095_U392
g23962 nand P3_U3908 P3_R1095_U161 ; P3_R1095_U393
g23963 nand P3_U3054 P3_R1095_U160 ; P3_R1095_U394
g23964 nand P3_R1095_U394 P3_R1095_U393 ; P3_R1095_U395
g23965 nand P3_U3053 P3_R1095_U395 P3_R1095_U89 ; P3_R1095_U396
g23966 nand P3_R1095_U15 P3_R1095_U90 P3_U3899 ; P3_R1095_U397
g23967 nand P3_U3899 P3_R1095_U90 ; P3_R1095_U398
g23968 nand P3_U3053 P3_R1095_U89 ; P3_R1095_U399
g23969 not P3_R1095_U135 ; P3_R1095_U400
g23970 nand P3_R1095_U308 P3_R1095_U400 ; P3_R1095_U401
g23971 nand P3_R1095_U135 P3_R1095_U163 ; P3_R1095_U402
g23972 nand P3_U3900 P3_R1095_U88 ; P3_R1095_U403
g23973 nand P3_U3052 P3_R1095_U85 ; P3_R1095_U404
g23974 nand P3_U3900 P3_R1095_U88 ; P3_R1095_U405
g23975 nand P3_U3052 P3_R1095_U85 ; P3_R1095_U406
g23976 nand P3_R1095_U406 P3_R1095_U405 ; P3_R1095_U407
g23977 nand P3_U3901 P3_R1095_U86 ; P3_R1095_U408
g23978 nand P3_U3056 P3_R1095_U50 ; P3_R1095_U409
g23979 nand P3_R1095_U315 P3_R1095_U91 ; P3_R1095_U410
g23980 nand P3_R1095_U164 P3_R1095_U303 ; P3_R1095_U411
g23981 nand P3_U3902 P3_R1095_U84 ; P3_R1095_U412
g23982 nand P3_U3057 P3_R1095_U83 ; P3_R1095_U413
g23983 not P3_R1095_U138 ; P3_R1095_U414
g23984 nand P3_R1095_U299 P3_R1095_U414 ; P3_R1095_U415
g23985 nand P3_R1095_U138 P3_R1095_U165 ; P3_R1095_U416
g23986 nand P3_U3903 P3_R1095_U82 ; P3_R1095_U417
g23987 nand P3_U3064 P3_R1095_U81 ; P3_R1095_U418
g23988 not P3_R1095_U139 ; P3_R1095_U419
g23989 nand P3_R1095_U295 P3_R1095_U419 ; P3_R1095_U420
g23990 nand P3_R1095_U139 P3_R1095_U166 ; P3_R1095_U421
g23991 nand P3_U3904 P3_R1095_U77 ; P3_R1095_U422
g23992 nand P3_U3065 P3_R1095_U74 ; P3_R1095_U423
g23993 nand P3_R1095_U423 P3_R1095_U422 ; P3_R1095_U424
g23994 nand P3_U3905 P3_R1095_U78 ; P3_R1095_U425
g23995 nand P3_U3060 P3_R1095_U75 ; P3_R1095_U426
g23996 nand P3_R1095_U325 P3_R1095_U92 ; P3_R1095_U427
g23997 nand P3_R1095_U167 P3_R1095_U317 ; P3_R1095_U428
g23998 nand P3_U3906 P3_R1095_U79 ; P3_R1095_U429
g23999 nand P3_U3074 P3_R1095_U76 ; P3_R1095_U430
g24000 nand P3_R1095_U326 P3_R1095_U169 ; P3_R1095_U431
g24001 nand P3_R1095_U285 P3_R1095_U168 ; P3_R1095_U432
g24002 nand P3_U3907 P3_R1095_U73 ; P3_R1095_U433
g24003 nand P3_U3075 P3_R1095_U72 ; P3_R1095_U434
g24004 not P3_R1095_U142 ; P3_R1095_U435
g24005 nand P3_R1095_U281 P3_R1095_U435 ; P3_R1095_U436
g24006 nand P3_R1095_U142 P3_R1095_U170 ; P3_R1095_U437
g24007 nand P3_U3392 P3_R1095_U31 ; P3_R1095_U438
g24008 nand P3_U3077 P3_R1095_U171 ; P3_R1095_U439
g24009 not P3_R1095_U143 ; P3_R1095_U440
g24010 nand P3_R1095_U200 P3_R1095_U440 ; P3_R1095_U441
g24011 nand P3_R1095_U143 P3_R1095_U172 ; P3_R1095_U442
g24012 nand P3_U3445 P3_R1095_U71 ; P3_R1095_U443
g24013 nand P3_U3080 P3_R1095_U70 ; P3_R1095_U444
g24014 not P3_R1095_U144 ; P3_R1095_U445
g24015 nand P3_R1095_U277 P3_R1095_U445 ; P3_R1095_U446
g24016 nand P3_R1095_U144 P3_R1095_U173 ; P3_R1095_U447
g24017 nand P3_U3443 P3_R1095_U69 ; P3_R1095_U448
g24018 nand P3_U3081 P3_R1095_U174 ; P3_R1095_U449
g24019 not P3_R1095_U145 ; P3_R1095_U450
g24020 nand P3_R1095_U275 P3_R1095_U450 ; P3_R1095_U451
g24021 nand P3_R1095_U145 P3_R1095_U175 ; P3_R1095_U452
g24022 nand P3_U3440 P3_R1095_U68 ; P3_R1095_U453
g24023 nand P3_U3068 P3_R1095_U67 ; P3_R1095_U454
g24024 not P3_R1095_U146 ; P3_R1095_U455
g24025 nand P3_R1095_U271 P3_R1095_U455 ; P3_R1095_U456
g24026 nand P3_R1095_U146 P3_R1095_U176 ; P3_R1095_U457
g24027 nand P3_U3437 P3_R1095_U63 ; P3_R1095_U458
g24028 nand P3_U3072 P3_R1095_U60 ; P3_R1095_U459
g24029 nand P3_R1095_U459 P3_R1095_U458 ; P3_R1095_U460
g24030 nand P3_U3434 P3_R1095_U64 ; P3_R1095_U461
g24031 nand P3_U3073 P3_R1095_U61 ; P3_R1095_U462
g24032 nand P3_R1095_U336 P3_R1095_U93 ; P3_R1095_U463
g24033 nand P3_R1095_U177 P3_R1095_U328 ; P3_R1095_U464
g24034 nand P3_U3431 P3_R1095_U65 ; P3_R1095_U465
g24035 nand P3_U3078 P3_R1095_U62 ; P3_R1095_U466
g24036 nand P3_R1095_U337 P3_R1095_U179 ; P3_R1095_U467
g24037 nand P3_R1095_U261 P3_R1095_U178 ; P3_R1095_U468
g24038 nand P3_U3428 P3_R1095_U59 ; P3_R1095_U469
g24039 nand P3_U3079 P3_R1095_U58 ; P3_R1095_U470
g24040 not P3_R1095_U149 ; P3_R1095_U471
g24041 nand P3_R1095_U257 P3_R1095_U471 ; P3_R1095_U472
g24042 nand P3_R1095_U149 P3_R1095_U180 ; P3_R1095_U473
g24043 nand P3_U3425 P3_R1095_U57 ; P3_R1095_U474
g24044 nand P3_U3071 P3_R1095_U56 ; P3_R1095_U475
g24045 not P3_R1095_U150 ; P3_R1095_U476
g24046 nand P3_R1095_U253 P3_R1095_U476 ; P3_R1095_U477
g24047 nand P3_R1095_U150 P3_R1095_U181 ; P3_R1095_U478
g24048 nand P3_U3422 P3_R1095_U53 ; P3_R1095_U479
g24049 nand P3_U3062 P3_R1095_U51 ; P3_R1095_U480
g24050 nand P3_R1095_U480 P3_R1095_U479 ; P3_R1095_U481
g24051 nand P3_U3419 P3_R1095_U54 ; P3_R1095_U482
g24052 nand P3_U3061 P3_R1095_U52 ; P3_R1095_U483
g24053 nand P3_R1095_U347 P3_R1095_U94 ; P3_R1095_U484
g24054 nand P3_R1095_U182 P3_R1095_U339 ; P3_R1095_U485
g24055 nand P3_R1212_U176 P3_R1212_U180 ; P3_R1212_U6
g24056 nand P3_R1212_U9 P3_R1212_U181 ; P3_R1212_U7
g24057 not P3_REG2_REG_0__SCAN_IN ; P3_R1212_U8
g24058 nand P3_R1212_U48 P3_REG2_REG_0__SCAN_IN ; P3_R1212_U9
g24059 not P3_REG2_REG_1__SCAN_IN ; P3_R1212_U10
g24060 not P3_U3391 ; P3_R1212_U11
g24061 not P3_REG2_REG_2__SCAN_IN ; P3_R1212_U12
g24062 not P3_U3394 ; P3_R1212_U13
g24063 not P3_REG2_REG_3__SCAN_IN ; P3_R1212_U14
g24064 not P3_U3397 ; P3_R1212_U15
g24065 not P3_REG2_REG_4__SCAN_IN ; P3_R1212_U16
g24066 not P3_U3400 ; P3_R1212_U17
g24067 not P3_REG2_REG_5__SCAN_IN ; P3_R1212_U18
g24068 not P3_U3403 ; P3_R1212_U19
g24069 not P3_REG2_REG_6__SCAN_IN ; P3_R1212_U20
g24070 not P3_U3406 ; P3_R1212_U21
g24071 not P3_REG2_REG_7__SCAN_IN ; P3_R1212_U22
g24072 not P3_U3409 ; P3_R1212_U23
g24073 not P3_REG2_REG_8__SCAN_IN ; P3_R1212_U24
g24074 not P3_U3412 ; P3_R1212_U25
g24075 not P3_REG2_REG_9__SCAN_IN ; P3_R1212_U26
g24076 not P3_U3415 ; P3_R1212_U27
g24077 not P3_REG2_REG_10__SCAN_IN ; P3_R1212_U28
g24078 not P3_U3418 ; P3_R1212_U29
g24079 not P3_REG2_REG_11__SCAN_IN ; P3_R1212_U30
g24080 not P3_U3421 ; P3_R1212_U31
g24081 not P3_REG2_REG_12__SCAN_IN ; P3_R1212_U32
g24082 not P3_U3424 ; P3_R1212_U33
g24083 not P3_REG2_REG_13__SCAN_IN ; P3_R1212_U34
g24084 not P3_U3427 ; P3_R1212_U35
g24085 not P3_REG2_REG_14__SCAN_IN ; P3_R1212_U36
g24086 not P3_U3430 ; P3_R1212_U37
g24087 nand P3_R1212_U159 P3_R1212_U158 ; P3_R1212_U38
g24088 not P3_REG2_REG_15__SCAN_IN ; P3_R1212_U39
g24089 not P3_U3433 ; P3_R1212_U40
g24090 not P3_REG2_REG_16__SCAN_IN ; P3_R1212_U41
g24091 not P3_U3436 ; P3_R1212_U42
g24092 not P3_REG2_REG_17__SCAN_IN ; P3_R1212_U43
g24093 not P3_U3439 ; P3_R1212_U44
g24094 not P3_REG2_REG_18__SCAN_IN ; P3_R1212_U45
g24095 not P3_U3442 ; P3_R1212_U46
g24096 nand P3_R1212_U171 P3_R1212_U170 ; P3_R1212_U47
g24097 not P3_U3386 ; P3_R1212_U48
g24098 nand P3_R1212_U186 P3_R1212_U185 ; P3_R1212_U49
g24099 nand P3_R1212_U191 P3_R1212_U190 ; P3_R1212_U50
g24100 nand P3_R1212_U196 P3_R1212_U195 ; P3_R1212_U51
g24101 nand P3_R1212_U201 P3_R1212_U200 ; P3_R1212_U52
g24102 nand P3_R1212_U206 P3_R1212_U205 ; P3_R1212_U53
g24103 nand P3_R1212_U211 P3_R1212_U210 ; P3_R1212_U54
g24104 nand P3_R1212_U216 P3_R1212_U215 ; P3_R1212_U55
g24105 nand P3_R1212_U221 P3_R1212_U220 ; P3_R1212_U56
g24106 nand P3_R1212_U226 P3_R1212_U225 ; P3_R1212_U57
g24107 nand P3_R1212_U236 P3_R1212_U235 ; P3_R1212_U58
g24108 nand P3_R1212_U241 P3_R1212_U240 ; P3_R1212_U59
g24109 nand P3_R1212_U246 P3_R1212_U245 ; P3_R1212_U60
g24110 nand P3_R1212_U251 P3_R1212_U250 ; P3_R1212_U61
g24111 nand P3_R1212_U256 P3_R1212_U255 ; P3_R1212_U62
g24112 nand P3_R1212_U261 P3_R1212_U260 ; P3_R1212_U63
g24113 nand P3_R1212_U266 P3_R1212_U265 ; P3_R1212_U64
g24114 nand P3_R1212_U271 P3_R1212_U270 ; P3_R1212_U65
g24115 nand P3_R1212_U276 P3_R1212_U275 ; P3_R1212_U66
g24116 nand P3_R1212_U183 P3_R1212_U182 ; P3_R1212_U67
g24117 nand P3_R1212_U188 P3_R1212_U187 ; P3_R1212_U68
g24118 nand P3_R1212_U193 P3_R1212_U192 ; P3_R1212_U69
g24119 nand P3_R1212_U198 P3_R1212_U197 ; P3_R1212_U70
g24120 nand P3_R1212_U203 P3_R1212_U202 ; P3_R1212_U71
g24121 nand P3_R1212_U208 P3_R1212_U207 ; P3_R1212_U72
g24122 nand P3_R1212_U213 P3_R1212_U212 ; P3_R1212_U73
g24123 nand P3_R1212_U218 P3_R1212_U217 ; P3_R1212_U74
g24124 nand P3_R1212_U223 P3_R1212_U222 ; P3_R1212_U75
g24125 and P3_R1212_U228 P3_R1212_U227 P3_R1212_U179 ; P3_R1212_U76
g24126 and P3_R1212_U175 P3_R1212_U231 ; P3_R1212_U77
g24127 nand P3_R1212_U233 P3_R1212_U232 ; P3_R1212_U78
g24128 nand P3_R1212_U238 P3_R1212_U237 ; P3_R1212_U79
g24129 nand P3_R1212_U243 P3_R1212_U242 ; P3_R1212_U80
g24130 nand P3_R1212_U248 P3_R1212_U247 ; P3_R1212_U81
g24131 nand P3_R1212_U253 P3_R1212_U252 ; P3_R1212_U82
g24132 nand P3_R1212_U258 P3_R1212_U257 ; P3_R1212_U83
g24133 nand P3_R1212_U263 P3_R1212_U262 ; P3_R1212_U84
g24134 nand P3_R1212_U268 P3_R1212_U267 ; P3_R1212_U85
g24135 nand P3_R1212_U273 P3_R1212_U272 ; P3_R1212_U86
g24136 nand P3_R1212_U135 P3_R1212_U134 ; P3_R1212_U87
g24137 nand P3_R1212_U131 P3_R1212_U130 ; P3_R1212_U88
g24138 nand P3_R1212_U127 P3_R1212_U126 ; P3_R1212_U89
g24139 nand P3_R1212_U123 P3_R1212_U122 ; P3_R1212_U90
g24140 nand P3_R1212_U119 P3_R1212_U118 ; P3_R1212_U91
g24141 nand P3_R1212_U115 P3_R1212_U114 ; P3_R1212_U92
g24142 nand P3_R1212_U111 P3_R1212_U110 ; P3_R1212_U93
g24143 nand P3_R1212_U107 P3_R1212_U106 ; P3_R1212_U94
g24144 not P3_REG2_REG_19__SCAN_IN ; P3_R1212_U95
g24145 not P3_U3379 ; P3_R1212_U96
g24146 nand P3_R1212_U167 P3_R1212_U166 ; P3_R1212_U97
g24147 nand P3_R1212_U163 P3_R1212_U162 ; P3_R1212_U98
g24148 nand P3_R1212_U155 P3_R1212_U154 ; P3_R1212_U99
g24149 nand P3_R1212_U151 P3_R1212_U150 ; P3_R1212_U100
g24150 nand P3_R1212_U147 P3_R1212_U146 ; P3_R1212_U101
g24151 nand P3_R1212_U143 P3_R1212_U142 ; P3_R1212_U102
g24152 nand P3_R1212_U139 P3_R1212_U138 ; P3_R1212_U103
g24153 not P3_R1212_U9 ; P3_R1212_U104
g24154 nand P3_R1212_U104 P3_REG2_REG_1__SCAN_IN ; P3_R1212_U105
g24155 nand P3_U3391 P3_R1212_U105 ; P3_R1212_U106
g24156 nand P3_R1212_U9 P3_R1212_U10 ; P3_R1212_U107
g24157 not P3_R1212_U94 ; P3_R1212_U108
g24158 nand P3_R1212_U13 P3_REG2_REG_2__SCAN_IN ; P3_R1212_U109
g24159 nand P3_R1212_U109 P3_R1212_U94 ; P3_R1212_U110
g24160 nand P3_U3394 P3_R1212_U12 ; P3_R1212_U111
g24161 not P3_R1212_U93 ; P3_R1212_U112
g24162 nand P3_R1212_U15 P3_REG2_REG_3__SCAN_IN ; P3_R1212_U113
g24163 nand P3_R1212_U113 P3_R1212_U93 ; P3_R1212_U114
g24164 nand P3_U3397 P3_R1212_U14 ; P3_R1212_U115
g24165 not P3_R1212_U92 ; P3_R1212_U116
g24166 nand P3_R1212_U17 P3_REG2_REG_4__SCAN_IN ; P3_R1212_U117
g24167 nand P3_R1212_U117 P3_R1212_U92 ; P3_R1212_U118
g24168 nand P3_U3400 P3_R1212_U16 ; P3_R1212_U119
g24169 not P3_R1212_U91 ; P3_R1212_U120
g24170 nand P3_R1212_U19 P3_REG2_REG_5__SCAN_IN ; P3_R1212_U121
g24171 nand P3_R1212_U121 P3_R1212_U91 ; P3_R1212_U122
g24172 nand P3_U3403 P3_R1212_U18 ; P3_R1212_U123
g24173 not P3_R1212_U90 ; P3_R1212_U124
g24174 nand P3_R1212_U21 P3_REG2_REG_6__SCAN_IN ; P3_R1212_U125
g24175 nand P3_R1212_U125 P3_R1212_U90 ; P3_R1212_U126
g24176 nand P3_U3406 P3_R1212_U20 ; P3_R1212_U127
g24177 not P3_R1212_U89 ; P3_R1212_U128
g24178 nand P3_R1212_U23 P3_REG2_REG_7__SCAN_IN ; P3_R1212_U129
g24179 nand P3_R1212_U129 P3_R1212_U89 ; P3_R1212_U130
g24180 nand P3_U3409 P3_R1212_U22 ; P3_R1212_U131
g24181 not P3_R1212_U88 ; P3_R1212_U132
g24182 nand P3_R1212_U25 P3_REG2_REG_8__SCAN_IN ; P3_R1212_U133
g24183 nand P3_R1212_U133 P3_R1212_U88 ; P3_R1212_U134
g24184 nand P3_U3412 P3_R1212_U24 ; P3_R1212_U135
g24185 not P3_R1212_U87 ; P3_R1212_U136
g24186 nand P3_R1212_U27 P3_REG2_REG_9__SCAN_IN ; P3_R1212_U137
g24187 nand P3_R1212_U137 P3_R1212_U87 ; P3_R1212_U138
g24188 nand P3_U3415 P3_R1212_U26 ; P3_R1212_U139
g24189 not P3_R1212_U103 ; P3_R1212_U140
g24190 nand P3_R1212_U29 P3_REG2_REG_10__SCAN_IN ; P3_R1212_U141
g24191 nand P3_R1212_U141 P3_R1212_U103 ; P3_R1212_U142
g24192 nand P3_U3418 P3_R1212_U28 ; P3_R1212_U143
g24193 not P3_R1212_U102 ; P3_R1212_U144
g24194 nand P3_R1212_U31 P3_REG2_REG_11__SCAN_IN ; P3_R1212_U145
g24195 nand P3_R1212_U145 P3_R1212_U102 ; P3_R1212_U146
g24196 nand P3_U3421 P3_R1212_U30 ; P3_R1212_U147
g24197 not P3_R1212_U101 ; P3_R1212_U148
g24198 nand P3_R1212_U33 P3_REG2_REG_12__SCAN_IN ; P3_R1212_U149
g24199 nand P3_R1212_U149 P3_R1212_U101 ; P3_R1212_U150
g24200 nand P3_U3424 P3_R1212_U32 ; P3_R1212_U151
g24201 not P3_R1212_U100 ; P3_R1212_U152
g24202 nand P3_R1212_U35 P3_REG2_REG_13__SCAN_IN ; P3_R1212_U153
g24203 nand P3_R1212_U153 P3_R1212_U100 ; P3_R1212_U154
g24204 nand P3_U3427 P3_R1212_U34 ; P3_R1212_U155
g24205 not P3_R1212_U99 ; P3_R1212_U156
g24206 nand P3_R1212_U37 P3_REG2_REG_14__SCAN_IN ; P3_R1212_U157
g24207 nand P3_R1212_U157 P3_R1212_U99 ; P3_R1212_U158
g24208 nand P3_U3430 P3_R1212_U36 ; P3_R1212_U159
g24209 not P3_R1212_U38 ; P3_R1212_U160
g24210 nand P3_R1212_U160 P3_REG2_REG_15__SCAN_IN ; P3_R1212_U161
g24211 nand P3_U3433 P3_R1212_U161 ; P3_R1212_U162
g24212 nand P3_R1212_U38 P3_R1212_U39 ; P3_R1212_U163
g24213 not P3_R1212_U98 ; P3_R1212_U164
g24214 nand P3_R1212_U42 P3_REG2_REG_16__SCAN_IN ; P3_R1212_U165
g24215 nand P3_R1212_U165 P3_R1212_U98 ; P3_R1212_U166
g24216 nand P3_U3436 P3_R1212_U41 ; P3_R1212_U167
g24217 not P3_R1212_U97 ; P3_R1212_U168
g24218 nand P3_R1212_U44 P3_REG2_REG_17__SCAN_IN ; P3_R1212_U169
g24219 nand P3_R1212_U169 P3_R1212_U97 ; P3_R1212_U170
g24220 nand P3_U3439 P3_R1212_U43 ; P3_R1212_U171
g24221 not P3_R1212_U47 ; P3_R1212_U172
g24222 nand P3_U3442 P3_R1212_U45 ; P3_R1212_U173
g24223 nand P3_R1212_U172 P3_R1212_U173 ; P3_R1212_U174
g24224 nand P3_R1212_U46 P3_REG2_REG_18__SCAN_IN ; P3_R1212_U175
g24225 nand P3_R1212_U77 P3_R1212_U174 ; P3_R1212_U176
g24226 nand P3_R1212_U46 P3_REG2_REG_18__SCAN_IN ; P3_R1212_U177
g24227 nand P3_R1212_U177 P3_R1212_U47 ; P3_R1212_U178
g24228 nand P3_U3442 P3_R1212_U45 ; P3_R1212_U179
g24229 nand P3_R1212_U76 P3_R1212_U178 ; P3_R1212_U180
g24230 nand P3_U3386 P3_R1212_U8 ; P3_R1212_U181
g24231 nand P3_R1212_U27 P3_REG2_REG_9__SCAN_IN ; P3_R1212_U182
g24232 nand P3_U3415 P3_R1212_U26 ; P3_R1212_U183
g24233 not P3_R1212_U67 ; P3_R1212_U184
g24234 nand P3_R1212_U136 P3_R1212_U184 ; P3_R1212_U185
g24235 nand P3_R1212_U67 P3_R1212_U87 ; P3_R1212_U186
g24236 nand P3_R1212_U25 P3_REG2_REG_8__SCAN_IN ; P3_R1212_U187
g24237 nand P3_U3412 P3_R1212_U24 ; P3_R1212_U188
g24238 not P3_R1212_U68 ; P3_R1212_U189
g24239 nand P3_R1212_U132 P3_R1212_U189 ; P3_R1212_U190
g24240 nand P3_R1212_U68 P3_R1212_U88 ; P3_R1212_U191
g24241 nand P3_R1212_U23 P3_REG2_REG_7__SCAN_IN ; P3_R1212_U192
g24242 nand P3_U3409 P3_R1212_U22 ; P3_R1212_U193
g24243 not P3_R1212_U69 ; P3_R1212_U194
g24244 nand P3_R1212_U128 P3_R1212_U194 ; P3_R1212_U195
g24245 nand P3_R1212_U69 P3_R1212_U89 ; P3_R1212_U196
g24246 nand P3_R1212_U21 P3_REG2_REG_6__SCAN_IN ; P3_R1212_U197
g24247 nand P3_U3406 P3_R1212_U20 ; P3_R1212_U198
g24248 not P3_R1212_U70 ; P3_R1212_U199
g24249 nand P3_R1212_U124 P3_R1212_U199 ; P3_R1212_U200
g24250 nand P3_R1212_U70 P3_R1212_U90 ; P3_R1212_U201
g24251 nand P3_R1212_U19 P3_REG2_REG_5__SCAN_IN ; P3_R1212_U202
g24252 nand P3_U3403 P3_R1212_U18 ; P3_R1212_U203
g24253 not P3_R1212_U71 ; P3_R1212_U204
g24254 nand P3_R1212_U120 P3_R1212_U204 ; P3_R1212_U205
g24255 nand P3_R1212_U71 P3_R1212_U91 ; P3_R1212_U206
g24256 nand P3_R1212_U17 P3_REG2_REG_4__SCAN_IN ; P3_R1212_U207
g24257 nand P3_U3400 P3_R1212_U16 ; P3_R1212_U208
g24258 not P3_R1212_U72 ; P3_R1212_U209
g24259 nand P3_R1212_U116 P3_R1212_U209 ; P3_R1212_U210
g24260 nand P3_R1212_U72 P3_R1212_U92 ; P3_R1212_U211
g24261 nand P3_R1212_U15 P3_REG2_REG_3__SCAN_IN ; P3_R1212_U212
g24262 nand P3_U3397 P3_R1212_U14 ; P3_R1212_U213
g24263 not P3_R1212_U73 ; P3_R1212_U214
g24264 nand P3_R1212_U112 P3_R1212_U214 ; P3_R1212_U215
g24265 nand P3_R1212_U73 P3_R1212_U93 ; P3_R1212_U216
g24266 nand P3_R1212_U13 P3_REG2_REG_2__SCAN_IN ; P3_R1212_U217
g24267 nand P3_U3394 P3_R1212_U12 ; P3_R1212_U218
g24268 not P3_R1212_U74 ; P3_R1212_U219
g24269 nand P3_R1212_U108 P3_R1212_U219 ; P3_R1212_U220
g24270 nand P3_R1212_U74 P3_R1212_U94 ; P3_R1212_U221
g24271 nand P3_R1212_U104 P3_R1212_U10 ; P3_R1212_U222
g24272 nand P3_R1212_U9 P3_REG2_REG_1__SCAN_IN ; P3_R1212_U223
g24273 not P3_R1212_U75 ; P3_R1212_U224
g24274 nand P3_R1212_U224 P3_U3391 ; P3_R1212_U225
g24275 nand P3_R1212_U75 P3_R1212_U11 ; P3_R1212_U226
g24276 nand P3_R1212_U96 P3_REG2_REG_19__SCAN_IN ; P3_R1212_U227
g24277 nand P3_U3379 P3_R1212_U95 ; P3_R1212_U228
g24278 nand P3_R1212_U96 P3_REG2_REG_19__SCAN_IN ; P3_R1212_U229
g24279 nand P3_U3379 P3_R1212_U95 ; P3_R1212_U230
g24280 nand P3_R1212_U230 P3_R1212_U229 ; P3_R1212_U231
g24281 nand P3_R1212_U46 P3_REG2_REG_18__SCAN_IN ; P3_R1212_U232
g24282 nand P3_U3442 P3_R1212_U45 ; P3_R1212_U233
g24283 not P3_R1212_U78 ; P3_R1212_U234
g24284 nand P3_R1212_U234 P3_R1212_U172 ; P3_R1212_U235
g24285 nand P3_R1212_U78 P3_R1212_U47 ; P3_R1212_U236
g24286 nand P3_R1212_U44 P3_REG2_REG_17__SCAN_IN ; P3_R1212_U237
g24287 nand P3_U3439 P3_R1212_U43 ; P3_R1212_U238
g24288 not P3_R1212_U79 ; P3_R1212_U239
g24289 nand P3_R1212_U168 P3_R1212_U239 ; P3_R1212_U240
g24290 nand P3_R1212_U79 P3_R1212_U97 ; P3_R1212_U241
g24291 nand P3_R1212_U42 P3_REG2_REG_16__SCAN_IN ; P3_R1212_U242
g24292 nand P3_U3436 P3_R1212_U41 ; P3_R1212_U243
g24293 not P3_R1212_U80 ; P3_R1212_U244
g24294 nand P3_R1212_U164 P3_R1212_U244 ; P3_R1212_U245
g24295 nand P3_R1212_U80 P3_R1212_U98 ; P3_R1212_U246
g24296 nand P3_U3433 P3_R1212_U39 ; P3_R1212_U247
g24297 nand P3_R1212_U40 P3_REG2_REG_15__SCAN_IN ; P3_R1212_U248
g24298 not P3_R1212_U81 ; P3_R1212_U249
g24299 nand P3_R1212_U249 P3_R1212_U160 ; P3_R1212_U250
g24300 nand P3_R1212_U81 P3_R1212_U38 ; P3_R1212_U251
g24301 nand P3_R1212_U37 P3_REG2_REG_14__SCAN_IN ; P3_R1212_U252
g24302 nand P3_U3430 P3_R1212_U36 ; P3_R1212_U253
g24303 not P3_R1212_U82 ; P3_R1212_U254
g24304 nand P3_R1212_U156 P3_R1212_U254 ; P3_R1212_U255
g24305 nand P3_R1212_U82 P3_R1212_U99 ; P3_R1212_U256
g24306 nand P3_R1212_U35 P3_REG2_REG_13__SCAN_IN ; P3_R1212_U257
g24307 nand P3_U3427 P3_R1212_U34 ; P3_R1212_U258
g24308 not P3_R1212_U83 ; P3_R1212_U259
g24309 nand P3_R1212_U152 P3_R1212_U259 ; P3_R1212_U260
g24310 nand P3_R1212_U83 P3_R1212_U100 ; P3_R1212_U261
g24311 nand P3_R1212_U33 P3_REG2_REG_12__SCAN_IN ; P3_R1212_U262
g24312 nand P3_U3424 P3_R1212_U32 ; P3_R1212_U263
g24313 not P3_R1212_U84 ; P3_R1212_U264
g24314 nand P3_R1212_U148 P3_R1212_U264 ; P3_R1212_U265
g24315 nand P3_R1212_U84 P3_R1212_U101 ; P3_R1212_U266
g24316 nand P3_R1212_U31 P3_REG2_REG_11__SCAN_IN ; P3_R1212_U267
g24317 nand P3_U3421 P3_R1212_U30 ; P3_R1212_U268
g24318 not P3_R1212_U85 ; P3_R1212_U269
g24319 nand P3_R1212_U144 P3_R1212_U269 ; P3_R1212_U270
g24320 nand P3_R1212_U85 P3_R1212_U102 ; P3_R1212_U271
g24321 nand P3_R1212_U29 P3_REG2_REG_10__SCAN_IN ; P3_R1212_U272
g24322 nand P3_U3418 P3_R1212_U28 ; P3_R1212_U273
g24323 not P3_R1212_U86 ; P3_R1212_U274
g24324 nand P3_R1212_U140 P3_R1212_U274 ; P3_R1212_U275
g24325 nand P3_R1212_U86 P3_R1212_U103 ; P3_R1212_U276
g24326 nand P3_R1209_U176 P3_R1209_U180 ; P3_R1209_U6
g24327 nand P3_R1209_U9 P3_R1209_U181 ; P3_R1209_U7
g24328 not P3_REG1_REG_0__SCAN_IN ; P3_R1209_U8
g24329 nand P3_R1209_U48 P3_REG1_REG_0__SCAN_IN ; P3_R1209_U9
g24330 not P3_REG1_REG_1__SCAN_IN ; P3_R1209_U10
g24331 not P3_U3391 ; P3_R1209_U11
g24332 not P3_REG1_REG_2__SCAN_IN ; P3_R1209_U12
g24333 not P3_U3394 ; P3_R1209_U13
g24334 not P3_REG1_REG_3__SCAN_IN ; P3_R1209_U14
g24335 not P3_U3397 ; P3_R1209_U15
g24336 not P3_REG1_REG_4__SCAN_IN ; P3_R1209_U16
g24337 not P3_U3400 ; P3_R1209_U17
g24338 not P3_REG1_REG_5__SCAN_IN ; P3_R1209_U18
g24339 not P3_U3403 ; P3_R1209_U19
g24340 not P3_REG1_REG_6__SCAN_IN ; P3_R1209_U20
g24341 not P3_U3406 ; P3_R1209_U21
g24342 not P3_REG1_REG_7__SCAN_IN ; P3_R1209_U22
g24343 not P3_U3409 ; P3_R1209_U23
g24344 not P3_REG1_REG_8__SCAN_IN ; P3_R1209_U24
g24345 not P3_U3412 ; P3_R1209_U25
g24346 not P3_REG1_REG_9__SCAN_IN ; P3_R1209_U26
g24347 not P3_U3415 ; P3_R1209_U27
g24348 not P3_REG1_REG_10__SCAN_IN ; P3_R1209_U28
g24349 not P3_U3418 ; P3_R1209_U29
g24350 not P3_REG1_REG_11__SCAN_IN ; P3_R1209_U30
g24351 not P3_U3421 ; P3_R1209_U31
g24352 not P3_REG1_REG_12__SCAN_IN ; P3_R1209_U32
g24353 not P3_U3424 ; P3_R1209_U33
g24354 not P3_REG1_REG_13__SCAN_IN ; P3_R1209_U34
g24355 not P3_U3427 ; P3_R1209_U35
g24356 not P3_REG1_REG_14__SCAN_IN ; P3_R1209_U36
g24357 not P3_U3430 ; P3_R1209_U37
g24358 nand P3_R1209_U159 P3_R1209_U158 ; P3_R1209_U38
g24359 not P3_REG1_REG_15__SCAN_IN ; P3_R1209_U39
g24360 not P3_U3433 ; P3_R1209_U40
g24361 not P3_REG1_REG_16__SCAN_IN ; P3_R1209_U41
g24362 not P3_U3436 ; P3_R1209_U42
g24363 not P3_REG1_REG_17__SCAN_IN ; P3_R1209_U43
g24364 not P3_U3439 ; P3_R1209_U44
g24365 not P3_REG1_REG_18__SCAN_IN ; P3_R1209_U45
g24366 not P3_U3442 ; P3_R1209_U46
g24367 nand P3_R1209_U171 P3_R1209_U170 ; P3_R1209_U47
g24368 not P3_U3386 ; P3_R1209_U48
g24369 nand P3_R1209_U186 P3_R1209_U185 ; P3_R1209_U49
g24370 nand P3_R1209_U191 P3_R1209_U190 ; P3_R1209_U50
g24371 nand P3_R1209_U196 P3_R1209_U195 ; P3_R1209_U51
g24372 nand P3_R1209_U201 P3_R1209_U200 ; P3_R1209_U52
g24373 nand P3_R1209_U206 P3_R1209_U205 ; P3_R1209_U53
g24374 nand P3_R1209_U211 P3_R1209_U210 ; P3_R1209_U54
g24375 nand P3_R1209_U216 P3_R1209_U215 ; P3_R1209_U55
g24376 nand P3_R1209_U221 P3_R1209_U220 ; P3_R1209_U56
g24377 nand P3_R1209_U226 P3_R1209_U225 ; P3_R1209_U57
g24378 nand P3_R1209_U236 P3_R1209_U235 ; P3_R1209_U58
g24379 nand P3_R1209_U241 P3_R1209_U240 ; P3_R1209_U59
g24380 nand P3_R1209_U246 P3_R1209_U245 ; P3_R1209_U60
g24381 nand P3_R1209_U251 P3_R1209_U250 ; P3_R1209_U61
g24382 nand P3_R1209_U256 P3_R1209_U255 ; P3_R1209_U62
g24383 nand P3_R1209_U261 P3_R1209_U260 ; P3_R1209_U63
g24384 nand P3_R1209_U266 P3_R1209_U265 ; P3_R1209_U64
g24385 nand P3_R1209_U271 P3_R1209_U270 ; P3_R1209_U65
g24386 nand P3_R1209_U276 P3_R1209_U275 ; P3_R1209_U66
g24387 nand P3_R1209_U183 P3_R1209_U182 ; P3_R1209_U67
g24388 nand P3_R1209_U188 P3_R1209_U187 ; P3_R1209_U68
g24389 nand P3_R1209_U193 P3_R1209_U192 ; P3_R1209_U69
g24390 nand P3_R1209_U198 P3_R1209_U197 ; P3_R1209_U70
g24391 nand P3_R1209_U203 P3_R1209_U202 ; P3_R1209_U71
g24392 nand P3_R1209_U208 P3_R1209_U207 ; P3_R1209_U72
g24393 nand P3_R1209_U213 P3_R1209_U212 ; P3_R1209_U73
g24394 nand P3_R1209_U218 P3_R1209_U217 ; P3_R1209_U74
g24395 nand P3_R1209_U223 P3_R1209_U222 ; P3_R1209_U75
g24396 and P3_R1209_U228 P3_R1209_U227 P3_R1209_U179 ; P3_R1209_U76
g24397 and P3_R1209_U175 P3_R1209_U231 ; P3_R1209_U77
g24398 nand P3_R1209_U233 P3_R1209_U232 ; P3_R1209_U78
g24399 nand P3_R1209_U238 P3_R1209_U237 ; P3_R1209_U79
g24400 nand P3_R1209_U243 P3_R1209_U242 ; P3_R1209_U80
g24401 nand P3_R1209_U248 P3_R1209_U247 ; P3_R1209_U81
g24402 nand P3_R1209_U253 P3_R1209_U252 ; P3_R1209_U82
g24403 nand P3_R1209_U258 P3_R1209_U257 ; P3_R1209_U83
g24404 nand P3_R1209_U263 P3_R1209_U262 ; P3_R1209_U84
g24405 nand P3_R1209_U268 P3_R1209_U267 ; P3_R1209_U85
g24406 nand P3_R1209_U273 P3_R1209_U272 ; P3_R1209_U86
g24407 nand P3_R1209_U135 P3_R1209_U134 ; P3_R1209_U87
g24408 nand P3_R1209_U131 P3_R1209_U130 ; P3_R1209_U88
g24409 nand P3_R1209_U127 P3_R1209_U126 ; P3_R1209_U89
g24410 nand P3_R1209_U123 P3_R1209_U122 ; P3_R1209_U90
g24411 nand P3_R1209_U119 P3_R1209_U118 ; P3_R1209_U91
g24412 nand P3_R1209_U115 P3_R1209_U114 ; P3_R1209_U92
g24413 nand P3_R1209_U111 P3_R1209_U110 ; P3_R1209_U93
g24414 nand P3_R1209_U107 P3_R1209_U106 ; P3_R1209_U94
g24415 not P3_REG1_REG_19__SCAN_IN ; P3_R1209_U95
g24416 not P3_U3379 ; P3_R1209_U96
g24417 nand P3_R1209_U167 P3_R1209_U166 ; P3_R1209_U97
g24418 nand P3_R1209_U163 P3_R1209_U162 ; P3_R1209_U98
g24419 nand P3_R1209_U155 P3_R1209_U154 ; P3_R1209_U99
g24420 nand P3_R1209_U151 P3_R1209_U150 ; P3_R1209_U100
g24421 nand P3_R1209_U147 P3_R1209_U146 ; P3_R1209_U101
g24422 nand P3_R1209_U143 P3_R1209_U142 ; P3_R1209_U102
g24423 nand P3_R1209_U139 P3_R1209_U138 ; P3_R1209_U103
g24424 not P3_R1209_U9 ; P3_R1209_U104
g24425 nand P3_R1209_U104 P3_REG1_REG_1__SCAN_IN ; P3_R1209_U105
g24426 nand P3_U3391 P3_R1209_U105 ; P3_R1209_U106
g24427 nand P3_R1209_U9 P3_R1209_U10 ; P3_R1209_U107
g24428 not P3_R1209_U94 ; P3_R1209_U108
g24429 nand P3_R1209_U13 P3_REG1_REG_2__SCAN_IN ; P3_R1209_U109
g24430 nand P3_R1209_U109 P3_R1209_U94 ; P3_R1209_U110
g24431 nand P3_U3394 P3_R1209_U12 ; P3_R1209_U111
g24432 not P3_R1209_U93 ; P3_R1209_U112
g24433 nand P3_R1209_U15 P3_REG1_REG_3__SCAN_IN ; P3_R1209_U113
g24434 nand P3_R1209_U113 P3_R1209_U93 ; P3_R1209_U114
g24435 nand P3_U3397 P3_R1209_U14 ; P3_R1209_U115
g24436 not P3_R1209_U92 ; P3_R1209_U116
g24437 nand P3_R1209_U17 P3_REG1_REG_4__SCAN_IN ; P3_R1209_U117
g24438 nand P3_R1209_U117 P3_R1209_U92 ; P3_R1209_U118
g24439 nand P3_U3400 P3_R1209_U16 ; P3_R1209_U119
g24440 not P3_R1209_U91 ; P3_R1209_U120
g24441 nand P3_R1209_U19 P3_REG1_REG_5__SCAN_IN ; P3_R1209_U121
g24442 nand P3_R1209_U121 P3_R1209_U91 ; P3_R1209_U122
g24443 nand P3_U3403 P3_R1209_U18 ; P3_R1209_U123
g24444 not P3_R1209_U90 ; P3_R1209_U124
g24445 nand P3_R1209_U21 P3_REG1_REG_6__SCAN_IN ; P3_R1209_U125
g24446 nand P3_R1209_U125 P3_R1209_U90 ; P3_R1209_U126
g24447 nand P3_U3406 P3_R1209_U20 ; P3_R1209_U127
g24448 not P3_R1209_U89 ; P3_R1209_U128
g24449 nand P3_R1209_U23 P3_REG1_REG_7__SCAN_IN ; P3_R1209_U129
g24450 nand P3_R1209_U129 P3_R1209_U89 ; P3_R1209_U130
g24451 nand P3_U3409 P3_R1209_U22 ; P3_R1209_U131
g24452 not P3_R1209_U88 ; P3_R1209_U132
g24453 nand P3_R1209_U25 P3_REG1_REG_8__SCAN_IN ; P3_R1209_U133
g24454 nand P3_R1209_U133 P3_R1209_U88 ; P3_R1209_U134
g24455 nand P3_U3412 P3_R1209_U24 ; P3_R1209_U135
g24456 not P3_R1209_U87 ; P3_R1209_U136
g24457 nand P3_R1209_U27 P3_REG1_REG_9__SCAN_IN ; P3_R1209_U137
g24458 nand P3_R1209_U137 P3_R1209_U87 ; P3_R1209_U138
g24459 nand P3_U3415 P3_R1209_U26 ; P3_R1209_U139
g24460 not P3_R1209_U103 ; P3_R1209_U140
g24461 nand P3_R1209_U29 P3_REG1_REG_10__SCAN_IN ; P3_R1209_U141
g24462 nand P3_R1209_U141 P3_R1209_U103 ; P3_R1209_U142
g24463 nand P3_U3418 P3_R1209_U28 ; P3_R1209_U143
g24464 not P3_R1209_U102 ; P3_R1209_U144
g24465 nand P3_R1209_U31 P3_REG1_REG_11__SCAN_IN ; P3_R1209_U145
g24466 nand P3_R1209_U145 P3_R1209_U102 ; P3_R1209_U146
g24467 nand P3_U3421 P3_R1209_U30 ; P3_R1209_U147
g24468 not P3_R1209_U101 ; P3_R1209_U148
g24469 nand P3_R1209_U33 P3_REG1_REG_12__SCAN_IN ; P3_R1209_U149
g24470 nand P3_R1209_U149 P3_R1209_U101 ; P3_R1209_U150
g24471 nand P3_U3424 P3_R1209_U32 ; P3_R1209_U151
g24472 not P3_R1209_U100 ; P3_R1209_U152
g24473 nand P3_R1209_U35 P3_REG1_REG_13__SCAN_IN ; P3_R1209_U153
g24474 nand P3_R1209_U153 P3_R1209_U100 ; P3_R1209_U154
g24475 nand P3_U3427 P3_R1209_U34 ; P3_R1209_U155
g24476 not P3_R1209_U99 ; P3_R1209_U156
g24477 nand P3_R1209_U37 P3_REG1_REG_14__SCAN_IN ; P3_R1209_U157
g24478 nand P3_R1209_U157 P3_R1209_U99 ; P3_R1209_U158
g24479 nand P3_U3430 P3_R1209_U36 ; P3_R1209_U159
g24480 not P3_R1209_U38 ; P3_R1209_U160
g24481 nand P3_R1209_U160 P3_REG1_REG_15__SCAN_IN ; P3_R1209_U161
g24482 nand P3_U3433 P3_R1209_U161 ; P3_R1209_U162
g24483 nand P3_R1209_U38 P3_R1209_U39 ; P3_R1209_U163
g24484 not P3_R1209_U98 ; P3_R1209_U164
g24485 nand P3_R1209_U42 P3_REG1_REG_16__SCAN_IN ; P3_R1209_U165
g24486 nand P3_R1209_U165 P3_R1209_U98 ; P3_R1209_U166
g24487 nand P3_U3436 P3_R1209_U41 ; P3_R1209_U167
g24488 not P3_R1209_U97 ; P3_R1209_U168
g24489 nand P3_R1209_U44 P3_REG1_REG_17__SCAN_IN ; P3_R1209_U169
g24490 nand P3_R1209_U169 P3_R1209_U97 ; P3_R1209_U170
g24491 nand P3_U3439 P3_R1209_U43 ; P3_R1209_U171
g24492 not P3_R1209_U47 ; P3_R1209_U172
g24493 nand P3_U3442 P3_R1209_U45 ; P3_R1209_U173
g24494 nand P3_R1209_U172 P3_R1209_U173 ; P3_R1209_U174
g24495 nand P3_R1209_U46 P3_REG1_REG_18__SCAN_IN ; P3_R1209_U175
g24496 nand P3_R1209_U77 P3_R1209_U174 ; P3_R1209_U176
g24497 nand P3_R1209_U46 P3_REG1_REG_18__SCAN_IN ; P3_R1209_U177
g24498 nand P3_R1209_U177 P3_R1209_U47 ; P3_R1209_U178
g24499 nand P3_U3442 P3_R1209_U45 ; P3_R1209_U179
g24500 nand P3_R1209_U76 P3_R1209_U178 ; P3_R1209_U180
g24501 nand P3_U3386 P3_R1209_U8 ; P3_R1209_U181
g24502 nand P3_R1209_U27 P3_REG1_REG_9__SCAN_IN ; P3_R1209_U182
g24503 nand P3_U3415 P3_R1209_U26 ; P3_R1209_U183
g24504 not P3_R1209_U67 ; P3_R1209_U184
g24505 nand P3_R1209_U136 P3_R1209_U184 ; P3_R1209_U185
g24506 nand P3_R1209_U67 P3_R1209_U87 ; P3_R1209_U186
g24507 nand P3_R1209_U25 P3_REG1_REG_8__SCAN_IN ; P3_R1209_U187
g24508 nand P3_U3412 P3_R1209_U24 ; P3_R1209_U188
g24509 not P3_R1209_U68 ; P3_R1209_U189
g24510 nand P3_R1209_U132 P3_R1209_U189 ; P3_R1209_U190
g24511 nand P3_R1209_U68 P3_R1209_U88 ; P3_R1209_U191
g24512 nand P3_R1209_U23 P3_REG1_REG_7__SCAN_IN ; P3_R1209_U192
g24513 nand P3_U3409 P3_R1209_U22 ; P3_R1209_U193
g24514 not P3_R1209_U69 ; P3_R1209_U194
g24515 nand P3_R1209_U128 P3_R1209_U194 ; P3_R1209_U195
g24516 nand P3_R1209_U69 P3_R1209_U89 ; P3_R1209_U196
g24517 nand P3_R1209_U21 P3_REG1_REG_6__SCAN_IN ; P3_R1209_U197
g24518 nand P3_U3406 P3_R1209_U20 ; P3_R1209_U198
g24519 not P3_R1209_U70 ; P3_R1209_U199
g24520 nand P3_R1209_U124 P3_R1209_U199 ; P3_R1209_U200
g24521 nand P3_R1209_U70 P3_R1209_U90 ; P3_R1209_U201
g24522 nand P3_R1209_U19 P3_REG1_REG_5__SCAN_IN ; P3_R1209_U202
g24523 nand P3_U3403 P3_R1209_U18 ; P3_R1209_U203
g24524 not P3_R1209_U71 ; P3_R1209_U204
g24525 nand P3_R1209_U120 P3_R1209_U204 ; P3_R1209_U205
g24526 nand P3_R1209_U71 P3_R1209_U91 ; P3_R1209_U206
g24527 nand P3_R1209_U17 P3_REG1_REG_4__SCAN_IN ; P3_R1209_U207
g24528 nand P3_U3400 P3_R1209_U16 ; P3_R1209_U208
g24529 not P3_R1209_U72 ; P3_R1209_U209
g24530 nand P3_R1209_U116 P3_R1209_U209 ; P3_R1209_U210
g24531 nand P3_R1209_U72 P3_R1209_U92 ; P3_R1209_U211
g24532 nand P3_R1209_U15 P3_REG1_REG_3__SCAN_IN ; P3_R1209_U212
g24533 nand P3_U3397 P3_R1209_U14 ; P3_R1209_U213
g24534 not P3_R1209_U73 ; P3_R1209_U214
g24535 nand P3_R1209_U112 P3_R1209_U214 ; P3_R1209_U215
g24536 nand P3_R1209_U73 P3_R1209_U93 ; P3_R1209_U216
g24537 nand P3_R1209_U13 P3_REG1_REG_2__SCAN_IN ; P3_R1209_U217
g24538 nand P3_U3394 P3_R1209_U12 ; P3_R1209_U218
g24539 not P3_R1209_U74 ; P3_R1209_U219
g24540 nand P3_R1209_U108 P3_R1209_U219 ; P3_R1209_U220
g24541 nand P3_R1209_U74 P3_R1209_U94 ; P3_R1209_U221
g24542 nand P3_R1209_U104 P3_R1209_U10 ; P3_R1209_U222
g24543 nand P3_R1209_U9 P3_REG1_REG_1__SCAN_IN ; P3_R1209_U223
g24544 not P3_R1209_U75 ; P3_R1209_U224
g24545 nand P3_R1209_U224 P3_U3391 ; P3_R1209_U225
g24546 nand P3_R1209_U75 P3_R1209_U11 ; P3_R1209_U226
g24547 nand P3_R1209_U96 P3_REG1_REG_19__SCAN_IN ; P3_R1209_U227
g24548 nand P3_U3379 P3_R1209_U95 ; P3_R1209_U228
g24549 nand P3_R1209_U96 P3_REG1_REG_19__SCAN_IN ; P3_R1209_U229
g24550 nand P3_U3379 P3_R1209_U95 ; P3_R1209_U230
g24551 nand P3_R1209_U230 P3_R1209_U229 ; P3_R1209_U231
g24552 nand P3_R1209_U46 P3_REG1_REG_18__SCAN_IN ; P3_R1209_U232
g24553 nand P3_U3442 P3_R1209_U45 ; P3_R1209_U233
g24554 not P3_R1209_U78 ; P3_R1209_U234
g24555 nand P3_R1209_U234 P3_R1209_U172 ; P3_R1209_U235
g24556 nand P3_R1209_U78 P3_R1209_U47 ; P3_R1209_U236
g24557 nand P3_R1209_U44 P3_REG1_REG_17__SCAN_IN ; P3_R1209_U237
g24558 nand P3_U3439 P3_R1209_U43 ; P3_R1209_U238
g24559 not P3_R1209_U79 ; P3_R1209_U239
g24560 nand P3_R1209_U168 P3_R1209_U239 ; P3_R1209_U240
g24561 nand P3_R1209_U79 P3_R1209_U97 ; P3_R1209_U241
g24562 nand P3_R1209_U42 P3_REG1_REG_16__SCAN_IN ; P3_R1209_U242
g24563 nand P3_U3436 P3_R1209_U41 ; P3_R1209_U243
g24564 not P3_R1209_U80 ; P3_R1209_U244
g24565 nand P3_R1209_U164 P3_R1209_U244 ; P3_R1209_U245
g24566 nand P3_R1209_U80 P3_R1209_U98 ; P3_R1209_U246
g24567 nand P3_U3433 P3_R1209_U39 ; P3_R1209_U247
g24568 nand P3_R1209_U40 P3_REG1_REG_15__SCAN_IN ; P3_R1209_U248
g24569 not P3_R1209_U81 ; P3_R1209_U249
g24570 nand P3_R1209_U249 P3_R1209_U160 ; P3_R1209_U250
g24571 nand P3_R1209_U81 P3_R1209_U38 ; P3_R1209_U251
g24572 nand P3_R1209_U37 P3_REG1_REG_14__SCAN_IN ; P3_R1209_U252
g24573 nand P3_U3430 P3_R1209_U36 ; P3_R1209_U253
g24574 not P3_R1209_U82 ; P3_R1209_U254
g24575 nand P3_R1209_U156 P3_R1209_U254 ; P3_R1209_U255
g24576 nand P3_R1209_U82 P3_R1209_U99 ; P3_R1209_U256
g24577 nand P3_R1209_U35 P3_REG1_REG_13__SCAN_IN ; P3_R1209_U257
g24578 nand P3_U3427 P3_R1209_U34 ; P3_R1209_U258
g24579 not P3_R1209_U83 ; P3_R1209_U259
g24580 nand P3_R1209_U152 P3_R1209_U259 ; P3_R1209_U260
g24581 nand P3_R1209_U83 P3_R1209_U100 ; P3_R1209_U261
g24582 nand P3_R1209_U33 P3_REG1_REG_12__SCAN_IN ; P3_R1209_U262
g24583 nand P3_U3424 P3_R1209_U32 ; P3_R1209_U263
g24584 not P3_R1209_U84 ; P3_R1209_U264
g24585 nand P3_R1209_U148 P3_R1209_U264 ; P3_R1209_U265
g24586 nand P3_R1209_U84 P3_R1209_U101 ; P3_R1209_U266
g24587 nand P3_R1209_U31 P3_REG1_REG_11__SCAN_IN ; P3_R1209_U267
g24588 nand P3_U3421 P3_R1209_U30 ; P3_R1209_U268
g24589 not P3_R1209_U85 ; P3_R1209_U269
g24590 nand P3_R1209_U144 P3_R1209_U269 ; P3_R1209_U270
g24591 nand P3_R1209_U85 P3_R1209_U102 ; P3_R1209_U271
g24592 nand P3_R1209_U29 P3_REG1_REG_10__SCAN_IN ; P3_R1209_U272
g24593 nand P3_U3418 P3_R1209_U28 ; P3_R1209_U273
g24594 not P3_R1209_U86 ; P3_R1209_U274
g24595 nand P3_R1209_U140 P3_R1209_U274 ; P3_R1209_U275
g24596 nand P3_R1209_U86 P3_R1209_U103 ; P3_R1209_U276
g24597 not P3_U3058 ; P3_R1300_U6
g24598 not P3_U3055 ; P3_R1300_U7
g24599 and P3_R1300_U10 P3_R1300_U9 ; P3_R1300_U8
g24600 nand P3_U3055 P3_R1300_U6 ; P3_R1300_U9
g24601 nand P3_U3058 P3_R1300_U7 ; P3_R1300_U10
g24602 and P3_R1200_U210 P3_R1200_U209 ; P3_R1200_U6
g24603 and P3_R1200_U189 P3_R1200_U245 ; P3_R1200_U7
g24604 and P3_R1200_U247 P3_R1200_U246 ; P3_R1200_U8
g24605 and P3_R1200_U190 P3_R1200_U262 ; P3_R1200_U9
g24606 and P3_R1200_U264 P3_R1200_U263 ; P3_R1200_U10
g24607 and P3_R1200_U191 P3_R1200_U286 ; P3_R1200_U11
g24608 and P3_R1200_U288 P3_R1200_U287 ; P3_R1200_U12
g24609 and P3_R1200_U208 P3_R1200_U194 P3_R1200_U213 ; P3_R1200_U13
g24610 and P3_R1200_U218 P3_R1200_U195 ; P3_R1200_U14
g24611 and P3_R1200_U392 P3_R1200_U391 ; P3_R1200_U15
g24612 nand P3_R1200_U342 P3_R1200_U345 ; P3_R1200_U16
g24613 nand P3_R1200_U331 P3_R1200_U334 ; P3_R1200_U17
g24614 nand P3_R1200_U320 P3_R1200_U323 ; P3_R1200_U18
g24615 nand P3_R1200_U312 P3_R1200_U314 ; P3_R1200_U19
g24616 nand P3_R1200_U162 P3_R1200_U183 P3_R1200_U351 ; P3_R1200_U20
g24617 nand P3_R1200_U241 P3_R1200_U243 ; P3_R1200_U21
g24618 nand P3_R1200_U233 P3_R1200_U236 ; P3_R1200_U22
g24619 nand P3_R1200_U225 P3_R1200_U227 ; P3_R1200_U23
g24620 nand P3_R1200_U172 P3_R1200_U348 ; P3_R1200_U24
g24621 not P3_U3069 ; P3_R1200_U25
g24622 nand P3_U3069 P3_R1200_U39 ; P3_R1200_U26
g24623 not P3_U3083 ; P3_R1200_U27
g24624 not P3_U3413 ; P3_R1200_U28
g24625 not P3_U3395 ; P3_R1200_U29
g24626 not P3_U3387 ; P3_R1200_U30
g24627 not P3_U3077 ; P3_R1200_U31
g24628 not P3_U3398 ; P3_R1200_U32
g24629 not P3_U3067 ; P3_R1200_U33
g24630 nand P3_U3067 P3_R1200_U29 ; P3_R1200_U34
g24631 not P3_U3063 ; P3_R1200_U35
g24632 not P3_U3404 ; P3_R1200_U36
g24633 not P3_U3407 ; P3_R1200_U37
g24634 not P3_U3401 ; P3_R1200_U38
g24635 not P3_U3410 ; P3_R1200_U39
g24636 not P3_U3070 ; P3_R1200_U40
g24637 not P3_U3066 ; P3_R1200_U41
g24638 not P3_U3059 ; P3_R1200_U42
g24639 nand P3_U3059 P3_R1200_U38 ; P3_R1200_U43
g24640 nand P3_R1200_U214 P3_R1200_U212 ; P3_R1200_U44
g24641 not P3_U3416 ; P3_R1200_U45
g24642 not P3_U3082 ; P3_R1200_U46
g24643 nand P3_R1200_U44 P3_R1200_U215 ; P3_R1200_U47
g24644 nand P3_R1200_U43 P3_R1200_U229 ; P3_R1200_U48
g24645 nand P3_R1200_U201 P3_R1200_U185 P3_R1200_U349 ; P3_R1200_U49
g24646 not P3_U3901 ; P3_R1200_U50
g24647 not P3_U3422 ; P3_R1200_U51
g24648 not P3_U3419 ; P3_R1200_U52
g24649 not P3_U3062 ; P3_R1200_U53
g24650 not P3_U3061 ; P3_R1200_U54
g24651 nand P3_U3082 P3_R1200_U45 ; P3_R1200_U55
g24652 not P3_U3425 ; P3_R1200_U56
g24653 not P3_U3071 ; P3_R1200_U57
g24654 not P3_U3428 ; P3_R1200_U58
g24655 not P3_U3079 ; P3_R1200_U59
g24656 not P3_U3437 ; P3_R1200_U60
g24657 not P3_U3434 ; P3_R1200_U61
g24658 not P3_U3431 ; P3_R1200_U62
g24659 not P3_U3072 ; P3_R1200_U63
g24660 not P3_U3073 ; P3_R1200_U64
g24661 not P3_U3078 ; P3_R1200_U65
g24662 nand P3_U3078 P3_R1200_U62 ; P3_R1200_U66
g24663 not P3_U3440 ; P3_R1200_U67
g24664 not P3_U3068 ; P3_R1200_U68
g24665 not P3_U3081 ; P3_R1200_U69
g24666 not P3_U3445 ; P3_R1200_U70
g24667 not P3_U3080 ; P3_R1200_U71
g24668 not P3_U3907 ; P3_R1200_U72
g24669 not P3_U3075 ; P3_R1200_U73
g24670 not P3_U3904 ; P3_R1200_U74
g24671 not P3_U3905 ; P3_R1200_U75
g24672 not P3_U3906 ; P3_R1200_U76
g24673 not P3_U3065 ; P3_R1200_U77
g24674 not P3_U3060 ; P3_R1200_U78
g24675 not P3_U3074 ; P3_R1200_U79
g24676 nand P3_U3074 P3_R1200_U76 ; P3_R1200_U80
g24677 not P3_U3903 ; P3_R1200_U81
g24678 not P3_U3064 ; P3_R1200_U82
g24679 not P3_U3902 ; P3_R1200_U83
g24680 not P3_U3057 ; P3_R1200_U84
g24681 not P3_U3900 ; P3_R1200_U85
g24682 not P3_U3056 ; P3_R1200_U86
g24683 nand P3_U3056 P3_R1200_U50 ; P3_R1200_U87
g24684 not P3_U3052 ; P3_R1200_U88
g24685 not P3_U3899 ; P3_R1200_U89
g24686 not P3_U3053 ; P3_R1200_U90
g24687 nand P3_R1200_U302 P3_R1200_U301 ; P3_R1200_U91
g24688 nand P3_R1200_U80 P3_R1200_U316 ; P3_R1200_U92
g24689 nand P3_R1200_U66 P3_R1200_U327 ; P3_R1200_U93
g24690 nand P3_R1200_U55 P3_R1200_U338 ; P3_R1200_U94
g24691 not P3_U3076 ; P3_R1200_U95
g24692 nand P3_R1200_U402 P3_R1200_U401 ; P3_R1200_U96
g24693 nand P3_R1200_U416 P3_R1200_U415 ; P3_R1200_U97
g24694 nand P3_R1200_U421 P3_R1200_U420 ; P3_R1200_U98
g24695 nand P3_R1200_U437 P3_R1200_U436 ; P3_R1200_U99
g24696 nand P3_R1200_U442 P3_R1200_U441 ; P3_R1200_U100
g24697 nand P3_R1200_U447 P3_R1200_U446 ; P3_R1200_U101
g24698 nand P3_R1200_U452 P3_R1200_U451 ; P3_R1200_U102
g24699 nand P3_R1200_U457 P3_R1200_U456 ; P3_R1200_U103
g24700 nand P3_R1200_U473 P3_R1200_U472 ; P3_R1200_U104
g24701 nand P3_R1200_U478 P3_R1200_U477 ; P3_R1200_U105
g24702 nand P3_R1200_U361 P3_R1200_U360 ; P3_R1200_U106
g24703 nand P3_R1200_U370 P3_R1200_U369 ; P3_R1200_U107
g24704 nand P3_R1200_U377 P3_R1200_U376 ; P3_R1200_U108
g24705 nand P3_R1200_U381 P3_R1200_U380 ; P3_R1200_U109
g24706 nand P3_R1200_U390 P3_R1200_U389 ; P3_R1200_U110
g24707 nand P3_R1200_U411 P3_R1200_U410 ; P3_R1200_U111
g24708 nand P3_R1200_U428 P3_R1200_U427 ; P3_R1200_U112
g24709 nand P3_R1200_U432 P3_R1200_U431 ; P3_R1200_U113
g24710 nand P3_R1200_U464 P3_R1200_U463 ; P3_R1200_U114
g24711 nand P3_R1200_U468 P3_R1200_U467 ; P3_R1200_U115
g24712 nand P3_R1200_U485 P3_R1200_U484 ; P3_R1200_U116
g24713 and P3_R1200_U352 P3_R1200_U193 ; P3_R1200_U117
g24714 and P3_R1200_U205 P3_R1200_U206 ; P3_R1200_U118
g24715 and P3_R1200_U14 P3_R1200_U13 ; P3_R1200_U119
g24716 and P3_R1200_U357 P3_R1200_U354 ; P3_R1200_U120
g24717 and P3_R1200_U363 P3_R1200_U362 P3_R1200_U26 ; P3_R1200_U121
g24718 and P3_R1200_U366 P3_R1200_U195 ; P3_R1200_U122
g24719 and P3_R1200_U235 P3_R1200_U6 ; P3_R1200_U123
g24720 and P3_R1200_U373 P3_R1200_U194 ; P3_R1200_U124
g24721 and P3_R1200_U383 P3_R1200_U382 P3_R1200_U34 ; P3_R1200_U125
g24722 and P3_R1200_U386 P3_R1200_U193 ; P3_R1200_U126
g24723 and P3_R1200_U222 P3_R1200_U7 ; P3_R1200_U127
g24724 and P3_R1200_U267 P3_R1200_U9 ; P3_R1200_U128
g24725 and P3_R1200_U291 P3_R1200_U11 ; P3_R1200_U129
g24726 and P3_R1200_U355 P3_R1200_U192 ; P3_R1200_U130
g24727 and P3_R1200_U306 P3_R1200_U307 ; P3_R1200_U131
g24728 and P3_R1200_U309 P3_R1200_U395 ; P3_R1200_U132
g24729 and P3_R1200_U306 P3_R1200_U307 ; P3_R1200_U133
g24730 and P3_R1200_U15 P3_R1200_U310 ; P3_R1200_U134
g24731 nand P3_R1200_U399 P3_R1200_U398 ; P3_R1200_U135
g24732 and P3_R1200_U404 P3_R1200_U403 P3_R1200_U87 ; P3_R1200_U136
g24733 and P3_R1200_U407 P3_R1200_U192 ; P3_R1200_U137
g24734 nand P3_R1200_U413 P3_R1200_U412 ; P3_R1200_U138
g24735 nand P3_R1200_U418 P3_R1200_U417 ; P3_R1200_U139
g24736 and P3_R1200_U322 P3_R1200_U12 ; P3_R1200_U140
g24737 and P3_R1200_U424 P3_R1200_U191 ; P3_R1200_U141
g24738 nand P3_R1200_U434 P3_R1200_U433 ; P3_R1200_U142
g24739 nand P3_R1200_U439 P3_R1200_U438 ; P3_R1200_U143
g24740 nand P3_R1200_U444 P3_R1200_U443 ; P3_R1200_U144
g24741 nand P3_R1200_U449 P3_R1200_U448 ; P3_R1200_U145
g24742 nand P3_R1200_U454 P3_R1200_U453 ; P3_R1200_U146
g24743 and P3_R1200_U333 P3_R1200_U10 ; P3_R1200_U147
g24744 and P3_R1200_U460 P3_R1200_U190 ; P3_R1200_U148
g24745 nand P3_R1200_U470 P3_R1200_U469 ; P3_R1200_U149
g24746 nand P3_R1200_U475 P3_R1200_U474 ; P3_R1200_U150
g24747 and P3_R1200_U344 P3_R1200_U8 ; P3_R1200_U151
g24748 and P3_R1200_U481 P3_R1200_U189 ; P3_R1200_U152
g24749 and P3_R1200_U359 P3_R1200_U358 ; P3_R1200_U153
g24750 nand P3_R1200_U120 P3_R1200_U356 ; P3_R1200_U154
g24751 and P3_R1200_U368 P3_R1200_U367 ; P3_R1200_U155
g24752 and P3_R1200_U375 P3_R1200_U374 ; P3_R1200_U156
g24753 and P3_R1200_U379 P3_R1200_U378 ; P3_R1200_U157
g24754 nand P3_R1200_U118 P3_R1200_U203 ; P3_R1200_U158
g24755 and P3_R1200_U388 P3_R1200_U387 ; P3_R1200_U159
g24756 not P3_U3908 ; P3_R1200_U160
g24757 not P3_U3054 ; P3_R1200_U161
g24758 and P3_R1200_U397 P3_R1200_U396 ; P3_R1200_U162
g24759 nand P3_R1200_U131 P3_R1200_U304 ; P3_R1200_U163
g24760 and P3_R1200_U409 P3_R1200_U408 ; P3_R1200_U164
g24761 nand P3_R1200_U298 P3_R1200_U297 ; P3_R1200_U165
g24762 nand P3_R1200_U294 P3_R1200_U293 ; P3_R1200_U166
g24763 and P3_R1200_U426 P3_R1200_U425 ; P3_R1200_U167
g24764 and P3_R1200_U430 P3_R1200_U429 ; P3_R1200_U168
g24765 nand P3_R1200_U284 P3_R1200_U283 ; P3_R1200_U169
g24766 nand P3_R1200_U280 P3_R1200_U279 ; P3_R1200_U170
g24767 not P3_U3392 ; P3_R1200_U171
g24768 nand P3_U3387 P3_R1200_U95 ; P3_R1200_U172
g24769 nand P3_R1200_U276 P3_R1200_U184 P3_R1200_U350 ; P3_R1200_U173
g24770 not P3_U3443 ; P3_R1200_U174
g24771 nand P3_R1200_U274 P3_R1200_U273 ; P3_R1200_U175
g24772 nand P3_R1200_U270 P3_R1200_U269 ; P3_R1200_U176
g24773 and P3_R1200_U462 P3_R1200_U461 ; P3_R1200_U177
g24774 and P3_R1200_U466 P3_R1200_U465 ; P3_R1200_U178
g24775 nand P3_R1200_U260 P3_R1200_U259 ; P3_R1200_U179
g24776 nand P3_R1200_U256 P3_R1200_U255 ; P3_R1200_U180
g24777 nand P3_R1200_U252 P3_R1200_U251 ; P3_R1200_U181
g24778 and P3_R1200_U483 P3_R1200_U482 ; P3_R1200_U182
g24779 nand P3_R1200_U132 P3_R1200_U163 ; P3_R1200_U183
g24780 nand P3_R1200_U175 P3_R1200_U174 ; P3_R1200_U184
g24781 nand P3_R1200_U172 P3_R1200_U171 ; P3_R1200_U185
g24782 not P3_R1200_U87 ; P3_R1200_U186
g24783 not P3_R1200_U34 ; P3_R1200_U187
g24784 not P3_R1200_U26 ; P3_R1200_U188
g24785 nand P3_U3419 P3_R1200_U54 ; P3_R1200_U189
g24786 nand P3_U3434 P3_R1200_U64 ; P3_R1200_U190
g24787 nand P3_U3905 P3_R1200_U78 ; P3_R1200_U191
g24788 nand P3_U3901 P3_R1200_U86 ; P3_R1200_U192
g24789 nand P3_U3395 P3_R1200_U33 ; P3_R1200_U193
g24790 nand P3_U3404 P3_R1200_U41 ; P3_R1200_U194
g24791 nand P3_U3410 P3_R1200_U25 ; P3_R1200_U195
g24792 not P3_R1200_U66 ; P3_R1200_U196
g24793 not P3_R1200_U80 ; P3_R1200_U197
g24794 not P3_R1200_U43 ; P3_R1200_U198
g24795 not P3_R1200_U55 ; P3_R1200_U199
g24796 not P3_R1200_U172 ; P3_R1200_U200
g24797 nand P3_U3077 P3_R1200_U172 ; P3_R1200_U201
g24798 not P3_R1200_U49 ; P3_R1200_U202
g24799 nand P3_R1200_U117 P3_R1200_U49 ; P3_R1200_U203
g24800 nand P3_R1200_U35 P3_R1200_U34 ; P3_R1200_U204
g24801 nand P3_R1200_U204 P3_R1200_U32 ; P3_R1200_U205
g24802 nand P3_U3063 P3_R1200_U187 ; P3_R1200_U206
g24803 not P3_R1200_U158 ; P3_R1200_U207
g24804 nand P3_U3407 P3_R1200_U40 ; P3_R1200_U208
g24805 nand P3_U3070 P3_R1200_U37 ; P3_R1200_U209
g24806 nand P3_U3066 P3_R1200_U36 ; P3_R1200_U210
g24807 nand P3_R1200_U198 P3_R1200_U194 ; P3_R1200_U211
g24808 nand P3_R1200_U6 P3_R1200_U211 ; P3_R1200_U212
g24809 nand P3_U3401 P3_R1200_U42 ; P3_R1200_U213
g24810 nand P3_U3407 P3_R1200_U40 ; P3_R1200_U214
g24811 nand P3_R1200_U13 P3_R1200_U158 ; P3_R1200_U215
g24812 not P3_R1200_U44 ; P3_R1200_U216
g24813 not P3_R1200_U47 ; P3_R1200_U217
g24814 nand P3_U3413 P3_R1200_U27 ; P3_R1200_U218
g24815 nand P3_R1200_U27 P3_R1200_U26 ; P3_R1200_U219
g24816 nand P3_U3083 P3_R1200_U188 ; P3_R1200_U220
g24817 not P3_R1200_U154 ; P3_R1200_U221
g24818 nand P3_U3416 P3_R1200_U46 ; P3_R1200_U222
g24819 nand P3_R1200_U222 P3_R1200_U55 ; P3_R1200_U223
g24820 nand P3_R1200_U217 P3_R1200_U26 ; P3_R1200_U224
g24821 nand P3_R1200_U122 P3_R1200_U224 ; P3_R1200_U225
g24822 nand P3_R1200_U47 P3_R1200_U195 ; P3_R1200_U226
g24823 nand P3_R1200_U121 P3_R1200_U226 ; P3_R1200_U227
g24824 nand P3_R1200_U26 P3_R1200_U195 ; P3_R1200_U228
g24825 nand P3_R1200_U213 P3_R1200_U158 ; P3_R1200_U229
g24826 not P3_R1200_U48 ; P3_R1200_U230
g24827 nand P3_U3066 P3_R1200_U36 ; P3_R1200_U231
g24828 nand P3_R1200_U230 P3_R1200_U231 ; P3_R1200_U232
g24829 nand P3_R1200_U124 P3_R1200_U232 ; P3_R1200_U233
g24830 nand P3_R1200_U48 P3_R1200_U194 ; P3_R1200_U234
g24831 nand P3_U3407 P3_R1200_U40 ; P3_R1200_U235
g24832 nand P3_R1200_U123 P3_R1200_U234 ; P3_R1200_U236
g24833 nand P3_U3066 P3_R1200_U36 ; P3_R1200_U237
g24834 nand P3_R1200_U194 P3_R1200_U237 ; P3_R1200_U238
g24835 nand P3_R1200_U213 P3_R1200_U43 ; P3_R1200_U239
g24836 nand P3_R1200_U202 P3_R1200_U34 ; P3_R1200_U240
g24837 nand P3_R1200_U126 P3_R1200_U240 ; P3_R1200_U241
g24838 nand P3_R1200_U49 P3_R1200_U193 ; P3_R1200_U242
g24839 nand P3_R1200_U125 P3_R1200_U242 ; P3_R1200_U243
g24840 nand P3_R1200_U193 P3_R1200_U34 ; P3_R1200_U244
g24841 nand P3_U3422 P3_R1200_U53 ; P3_R1200_U245
g24842 nand P3_U3062 P3_R1200_U51 ; P3_R1200_U246
g24843 nand P3_U3061 P3_R1200_U52 ; P3_R1200_U247
g24844 nand P3_R1200_U199 P3_R1200_U7 ; P3_R1200_U248
g24845 nand P3_R1200_U8 P3_R1200_U248 ; P3_R1200_U249
g24846 nand P3_U3422 P3_R1200_U53 ; P3_R1200_U250
g24847 nand P3_R1200_U127 P3_R1200_U154 ; P3_R1200_U251
g24848 nand P3_R1200_U250 P3_R1200_U249 ; P3_R1200_U252
g24849 not P3_R1200_U181 ; P3_R1200_U253
g24850 nand P3_U3425 P3_R1200_U57 ; P3_R1200_U254
g24851 nand P3_R1200_U254 P3_R1200_U181 ; P3_R1200_U255
g24852 nand P3_U3071 P3_R1200_U56 ; P3_R1200_U256
g24853 not P3_R1200_U180 ; P3_R1200_U257
g24854 nand P3_U3428 P3_R1200_U59 ; P3_R1200_U258
g24855 nand P3_R1200_U258 P3_R1200_U180 ; P3_R1200_U259
g24856 nand P3_U3079 P3_R1200_U58 ; P3_R1200_U260
g24857 not P3_R1200_U179 ; P3_R1200_U261
g24858 nand P3_U3437 P3_R1200_U63 ; P3_R1200_U262
g24859 nand P3_U3072 P3_R1200_U60 ; P3_R1200_U263
g24860 nand P3_U3073 P3_R1200_U61 ; P3_R1200_U264
g24861 nand P3_R1200_U196 P3_R1200_U9 ; P3_R1200_U265
g24862 nand P3_R1200_U10 P3_R1200_U265 ; P3_R1200_U266
g24863 nand P3_U3431 P3_R1200_U65 ; P3_R1200_U267
g24864 nand P3_U3437 P3_R1200_U63 ; P3_R1200_U268
g24865 nand P3_R1200_U128 P3_R1200_U179 ; P3_R1200_U269
g24866 nand P3_R1200_U268 P3_R1200_U266 ; P3_R1200_U270
g24867 not P3_R1200_U176 ; P3_R1200_U271
g24868 nand P3_U3440 P3_R1200_U68 ; P3_R1200_U272
g24869 nand P3_R1200_U272 P3_R1200_U176 ; P3_R1200_U273
g24870 nand P3_U3068 P3_R1200_U67 ; P3_R1200_U274
g24871 not P3_R1200_U175 ; P3_R1200_U275
g24872 nand P3_U3081 P3_R1200_U175 ; P3_R1200_U276
g24873 not P3_R1200_U173 ; P3_R1200_U277
g24874 nand P3_U3445 P3_R1200_U71 ; P3_R1200_U278
g24875 nand P3_R1200_U278 P3_R1200_U173 ; P3_R1200_U279
g24876 nand P3_U3080 P3_R1200_U70 ; P3_R1200_U280
g24877 not P3_R1200_U170 ; P3_R1200_U281
g24878 nand P3_U3907 P3_R1200_U73 ; P3_R1200_U282
g24879 nand P3_R1200_U282 P3_R1200_U170 ; P3_R1200_U283
g24880 nand P3_U3075 P3_R1200_U72 ; P3_R1200_U284
g24881 not P3_R1200_U169 ; P3_R1200_U285
g24882 nand P3_U3904 P3_R1200_U77 ; P3_R1200_U286
g24883 nand P3_U3065 P3_R1200_U74 ; P3_R1200_U287
g24884 nand P3_U3060 P3_R1200_U75 ; P3_R1200_U288
g24885 nand P3_R1200_U197 P3_R1200_U11 ; P3_R1200_U289
g24886 nand P3_R1200_U12 P3_R1200_U289 ; P3_R1200_U290
g24887 nand P3_U3906 P3_R1200_U79 ; P3_R1200_U291
g24888 nand P3_U3904 P3_R1200_U77 ; P3_R1200_U292
g24889 nand P3_R1200_U129 P3_R1200_U169 ; P3_R1200_U293
g24890 nand P3_R1200_U292 P3_R1200_U290 ; P3_R1200_U294
g24891 not P3_R1200_U166 ; P3_R1200_U295
g24892 nand P3_U3903 P3_R1200_U82 ; P3_R1200_U296
g24893 nand P3_R1200_U296 P3_R1200_U166 ; P3_R1200_U297
g24894 nand P3_U3064 P3_R1200_U81 ; P3_R1200_U298
g24895 not P3_R1200_U165 ; P3_R1200_U299
g24896 nand P3_U3902 P3_R1200_U84 ; P3_R1200_U300
g24897 nand P3_R1200_U300 P3_R1200_U165 ; P3_R1200_U301
g24898 nand P3_U3057 P3_R1200_U83 ; P3_R1200_U302
g24899 not P3_R1200_U91 ; P3_R1200_U303
g24900 nand P3_R1200_U130 P3_R1200_U91 ; P3_R1200_U304
g24901 nand P3_R1200_U88 P3_R1200_U87 ; P3_R1200_U305
g24902 nand P3_R1200_U305 P3_R1200_U85 ; P3_R1200_U306
g24903 nand P3_U3052 P3_R1200_U186 ; P3_R1200_U307
g24904 not P3_R1200_U163 ; P3_R1200_U308
g24905 nand P3_U3899 P3_R1200_U90 ; P3_R1200_U309
g24906 nand P3_U3053 P3_R1200_U89 ; P3_R1200_U310
g24907 nand P3_R1200_U303 P3_R1200_U87 ; P3_R1200_U311
g24908 nand P3_R1200_U137 P3_R1200_U311 ; P3_R1200_U312
g24909 nand P3_R1200_U91 P3_R1200_U192 ; P3_R1200_U313
g24910 nand P3_R1200_U136 P3_R1200_U313 ; P3_R1200_U314
g24911 nand P3_R1200_U192 P3_R1200_U87 ; P3_R1200_U315
g24912 nand P3_R1200_U291 P3_R1200_U169 ; P3_R1200_U316
g24913 not P3_R1200_U92 ; P3_R1200_U317
g24914 nand P3_U3060 P3_R1200_U75 ; P3_R1200_U318
g24915 nand P3_R1200_U317 P3_R1200_U318 ; P3_R1200_U319
g24916 nand P3_R1200_U141 P3_R1200_U319 ; P3_R1200_U320
g24917 nand P3_R1200_U92 P3_R1200_U191 ; P3_R1200_U321
g24918 nand P3_U3904 P3_R1200_U77 ; P3_R1200_U322
g24919 nand P3_R1200_U140 P3_R1200_U321 ; P3_R1200_U323
g24920 nand P3_U3060 P3_R1200_U75 ; P3_R1200_U324
g24921 nand P3_R1200_U191 P3_R1200_U324 ; P3_R1200_U325
g24922 nand P3_R1200_U291 P3_R1200_U80 ; P3_R1200_U326
g24923 nand P3_R1200_U267 P3_R1200_U179 ; P3_R1200_U327
g24924 not P3_R1200_U93 ; P3_R1200_U328
g24925 nand P3_U3073 P3_R1200_U61 ; P3_R1200_U329
g24926 nand P3_R1200_U328 P3_R1200_U329 ; P3_R1200_U330
g24927 nand P3_R1200_U148 P3_R1200_U330 ; P3_R1200_U331
g24928 nand P3_R1200_U93 P3_R1200_U190 ; P3_R1200_U332
g24929 nand P3_U3437 P3_R1200_U63 ; P3_R1200_U333
g24930 nand P3_R1200_U147 P3_R1200_U332 ; P3_R1200_U334
g24931 nand P3_U3073 P3_R1200_U61 ; P3_R1200_U335
g24932 nand P3_R1200_U190 P3_R1200_U335 ; P3_R1200_U336
g24933 nand P3_R1200_U267 P3_R1200_U66 ; P3_R1200_U337
g24934 nand P3_R1200_U222 P3_R1200_U154 ; P3_R1200_U338
g24935 not P3_R1200_U94 ; P3_R1200_U339
g24936 nand P3_U3061 P3_R1200_U52 ; P3_R1200_U340
g24937 nand P3_R1200_U339 P3_R1200_U340 ; P3_R1200_U341
g24938 nand P3_R1200_U152 P3_R1200_U341 ; P3_R1200_U342
g24939 nand P3_R1200_U94 P3_R1200_U189 ; P3_R1200_U343
g24940 nand P3_U3422 P3_R1200_U53 ; P3_R1200_U344
g24941 nand P3_R1200_U151 P3_R1200_U343 ; P3_R1200_U345
g24942 nand P3_U3061 P3_R1200_U52 ; P3_R1200_U346
g24943 nand P3_R1200_U189 P3_R1200_U346 ; P3_R1200_U347
g24944 nand P3_U3076 P3_R1200_U30 ; P3_R1200_U348
g24945 nand P3_U3077 P3_R1200_U171 ; P3_R1200_U349
g24946 nand P3_U3081 P3_R1200_U174 ; P3_R1200_U350
g24947 nand P3_R1200_U133 P3_R1200_U304 P3_R1200_U134 ; P3_R1200_U351
g24948 nand P3_U3398 P3_R1200_U35 ; P3_R1200_U352
g24949 nand P3_U3413 P3_R1200_U220 ; P3_R1200_U353
g24950 nand P3_R1200_U353 P3_R1200_U219 ; P3_R1200_U354
g24951 nand P3_U3900 P3_R1200_U88 ; P3_R1200_U355
g24952 nand P3_R1200_U119 P3_R1200_U158 ; P3_R1200_U356
g24953 nand P3_R1200_U216 P3_R1200_U14 ; P3_R1200_U357
g24954 nand P3_U3416 P3_R1200_U46 ; P3_R1200_U358
g24955 nand P3_U3082 P3_R1200_U45 ; P3_R1200_U359
g24956 nand P3_R1200_U223 P3_R1200_U154 ; P3_R1200_U360
g24957 nand P3_R1200_U221 P3_R1200_U153 ; P3_R1200_U361
g24958 nand P3_U3413 P3_R1200_U27 ; P3_R1200_U362
g24959 nand P3_U3083 P3_R1200_U28 ; P3_R1200_U363
g24960 nand P3_U3413 P3_R1200_U27 ; P3_R1200_U364
g24961 nand P3_U3083 P3_R1200_U28 ; P3_R1200_U365
g24962 nand P3_R1200_U365 P3_R1200_U364 ; P3_R1200_U366
g24963 nand P3_U3410 P3_R1200_U25 ; P3_R1200_U367
g24964 nand P3_U3069 P3_R1200_U39 ; P3_R1200_U368
g24965 nand P3_R1200_U228 P3_R1200_U47 ; P3_R1200_U369
g24966 nand P3_R1200_U155 P3_R1200_U217 ; P3_R1200_U370
g24967 nand P3_U3407 P3_R1200_U40 ; P3_R1200_U371
g24968 nand P3_U3070 P3_R1200_U37 ; P3_R1200_U372
g24969 nand P3_R1200_U372 P3_R1200_U371 ; P3_R1200_U373
g24970 nand P3_U3404 P3_R1200_U41 ; P3_R1200_U374
g24971 nand P3_U3066 P3_R1200_U36 ; P3_R1200_U375
g24972 nand P3_R1200_U238 P3_R1200_U48 ; P3_R1200_U376
g24973 nand P3_R1200_U156 P3_R1200_U230 ; P3_R1200_U377
g24974 nand P3_U3401 P3_R1200_U42 ; P3_R1200_U378
g24975 nand P3_U3059 P3_R1200_U38 ; P3_R1200_U379
g24976 nand P3_R1200_U239 P3_R1200_U158 ; P3_R1200_U380
g24977 nand P3_R1200_U207 P3_R1200_U157 ; P3_R1200_U381
g24978 nand P3_U3398 P3_R1200_U35 ; P3_R1200_U382
g24979 nand P3_U3063 P3_R1200_U32 ; P3_R1200_U383
g24980 nand P3_U3398 P3_R1200_U35 ; P3_R1200_U384
g24981 nand P3_U3063 P3_R1200_U32 ; P3_R1200_U385
g24982 nand P3_R1200_U385 P3_R1200_U384 ; P3_R1200_U386
g24983 nand P3_U3395 P3_R1200_U33 ; P3_R1200_U387
g24984 nand P3_U3067 P3_R1200_U29 ; P3_R1200_U388
g24985 nand P3_R1200_U244 P3_R1200_U49 ; P3_R1200_U389
g24986 nand P3_R1200_U159 P3_R1200_U202 ; P3_R1200_U390
g24987 nand P3_U3908 P3_R1200_U161 ; P3_R1200_U391
g24988 nand P3_U3054 P3_R1200_U160 ; P3_R1200_U392
g24989 nand P3_U3908 P3_R1200_U161 ; P3_R1200_U393
g24990 nand P3_U3054 P3_R1200_U160 ; P3_R1200_U394
g24991 nand P3_R1200_U394 P3_R1200_U393 ; P3_R1200_U395
g24992 nand P3_U3053 P3_R1200_U395 P3_R1200_U89 ; P3_R1200_U396
g24993 nand P3_R1200_U15 P3_R1200_U90 P3_U3899 ; P3_R1200_U397
g24994 nand P3_U3899 P3_R1200_U90 ; P3_R1200_U398
g24995 nand P3_U3053 P3_R1200_U89 ; P3_R1200_U399
g24996 not P3_R1200_U135 ; P3_R1200_U400
g24997 nand P3_R1200_U308 P3_R1200_U400 ; P3_R1200_U401
g24998 nand P3_R1200_U135 P3_R1200_U163 ; P3_R1200_U402
g24999 nand P3_U3900 P3_R1200_U88 ; P3_R1200_U403
g25000 nand P3_U3052 P3_R1200_U85 ; P3_R1200_U404
g25001 nand P3_U3900 P3_R1200_U88 ; P3_R1200_U405
g25002 nand P3_U3052 P3_R1200_U85 ; P3_R1200_U406
g25003 nand P3_R1200_U406 P3_R1200_U405 ; P3_R1200_U407
g25004 nand P3_U3901 P3_R1200_U86 ; P3_R1200_U408
g25005 nand P3_U3056 P3_R1200_U50 ; P3_R1200_U409
g25006 nand P3_R1200_U315 P3_R1200_U91 ; P3_R1200_U410
g25007 nand P3_R1200_U164 P3_R1200_U303 ; P3_R1200_U411
g25008 nand P3_U3902 P3_R1200_U84 ; P3_R1200_U412
g25009 nand P3_U3057 P3_R1200_U83 ; P3_R1200_U413
g25010 not P3_R1200_U138 ; P3_R1200_U414
g25011 nand P3_R1200_U299 P3_R1200_U414 ; P3_R1200_U415
g25012 nand P3_R1200_U138 P3_R1200_U165 ; P3_R1200_U416
g25013 nand P3_U3903 P3_R1200_U82 ; P3_R1200_U417
g25014 nand P3_U3064 P3_R1200_U81 ; P3_R1200_U418
g25015 not P3_R1200_U139 ; P3_R1200_U419
g25016 nand P3_R1200_U295 P3_R1200_U419 ; P3_R1200_U420
g25017 nand P3_R1200_U139 P3_R1200_U166 ; P3_R1200_U421
g25018 nand P3_U3904 P3_R1200_U77 ; P3_R1200_U422
g25019 nand P3_U3065 P3_R1200_U74 ; P3_R1200_U423
g25020 nand P3_R1200_U423 P3_R1200_U422 ; P3_R1200_U424
g25021 nand P3_U3905 P3_R1200_U78 ; P3_R1200_U425
g25022 nand P3_U3060 P3_R1200_U75 ; P3_R1200_U426
g25023 nand P3_R1200_U325 P3_R1200_U92 ; P3_R1200_U427
g25024 nand P3_R1200_U167 P3_R1200_U317 ; P3_R1200_U428
g25025 nand P3_U3906 P3_R1200_U79 ; P3_R1200_U429
g25026 nand P3_U3074 P3_R1200_U76 ; P3_R1200_U430
g25027 nand P3_R1200_U326 P3_R1200_U169 ; P3_R1200_U431
g25028 nand P3_R1200_U285 P3_R1200_U168 ; P3_R1200_U432
g25029 nand P3_U3907 P3_R1200_U73 ; P3_R1200_U433
g25030 nand P3_U3075 P3_R1200_U72 ; P3_R1200_U434
g25031 not P3_R1200_U142 ; P3_R1200_U435
g25032 nand P3_R1200_U281 P3_R1200_U435 ; P3_R1200_U436
g25033 nand P3_R1200_U142 P3_R1200_U170 ; P3_R1200_U437
g25034 nand P3_U3392 P3_R1200_U31 ; P3_R1200_U438
g25035 nand P3_U3077 P3_R1200_U171 ; P3_R1200_U439
g25036 not P3_R1200_U143 ; P3_R1200_U440
g25037 nand P3_R1200_U200 P3_R1200_U440 ; P3_R1200_U441
g25038 nand P3_R1200_U143 P3_R1200_U172 ; P3_R1200_U442
g25039 nand P3_U3445 P3_R1200_U71 ; P3_R1200_U443
g25040 nand P3_U3080 P3_R1200_U70 ; P3_R1200_U444
g25041 not P3_R1200_U144 ; P3_R1200_U445
g25042 nand P3_R1200_U277 P3_R1200_U445 ; P3_R1200_U446
g25043 nand P3_R1200_U144 P3_R1200_U173 ; P3_R1200_U447
g25044 nand P3_U3443 P3_R1200_U69 ; P3_R1200_U448
g25045 nand P3_U3081 P3_R1200_U174 ; P3_R1200_U449
g25046 not P3_R1200_U145 ; P3_R1200_U450
g25047 nand P3_R1200_U275 P3_R1200_U450 ; P3_R1200_U451
g25048 nand P3_R1200_U145 P3_R1200_U175 ; P3_R1200_U452
g25049 nand P3_U3440 P3_R1200_U68 ; P3_R1200_U453
g25050 nand P3_U3068 P3_R1200_U67 ; P3_R1200_U454
g25051 not P3_R1200_U146 ; P3_R1200_U455
g25052 nand P3_R1200_U271 P3_R1200_U455 ; P3_R1200_U456
g25053 nand P3_R1200_U146 P3_R1200_U176 ; P3_R1200_U457
g25054 nand P3_U3437 P3_R1200_U63 ; P3_R1200_U458
g25055 nand P3_U3072 P3_R1200_U60 ; P3_R1200_U459
g25056 nand P3_R1200_U459 P3_R1200_U458 ; P3_R1200_U460
g25057 nand P3_U3434 P3_R1200_U64 ; P3_R1200_U461
g25058 nand P3_U3073 P3_R1200_U61 ; P3_R1200_U462
g25059 nand P3_R1200_U336 P3_R1200_U93 ; P3_R1200_U463
g25060 nand P3_R1200_U177 P3_R1200_U328 ; P3_R1200_U464
g25061 nand P3_U3431 P3_R1200_U65 ; P3_R1200_U465
g25062 nand P3_U3078 P3_R1200_U62 ; P3_R1200_U466
g25063 nand P3_R1200_U337 P3_R1200_U179 ; P3_R1200_U467
g25064 nand P3_R1200_U261 P3_R1200_U178 ; P3_R1200_U468
g25065 nand P3_U3428 P3_R1200_U59 ; P3_R1200_U469
g25066 nand P3_U3079 P3_R1200_U58 ; P3_R1200_U470
g25067 not P3_R1200_U149 ; P3_R1200_U471
g25068 nand P3_R1200_U257 P3_R1200_U471 ; P3_R1200_U472
g25069 nand P3_R1200_U149 P3_R1200_U180 ; P3_R1200_U473
g25070 nand P3_U3425 P3_R1200_U57 ; P3_R1200_U474
g25071 nand P3_U3071 P3_R1200_U56 ; P3_R1200_U475
g25072 not P3_R1200_U150 ; P3_R1200_U476
g25073 nand P3_R1200_U253 P3_R1200_U476 ; P3_R1200_U477
g25074 nand P3_R1200_U150 P3_R1200_U181 ; P3_R1200_U478
g25075 nand P3_U3422 P3_R1200_U53 ; P3_R1200_U479
g25076 nand P3_U3062 P3_R1200_U51 ; P3_R1200_U480
g25077 nand P3_R1200_U480 P3_R1200_U479 ; P3_R1200_U481
g25078 nand P3_U3419 P3_R1200_U54 ; P3_R1200_U482
g25079 nand P3_U3061 P3_R1200_U52 ; P3_R1200_U483
g25080 nand P3_R1200_U347 P3_R1200_U94 ; P3_R1200_U484
g25081 nand P3_R1200_U182 P3_R1200_U339 ; P3_R1200_U485
g25082 and P3_R1179_U210 P3_R1179_U209 ; P3_R1179_U6
g25083 and P3_R1179_U189 P3_R1179_U245 ; P3_R1179_U7
g25084 and P3_R1179_U247 P3_R1179_U246 ; P3_R1179_U8
g25085 and P3_R1179_U190 P3_R1179_U262 ; P3_R1179_U9
g25086 and P3_R1179_U264 P3_R1179_U263 ; P3_R1179_U10
g25087 and P3_R1179_U191 P3_R1179_U286 ; P3_R1179_U11
g25088 and P3_R1179_U288 P3_R1179_U287 ; P3_R1179_U12
g25089 and P3_R1179_U208 P3_R1179_U194 P3_R1179_U213 ; P3_R1179_U13
g25090 and P3_R1179_U218 P3_R1179_U195 ; P3_R1179_U14
g25091 and P3_R1179_U392 P3_R1179_U391 ; P3_R1179_U15
g25092 nand P3_R1179_U342 P3_R1179_U345 ; P3_R1179_U16
g25093 nand P3_R1179_U331 P3_R1179_U334 ; P3_R1179_U17
g25094 nand P3_R1179_U320 P3_R1179_U323 ; P3_R1179_U18
g25095 nand P3_R1179_U312 P3_R1179_U314 ; P3_R1179_U19
g25096 nand P3_R1179_U162 P3_R1179_U183 P3_R1179_U351 ; P3_R1179_U20
g25097 nand P3_R1179_U241 P3_R1179_U243 ; P3_R1179_U21
g25098 nand P3_R1179_U233 P3_R1179_U236 ; P3_R1179_U22
g25099 nand P3_R1179_U225 P3_R1179_U227 ; P3_R1179_U23
g25100 nand P3_R1179_U172 P3_R1179_U348 ; P3_R1179_U24
g25101 not P3_U3069 ; P3_R1179_U25
g25102 nand P3_U3069 P3_R1179_U39 ; P3_R1179_U26
g25103 not P3_U3083 ; P3_R1179_U27
g25104 not P3_U3413 ; P3_R1179_U28
g25105 not P3_U3395 ; P3_R1179_U29
g25106 not P3_U3387 ; P3_R1179_U30
g25107 not P3_U3077 ; P3_R1179_U31
g25108 not P3_U3398 ; P3_R1179_U32
g25109 not P3_U3067 ; P3_R1179_U33
g25110 nand P3_U3067 P3_R1179_U29 ; P3_R1179_U34
g25111 not P3_U3063 ; P3_R1179_U35
g25112 not P3_U3404 ; P3_R1179_U36
g25113 not P3_U3407 ; P3_R1179_U37
g25114 not P3_U3401 ; P3_R1179_U38
g25115 not P3_U3410 ; P3_R1179_U39
g25116 not P3_U3070 ; P3_R1179_U40
g25117 not P3_U3066 ; P3_R1179_U41
g25118 not P3_U3059 ; P3_R1179_U42
g25119 nand P3_U3059 P3_R1179_U38 ; P3_R1179_U43
g25120 nand P3_R1179_U214 P3_R1179_U212 ; P3_R1179_U44
g25121 not P3_U3416 ; P3_R1179_U45
g25122 not P3_U3082 ; P3_R1179_U46
g25123 nand P3_R1179_U44 P3_R1179_U215 ; P3_R1179_U47
g25124 nand P3_R1179_U43 P3_R1179_U229 ; P3_R1179_U48
g25125 nand P3_R1179_U201 P3_R1179_U185 P3_R1179_U349 ; P3_R1179_U49
g25126 not P3_U3901 ; P3_R1179_U50
g25127 not P3_U3422 ; P3_R1179_U51
g25128 not P3_U3419 ; P3_R1179_U52
g25129 not P3_U3062 ; P3_R1179_U53
g25130 not P3_U3061 ; P3_R1179_U54
g25131 nand P3_U3082 P3_R1179_U45 ; P3_R1179_U55
g25132 not P3_U3425 ; P3_R1179_U56
g25133 not P3_U3071 ; P3_R1179_U57
g25134 not P3_U3428 ; P3_R1179_U58
g25135 not P3_U3079 ; P3_R1179_U59
g25136 not P3_U3437 ; P3_R1179_U60
g25137 not P3_U3434 ; P3_R1179_U61
g25138 not P3_U3431 ; P3_R1179_U62
g25139 not P3_U3072 ; P3_R1179_U63
g25140 not P3_U3073 ; P3_R1179_U64
g25141 not P3_U3078 ; P3_R1179_U65
g25142 nand P3_U3078 P3_R1179_U62 ; P3_R1179_U66
g25143 not P3_U3440 ; P3_R1179_U67
g25144 not P3_U3068 ; P3_R1179_U68
g25145 not P3_U3081 ; P3_R1179_U69
g25146 not P3_U3445 ; P3_R1179_U70
g25147 not P3_U3080 ; P3_R1179_U71
g25148 not P3_U3907 ; P3_R1179_U72
g25149 not P3_U3075 ; P3_R1179_U73
g25150 not P3_U3904 ; P3_R1179_U74
g25151 not P3_U3905 ; P3_R1179_U75
g25152 not P3_U3906 ; P3_R1179_U76
g25153 not P3_U3065 ; P3_R1179_U77
g25154 not P3_U3060 ; P3_R1179_U78
g25155 not P3_U3074 ; P3_R1179_U79
g25156 nand P3_U3074 P3_R1179_U76 ; P3_R1179_U80
g25157 not P3_U3903 ; P3_R1179_U81
g25158 not P3_U3064 ; P3_R1179_U82
g25159 not P3_U3902 ; P3_R1179_U83
g25160 not P3_U3057 ; P3_R1179_U84
g25161 not P3_U3900 ; P3_R1179_U85
g25162 not P3_U3056 ; P3_R1179_U86
g25163 nand P3_U3056 P3_R1179_U50 ; P3_R1179_U87
g25164 not P3_U3052 ; P3_R1179_U88
g25165 not P3_U3899 ; P3_R1179_U89
g25166 not P3_U3053 ; P3_R1179_U90
g25167 nand P3_R1179_U302 P3_R1179_U301 ; P3_R1179_U91
g25168 nand P3_R1179_U80 P3_R1179_U316 ; P3_R1179_U92
g25169 nand P3_R1179_U66 P3_R1179_U327 ; P3_R1179_U93
g25170 nand P3_R1179_U55 P3_R1179_U338 ; P3_R1179_U94
g25171 not P3_U3076 ; P3_R1179_U95
g25172 nand P3_R1179_U402 P3_R1179_U401 ; P3_R1179_U96
g25173 nand P3_R1179_U416 P3_R1179_U415 ; P3_R1179_U97
g25174 nand P3_R1179_U421 P3_R1179_U420 ; P3_R1179_U98
g25175 nand P3_R1179_U437 P3_R1179_U436 ; P3_R1179_U99
g25176 nand P3_R1179_U442 P3_R1179_U441 ; P3_R1179_U100
g25177 nand P3_R1179_U447 P3_R1179_U446 ; P3_R1179_U101
g25178 nand P3_R1179_U452 P3_R1179_U451 ; P3_R1179_U102
g25179 nand P3_R1179_U457 P3_R1179_U456 ; P3_R1179_U103
g25180 nand P3_R1179_U473 P3_R1179_U472 ; P3_R1179_U104
g25181 nand P3_R1179_U478 P3_R1179_U477 ; P3_R1179_U105
g25182 nand P3_R1179_U361 P3_R1179_U360 ; P3_R1179_U106
g25183 nand P3_R1179_U370 P3_R1179_U369 ; P3_R1179_U107
g25184 nand P3_R1179_U377 P3_R1179_U376 ; P3_R1179_U108
g25185 nand P3_R1179_U381 P3_R1179_U380 ; P3_R1179_U109
g25186 nand P3_R1179_U390 P3_R1179_U389 ; P3_R1179_U110
g25187 nand P3_R1179_U411 P3_R1179_U410 ; P3_R1179_U111
g25188 nand P3_R1179_U428 P3_R1179_U427 ; P3_R1179_U112
g25189 nand P3_R1179_U432 P3_R1179_U431 ; P3_R1179_U113
g25190 nand P3_R1179_U464 P3_R1179_U463 ; P3_R1179_U114
g25191 nand P3_R1179_U468 P3_R1179_U467 ; P3_R1179_U115
g25192 nand P3_R1179_U485 P3_R1179_U484 ; P3_R1179_U116
g25193 and P3_R1179_U352 P3_R1179_U193 ; P3_R1179_U117
g25194 and P3_R1179_U205 P3_R1179_U206 ; P3_R1179_U118
g25195 and P3_R1179_U14 P3_R1179_U13 ; P3_R1179_U119
g25196 and P3_R1179_U357 P3_R1179_U354 ; P3_R1179_U120
g25197 and P3_R1179_U363 P3_R1179_U362 P3_R1179_U26 ; P3_R1179_U121
g25198 and P3_R1179_U366 P3_R1179_U195 ; P3_R1179_U122
g25199 and P3_R1179_U235 P3_R1179_U6 ; P3_R1179_U123
g25200 and P3_R1179_U373 P3_R1179_U194 ; P3_R1179_U124
g25201 and P3_R1179_U383 P3_R1179_U382 P3_R1179_U34 ; P3_R1179_U125
g25202 and P3_R1179_U386 P3_R1179_U193 ; P3_R1179_U126
g25203 and P3_R1179_U222 P3_R1179_U7 ; P3_R1179_U127
g25204 and P3_R1179_U267 P3_R1179_U9 ; P3_R1179_U128
g25205 and P3_R1179_U291 P3_R1179_U11 ; P3_R1179_U129
g25206 and P3_R1179_U355 P3_R1179_U192 ; P3_R1179_U130
g25207 and P3_R1179_U306 P3_R1179_U307 ; P3_R1179_U131
g25208 and P3_R1179_U309 P3_R1179_U395 ; P3_R1179_U132
g25209 and P3_R1179_U306 P3_R1179_U307 ; P3_R1179_U133
g25210 and P3_R1179_U15 P3_R1179_U310 ; P3_R1179_U134
g25211 nand P3_R1179_U399 P3_R1179_U398 ; P3_R1179_U135
g25212 and P3_R1179_U404 P3_R1179_U403 P3_R1179_U87 ; P3_R1179_U136
g25213 and P3_R1179_U407 P3_R1179_U192 ; P3_R1179_U137
g25214 nand P3_R1179_U413 P3_R1179_U412 ; P3_R1179_U138
g25215 nand P3_R1179_U418 P3_R1179_U417 ; P3_R1179_U139
g25216 and P3_R1179_U322 P3_R1179_U12 ; P3_R1179_U140
g25217 and P3_R1179_U424 P3_R1179_U191 ; P3_R1179_U141
g25218 nand P3_R1179_U434 P3_R1179_U433 ; P3_R1179_U142
g25219 nand P3_R1179_U439 P3_R1179_U438 ; P3_R1179_U143
g25220 nand P3_R1179_U444 P3_R1179_U443 ; P3_R1179_U144
g25221 nand P3_R1179_U449 P3_R1179_U448 ; P3_R1179_U145
g25222 nand P3_R1179_U454 P3_R1179_U453 ; P3_R1179_U146
g25223 and P3_R1179_U333 P3_R1179_U10 ; P3_R1179_U147
g25224 and P3_R1179_U460 P3_R1179_U190 ; P3_R1179_U148
g25225 nand P3_R1179_U470 P3_R1179_U469 ; P3_R1179_U149
g25226 nand P3_R1179_U475 P3_R1179_U474 ; P3_R1179_U150
g25227 and P3_R1179_U344 P3_R1179_U8 ; P3_R1179_U151
g25228 and P3_R1179_U481 P3_R1179_U189 ; P3_R1179_U152
g25229 and P3_R1179_U359 P3_R1179_U358 ; P3_R1179_U153
g25230 nand P3_R1179_U120 P3_R1179_U356 ; P3_R1179_U154
g25231 and P3_R1179_U368 P3_R1179_U367 ; P3_R1179_U155
g25232 and P3_R1179_U375 P3_R1179_U374 ; P3_R1179_U156
g25233 and P3_R1179_U379 P3_R1179_U378 ; P3_R1179_U157
g25234 nand P3_R1179_U118 P3_R1179_U203 ; P3_R1179_U158
g25235 and P3_R1179_U388 P3_R1179_U387 ; P3_R1179_U159
g25236 not P3_U3908 ; P3_R1179_U160
g25237 not P3_U3054 ; P3_R1179_U161
g25238 and P3_R1179_U397 P3_R1179_U396 ; P3_R1179_U162
g25239 nand P3_R1179_U131 P3_R1179_U304 ; P3_R1179_U163
g25240 and P3_R1179_U409 P3_R1179_U408 ; P3_R1179_U164
g25241 nand P3_R1179_U298 P3_R1179_U297 ; P3_R1179_U165
g25242 nand P3_R1179_U294 P3_R1179_U293 ; P3_R1179_U166
g25243 and P3_R1179_U426 P3_R1179_U425 ; P3_R1179_U167
g25244 and P3_R1179_U430 P3_R1179_U429 ; P3_R1179_U168
g25245 nand P3_R1179_U284 P3_R1179_U283 ; P3_R1179_U169
g25246 nand P3_R1179_U280 P3_R1179_U279 ; P3_R1179_U170
g25247 not P3_U3392 ; P3_R1179_U171
g25248 nand P3_U3387 P3_R1179_U95 ; P3_R1179_U172
g25249 nand P3_R1179_U276 P3_R1179_U184 P3_R1179_U350 ; P3_R1179_U173
g25250 not P3_U3443 ; P3_R1179_U174
g25251 nand P3_R1179_U274 P3_R1179_U273 ; P3_R1179_U175
g25252 nand P3_R1179_U270 P3_R1179_U269 ; P3_R1179_U176
g25253 and P3_R1179_U462 P3_R1179_U461 ; P3_R1179_U177
g25254 and P3_R1179_U466 P3_R1179_U465 ; P3_R1179_U178
g25255 nand P3_R1179_U260 P3_R1179_U259 ; P3_R1179_U179
g25256 nand P3_R1179_U256 P3_R1179_U255 ; P3_R1179_U180
g25257 nand P3_R1179_U252 P3_R1179_U251 ; P3_R1179_U181
g25258 and P3_R1179_U483 P3_R1179_U482 ; P3_R1179_U182
g25259 nand P3_R1179_U132 P3_R1179_U163 ; P3_R1179_U183
g25260 nand P3_R1179_U175 P3_R1179_U174 ; P3_R1179_U184
g25261 nand P3_R1179_U172 P3_R1179_U171 ; P3_R1179_U185
g25262 not P3_R1179_U87 ; P3_R1179_U186
g25263 not P3_R1179_U34 ; P3_R1179_U187
g25264 not P3_R1179_U26 ; P3_R1179_U188
g25265 nand P3_U3419 P3_R1179_U54 ; P3_R1179_U189
g25266 nand P3_U3434 P3_R1179_U64 ; P3_R1179_U190
g25267 nand P3_U3905 P3_R1179_U78 ; P3_R1179_U191
g25268 nand P3_U3901 P3_R1179_U86 ; P3_R1179_U192
g25269 nand P3_U3395 P3_R1179_U33 ; P3_R1179_U193
g25270 nand P3_U3404 P3_R1179_U41 ; P3_R1179_U194
g25271 nand P3_U3410 P3_R1179_U25 ; P3_R1179_U195
g25272 not P3_R1179_U66 ; P3_R1179_U196
g25273 not P3_R1179_U80 ; P3_R1179_U197
g25274 not P3_R1179_U43 ; P3_R1179_U198
g25275 not P3_R1179_U55 ; P3_R1179_U199
g25276 not P3_R1179_U172 ; P3_R1179_U200
g25277 nand P3_U3077 P3_R1179_U172 ; P3_R1179_U201
g25278 not P3_R1179_U49 ; P3_R1179_U202
g25279 nand P3_R1179_U117 P3_R1179_U49 ; P3_R1179_U203
g25280 nand P3_R1179_U35 P3_R1179_U34 ; P3_R1179_U204
g25281 nand P3_R1179_U204 P3_R1179_U32 ; P3_R1179_U205
g25282 nand P3_U3063 P3_R1179_U187 ; P3_R1179_U206
g25283 not P3_R1179_U158 ; P3_R1179_U207
g25284 nand P3_U3407 P3_R1179_U40 ; P3_R1179_U208
g25285 nand P3_U3070 P3_R1179_U37 ; P3_R1179_U209
g25286 nand P3_U3066 P3_R1179_U36 ; P3_R1179_U210
g25287 nand P3_R1179_U198 P3_R1179_U194 ; P3_R1179_U211
g25288 nand P3_R1179_U6 P3_R1179_U211 ; P3_R1179_U212
g25289 nand P3_U3401 P3_R1179_U42 ; P3_R1179_U213
g25290 nand P3_U3407 P3_R1179_U40 ; P3_R1179_U214
g25291 nand P3_R1179_U13 P3_R1179_U158 ; P3_R1179_U215
g25292 not P3_R1179_U44 ; P3_R1179_U216
g25293 not P3_R1179_U47 ; P3_R1179_U217
g25294 nand P3_U3413 P3_R1179_U27 ; P3_R1179_U218
g25295 nand P3_R1179_U27 P3_R1179_U26 ; P3_R1179_U219
g25296 nand P3_U3083 P3_R1179_U188 ; P3_R1179_U220
g25297 not P3_R1179_U154 ; P3_R1179_U221
g25298 nand P3_U3416 P3_R1179_U46 ; P3_R1179_U222
g25299 nand P3_R1179_U222 P3_R1179_U55 ; P3_R1179_U223
g25300 nand P3_R1179_U217 P3_R1179_U26 ; P3_R1179_U224
g25301 nand P3_R1179_U122 P3_R1179_U224 ; P3_R1179_U225
g25302 nand P3_R1179_U47 P3_R1179_U195 ; P3_R1179_U226
g25303 nand P3_R1179_U121 P3_R1179_U226 ; P3_R1179_U227
g25304 nand P3_R1179_U26 P3_R1179_U195 ; P3_R1179_U228
g25305 nand P3_R1179_U213 P3_R1179_U158 ; P3_R1179_U229
g25306 not P3_R1179_U48 ; P3_R1179_U230
g25307 nand P3_U3066 P3_R1179_U36 ; P3_R1179_U231
g25308 nand P3_R1179_U230 P3_R1179_U231 ; P3_R1179_U232
g25309 nand P3_R1179_U124 P3_R1179_U232 ; P3_R1179_U233
g25310 nand P3_R1179_U48 P3_R1179_U194 ; P3_R1179_U234
g25311 nand P3_U3407 P3_R1179_U40 ; P3_R1179_U235
g25312 nand P3_R1179_U123 P3_R1179_U234 ; P3_R1179_U236
g25313 nand P3_U3066 P3_R1179_U36 ; P3_R1179_U237
g25314 nand P3_R1179_U194 P3_R1179_U237 ; P3_R1179_U238
g25315 nand P3_R1179_U213 P3_R1179_U43 ; P3_R1179_U239
g25316 nand P3_R1179_U202 P3_R1179_U34 ; P3_R1179_U240
g25317 nand P3_R1179_U126 P3_R1179_U240 ; P3_R1179_U241
g25318 nand P3_R1179_U49 P3_R1179_U193 ; P3_R1179_U242
g25319 nand P3_R1179_U125 P3_R1179_U242 ; P3_R1179_U243
g25320 nand P3_R1179_U193 P3_R1179_U34 ; P3_R1179_U244
g25321 nand P3_U3422 P3_R1179_U53 ; P3_R1179_U245
g25322 nand P3_U3062 P3_R1179_U51 ; P3_R1179_U246
g25323 nand P3_U3061 P3_R1179_U52 ; P3_R1179_U247
g25324 nand P3_R1179_U199 P3_R1179_U7 ; P3_R1179_U248
g25325 nand P3_R1179_U8 P3_R1179_U248 ; P3_R1179_U249
g25326 nand P3_U3422 P3_R1179_U53 ; P3_R1179_U250
g25327 nand P3_R1179_U127 P3_R1179_U154 ; P3_R1179_U251
g25328 nand P3_R1179_U250 P3_R1179_U249 ; P3_R1179_U252
g25329 not P3_R1179_U181 ; P3_R1179_U253
g25330 nand P3_U3425 P3_R1179_U57 ; P3_R1179_U254
g25331 nand P3_R1179_U254 P3_R1179_U181 ; P3_R1179_U255
g25332 nand P3_U3071 P3_R1179_U56 ; P3_R1179_U256
g25333 not P3_R1179_U180 ; P3_R1179_U257
g25334 nand P3_U3428 P3_R1179_U59 ; P3_R1179_U258
g25335 nand P3_R1179_U258 P3_R1179_U180 ; P3_R1179_U259
g25336 nand P3_U3079 P3_R1179_U58 ; P3_R1179_U260
g25337 not P3_R1179_U179 ; P3_R1179_U261
g25338 nand P3_U3437 P3_R1179_U63 ; P3_R1179_U262
g25339 nand P3_U3072 P3_R1179_U60 ; P3_R1179_U263
g25340 nand P3_U3073 P3_R1179_U61 ; P3_R1179_U264
g25341 nand P3_R1179_U196 P3_R1179_U9 ; P3_R1179_U265
g25342 nand P3_R1179_U10 P3_R1179_U265 ; P3_R1179_U266
g25343 nand P3_U3431 P3_R1179_U65 ; P3_R1179_U267
g25344 nand P3_U3437 P3_R1179_U63 ; P3_R1179_U268
g25345 nand P3_R1179_U128 P3_R1179_U179 ; P3_R1179_U269
g25346 nand P3_R1179_U268 P3_R1179_U266 ; P3_R1179_U270
g25347 not P3_R1179_U176 ; P3_R1179_U271
g25348 nand P3_U3440 P3_R1179_U68 ; P3_R1179_U272
g25349 nand P3_R1179_U272 P3_R1179_U176 ; P3_R1179_U273
g25350 nand P3_U3068 P3_R1179_U67 ; P3_R1179_U274
g25351 not P3_R1179_U175 ; P3_R1179_U275
g25352 nand P3_U3081 P3_R1179_U175 ; P3_R1179_U276
g25353 not P3_R1179_U173 ; P3_R1179_U277
g25354 nand P3_U3445 P3_R1179_U71 ; P3_R1179_U278
g25355 nand P3_R1179_U278 P3_R1179_U173 ; P3_R1179_U279
g25356 nand P3_U3080 P3_R1179_U70 ; P3_R1179_U280
g25357 not P3_R1179_U170 ; P3_R1179_U281
g25358 nand P3_U3907 P3_R1179_U73 ; P3_R1179_U282
g25359 nand P3_R1179_U282 P3_R1179_U170 ; P3_R1179_U283
g25360 nand P3_U3075 P3_R1179_U72 ; P3_R1179_U284
g25361 not P3_R1179_U169 ; P3_R1179_U285
g25362 nand P3_U3904 P3_R1179_U77 ; P3_R1179_U286
g25363 nand P3_U3065 P3_R1179_U74 ; P3_R1179_U287
g25364 nand P3_U3060 P3_R1179_U75 ; P3_R1179_U288
g25365 nand P3_R1179_U197 P3_R1179_U11 ; P3_R1179_U289
g25366 nand P3_R1179_U12 P3_R1179_U289 ; P3_R1179_U290
g25367 nand P3_U3906 P3_R1179_U79 ; P3_R1179_U291
g25368 nand P3_U3904 P3_R1179_U77 ; P3_R1179_U292
g25369 nand P3_R1179_U129 P3_R1179_U169 ; P3_R1179_U293
g25370 nand P3_R1179_U292 P3_R1179_U290 ; P3_R1179_U294
g25371 not P3_R1179_U166 ; P3_R1179_U295
g25372 nand P3_U3903 P3_R1179_U82 ; P3_R1179_U296
g25373 nand P3_R1179_U296 P3_R1179_U166 ; P3_R1179_U297
g25374 nand P3_U3064 P3_R1179_U81 ; P3_R1179_U298
g25375 not P3_R1179_U165 ; P3_R1179_U299
g25376 nand P3_U3902 P3_R1179_U84 ; P3_R1179_U300
g25377 nand P3_R1179_U300 P3_R1179_U165 ; P3_R1179_U301
g25378 nand P3_U3057 P3_R1179_U83 ; P3_R1179_U302
g25379 not P3_R1179_U91 ; P3_R1179_U303
g25380 nand P3_R1179_U130 P3_R1179_U91 ; P3_R1179_U304
g25381 nand P3_R1179_U88 P3_R1179_U87 ; P3_R1179_U305
g25382 nand P3_R1179_U305 P3_R1179_U85 ; P3_R1179_U306
g25383 nand P3_U3052 P3_R1179_U186 ; P3_R1179_U307
g25384 not P3_R1179_U163 ; P3_R1179_U308
g25385 nand P3_U3899 P3_R1179_U90 ; P3_R1179_U309
g25386 nand P3_U3053 P3_R1179_U89 ; P3_R1179_U310
g25387 nand P3_R1179_U303 P3_R1179_U87 ; P3_R1179_U311
g25388 nand P3_R1179_U137 P3_R1179_U311 ; P3_R1179_U312
g25389 nand P3_R1179_U91 P3_R1179_U192 ; P3_R1179_U313
g25390 nand P3_R1179_U136 P3_R1179_U313 ; P3_R1179_U314
g25391 nand P3_R1179_U192 P3_R1179_U87 ; P3_R1179_U315
g25392 nand P3_R1179_U291 P3_R1179_U169 ; P3_R1179_U316
g25393 not P3_R1179_U92 ; P3_R1179_U317
g25394 nand P3_U3060 P3_R1179_U75 ; P3_R1179_U318
g25395 nand P3_R1179_U317 P3_R1179_U318 ; P3_R1179_U319
g25396 nand P3_R1179_U141 P3_R1179_U319 ; P3_R1179_U320
g25397 nand P3_R1179_U92 P3_R1179_U191 ; P3_R1179_U321
g25398 nand P3_U3904 P3_R1179_U77 ; P3_R1179_U322
g25399 nand P3_R1179_U140 P3_R1179_U321 ; P3_R1179_U323
g25400 nand P3_U3060 P3_R1179_U75 ; P3_R1179_U324
g25401 nand P3_R1179_U191 P3_R1179_U324 ; P3_R1179_U325
g25402 nand P3_R1179_U291 P3_R1179_U80 ; P3_R1179_U326
g25403 nand P3_R1179_U267 P3_R1179_U179 ; P3_R1179_U327
g25404 not P3_R1179_U93 ; P3_R1179_U328
g25405 nand P3_U3073 P3_R1179_U61 ; P3_R1179_U329
g25406 nand P3_R1179_U328 P3_R1179_U329 ; P3_R1179_U330
g25407 nand P3_R1179_U148 P3_R1179_U330 ; P3_R1179_U331
g25408 nand P3_R1179_U93 P3_R1179_U190 ; P3_R1179_U332
g25409 nand P3_U3437 P3_R1179_U63 ; P3_R1179_U333
g25410 nand P3_R1179_U147 P3_R1179_U332 ; P3_R1179_U334
g25411 nand P3_U3073 P3_R1179_U61 ; P3_R1179_U335
g25412 nand P3_R1179_U190 P3_R1179_U335 ; P3_R1179_U336
g25413 nand P3_R1179_U267 P3_R1179_U66 ; P3_R1179_U337
g25414 nand P3_R1179_U222 P3_R1179_U154 ; P3_R1179_U338
g25415 not P3_R1179_U94 ; P3_R1179_U339
g25416 nand P3_U3061 P3_R1179_U52 ; P3_R1179_U340
g25417 nand P3_R1179_U339 P3_R1179_U340 ; P3_R1179_U341
g25418 nand P3_R1179_U152 P3_R1179_U341 ; P3_R1179_U342
g25419 nand P3_R1179_U94 P3_R1179_U189 ; P3_R1179_U343
g25420 nand P3_U3422 P3_R1179_U53 ; P3_R1179_U344
g25421 nand P3_R1179_U151 P3_R1179_U343 ; P3_R1179_U345
g25422 nand P3_U3061 P3_R1179_U52 ; P3_R1179_U346
g25423 nand P3_R1179_U189 P3_R1179_U346 ; P3_R1179_U347
g25424 nand P3_U3076 P3_R1179_U30 ; P3_R1179_U348
g25425 nand P3_U3077 P3_R1179_U171 ; P3_R1179_U349
g25426 nand P3_U3081 P3_R1179_U174 ; P3_R1179_U350
g25427 nand P3_R1179_U133 P3_R1179_U304 P3_R1179_U134 ; P3_R1179_U351
g25428 nand P3_U3398 P3_R1179_U35 ; P3_R1179_U352
g25429 nand P3_U3413 P3_R1179_U220 ; P3_R1179_U353
g25430 nand P3_R1179_U353 P3_R1179_U219 ; P3_R1179_U354
g25431 nand P3_U3900 P3_R1179_U88 ; P3_R1179_U355
g25432 nand P3_R1179_U119 P3_R1179_U158 ; P3_R1179_U356
g25433 nand P3_R1179_U216 P3_R1179_U14 ; P3_R1179_U357
g25434 nand P3_U3416 P3_R1179_U46 ; P3_R1179_U358
g25435 nand P3_U3082 P3_R1179_U45 ; P3_R1179_U359
g25436 nand P3_R1179_U223 P3_R1179_U154 ; P3_R1179_U360
g25437 nand P3_R1179_U221 P3_R1179_U153 ; P3_R1179_U361
g25438 nand P3_U3413 P3_R1179_U27 ; P3_R1179_U362
g25439 nand P3_U3083 P3_R1179_U28 ; P3_R1179_U363
g25440 nand P3_U3413 P3_R1179_U27 ; P3_R1179_U364
g25441 nand P3_U3083 P3_R1179_U28 ; P3_R1179_U365
g25442 nand P3_R1179_U365 P3_R1179_U364 ; P3_R1179_U366
g25443 nand P3_U3410 P3_R1179_U25 ; P3_R1179_U367
g25444 nand P3_U3069 P3_R1179_U39 ; P3_R1179_U368
g25445 nand P3_R1179_U228 P3_R1179_U47 ; P3_R1179_U369
g25446 nand P3_R1179_U155 P3_R1179_U217 ; P3_R1179_U370
g25447 nand P3_U3407 P3_R1179_U40 ; P3_R1179_U371
g25448 nand P3_U3070 P3_R1179_U37 ; P3_R1179_U372
g25449 nand P3_R1179_U372 P3_R1179_U371 ; P3_R1179_U373
g25450 nand P3_U3404 P3_R1179_U41 ; P3_R1179_U374
g25451 nand P3_U3066 P3_R1179_U36 ; P3_R1179_U375
g25452 nand P3_R1179_U238 P3_R1179_U48 ; P3_R1179_U376
g25453 nand P3_R1179_U156 P3_R1179_U230 ; P3_R1179_U377
g25454 nand P3_U3401 P3_R1179_U42 ; P3_R1179_U378
g25455 nand P3_U3059 P3_R1179_U38 ; P3_R1179_U379
g25456 nand P3_R1179_U239 P3_R1179_U158 ; P3_R1179_U380
g25457 nand P3_R1179_U207 P3_R1179_U157 ; P3_R1179_U381
g25458 nand P3_U3398 P3_R1179_U35 ; P3_R1179_U382
g25459 nand P3_U3063 P3_R1179_U32 ; P3_R1179_U383
g25460 nand P3_U3398 P3_R1179_U35 ; P3_R1179_U384
g25461 nand P3_U3063 P3_R1179_U32 ; P3_R1179_U385
g25462 nand P3_R1179_U385 P3_R1179_U384 ; P3_R1179_U386
g25463 nand P3_U3395 P3_R1179_U33 ; P3_R1179_U387
g25464 nand P3_U3067 P3_R1179_U29 ; P3_R1179_U388
g25465 nand P3_R1179_U244 P3_R1179_U49 ; P3_R1179_U389
g25466 nand P3_R1179_U159 P3_R1179_U202 ; P3_R1179_U390
g25467 nand P3_U3908 P3_R1179_U161 ; P3_R1179_U391
g25468 nand P3_U3054 P3_R1179_U160 ; P3_R1179_U392
g25469 nand P3_U3908 P3_R1179_U161 ; P3_R1179_U393
g25470 nand P3_U3054 P3_R1179_U160 ; P3_R1179_U394
g25471 nand P3_R1179_U394 P3_R1179_U393 ; P3_R1179_U395
g25472 nand P3_U3053 P3_R1179_U395 P3_R1179_U89 ; P3_R1179_U396
g25473 nand P3_R1179_U15 P3_R1179_U90 P3_U3899 ; P3_R1179_U397
g25474 nand P3_U3899 P3_R1179_U90 ; P3_R1179_U398
g25475 nand P3_U3053 P3_R1179_U89 ; P3_R1179_U399
g25476 not P3_R1179_U135 ; P3_R1179_U400
g25477 nand P3_R1179_U308 P3_R1179_U400 ; P3_R1179_U401
g25478 nand P3_R1179_U135 P3_R1179_U163 ; P3_R1179_U402
g25479 nand P3_U3900 P3_R1179_U88 ; P3_R1179_U403
g25480 nand P3_U3052 P3_R1179_U85 ; P3_R1179_U404
g25481 nand P3_U3900 P3_R1179_U88 ; P3_R1179_U405
g25482 nand P3_U3052 P3_R1179_U85 ; P3_R1179_U406
g25483 nand P3_R1179_U406 P3_R1179_U405 ; P3_R1179_U407
g25484 nand P3_U3901 P3_R1179_U86 ; P3_R1179_U408
g25485 nand P3_U3056 P3_R1179_U50 ; P3_R1179_U409
g25486 nand P3_R1179_U315 P3_R1179_U91 ; P3_R1179_U410
g25487 nand P3_R1179_U164 P3_R1179_U303 ; P3_R1179_U411
g25488 nand P3_U3902 P3_R1179_U84 ; P3_R1179_U412
g25489 nand P3_U3057 P3_R1179_U83 ; P3_R1179_U413
g25490 not P3_R1179_U138 ; P3_R1179_U414
g25491 nand P3_R1179_U299 P3_R1179_U414 ; P3_R1179_U415
g25492 nand P3_R1179_U138 P3_R1179_U165 ; P3_R1179_U416
g25493 nand P3_U3903 P3_R1179_U82 ; P3_R1179_U417
g25494 nand P3_U3064 P3_R1179_U81 ; P3_R1179_U418
g25495 not P3_R1179_U139 ; P3_R1179_U419
g25496 nand P3_R1179_U295 P3_R1179_U419 ; P3_R1179_U420
g25497 nand P3_R1179_U139 P3_R1179_U166 ; P3_R1179_U421
g25498 nand P3_U3904 P3_R1179_U77 ; P3_R1179_U422
g25499 nand P3_U3065 P3_R1179_U74 ; P3_R1179_U423
g25500 nand P3_R1179_U423 P3_R1179_U422 ; P3_R1179_U424
g25501 nand P3_U3905 P3_R1179_U78 ; P3_R1179_U425
g25502 nand P3_U3060 P3_R1179_U75 ; P3_R1179_U426
g25503 nand P3_R1179_U325 P3_R1179_U92 ; P3_R1179_U427
g25504 nand P3_R1179_U167 P3_R1179_U317 ; P3_R1179_U428
g25505 nand P3_U3906 P3_R1179_U79 ; P3_R1179_U429
g25506 nand P3_U3074 P3_R1179_U76 ; P3_R1179_U430
g25507 nand P3_R1179_U326 P3_R1179_U169 ; P3_R1179_U431
g25508 nand P3_R1179_U285 P3_R1179_U168 ; P3_R1179_U432
g25509 nand P3_U3907 P3_R1179_U73 ; P3_R1179_U433
g25510 nand P3_U3075 P3_R1179_U72 ; P3_R1179_U434
g25511 not P3_R1179_U142 ; P3_R1179_U435
g25512 nand P3_R1179_U281 P3_R1179_U435 ; P3_R1179_U436
g25513 nand P3_R1179_U142 P3_R1179_U170 ; P3_R1179_U437
g25514 nand P3_U3392 P3_R1179_U31 ; P3_R1179_U438
g25515 nand P3_U3077 P3_R1179_U171 ; P3_R1179_U439
g25516 not P3_R1179_U143 ; P3_R1179_U440
g25517 nand P3_R1179_U200 P3_R1179_U440 ; P3_R1179_U441
g25518 nand P3_R1179_U143 P3_R1179_U172 ; P3_R1179_U442
g25519 nand P3_U3445 P3_R1179_U71 ; P3_R1179_U443
g25520 nand P3_U3080 P3_R1179_U70 ; P3_R1179_U444
g25521 not P3_R1179_U144 ; P3_R1179_U445
g25522 nand P3_R1179_U277 P3_R1179_U445 ; P3_R1179_U446
g25523 nand P3_R1179_U144 P3_R1179_U173 ; P3_R1179_U447
g25524 nand P3_U3443 P3_R1179_U69 ; P3_R1179_U448
g25525 nand P3_U3081 P3_R1179_U174 ; P3_R1179_U449
g25526 not P3_R1179_U145 ; P3_R1179_U450
g25527 nand P3_R1179_U275 P3_R1179_U450 ; P3_R1179_U451
g25528 nand P3_R1179_U145 P3_R1179_U175 ; P3_R1179_U452
g25529 nand P3_U3440 P3_R1179_U68 ; P3_R1179_U453
g25530 nand P3_U3068 P3_R1179_U67 ; P3_R1179_U454
g25531 not P3_R1179_U146 ; P3_R1179_U455
g25532 nand P3_R1179_U271 P3_R1179_U455 ; P3_R1179_U456
g25533 nand P3_R1179_U146 P3_R1179_U176 ; P3_R1179_U457
g25534 nand P3_U3437 P3_R1179_U63 ; P3_R1179_U458
g25535 nand P3_U3072 P3_R1179_U60 ; P3_R1179_U459
g25536 nand P3_R1179_U459 P3_R1179_U458 ; P3_R1179_U460
g25537 nand P3_U3434 P3_R1179_U64 ; P3_R1179_U461
g25538 nand P3_U3073 P3_R1179_U61 ; P3_R1179_U462
g25539 nand P3_R1179_U336 P3_R1179_U93 ; P3_R1179_U463
g25540 nand P3_R1179_U177 P3_R1179_U328 ; P3_R1179_U464
g25541 nand P3_U3431 P3_R1179_U65 ; P3_R1179_U465
g25542 nand P3_U3078 P3_R1179_U62 ; P3_R1179_U466
g25543 nand P3_R1179_U337 P3_R1179_U179 ; P3_R1179_U467
g25544 nand P3_R1179_U261 P3_R1179_U178 ; P3_R1179_U468
g25545 nand P3_U3428 P3_R1179_U59 ; P3_R1179_U469
g25546 nand P3_U3079 P3_R1179_U58 ; P3_R1179_U470
g25547 not P3_R1179_U149 ; P3_R1179_U471
g25548 nand P3_R1179_U257 P3_R1179_U471 ; P3_R1179_U472
g25549 nand P3_R1179_U149 P3_R1179_U180 ; P3_R1179_U473
g25550 nand P3_U3425 P3_R1179_U57 ; P3_R1179_U474
g25551 nand P3_U3071 P3_R1179_U56 ; P3_R1179_U475
g25552 not P3_R1179_U150 ; P3_R1179_U476
g25553 nand P3_R1179_U253 P3_R1179_U476 ; P3_R1179_U477
g25554 nand P3_R1179_U150 P3_R1179_U181 ; P3_R1179_U478
g25555 nand P3_U3422 P3_R1179_U53 ; P3_R1179_U479
g25556 nand P3_U3062 P3_R1179_U51 ; P3_R1179_U480
g25557 nand P3_R1179_U480 P3_R1179_U479 ; P3_R1179_U481
g25558 nand P3_U3419 P3_R1179_U54 ; P3_R1179_U482
g25559 nand P3_U3061 P3_R1179_U52 ; P3_R1179_U483
g25560 nand P3_R1179_U347 P3_R1179_U94 ; P3_R1179_U484
g25561 nand P3_R1179_U182 P3_R1179_U339 ; P3_R1179_U485
g25562 and P3_R1269_U107 P3_R1269_U108 ; P3_R1269_U6
g25563 and P3_R1269_U118 P3_R1269_U117 ; P3_R1269_U7
g25564 and P3_R1269_U142 P3_R1269_U141 ; P3_R1269_U8
g25565 and P3_R1269_U200 P3_R1269_U199 ; P3_R1269_U9
g25566 and P3_R1269_U202 P3_R1269_U201 ; P3_R1269_U10
g25567 nand P3_R1269_U10 P3_R1269_U194 P3_R1269_U196 ; P3_R1269_U11
g25568 not P3_U3116 ; P3_R1269_U12
g25569 not P3_U3094 ; P3_R1269_U13
g25570 not P3_U3095 ; P3_R1269_U14
g25571 not P3_U3130 ; P3_R1269_U15
g25572 not P3_U3136 ; P3_R1269_U16
g25573 not P3_U3135 ; P3_R1269_U17
g25574 not P3_U3106 ; P3_R1269_U18
g25575 not P3_U3107 ; P3_R1269_U19
g25576 not P3_U3112 ; P3_R1269_U20
g25577 not P3_U3113 ; P3_R1269_U21
g25578 not P3_U3114 ; P3_R1269_U22
g25579 not P3_U3142 ; P3_R1269_U23
g25580 not P3_U3141 ; P3_R1269_U24
g25581 not P3_U3146 ; P3_R1269_U25
g25582 not P3_U3145 ; P3_R1269_U26
g25583 not P3_U3144 ; P3_R1269_U27
g25584 not P3_U3143 ; P3_R1269_U28
g25585 not P3_U3111 ; P3_R1269_U29
g25586 not P3_U3109 ; P3_R1269_U30
g25587 not P3_U3110 ; P3_R1269_U31
g25588 not P3_U3108 ; P3_R1269_U32
g25589 not P3_U3140 ; P3_R1269_U33
g25590 not P3_U3139 ; P3_R1269_U34
g25591 not P3_U3138 ; P3_R1269_U35
g25592 not P3_U3137 ; P3_R1269_U36
g25593 not P3_U3101 ; P3_R1269_U37
g25594 not P3_U3100 ; P3_R1269_U38
g25595 not P3_U3104 ; P3_R1269_U39
g25596 not P3_U3105 ; P3_R1269_U40
g25597 not P3_U3103 ; P3_R1269_U41
g25598 not P3_U3102 ; P3_R1269_U42
g25599 not P3_U3134 ; P3_R1269_U43
g25600 not P3_U3133 ; P3_R1269_U44
g25601 not P3_U3132 ; P3_R1269_U45
g25602 not P3_U3131 ; P3_R1269_U46
g25603 not P3_U3099 ; P3_R1269_U47
g25604 not P3_U3098 ; P3_R1269_U48
g25605 nand P3_R1269_U157 P3_R1269_U156 ; P3_R1269_U49
g25606 not P3_U3129 ; P3_R1269_U50
g25607 not P3_U3096 ; P3_R1269_U51
g25608 not P3_U3123 ; P3_R1269_U52
g25609 not P3_U3124 ; P3_R1269_U53
g25610 not P3_U3128 ; P3_R1269_U54
g25611 not P3_U3127 ; P3_R1269_U55
g25612 not P3_U3126 ; P3_R1269_U56
g25613 not P3_U3125 ; P3_R1269_U57
g25614 not P3_U3087 ; P3_R1269_U58
g25615 not P3_U3089 ; P3_R1269_U59
g25616 not P3_U3088 ; P3_R1269_U60
g25617 not P3_U3086 ; P3_R1269_U61
g25618 not P3_U3093 ; P3_R1269_U62
g25619 not P3_U3092 ; P3_R1269_U63
g25620 not P3_U3090 ; P3_R1269_U64
g25621 not P3_U3091 ; P3_R1269_U65
g25622 not P3_U3120 ; P3_R1269_U66
g25623 not P3_U3119 ; P3_R1269_U67
g25624 nand P3_R1269_U178 P3_R1269_U177 ; P3_R1269_U68
g25625 not P3_U3121 ; P3_R1269_U69
g25626 not P3_U3122 ; P3_R1269_U70
g25627 not P3_U3118 ; P3_R1269_U71
g25628 not P3_U3149 ; P3_R1269_U72
g25629 and P3_R1269_U111 P3_R1269_U110 ; P3_R1269_U73
g25630 and P3_R1269_U7 P3_R1269_U124 ; P3_R1269_U74
g25631 and P3_U3111 P3_R1269_U28 ; P3_R1269_U75
g25632 and P3_U3110 P3_R1269_U23 ; P3_R1269_U76
g25633 and P3_R1269_U126 P3_R1269_U127 P3_R1269_U78 ; P3_R1269_U77
g25634 and P3_R1269_U130 P3_R1269_U129 ; P3_R1269_U78
g25635 and P3_R1269_U6 P3_R1269_U80 ; P3_R1269_U79
g25636 and P3_R1269_U138 P3_R1269_U139 ; P3_R1269_U80
g25637 and P3_U3104 P3_R1269_U16 ; P3_R1269_U81
g25638 and P3_U3105 P3_R1269_U36 ; P3_R1269_U82
g25639 and P3_R1269_U143 P3_R1269_U144 P3_R1269_U85 ; P3_R1269_U83
g25640 and P3_R1269_U146 P3_R1269_U145 ; P3_R1269_U84
g25641 and P3_R1269_U84 P3_R1269_U8 ; P3_R1269_U85
g25642 and P3_U3134 P3_R1269_U42 ; P3_R1269_U86
g25643 and P3_U3133 P3_R1269_U37 ; P3_R1269_U87
g25644 and P3_R1269_U148 P3_R1269_U150 P3_R1269_U89 ; P3_R1269_U88
g25645 and P3_R1269_U152 P3_R1269_U151 ; P3_R1269_U89
g25646 and P3_R1269_U104 P3_R1269_U103 ; P3_R1269_U90
g25647 and P3_R1269_U162 P3_R1269_U161 ; P3_R1269_U91
g25648 and P3_U3128 P3_R1269_U51 ; P3_R1269_U92
g25649 and P3_R1269_U170 P3_R1269_U169 P3_R1269_U171 P3_R1269_U165 ; P3_R1269_U93
g25650 and P3_R1269_U175 P3_R1269_U174 ; P3_R1269_U94
g25651 and P3_R1269_U172 P3_R1269_U94 P3_R1269_U173 P3_R1269_U96 P3_R1269_U176 ; P3_R1269_U95
g25652 and P3_R1269_U193 P3_R1269_U191 P3_R1269_U192 ; P3_R1269_U96
g25653 and P3_U3120 P3_R1269_U60 ; P3_R1269_U97
g25654 and P3_R1269_U174 P3_R1269_U175 ; P3_R1269_U98
g25655 and P3_R1269_U198 P3_R1269_U186 ; P3_R1269_U99
g25656 not P3_U3084 ; P3_R1269_U100
g25657 not P3_U3085 ; P3_R1269_U101
g25658 nand P3_R1269_U187 P3_R1269_U195 ; P3_R1269_U102
g25659 nand P3_U3094 P3_R1269_U56 ; P3_R1269_U103
g25660 nand P3_U3095 P3_R1269_U55 ; P3_R1269_U104
g25661 nand P3_U3130 P3_R1269_U48 ; P3_R1269_U105
g25662 nand P3_U3106 P3_R1269_U35 ; P3_R1269_U106
g25663 nand P3_U3135 P3_R1269_U41 ; P3_R1269_U107
g25664 nand P3_U3136 P3_R1269_U39 ; P3_R1269_U108
g25665 nand P3_U3107 P3_R1269_U34 ; P3_R1269_U109
g25666 nand P3_U3112 P3_R1269_U27 ; P3_R1269_U110
g25667 nand P3_U3113 P3_R1269_U26 ; P3_R1269_U111
g25668 nand P3_U3147 P3_U3148 ; P3_R1269_U112
g25669 nand P3_U3115 P3_R1269_U112 ; P3_R1269_U113
g25670 or P3_U3147 P3_U3148 ; P3_R1269_U114
g25671 nand P3_U3114 P3_R1269_U25 ; P3_R1269_U115
g25672 nand P3_R1269_U111 P3_R1269_U110 P3_R1269_U113 P3_R1269_U115 P3_R1269_U114 ; P3_R1269_U116
g25673 nand P3_U3142 P3_R1269_U31 ; P3_R1269_U117
g25674 nand P3_U3141 P3_R1269_U30 ; P3_R1269_U118
g25675 nand P3_U3146 P3_R1269_U22 ; P3_R1269_U119
g25676 nand P3_U3145 P3_R1269_U21 ; P3_R1269_U120
g25677 nand P3_R1269_U120 P3_R1269_U119 ; P3_R1269_U121
g25678 nand P3_R1269_U73 P3_R1269_U121 ; P3_R1269_U122
g25679 nand P3_U3144 P3_R1269_U20 ; P3_R1269_U123
g25680 nand P3_U3143 P3_R1269_U29 ; P3_R1269_U124
g25681 nand P3_R1269_U122 P3_R1269_U123 P3_R1269_U116 P3_R1269_U74 ; P3_R1269_U125
g25682 nand P3_R1269_U75 P3_R1269_U7 ; P3_R1269_U126
g25683 nand P3_U3109 P3_R1269_U24 ; P3_R1269_U127
g25684 nand P3_U3141 P3_R1269_U30 ; P3_R1269_U128
g25685 nand P3_R1269_U76 P3_R1269_U128 ; P3_R1269_U129
g25686 nand P3_U3108 P3_R1269_U33 ; P3_R1269_U130
g25687 nand P3_R1269_U125 P3_R1269_U77 ; P3_R1269_U131
g25688 nand P3_U3140 P3_R1269_U32 ; P3_R1269_U132
g25689 nand P3_R1269_U132 P3_R1269_U131 ; P3_R1269_U133
g25690 nand P3_R1269_U133 P3_R1269_U109 ; P3_R1269_U134
g25691 nand P3_U3139 P3_R1269_U19 ; P3_R1269_U135
g25692 nand P3_R1269_U135 P3_R1269_U134 ; P3_R1269_U136
g25693 nand P3_R1269_U136 P3_R1269_U106 ; P3_R1269_U137
g25694 nand P3_U3138 P3_R1269_U18 ; P3_R1269_U138
g25695 nand P3_U3137 P3_R1269_U40 ; P3_R1269_U139
g25696 nand P3_R1269_U137 P3_R1269_U79 ; P3_R1269_U140
g25697 nand P3_U3101 P3_R1269_U44 ; P3_R1269_U141
g25698 nand P3_U3100 P3_R1269_U45 ; P3_R1269_U142
g25699 nand P3_R1269_U81 P3_R1269_U107 ; P3_R1269_U143
g25700 nand P3_R1269_U82 P3_R1269_U6 ; P3_R1269_U144
g25701 nand P3_U3103 P3_R1269_U17 ; P3_R1269_U145
g25702 nand P3_U3102 P3_R1269_U43 ; P3_R1269_U146
g25703 nand P3_R1269_U140 P3_R1269_U83 ; P3_R1269_U147
g25704 nand P3_R1269_U86 P3_R1269_U8 ; P3_R1269_U148
g25705 nand P3_U3100 P3_R1269_U45 ; P3_R1269_U149
g25706 nand P3_R1269_U87 P3_R1269_U149 ; P3_R1269_U150
g25707 nand P3_U3132 P3_R1269_U38 ; P3_R1269_U151
g25708 nand P3_U3131 P3_R1269_U47 ; P3_R1269_U152
g25709 nand P3_R1269_U147 P3_R1269_U88 ; P3_R1269_U153
g25710 nand P3_U3099 P3_R1269_U46 ; P3_R1269_U154
g25711 nand P3_R1269_U154 P3_R1269_U153 ; P3_R1269_U155
g25712 nand P3_R1269_U155 P3_R1269_U105 ; P3_R1269_U156
g25713 nand P3_U3098 P3_R1269_U15 ; P3_R1269_U157
g25714 not P3_R1269_U49 ; P3_R1269_U158
g25715 nand P3_U3129 P3_R1269_U158 ; P3_R1269_U159
g25716 nand P3_U3097 P3_R1269_U159 ; P3_R1269_U160
g25717 nand P3_R1269_U49 P3_R1269_U50 ; P3_R1269_U161
g25718 nand P3_U3096 P3_R1269_U54 ; P3_R1269_U162
g25719 nand P3_R1269_U90 P3_R1269_U160 P3_R1269_U91 ; P3_R1269_U163
g25720 nand P3_U3123 P3_R1269_U65 ; P3_R1269_U164
g25721 nand P3_U3124 P3_R1269_U63 ; P3_R1269_U165
g25722 nand P3_R1269_U92 P3_R1269_U104 ; P3_R1269_U166
g25723 nand P3_U3127 P3_R1269_U14 ; P3_R1269_U167
g25724 nand P3_R1269_U167 P3_R1269_U166 ; P3_R1269_U168
g25725 nand P3_R1269_U168 P3_R1269_U103 ; P3_R1269_U169
g25726 nand P3_U3126 P3_R1269_U13 ; P3_R1269_U170
g25727 nand P3_U3125 P3_R1269_U62 ; P3_R1269_U171
g25728 nand P3_R1269_U93 P3_R1269_U163 P3_R1269_U164 ; P3_R1269_U172
g25729 nand P3_U3087 P3_R1269_U67 ; P3_R1269_U173
g25730 nand P3_U3089 P3_R1269_U69 ; P3_R1269_U174
g25731 nand P3_U3088 P3_R1269_U66 ; P3_R1269_U175
g25732 nand P3_U3086 P3_R1269_U71 ; P3_R1269_U176
g25733 nand P3_R1269_U97 P3_R1269_U173 ; P3_R1269_U177
g25734 nand P3_U3119 P3_R1269_U58 ; P3_R1269_U178
g25735 not P3_R1269_U68 ; P3_R1269_U179
g25736 nand P3_U3121 P3_R1269_U59 ; P3_R1269_U180
g25737 nand P3_U3122 P3_R1269_U64 ; P3_R1269_U181
g25738 nand P3_R1269_U181 P3_R1269_U180 ; P3_R1269_U182
g25739 nand P3_R1269_U179 P3_R1269_U71 ; P3_R1269_U183
g25740 nand P3_R1269_U183 P3_R1269_U61 ; P3_R1269_U184
g25741 nand P3_R1269_U98 P3_R1269_U182 P3_R1269_U173 P3_R1269_U176 ; P3_R1269_U185
g25742 nand P3_U3118 P3_R1269_U68 ; P3_R1269_U186
g25743 nand P3_R1269_U9 P3_R1269_U101 ; P3_R1269_U187
g25744 nand P3_U3093 P3_R1269_U57 ; P3_R1269_U188
g25745 nand P3_U3092 P3_R1269_U53 ; P3_R1269_U189
g25746 nand P3_R1269_U189 P3_R1269_U188 ; P3_R1269_U190
g25747 nand P3_R1269_U165 P3_R1269_U190 P3_R1269_U164 ; P3_R1269_U191
g25748 nand P3_U3090 P3_R1269_U70 ; P3_R1269_U192
g25749 nand P3_U3091 P3_R1269_U52 ; P3_R1269_U193
g25750 nand P3_R1269_U102 P3_R1269_U95 ; P3_R1269_U194
g25751 nand P3_U3117 P3_R1269_U9 ; P3_R1269_U195
g25752 nand P3_R1269_U197 P3_R1269_U102 ; P3_R1269_U196
g25753 nand P3_R1269_U185 P3_R1269_U184 P3_R1269_U99 ; P3_R1269_U197
g25754 nand P3_U3117 P3_R1269_U101 ; P3_R1269_U198
g25755 nand P3_U3084 P3_R1269_U12 ; P3_R1269_U199
g25756 nand P3_U3116 P3_R1269_U100 ; P3_R1269_U200
g25757 nand P3_U3116 P3_R1269_U72 P3_R1269_U100 ; P3_R1269_U201
g25758 nand P3_U3149 P3_R1269_U12 P3_U3084 ; P3_R1269_U202
g25759 and P3_R1110_U179 P3_R1110_U178 ; P3_R1110_U4
g25760 and P3_R1110_U197 P3_R1110_U196 ; P3_R1110_U5
g25761 and P3_R1110_U237 P3_R1110_U236 ; P3_R1110_U6
g25762 and P3_R1110_U246 P3_R1110_U245 ; P3_R1110_U7
g25763 and P3_R1110_U264 P3_R1110_U263 ; P3_R1110_U8
g25764 and P3_R1110_U272 P3_R1110_U271 ; P3_R1110_U9
g25765 and P3_R1110_U351 P3_R1110_U348 ; P3_R1110_U10
g25766 and P3_R1110_U344 P3_R1110_U341 ; P3_R1110_U11
g25767 and P3_R1110_U335 P3_R1110_U332 ; P3_R1110_U12
g25768 and P3_R1110_U326 P3_R1110_U323 ; P3_R1110_U13
g25769 and P3_R1110_U320 P3_R1110_U318 ; P3_R1110_U14
g25770 and P3_R1110_U313 P3_R1110_U310 ; P3_R1110_U15
g25771 and P3_R1110_U235 P3_R1110_U232 ; P3_R1110_U16
g25772 and P3_R1110_U227 P3_R1110_U224 ; P3_R1110_U17
g25773 and P3_R1110_U213 P3_R1110_U210 ; P3_R1110_U18
g25774 not P3_U3407 ; P3_R1110_U19
g25775 not P3_U3070 ; P3_R1110_U20
g25776 not P3_U3069 ; P3_R1110_U21
g25777 nand P3_U3070 P3_U3407 ; P3_R1110_U22
g25778 not P3_U3410 ; P3_R1110_U23
g25779 not P3_U3401 ; P3_R1110_U24
g25780 not P3_U3059 ; P3_R1110_U25
g25781 not P3_U3066 ; P3_R1110_U26
g25782 not P3_U3395 ; P3_R1110_U27
g25783 not P3_U3067 ; P3_R1110_U28
g25784 not P3_U3387 ; P3_R1110_U29
g25785 not P3_U3076 ; P3_R1110_U30
g25786 nand P3_U3076 P3_U3387 ; P3_R1110_U31
g25787 not P3_U3398 ; P3_R1110_U32
g25788 not P3_U3063 ; P3_R1110_U33
g25789 nand P3_U3059 P3_U3401 ; P3_R1110_U34
g25790 not P3_U3404 ; P3_R1110_U35
g25791 not P3_U3413 ; P3_R1110_U36
g25792 not P3_U3083 ; P3_R1110_U37
g25793 not P3_U3082 ; P3_R1110_U38
g25794 not P3_U3416 ; P3_R1110_U39
g25795 nand P3_R1110_U61 P3_R1110_U205 ; P3_R1110_U40
g25796 nand P3_R1110_U117 P3_R1110_U193 ; P3_R1110_U41
g25797 nand P3_R1110_U182 P3_R1110_U183 ; P3_R1110_U42
g25798 nand P3_U3392 P3_U3077 ; P3_R1110_U43
g25799 nand P3_R1110_U122 P3_R1110_U219 ; P3_R1110_U44
g25800 nand P3_R1110_U216 P3_R1110_U215 ; P3_R1110_U45
g25801 not P3_U3900 ; P3_R1110_U46
g25802 not P3_U3052 ; P3_R1110_U47
g25803 not P3_U3056 ; P3_R1110_U48
g25804 not P3_U3901 ; P3_R1110_U49
g25805 not P3_U3902 ; P3_R1110_U50
g25806 not P3_U3057 ; P3_R1110_U51
g25807 not P3_U3903 ; P3_R1110_U52
g25808 not P3_U3064 ; P3_R1110_U53
g25809 not P3_U3906 ; P3_R1110_U54
g25810 not P3_U3074 ; P3_R1110_U55
g25811 not P3_U3437 ; P3_R1110_U56
g25812 not P3_U3072 ; P3_R1110_U57
g25813 not P3_U3068 ; P3_R1110_U58
g25814 nand P3_U3072 P3_U3437 ; P3_R1110_U59
g25815 not P3_U3440 ; P3_R1110_U60
g25816 nand P3_U3083 P3_U3413 ; P3_R1110_U61
g25817 not P3_U3419 ; P3_R1110_U62
g25818 not P3_U3061 ; P3_R1110_U63
g25819 not P3_U3425 ; P3_R1110_U64
g25820 not P3_U3071 ; P3_R1110_U65
g25821 not P3_U3422 ; P3_R1110_U66
g25822 not P3_U3062 ; P3_R1110_U67
g25823 nand P3_U3062 P3_U3422 ; P3_R1110_U68
g25824 not P3_U3428 ; P3_R1110_U69
g25825 not P3_U3079 ; P3_R1110_U70
g25826 not P3_U3431 ; P3_R1110_U71
g25827 not P3_U3078 ; P3_R1110_U72
g25828 not P3_U3434 ; P3_R1110_U73
g25829 not P3_U3073 ; P3_R1110_U74
g25830 not P3_U3443 ; P3_R1110_U75
g25831 not P3_U3081 ; P3_R1110_U76
g25832 nand P3_U3081 P3_U3443 ; P3_R1110_U77
g25833 not P3_U3445 ; P3_R1110_U78
g25834 not P3_U3080 ; P3_R1110_U79
g25835 nand P3_U3080 P3_U3445 ; P3_R1110_U80
g25836 not P3_U3907 ; P3_R1110_U81
g25837 not P3_U3905 ; P3_R1110_U82
g25838 not P3_U3060 ; P3_R1110_U83
g25839 not P3_U3904 ; P3_R1110_U84
g25840 not P3_U3065 ; P3_R1110_U85
g25841 nand P3_U3901 P3_U3056 ; P3_R1110_U86
g25842 not P3_U3053 ; P3_R1110_U87
g25843 not P3_U3899 ; P3_R1110_U88
g25844 nand P3_R1110_U306 P3_R1110_U176 ; P3_R1110_U89
g25845 not P3_U3075 ; P3_R1110_U90
g25846 nand P3_R1110_U77 P3_R1110_U315 ; P3_R1110_U91
g25847 nand P3_R1110_U261 P3_R1110_U260 ; P3_R1110_U92
g25848 nand P3_R1110_U68 P3_R1110_U337 ; P3_R1110_U93
g25849 nand P3_R1110_U457 P3_R1110_U456 ; P3_R1110_U94
g25850 nand P3_R1110_U504 P3_R1110_U503 ; P3_R1110_U95
g25851 nand P3_R1110_U375 P3_R1110_U374 ; P3_R1110_U96
g25852 nand P3_R1110_U380 P3_R1110_U379 ; P3_R1110_U97
g25853 nand P3_R1110_U387 P3_R1110_U386 ; P3_R1110_U98
g25854 nand P3_R1110_U394 P3_R1110_U393 ; P3_R1110_U99
g25855 nand P3_R1110_U399 P3_R1110_U398 ; P3_R1110_U100
g25856 nand P3_R1110_U408 P3_R1110_U407 ; P3_R1110_U101
g25857 nand P3_R1110_U415 P3_R1110_U414 ; P3_R1110_U102
g25858 nand P3_R1110_U422 P3_R1110_U421 ; P3_R1110_U103
g25859 nand P3_R1110_U429 P3_R1110_U428 ; P3_R1110_U104
g25860 nand P3_R1110_U434 P3_R1110_U433 ; P3_R1110_U105
g25861 nand P3_R1110_U441 P3_R1110_U440 ; P3_R1110_U106
g25862 nand P3_R1110_U448 P3_R1110_U447 ; P3_R1110_U107
g25863 nand P3_R1110_U462 P3_R1110_U461 ; P3_R1110_U108
g25864 nand P3_R1110_U467 P3_R1110_U466 ; P3_R1110_U109
g25865 nand P3_R1110_U474 P3_R1110_U473 ; P3_R1110_U110
g25866 nand P3_R1110_U481 P3_R1110_U480 ; P3_R1110_U111
g25867 nand P3_R1110_U488 P3_R1110_U487 ; P3_R1110_U112
g25868 nand P3_R1110_U495 P3_R1110_U494 ; P3_R1110_U113
g25869 nand P3_R1110_U500 P3_R1110_U499 ; P3_R1110_U114
g25870 and P3_R1110_U189 P3_R1110_U187 ; P3_R1110_U115
g25871 and P3_R1110_U4 P3_R1110_U180 ; P3_R1110_U116
g25872 and P3_R1110_U194 P3_R1110_U192 ; P3_R1110_U117
g25873 and P3_R1110_U201 P3_R1110_U200 ; P3_R1110_U118
g25874 and P3_R1110_U382 P3_R1110_U381 P3_R1110_U22 ; P3_R1110_U119
g25875 and P3_R1110_U212 P3_R1110_U5 ; P3_R1110_U120
g25876 and P3_R1110_U181 P3_R1110_U180 ; P3_R1110_U121
g25877 and P3_R1110_U220 P3_R1110_U218 ; P3_R1110_U122
g25878 and P3_R1110_U389 P3_R1110_U388 P3_R1110_U34 ; P3_R1110_U123
g25879 and P3_R1110_U226 P3_R1110_U4 ; P3_R1110_U124
g25880 and P3_R1110_U234 P3_R1110_U181 ; P3_R1110_U125
g25881 and P3_R1110_U204 P3_R1110_U6 ; P3_R1110_U126
g25882 and P3_R1110_U239 P3_R1110_U171 ; P3_R1110_U127
g25883 and P3_R1110_U250 P3_R1110_U7 ; P3_R1110_U128
g25884 and P3_R1110_U248 P3_R1110_U172 ; P3_R1110_U129
g25885 and P3_R1110_U268 P3_R1110_U267 ; P3_R1110_U130
g25886 and P3_R1110_U9 P3_R1110_U282 P3_R1110_U273 ; P3_R1110_U131
g25887 and P3_R1110_U285 P3_R1110_U280 ; P3_R1110_U132
g25888 and P3_R1110_U301 P3_R1110_U298 ; P3_R1110_U133
g25889 and P3_R1110_U368 P3_R1110_U302 ; P3_R1110_U134
g25890 and P3_R1110_U160 P3_R1110_U278 ; P3_R1110_U135
g25891 and P3_R1110_U455 P3_R1110_U454 P3_R1110_U80 ; P3_R1110_U136
g25892 and P3_R1110_U325 P3_R1110_U9 ; P3_R1110_U137
g25893 and P3_R1110_U469 P3_R1110_U468 P3_R1110_U59 ; P3_R1110_U138
g25894 and P3_R1110_U334 P3_R1110_U8 ; P3_R1110_U139
g25895 and P3_R1110_U490 P3_R1110_U489 P3_R1110_U172 ; P3_R1110_U140
g25896 and P3_R1110_U343 P3_R1110_U7 ; P3_R1110_U141
g25897 and P3_R1110_U502 P3_R1110_U501 P3_R1110_U171 ; P3_R1110_U142
g25898 and P3_R1110_U350 P3_R1110_U6 ; P3_R1110_U143
g25899 nand P3_R1110_U118 P3_R1110_U202 ; P3_R1110_U144
g25900 nand P3_R1110_U217 P3_R1110_U229 ; P3_R1110_U145
g25901 not P3_U3054 ; P3_R1110_U146
g25902 not P3_U3908 ; P3_R1110_U147
g25903 and P3_R1110_U403 P3_R1110_U402 ; P3_R1110_U148
g25904 nand P3_R1110_U304 P3_R1110_U169 P3_R1110_U364 ; P3_R1110_U149
g25905 and P3_R1110_U410 P3_R1110_U409 ; P3_R1110_U150
g25906 nand P3_R1110_U370 P3_R1110_U369 P3_R1110_U134 ; P3_R1110_U151
g25907 and P3_R1110_U417 P3_R1110_U416 ; P3_R1110_U152
g25908 nand P3_R1110_U365 P3_R1110_U299 P3_R1110_U86 ; P3_R1110_U153
g25909 and P3_R1110_U424 P3_R1110_U423 ; P3_R1110_U154
g25910 nand P3_R1110_U293 P3_R1110_U292 ; P3_R1110_U155
g25911 and P3_R1110_U436 P3_R1110_U435 ; P3_R1110_U156
g25912 nand P3_R1110_U289 P3_R1110_U288 ; P3_R1110_U157
g25913 and P3_R1110_U443 P3_R1110_U442 ; P3_R1110_U158
g25914 nand P3_R1110_U132 P3_R1110_U284 ; P3_R1110_U159
g25915 and P3_R1110_U450 P3_R1110_U449 ; P3_R1110_U160
g25916 nand P3_R1110_U43 P3_R1110_U327 ; P3_R1110_U161
g25917 nand P3_R1110_U130 P3_R1110_U269 ; P3_R1110_U162
g25918 and P3_R1110_U476 P3_R1110_U475 ; P3_R1110_U163
g25919 nand P3_R1110_U257 P3_R1110_U256 ; P3_R1110_U164
g25920 and P3_R1110_U483 P3_R1110_U482 ; P3_R1110_U165
g25921 nand P3_R1110_U253 P3_R1110_U252 ; P3_R1110_U166
g25922 nand P3_R1110_U243 P3_R1110_U242 ; P3_R1110_U167
g25923 nand P3_R1110_U367 P3_R1110_U366 ; P3_R1110_U168
g25924 nand P3_U3053 P3_R1110_U151 ; P3_R1110_U169
g25925 not P3_R1110_U34 ; P3_R1110_U170
g25926 nand P3_U3416 P3_U3082 ; P3_R1110_U171
g25927 nand P3_U3071 P3_U3425 ; P3_R1110_U172
g25928 nand P3_U3057 P3_U3902 ; P3_R1110_U173
g25929 not P3_R1110_U68 ; P3_R1110_U174
g25930 not P3_R1110_U77 ; P3_R1110_U175
g25931 nand P3_U3064 P3_U3903 ; P3_R1110_U176
g25932 not P3_R1110_U61 ; P3_R1110_U177
g25933 or P3_U3066 P3_U3404 ; P3_R1110_U178
g25934 or P3_U3059 P3_U3401 ; P3_R1110_U179
g25935 or P3_U3398 P3_U3063 ; P3_R1110_U180
g25936 or P3_U3395 P3_U3067 ; P3_R1110_U181
g25937 not P3_R1110_U31 ; P3_R1110_U182
g25938 or P3_U3392 P3_U3077 ; P3_R1110_U183
g25939 not P3_R1110_U42 ; P3_R1110_U184
g25940 not P3_R1110_U43 ; P3_R1110_U185
g25941 nand P3_R1110_U42 P3_R1110_U43 ; P3_R1110_U186
g25942 nand P3_U3067 P3_U3395 ; P3_R1110_U187
g25943 nand P3_R1110_U186 P3_R1110_U181 ; P3_R1110_U188
g25944 nand P3_U3063 P3_U3398 ; P3_R1110_U189
g25945 nand P3_R1110_U115 P3_R1110_U188 ; P3_R1110_U190
g25946 nand P3_R1110_U35 P3_R1110_U34 ; P3_R1110_U191
g25947 nand P3_U3066 P3_R1110_U191 ; P3_R1110_U192
g25948 nand P3_R1110_U116 P3_R1110_U190 ; P3_R1110_U193
g25949 nand P3_U3404 P3_R1110_U170 ; P3_R1110_U194
g25950 not P3_R1110_U41 ; P3_R1110_U195
g25951 or P3_U3069 P3_U3410 ; P3_R1110_U196
g25952 or P3_U3070 P3_U3407 ; P3_R1110_U197
g25953 not P3_R1110_U22 ; P3_R1110_U198
g25954 nand P3_R1110_U23 P3_R1110_U22 ; P3_R1110_U199
g25955 nand P3_U3069 P3_R1110_U199 ; P3_R1110_U200
g25956 nand P3_U3410 P3_R1110_U198 ; P3_R1110_U201
g25957 nand P3_R1110_U5 P3_R1110_U41 ; P3_R1110_U202
g25958 not P3_R1110_U144 ; P3_R1110_U203
g25959 or P3_U3413 P3_U3083 ; P3_R1110_U204
g25960 nand P3_R1110_U204 P3_R1110_U144 ; P3_R1110_U205
g25961 not P3_R1110_U40 ; P3_R1110_U206
g25962 or P3_U3082 P3_U3416 ; P3_R1110_U207
g25963 or P3_U3407 P3_U3070 ; P3_R1110_U208
g25964 nand P3_R1110_U208 P3_R1110_U41 ; P3_R1110_U209
g25965 nand P3_R1110_U119 P3_R1110_U209 ; P3_R1110_U210
g25966 nand P3_R1110_U195 P3_R1110_U22 ; P3_R1110_U211
g25967 nand P3_U3410 P3_U3069 ; P3_R1110_U212
g25968 nand P3_R1110_U120 P3_R1110_U211 ; P3_R1110_U213
g25969 or P3_U3070 P3_U3407 ; P3_R1110_U214
g25970 nand P3_R1110_U185 P3_R1110_U181 ; P3_R1110_U215
g25971 nand P3_U3067 P3_U3395 ; P3_R1110_U216
g25972 not P3_R1110_U45 ; P3_R1110_U217
g25973 nand P3_R1110_U121 P3_R1110_U184 ; P3_R1110_U218
g25974 nand P3_R1110_U45 P3_R1110_U180 ; P3_R1110_U219
g25975 nand P3_U3063 P3_U3398 ; P3_R1110_U220
g25976 not P3_R1110_U44 ; P3_R1110_U221
g25977 or P3_U3401 P3_U3059 ; P3_R1110_U222
g25978 nand P3_R1110_U222 P3_R1110_U44 ; P3_R1110_U223
g25979 nand P3_R1110_U123 P3_R1110_U223 ; P3_R1110_U224
g25980 nand P3_R1110_U221 P3_R1110_U34 ; P3_R1110_U225
g25981 nand P3_U3404 P3_U3066 ; P3_R1110_U226
g25982 nand P3_R1110_U124 P3_R1110_U225 ; P3_R1110_U227
g25983 or P3_U3059 P3_U3401 ; P3_R1110_U228
g25984 nand P3_R1110_U184 P3_R1110_U181 ; P3_R1110_U229
g25985 not P3_R1110_U145 ; P3_R1110_U230
g25986 nand P3_U3063 P3_U3398 ; P3_R1110_U231
g25987 nand P3_R1110_U401 P3_R1110_U400 P3_R1110_U43 P3_R1110_U42 ; P3_R1110_U232
g25988 nand P3_R1110_U43 P3_R1110_U42 ; P3_R1110_U233
g25989 nand P3_U3067 P3_U3395 ; P3_R1110_U234
g25990 nand P3_R1110_U125 P3_R1110_U233 ; P3_R1110_U235
g25991 or P3_U3082 P3_U3416 ; P3_R1110_U236
g25992 or P3_U3061 P3_U3419 ; P3_R1110_U237
g25993 nand P3_R1110_U177 P3_R1110_U6 ; P3_R1110_U238
g25994 nand P3_U3061 P3_U3419 ; P3_R1110_U239
g25995 nand P3_R1110_U127 P3_R1110_U238 ; P3_R1110_U240
g25996 or P3_U3419 P3_U3061 ; P3_R1110_U241
g25997 nand P3_R1110_U126 P3_R1110_U144 ; P3_R1110_U242
g25998 nand P3_R1110_U241 P3_R1110_U240 ; P3_R1110_U243
g25999 not P3_R1110_U167 ; P3_R1110_U244
g26000 or P3_U3079 P3_U3428 ; P3_R1110_U245
g26001 or P3_U3071 P3_U3425 ; P3_R1110_U246
g26002 nand P3_R1110_U174 P3_R1110_U7 ; P3_R1110_U247
g26003 nand P3_U3079 P3_U3428 ; P3_R1110_U248
g26004 nand P3_R1110_U129 P3_R1110_U247 ; P3_R1110_U249
g26005 or P3_U3422 P3_U3062 ; P3_R1110_U250
g26006 or P3_U3428 P3_U3079 ; P3_R1110_U251
g26007 nand P3_R1110_U128 P3_R1110_U167 ; P3_R1110_U252
g26008 nand P3_R1110_U251 P3_R1110_U249 ; P3_R1110_U253
g26009 not P3_R1110_U166 ; P3_R1110_U254
g26010 or P3_U3431 P3_U3078 ; P3_R1110_U255
g26011 nand P3_R1110_U255 P3_R1110_U166 ; P3_R1110_U256
g26012 nand P3_U3078 P3_U3431 ; P3_R1110_U257
g26013 not P3_R1110_U164 ; P3_R1110_U258
g26014 or P3_U3434 P3_U3073 ; P3_R1110_U259
g26015 nand P3_R1110_U259 P3_R1110_U164 ; P3_R1110_U260
g26016 nand P3_U3073 P3_U3434 ; P3_R1110_U261
g26017 not P3_R1110_U92 ; P3_R1110_U262
g26018 or P3_U3068 P3_U3440 ; P3_R1110_U263
g26019 or P3_U3072 P3_U3437 ; P3_R1110_U264
g26020 not P3_R1110_U59 ; P3_R1110_U265
g26021 nand P3_R1110_U60 P3_R1110_U59 ; P3_R1110_U266
g26022 nand P3_U3068 P3_R1110_U266 ; P3_R1110_U267
g26023 nand P3_U3440 P3_R1110_U265 ; P3_R1110_U268
g26024 nand P3_R1110_U8 P3_R1110_U92 ; P3_R1110_U269
g26025 not P3_R1110_U162 ; P3_R1110_U270
g26026 or P3_U3075 P3_U3907 ; P3_R1110_U271
g26027 or P3_U3080 P3_U3445 ; P3_R1110_U272
g26028 or P3_U3074 P3_U3906 ; P3_R1110_U273
g26029 not P3_R1110_U80 ; P3_R1110_U274
g26030 nand P3_U3907 P3_R1110_U274 ; P3_R1110_U275
g26031 nand P3_R1110_U275 P3_R1110_U90 ; P3_R1110_U276
g26032 nand P3_R1110_U80 P3_R1110_U81 ; P3_R1110_U277
g26033 nand P3_R1110_U277 P3_R1110_U276 ; P3_R1110_U278
g26034 nand P3_R1110_U175 P3_R1110_U9 ; P3_R1110_U279
g26035 nand P3_U3074 P3_U3906 ; P3_R1110_U280
g26036 nand P3_R1110_U278 P3_R1110_U279 ; P3_R1110_U281
g26037 or P3_U3443 P3_U3081 ; P3_R1110_U282
g26038 or P3_U3906 P3_U3074 ; P3_R1110_U283
g26039 nand P3_R1110_U162 P3_R1110_U131 ; P3_R1110_U284
g26040 nand P3_R1110_U283 P3_R1110_U281 ; P3_R1110_U285
g26041 not P3_R1110_U159 ; P3_R1110_U286
g26042 or P3_U3905 P3_U3060 ; P3_R1110_U287
g26043 nand P3_R1110_U287 P3_R1110_U159 ; P3_R1110_U288
g26044 nand P3_U3060 P3_U3905 ; P3_R1110_U289
g26045 not P3_R1110_U157 ; P3_R1110_U290
g26046 or P3_U3904 P3_U3065 ; P3_R1110_U291
g26047 nand P3_R1110_U291 P3_R1110_U157 ; P3_R1110_U292
g26048 nand P3_U3065 P3_U3904 ; P3_R1110_U293
g26049 not P3_R1110_U155 ; P3_R1110_U294
g26050 or P3_U3057 P3_U3902 ; P3_R1110_U295
g26051 nand P3_R1110_U176 P3_R1110_U173 ; P3_R1110_U296
g26052 not P3_R1110_U86 ; P3_R1110_U297
g26053 or P3_U3903 P3_U3064 ; P3_R1110_U298
g26054 nand P3_R1110_U155 P3_R1110_U298 P3_R1110_U168 ; P3_R1110_U299
g26055 not P3_R1110_U153 ; P3_R1110_U300
g26056 or P3_U3900 P3_U3052 ; P3_R1110_U301
g26057 nand P3_U3052 P3_U3900 ; P3_R1110_U302
g26058 not P3_R1110_U151 ; P3_R1110_U303
g26059 nand P3_U3899 P3_R1110_U151 ; P3_R1110_U304
g26060 not P3_R1110_U149 ; P3_R1110_U305
g26061 nand P3_R1110_U298 P3_R1110_U155 ; P3_R1110_U306
g26062 not P3_R1110_U89 ; P3_R1110_U307
g26063 or P3_U3902 P3_U3057 ; P3_R1110_U308
g26064 nand P3_R1110_U308 P3_R1110_U89 ; P3_R1110_U309
g26065 nand P3_R1110_U309 P3_R1110_U173 P3_R1110_U154 ; P3_R1110_U310
g26066 nand P3_R1110_U307 P3_R1110_U173 ; P3_R1110_U311
g26067 nand P3_U3901 P3_U3056 ; P3_R1110_U312
g26068 nand P3_R1110_U311 P3_R1110_U312 P3_R1110_U168 ; P3_R1110_U313
g26069 or P3_U3057 P3_U3902 ; P3_R1110_U314
g26070 nand P3_R1110_U282 P3_R1110_U162 ; P3_R1110_U315
g26071 not P3_R1110_U91 ; P3_R1110_U316
g26072 nand P3_R1110_U9 P3_R1110_U91 ; P3_R1110_U317
g26073 nand P3_R1110_U135 P3_R1110_U317 ; P3_R1110_U318
g26074 nand P3_R1110_U317 P3_R1110_U278 ; P3_R1110_U319
g26075 nand P3_R1110_U453 P3_R1110_U319 ; P3_R1110_U320
g26076 or P3_U3445 P3_U3080 ; P3_R1110_U321
g26077 nand P3_R1110_U321 P3_R1110_U91 ; P3_R1110_U322
g26078 nand P3_R1110_U136 P3_R1110_U322 ; P3_R1110_U323
g26079 nand P3_R1110_U316 P3_R1110_U80 ; P3_R1110_U324
g26080 nand P3_U3075 P3_U3907 ; P3_R1110_U325
g26081 nand P3_R1110_U137 P3_R1110_U324 ; P3_R1110_U326
g26082 or P3_U3392 P3_U3077 ; P3_R1110_U327
g26083 not P3_R1110_U161 ; P3_R1110_U328
g26084 or P3_U3080 P3_U3445 ; P3_R1110_U329
g26085 or P3_U3437 P3_U3072 ; P3_R1110_U330
g26086 nand P3_R1110_U330 P3_R1110_U92 ; P3_R1110_U331
g26087 nand P3_R1110_U138 P3_R1110_U331 ; P3_R1110_U332
g26088 nand P3_R1110_U262 P3_R1110_U59 ; P3_R1110_U333
g26089 nand P3_U3440 P3_U3068 ; P3_R1110_U334
g26090 nand P3_R1110_U139 P3_R1110_U333 ; P3_R1110_U335
g26091 or P3_U3072 P3_U3437 ; P3_R1110_U336
g26092 nand P3_R1110_U250 P3_R1110_U167 ; P3_R1110_U337
g26093 not P3_R1110_U93 ; P3_R1110_U338
g26094 or P3_U3425 P3_U3071 ; P3_R1110_U339
g26095 nand P3_R1110_U339 P3_R1110_U93 ; P3_R1110_U340
g26096 nand P3_R1110_U140 P3_R1110_U340 ; P3_R1110_U341
g26097 nand P3_R1110_U338 P3_R1110_U172 ; P3_R1110_U342
g26098 nand P3_U3079 P3_U3428 ; P3_R1110_U343
g26099 nand P3_R1110_U141 P3_R1110_U342 ; P3_R1110_U344
g26100 or P3_U3071 P3_U3425 ; P3_R1110_U345
g26101 or P3_U3416 P3_U3082 ; P3_R1110_U346
g26102 nand P3_R1110_U346 P3_R1110_U40 ; P3_R1110_U347
g26103 nand P3_R1110_U142 P3_R1110_U347 ; P3_R1110_U348
g26104 nand P3_R1110_U206 P3_R1110_U171 ; P3_R1110_U349
g26105 nand P3_U3061 P3_U3419 ; P3_R1110_U350
g26106 nand P3_R1110_U143 P3_R1110_U349 ; P3_R1110_U351
g26107 nand P3_R1110_U207 P3_R1110_U171 ; P3_R1110_U352
g26108 nand P3_R1110_U204 P3_R1110_U61 ; P3_R1110_U353
g26109 nand P3_R1110_U214 P3_R1110_U22 ; P3_R1110_U354
g26110 nand P3_R1110_U228 P3_R1110_U34 ; P3_R1110_U355
g26111 nand P3_R1110_U231 P3_R1110_U180 ; P3_R1110_U356
g26112 nand P3_R1110_U314 P3_R1110_U173 ; P3_R1110_U357
g26113 nand P3_R1110_U298 P3_R1110_U176 ; P3_R1110_U358
g26114 nand P3_R1110_U329 P3_R1110_U80 ; P3_R1110_U359
g26115 nand P3_R1110_U282 P3_R1110_U77 ; P3_R1110_U360
g26116 nand P3_R1110_U336 P3_R1110_U59 ; P3_R1110_U361
g26117 nand P3_R1110_U345 P3_R1110_U172 ; P3_R1110_U362
g26118 nand P3_R1110_U250 P3_R1110_U68 ; P3_R1110_U363
g26119 nand P3_U3899 P3_U3053 ; P3_R1110_U364
g26120 nand P3_R1110_U296 P3_R1110_U168 ; P3_R1110_U365
g26121 nand P3_U3056 P3_R1110_U295 ; P3_R1110_U366
g26122 nand P3_U3901 P3_R1110_U295 ; P3_R1110_U367
g26123 nand P3_R1110_U296 P3_R1110_U168 P3_R1110_U301 ; P3_R1110_U368
g26124 nand P3_R1110_U155 P3_R1110_U168 P3_R1110_U133 ; P3_R1110_U369
g26125 nand P3_R1110_U297 P3_R1110_U301 ; P3_R1110_U370
g26126 nand P3_U3082 P3_R1110_U39 ; P3_R1110_U371
g26127 nand P3_U3416 P3_R1110_U38 ; P3_R1110_U372
g26128 nand P3_R1110_U372 P3_R1110_U371 ; P3_R1110_U373
g26129 nand P3_R1110_U352 P3_R1110_U40 ; P3_R1110_U374
g26130 nand P3_R1110_U373 P3_R1110_U206 ; P3_R1110_U375
g26131 nand P3_U3083 P3_R1110_U36 ; P3_R1110_U376
g26132 nand P3_U3413 P3_R1110_U37 ; P3_R1110_U377
g26133 nand P3_R1110_U377 P3_R1110_U376 ; P3_R1110_U378
g26134 nand P3_R1110_U353 P3_R1110_U144 ; P3_R1110_U379
g26135 nand P3_R1110_U203 P3_R1110_U378 ; P3_R1110_U380
g26136 nand P3_U3069 P3_R1110_U23 ; P3_R1110_U381
g26137 nand P3_U3410 P3_R1110_U21 ; P3_R1110_U382
g26138 nand P3_U3070 P3_R1110_U19 ; P3_R1110_U383
g26139 nand P3_U3407 P3_R1110_U20 ; P3_R1110_U384
g26140 nand P3_R1110_U384 P3_R1110_U383 ; P3_R1110_U385
g26141 nand P3_R1110_U354 P3_R1110_U41 ; P3_R1110_U386
g26142 nand P3_R1110_U385 P3_R1110_U195 ; P3_R1110_U387
g26143 nand P3_U3066 P3_R1110_U35 ; P3_R1110_U388
g26144 nand P3_U3404 P3_R1110_U26 ; P3_R1110_U389
g26145 nand P3_U3059 P3_R1110_U24 ; P3_R1110_U390
g26146 nand P3_U3401 P3_R1110_U25 ; P3_R1110_U391
g26147 nand P3_R1110_U391 P3_R1110_U390 ; P3_R1110_U392
g26148 nand P3_R1110_U355 P3_R1110_U44 ; P3_R1110_U393
g26149 nand P3_R1110_U392 P3_R1110_U221 ; P3_R1110_U394
g26150 nand P3_U3063 P3_R1110_U32 ; P3_R1110_U395
g26151 nand P3_U3398 P3_R1110_U33 ; P3_R1110_U396
g26152 nand P3_R1110_U396 P3_R1110_U395 ; P3_R1110_U397
g26153 nand P3_R1110_U356 P3_R1110_U145 ; P3_R1110_U398
g26154 nand P3_R1110_U230 P3_R1110_U397 ; P3_R1110_U399
g26155 nand P3_U3067 P3_R1110_U27 ; P3_R1110_U400
g26156 nand P3_U3395 P3_R1110_U28 ; P3_R1110_U401
g26157 nand P3_U3054 P3_R1110_U147 ; P3_R1110_U402
g26158 nand P3_U3908 P3_R1110_U146 ; P3_R1110_U403
g26159 nand P3_U3054 P3_R1110_U147 ; P3_R1110_U404
g26160 nand P3_U3908 P3_R1110_U146 ; P3_R1110_U405
g26161 nand P3_R1110_U405 P3_R1110_U404 ; P3_R1110_U406
g26162 nand P3_R1110_U148 P3_R1110_U149 ; P3_R1110_U407
g26163 nand P3_R1110_U305 P3_R1110_U406 ; P3_R1110_U408
g26164 nand P3_U3053 P3_R1110_U88 ; P3_R1110_U409
g26165 nand P3_U3899 P3_R1110_U87 ; P3_R1110_U410
g26166 nand P3_U3053 P3_R1110_U88 ; P3_R1110_U411
g26167 nand P3_U3899 P3_R1110_U87 ; P3_R1110_U412
g26168 nand P3_R1110_U412 P3_R1110_U411 ; P3_R1110_U413
g26169 nand P3_R1110_U150 P3_R1110_U151 ; P3_R1110_U414
g26170 nand P3_R1110_U303 P3_R1110_U413 ; P3_R1110_U415
g26171 nand P3_U3052 P3_R1110_U46 ; P3_R1110_U416
g26172 nand P3_U3900 P3_R1110_U47 ; P3_R1110_U417
g26173 nand P3_U3052 P3_R1110_U46 ; P3_R1110_U418
g26174 nand P3_U3900 P3_R1110_U47 ; P3_R1110_U419
g26175 nand P3_R1110_U419 P3_R1110_U418 ; P3_R1110_U420
g26176 nand P3_R1110_U152 P3_R1110_U153 ; P3_R1110_U421
g26177 nand P3_R1110_U300 P3_R1110_U420 ; P3_R1110_U422
g26178 nand P3_U3056 P3_R1110_U49 ; P3_R1110_U423
g26179 nand P3_U3901 P3_R1110_U48 ; P3_R1110_U424
g26180 nand P3_U3057 P3_R1110_U50 ; P3_R1110_U425
g26181 nand P3_U3902 P3_R1110_U51 ; P3_R1110_U426
g26182 nand P3_R1110_U426 P3_R1110_U425 ; P3_R1110_U427
g26183 nand P3_R1110_U357 P3_R1110_U89 ; P3_R1110_U428
g26184 nand P3_R1110_U427 P3_R1110_U307 ; P3_R1110_U429
g26185 nand P3_U3064 P3_R1110_U52 ; P3_R1110_U430
g26186 nand P3_U3903 P3_R1110_U53 ; P3_R1110_U431
g26187 nand P3_R1110_U431 P3_R1110_U430 ; P3_R1110_U432
g26188 nand P3_R1110_U358 P3_R1110_U155 ; P3_R1110_U433
g26189 nand P3_R1110_U294 P3_R1110_U432 ; P3_R1110_U434
g26190 nand P3_U3065 P3_R1110_U84 ; P3_R1110_U435
g26191 nand P3_U3904 P3_R1110_U85 ; P3_R1110_U436
g26192 nand P3_U3065 P3_R1110_U84 ; P3_R1110_U437
g26193 nand P3_U3904 P3_R1110_U85 ; P3_R1110_U438
g26194 nand P3_R1110_U438 P3_R1110_U437 ; P3_R1110_U439
g26195 nand P3_R1110_U156 P3_R1110_U157 ; P3_R1110_U440
g26196 nand P3_R1110_U290 P3_R1110_U439 ; P3_R1110_U441
g26197 nand P3_U3060 P3_R1110_U82 ; P3_R1110_U442
g26198 nand P3_U3905 P3_R1110_U83 ; P3_R1110_U443
g26199 nand P3_U3060 P3_R1110_U82 ; P3_R1110_U444
g26200 nand P3_U3905 P3_R1110_U83 ; P3_R1110_U445
g26201 nand P3_R1110_U445 P3_R1110_U444 ; P3_R1110_U446
g26202 nand P3_R1110_U158 P3_R1110_U159 ; P3_R1110_U447
g26203 nand P3_R1110_U286 P3_R1110_U446 ; P3_R1110_U448
g26204 nand P3_U3074 P3_R1110_U54 ; P3_R1110_U449
g26205 nand P3_U3906 P3_R1110_U55 ; P3_R1110_U450
g26206 nand P3_U3074 P3_R1110_U54 ; P3_R1110_U451
g26207 nand P3_U3906 P3_R1110_U55 ; P3_R1110_U452
g26208 nand P3_R1110_U452 P3_R1110_U451 ; P3_R1110_U453
g26209 nand P3_U3075 P3_R1110_U81 ; P3_R1110_U454
g26210 nand P3_U3907 P3_R1110_U90 ; P3_R1110_U455
g26211 nand P3_R1110_U182 P3_R1110_U161 ; P3_R1110_U456
g26212 nand P3_R1110_U328 P3_R1110_U31 ; P3_R1110_U457
g26213 nand P3_U3080 P3_R1110_U78 ; P3_R1110_U458
g26214 nand P3_U3445 P3_R1110_U79 ; P3_R1110_U459
g26215 nand P3_R1110_U459 P3_R1110_U458 ; P3_R1110_U460
g26216 nand P3_R1110_U359 P3_R1110_U91 ; P3_R1110_U461
g26217 nand P3_R1110_U460 P3_R1110_U316 ; P3_R1110_U462
g26218 nand P3_U3081 P3_R1110_U75 ; P3_R1110_U463
g26219 nand P3_U3443 P3_R1110_U76 ; P3_R1110_U464
g26220 nand P3_R1110_U464 P3_R1110_U463 ; P3_R1110_U465
g26221 nand P3_R1110_U360 P3_R1110_U162 ; P3_R1110_U466
g26222 nand P3_R1110_U270 P3_R1110_U465 ; P3_R1110_U467
g26223 nand P3_U3068 P3_R1110_U60 ; P3_R1110_U468
g26224 nand P3_U3440 P3_R1110_U58 ; P3_R1110_U469
g26225 nand P3_U3072 P3_R1110_U56 ; P3_R1110_U470
g26226 nand P3_U3437 P3_R1110_U57 ; P3_R1110_U471
g26227 nand P3_R1110_U471 P3_R1110_U470 ; P3_R1110_U472
g26228 nand P3_R1110_U361 P3_R1110_U92 ; P3_R1110_U473
g26229 nand P3_R1110_U472 P3_R1110_U262 ; P3_R1110_U474
g26230 nand P3_U3073 P3_R1110_U73 ; P3_R1110_U475
g26231 nand P3_U3434 P3_R1110_U74 ; P3_R1110_U476
g26232 nand P3_U3073 P3_R1110_U73 ; P3_R1110_U477
g26233 nand P3_U3434 P3_R1110_U74 ; P3_R1110_U478
g26234 nand P3_R1110_U478 P3_R1110_U477 ; P3_R1110_U479
g26235 nand P3_R1110_U163 P3_R1110_U164 ; P3_R1110_U480
g26236 nand P3_R1110_U258 P3_R1110_U479 ; P3_R1110_U481
g26237 nand P3_U3078 P3_R1110_U71 ; P3_R1110_U482
g26238 nand P3_U3431 P3_R1110_U72 ; P3_R1110_U483
g26239 nand P3_U3078 P3_R1110_U71 ; P3_R1110_U484
g26240 nand P3_U3431 P3_R1110_U72 ; P3_R1110_U485
g26241 nand P3_R1110_U485 P3_R1110_U484 ; P3_R1110_U486
g26242 nand P3_R1110_U165 P3_R1110_U166 ; P3_R1110_U487
g26243 nand P3_R1110_U254 P3_R1110_U486 ; P3_R1110_U488
g26244 nand P3_U3079 P3_R1110_U69 ; P3_R1110_U489
g26245 nand P3_U3428 P3_R1110_U70 ; P3_R1110_U490
g26246 nand P3_U3071 P3_R1110_U64 ; P3_R1110_U491
g26247 nand P3_U3425 P3_R1110_U65 ; P3_R1110_U492
g26248 nand P3_R1110_U492 P3_R1110_U491 ; P3_R1110_U493
g26249 nand P3_R1110_U362 P3_R1110_U93 ; P3_R1110_U494
g26250 nand P3_R1110_U493 P3_R1110_U338 ; P3_R1110_U495
g26251 nand P3_U3062 P3_R1110_U66 ; P3_R1110_U496
g26252 nand P3_U3422 P3_R1110_U67 ; P3_R1110_U497
g26253 nand P3_R1110_U497 P3_R1110_U496 ; P3_R1110_U498
g26254 nand P3_R1110_U363 P3_R1110_U167 ; P3_R1110_U499
g26255 nand P3_R1110_U244 P3_R1110_U498 ; P3_R1110_U500
g26256 nand P3_U3061 P3_R1110_U62 ; P3_R1110_U501
g26257 nand P3_U3419 P3_R1110_U63 ; P3_R1110_U502
g26258 nand P3_U3076 P3_R1110_U29 ; P3_R1110_U503
g26259 nand P3_U3387 P3_R1110_U30 ; P3_R1110_U504
g26260 and P3_U3058 P3_R1297_U7 ; P3_R1297_U6
g26261 not P3_U3055 ; P3_R1297_U7
g26262 and P3_R1077_U179 P3_R1077_U178 ; P3_R1077_U4
g26263 and P3_R1077_U197 P3_R1077_U196 ; P3_R1077_U5
g26264 and P3_R1077_U237 P3_R1077_U236 ; P3_R1077_U6
g26265 and P3_R1077_U246 P3_R1077_U245 ; P3_R1077_U7
g26266 and P3_R1077_U264 P3_R1077_U263 ; P3_R1077_U8
g26267 and P3_R1077_U272 P3_R1077_U271 ; P3_R1077_U9
g26268 and P3_R1077_U351 P3_R1077_U348 ; P3_R1077_U10
g26269 and P3_R1077_U344 P3_R1077_U341 ; P3_R1077_U11
g26270 and P3_R1077_U335 P3_R1077_U332 ; P3_R1077_U12
g26271 and P3_R1077_U326 P3_R1077_U323 ; P3_R1077_U13
g26272 and P3_R1077_U320 P3_R1077_U318 ; P3_R1077_U14
g26273 and P3_R1077_U313 P3_R1077_U310 ; P3_R1077_U15
g26274 and P3_R1077_U235 P3_R1077_U232 ; P3_R1077_U16
g26275 and P3_R1077_U227 P3_R1077_U224 ; P3_R1077_U17
g26276 and P3_R1077_U213 P3_R1077_U210 ; P3_R1077_U18
g26277 not P3_U3407 ; P3_R1077_U19
g26278 not P3_U3070 ; P3_R1077_U20
g26279 not P3_U3069 ; P3_R1077_U21
g26280 nand P3_U3070 P3_U3407 ; P3_R1077_U22
g26281 not P3_U3410 ; P3_R1077_U23
g26282 not P3_U3401 ; P3_R1077_U24
g26283 not P3_U3059 ; P3_R1077_U25
g26284 not P3_U3066 ; P3_R1077_U26
g26285 not P3_U3395 ; P3_R1077_U27
g26286 not P3_U3067 ; P3_R1077_U28
g26287 not P3_U3387 ; P3_R1077_U29
g26288 not P3_U3076 ; P3_R1077_U30
g26289 nand P3_U3076 P3_U3387 ; P3_R1077_U31
g26290 not P3_U3398 ; P3_R1077_U32
g26291 not P3_U3063 ; P3_R1077_U33
g26292 nand P3_U3059 P3_U3401 ; P3_R1077_U34
g26293 not P3_U3404 ; P3_R1077_U35
g26294 not P3_U3413 ; P3_R1077_U36
g26295 not P3_U3083 ; P3_R1077_U37
g26296 not P3_U3082 ; P3_R1077_U38
g26297 not P3_U3416 ; P3_R1077_U39
g26298 nand P3_R1077_U61 P3_R1077_U205 ; P3_R1077_U40
g26299 nand P3_R1077_U117 P3_R1077_U193 ; P3_R1077_U41
g26300 nand P3_R1077_U182 P3_R1077_U183 ; P3_R1077_U42
g26301 nand P3_U3392 P3_U3077 ; P3_R1077_U43
g26302 nand P3_R1077_U122 P3_R1077_U219 ; P3_R1077_U44
g26303 nand P3_R1077_U216 P3_R1077_U215 ; P3_R1077_U45
g26304 not P3_U3900 ; P3_R1077_U46
g26305 not P3_U3052 ; P3_R1077_U47
g26306 not P3_U3056 ; P3_R1077_U48
g26307 not P3_U3901 ; P3_R1077_U49
g26308 not P3_U3902 ; P3_R1077_U50
g26309 not P3_U3057 ; P3_R1077_U51
g26310 not P3_U3903 ; P3_R1077_U52
g26311 not P3_U3064 ; P3_R1077_U53
g26312 not P3_U3906 ; P3_R1077_U54
g26313 not P3_U3074 ; P3_R1077_U55
g26314 not P3_U3437 ; P3_R1077_U56
g26315 not P3_U3072 ; P3_R1077_U57
g26316 not P3_U3068 ; P3_R1077_U58
g26317 nand P3_U3072 P3_U3437 ; P3_R1077_U59
g26318 not P3_U3440 ; P3_R1077_U60
g26319 nand P3_U3083 P3_U3413 ; P3_R1077_U61
g26320 not P3_U3419 ; P3_R1077_U62
g26321 not P3_U3061 ; P3_R1077_U63
g26322 not P3_U3425 ; P3_R1077_U64
g26323 not P3_U3071 ; P3_R1077_U65
g26324 not P3_U3422 ; P3_R1077_U66
g26325 not P3_U3062 ; P3_R1077_U67
g26326 nand P3_U3062 P3_U3422 ; P3_R1077_U68
g26327 not P3_U3428 ; P3_R1077_U69
g26328 not P3_U3079 ; P3_R1077_U70
g26329 not P3_U3431 ; P3_R1077_U71
g26330 not P3_U3078 ; P3_R1077_U72
g26331 not P3_U3434 ; P3_R1077_U73
g26332 not P3_U3073 ; P3_R1077_U74
g26333 not P3_U3443 ; P3_R1077_U75
g26334 not P3_U3081 ; P3_R1077_U76
g26335 nand P3_U3081 P3_U3443 ; P3_R1077_U77
g26336 not P3_U3445 ; P3_R1077_U78
g26337 not P3_U3080 ; P3_R1077_U79
g26338 nand P3_U3080 P3_U3445 ; P3_R1077_U80
g26339 not P3_U3907 ; P3_R1077_U81
g26340 not P3_U3905 ; P3_R1077_U82
g26341 not P3_U3060 ; P3_R1077_U83
g26342 not P3_U3904 ; P3_R1077_U84
g26343 not P3_U3065 ; P3_R1077_U85
g26344 nand P3_U3901 P3_U3056 ; P3_R1077_U86
g26345 not P3_U3053 ; P3_R1077_U87
g26346 not P3_U3899 ; P3_R1077_U88
g26347 nand P3_R1077_U306 P3_R1077_U176 ; P3_R1077_U89
g26348 not P3_U3075 ; P3_R1077_U90
g26349 nand P3_R1077_U77 P3_R1077_U315 ; P3_R1077_U91
g26350 nand P3_R1077_U261 P3_R1077_U260 ; P3_R1077_U92
g26351 nand P3_R1077_U68 P3_R1077_U337 ; P3_R1077_U93
g26352 nand P3_R1077_U457 P3_R1077_U456 ; P3_R1077_U94
g26353 nand P3_R1077_U504 P3_R1077_U503 ; P3_R1077_U95
g26354 nand P3_R1077_U375 P3_R1077_U374 ; P3_R1077_U96
g26355 nand P3_R1077_U380 P3_R1077_U379 ; P3_R1077_U97
g26356 nand P3_R1077_U387 P3_R1077_U386 ; P3_R1077_U98
g26357 nand P3_R1077_U394 P3_R1077_U393 ; P3_R1077_U99
g26358 nand P3_R1077_U399 P3_R1077_U398 ; P3_R1077_U100
g26359 nand P3_R1077_U408 P3_R1077_U407 ; P3_R1077_U101
g26360 nand P3_R1077_U415 P3_R1077_U414 ; P3_R1077_U102
g26361 nand P3_R1077_U422 P3_R1077_U421 ; P3_R1077_U103
g26362 nand P3_R1077_U429 P3_R1077_U428 ; P3_R1077_U104
g26363 nand P3_R1077_U434 P3_R1077_U433 ; P3_R1077_U105
g26364 nand P3_R1077_U441 P3_R1077_U440 ; P3_R1077_U106
g26365 nand P3_R1077_U448 P3_R1077_U447 ; P3_R1077_U107
g26366 nand P3_R1077_U462 P3_R1077_U461 ; P3_R1077_U108
g26367 nand P3_R1077_U467 P3_R1077_U466 ; P3_R1077_U109
g26368 nand P3_R1077_U474 P3_R1077_U473 ; P3_R1077_U110
g26369 nand P3_R1077_U481 P3_R1077_U480 ; P3_R1077_U111
g26370 nand P3_R1077_U488 P3_R1077_U487 ; P3_R1077_U112
g26371 nand P3_R1077_U495 P3_R1077_U494 ; P3_R1077_U113
g26372 nand P3_R1077_U500 P3_R1077_U499 ; P3_R1077_U114
g26373 and P3_R1077_U189 P3_R1077_U187 ; P3_R1077_U115
g26374 and P3_R1077_U4 P3_R1077_U180 ; P3_R1077_U116
g26375 and P3_R1077_U194 P3_R1077_U192 ; P3_R1077_U117
g26376 and P3_R1077_U201 P3_R1077_U200 ; P3_R1077_U118
g26377 and P3_R1077_U382 P3_R1077_U381 P3_R1077_U22 ; P3_R1077_U119
g26378 and P3_R1077_U212 P3_R1077_U5 ; P3_R1077_U120
g26379 and P3_R1077_U181 P3_R1077_U180 ; P3_R1077_U121
g26380 and P3_R1077_U220 P3_R1077_U218 ; P3_R1077_U122
g26381 and P3_R1077_U389 P3_R1077_U388 P3_R1077_U34 ; P3_R1077_U123
g26382 and P3_R1077_U226 P3_R1077_U4 ; P3_R1077_U124
g26383 and P3_R1077_U234 P3_R1077_U181 ; P3_R1077_U125
g26384 and P3_R1077_U204 P3_R1077_U6 ; P3_R1077_U126
g26385 and P3_R1077_U239 P3_R1077_U171 ; P3_R1077_U127
g26386 and P3_R1077_U250 P3_R1077_U7 ; P3_R1077_U128
g26387 and P3_R1077_U248 P3_R1077_U172 ; P3_R1077_U129
g26388 and P3_R1077_U268 P3_R1077_U267 ; P3_R1077_U130
g26389 and P3_R1077_U9 P3_R1077_U282 P3_R1077_U273 ; P3_R1077_U131
g26390 and P3_R1077_U285 P3_R1077_U280 ; P3_R1077_U132
g26391 and P3_R1077_U301 P3_R1077_U298 ; P3_R1077_U133
g26392 and P3_R1077_U368 P3_R1077_U302 ; P3_R1077_U134
g26393 and P3_R1077_U160 P3_R1077_U278 ; P3_R1077_U135
g26394 and P3_R1077_U455 P3_R1077_U454 P3_R1077_U80 ; P3_R1077_U136
g26395 and P3_R1077_U325 P3_R1077_U9 ; P3_R1077_U137
g26396 and P3_R1077_U469 P3_R1077_U468 P3_R1077_U59 ; P3_R1077_U138
g26397 and P3_R1077_U334 P3_R1077_U8 ; P3_R1077_U139
g26398 and P3_R1077_U490 P3_R1077_U489 P3_R1077_U172 ; P3_R1077_U140
g26399 and P3_R1077_U343 P3_R1077_U7 ; P3_R1077_U141
g26400 and P3_R1077_U502 P3_R1077_U501 P3_R1077_U171 ; P3_R1077_U142
g26401 and P3_R1077_U350 P3_R1077_U6 ; P3_R1077_U143
g26402 nand P3_R1077_U118 P3_R1077_U202 ; P3_R1077_U144
g26403 nand P3_R1077_U217 P3_R1077_U229 ; P3_R1077_U145
g26404 not P3_U3054 ; P3_R1077_U146
g26405 not P3_U3908 ; P3_R1077_U147
g26406 and P3_R1077_U403 P3_R1077_U402 ; P3_R1077_U148
g26407 nand P3_R1077_U304 P3_R1077_U169 P3_R1077_U364 ; P3_R1077_U149
g26408 and P3_R1077_U410 P3_R1077_U409 ; P3_R1077_U150
g26409 nand P3_R1077_U370 P3_R1077_U369 P3_R1077_U134 ; P3_R1077_U151
g26410 and P3_R1077_U417 P3_R1077_U416 ; P3_R1077_U152
g26411 nand P3_R1077_U365 P3_R1077_U299 P3_R1077_U86 ; P3_R1077_U153
g26412 and P3_R1077_U424 P3_R1077_U423 ; P3_R1077_U154
g26413 nand P3_R1077_U293 P3_R1077_U292 ; P3_R1077_U155
g26414 and P3_R1077_U436 P3_R1077_U435 ; P3_R1077_U156
g26415 nand P3_R1077_U289 P3_R1077_U288 ; P3_R1077_U157
g26416 and P3_R1077_U443 P3_R1077_U442 ; P3_R1077_U158
g26417 nand P3_R1077_U132 P3_R1077_U284 ; P3_R1077_U159
g26418 and P3_R1077_U450 P3_R1077_U449 ; P3_R1077_U160
g26419 nand P3_R1077_U43 P3_R1077_U327 ; P3_R1077_U161
g26420 nand P3_R1077_U130 P3_R1077_U269 ; P3_R1077_U162
g26421 and P3_R1077_U476 P3_R1077_U475 ; P3_R1077_U163
g26422 nand P3_R1077_U257 P3_R1077_U256 ; P3_R1077_U164
g26423 and P3_R1077_U483 P3_R1077_U482 ; P3_R1077_U165
g26424 nand P3_R1077_U253 P3_R1077_U252 ; P3_R1077_U166
g26425 nand P3_R1077_U243 P3_R1077_U242 ; P3_R1077_U167
g26426 nand P3_R1077_U367 P3_R1077_U366 ; P3_R1077_U168
g26427 nand P3_U3053 P3_R1077_U151 ; P3_R1077_U169
g26428 not P3_R1077_U34 ; P3_R1077_U170
g26429 nand P3_U3416 P3_U3082 ; P3_R1077_U171
g26430 nand P3_U3071 P3_U3425 ; P3_R1077_U172
g26431 nand P3_U3057 P3_U3902 ; P3_R1077_U173
g26432 not P3_R1077_U68 ; P3_R1077_U174
g26433 not P3_R1077_U77 ; P3_R1077_U175
g26434 nand P3_U3064 P3_U3903 ; P3_R1077_U176
g26435 not P3_R1077_U61 ; P3_R1077_U177
g26436 or P3_U3066 P3_U3404 ; P3_R1077_U178
g26437 or P3_U3059 P3_U3401 ; P3_R1077_U179
g26438 or P3_U3398 P3_U3063 ; P3_R1077_U180
g26439 or P3_U3395 P3_U3067 ; P3_R1077_U181
g26440 not P3_R1077_U31 ; P3_R1077_U182
g26441 or P3_U3392 P3_U3077 ; P3_R1077_U183
g26442 not P3_R1077_U42 ; P3_R1077_U184
g26443 not P3_R1077_U43 ; P3_R1077_U185
g26444 nand P3_R1077_U42 P3_R1077_U43 ; P3_R1077_U186
g26445 nand P3_U3067 P3_U3395 ; P3_R1077_U187
g26446 nand P3_R1077_U186 P3_R1077_U181 ; P3_R1077_U188
g26447 nand P3_U3063 P3_U3398 ; P3_R1077_U189
g26448 nand P3_R1077_U115 P3_R1077_U188 ; P3_R1077_U190
g26449 nand P3_R1077_U35 P3_R1077_U34 ; P3_R1077_U191
g26450 nand P3_U3066 P3_R1077_U191 ; P3_R1077_U192
g26451 nand P3_R1077_U116 P3_R1077_U190 ; P3_R1077_U193
g26452 nand P3_U3404 P3_R1077_U170 ; P3_R1077_U194
g26453 not P3_R1077_U41 ; P3_R1077_U195
g26454 or P3_U3069 P3_U3410 ; P3_R1077_U196
g26455 or P3_U3070 P3_U3407 ; P3_R1077_U197
g26456 not P3_R1077_U22 ; P3_R1077_U198
g26457 nand P3_R1077_U23 P3_R1077_U22 ; P3_R1077_U199
g26458 nand P3_U3069 P3_R1077_U199 ; P3_R1077_U200
g26459 nand P3_U3410 P3_R1077_U198 ; P3_R1077_U201
g26460 nand P3_R1077_U5 P3_R1077_U41 ; P3_R1077_U202
g26461 not P3_R1077_U144 ; P3_R1077_U203
g26462 or P3_U3413 P3_U3083 ; P3_R1077_U204
g26463 nand P3_R1077_U204 P3_R1077_U144 ; P3_R1077_U205
g26464 not P3_R1077_U40 ; P3_R1077_U206
g26465 or P3_U3082 P3_U3416 ; P3_R1077_U207
g26466 or P3_U3407 P3_U3070 ; P3_R1077_U208
g26467 nand P3_R1077_U208 P3_R1077_U41 ; P3_R1077_U209
g26468 nand P3_R1077_U119 P3_R1077_U209 ; P3_R1077_U210
g26469 nand P3_R1077_U195 P3_R1077_U22 ; P3_R1077_U211
g26470 nand P3_U3410 P3_U3069 ; P3_R1077_U212
g26471 nand P3_R1077_U120 P3_R1077_U211 ; P3_R1077_U213
g26472 or P3_U3070 P3_U3407 ; P3_R1077_U214
g26473 nand P3_R1077_U185 P3_R1077_U181 ; P3_R1077_U215
g26474 nand P3_U3067 P3_U3395 ; P3_R1077_U216
g26475 not P3_R1077_U45 ; P3_R1077_U217
g26476 nand P3_R1077_U121 P3_R1077_U184 ; P3_R1077_U218
g26477 nand P3_R1077_U45 P3_R1077_U180 ; P3_R1077_U219
g26478 nand P3_U3063 P3_U3398 ; P3_R1077_U220
g26479 not P3_R1077_U44 ; P3_R1077_U221
g26480 or P3_U3401 P3_U3059 ; P3_R1077_U222
g26481 nand P3_R1077_U222 P3_R1077_U44 ; P3_R1077_U223
g26482 nand P3_R1077_U123 P3_R1077_U223 ; P3_R1077_U224
g26483 nand P3_R1077_U221 P3_R1077_U34 ; P3_R1077_U225
g26484 nand P3_U3404 P3_U3066 ; P3_R1077_U226
g26485 nand P3_R1077_U124 P3_R1077_U225 ; P3_R1077_U227
g26486 or P3_U3059 P3_U3401 ; P3_R1077_U228
g26487 nand P3_R1077_U184 P3_R1077_U181 ; P3_R1077_U229
g26488 not P3_R1077_U145 ; P3_R1077_U230
g26489 nand P3_U3063 P3_U3398 ; P3_R1077_U231
g26490 nand P3_R1077_U401 P3_R1077_U400 P3_R1077_U43 P3_R1077_U42 ; P3_R1077_U232
g26491 nand P3_R1077_U43 P3_R1077_U42 ; P3_R1077_U233
g26492 nand P3_U3067 P3_U3395 ; P3_R1077_U234
g26493 nand P3_R1077_U125 P3_R1077_U233 ; P3_R1077_U235
g26494 or P3_U3082 P3_U3416 ; P3_R1077_U236
g26495 or P3_U3061 P3_U3419 ; P3_R1077_U237
g26496 nand P3_R1077_U177 P3_R1077_U6 ; P3_R1077_U238
g26497 nand P3_U3061 P3_U3419 ; P3_R1077_U239
g26498 nand P3_R1077_U127 P3_R1077_U238 ; P3_R1077_U240
g26499 or P3_U3419 P3_U3061 ; P3_R1077_U241
g26500 nand P3_R1077_U126 P3_R1077_U144 ; P3_R1077_U242
g26501 nand P3_R1077_U241 P3_R1077_U240 ; P3_R1077_U243
g26502 not P3_R1077_U167 ; P3_R1077_U244
g26503 or P3_U3079 P3_U3428 ; P3_R1077_U245
g26504 or P3_U3071 P3_U3425 ; P3_R1077_U246
g26505 nand P3_R1077_U174 P3_R1077_U7 ; P3_R1077_U247
g26506 nand P3_U3079 P3_U3428 ; P3_R1077_U248
g26507 nand P3_R1077_U129 P3_R1077_U247 ; P3_R1077_U249
g26508 or P3_U3422 P3_U3062 ; P3_R1077_U250
g26509 or P3_U3428 P3_U3079 ; P3_R1077_U251
g26510 nand P3_R1077_U128 P3_R1077_U167 ; P3_R1077_U252
g26511 nand P3_R1077_U251 P3_R1077_U249 ; P3_R1077_U253
g26512 not P3_R1077_U166 ; P3_R1077_U254
g26513 or P3_U3431 P3_U3078 ; P3_R1077_U255
g26514 nand P3_R1077_U255 P3_R1077_U166 ; P3_R1077_U256
g26515 nand P3_U3078 P3_U3431 ; P3_R1077_U257
g26516 not P3_R1077_U164 ; P3_R1077_U258
g26517 or P3_U3434 P3_U3073 ; P3_R1077_U259
g26518 nand P3_R1077_U259 P3_R1077_U164 ; P3_R1077_U260
g26519 nand P3_U3073 P3_U3434 ; P3_R1077_U261
g26520 not P3_R1077_U92 ; P3_R1077_U262
g26521 or P3_U3068 P3_U3440 ; P3_R1077_U263
g26522 or P3_U3072 P3_U3437 ; P3_R1077_U264
g26523 not P3_R1077_U59 ; P3_R1077_U265
g26524 nand P3_R1077_U60 P3_R1077_U59 ; P3_R1077_U266
g26525 nand P3_U3068 P3_R1077_U266 ; P3_R1077_U267
g26526 nand P3_U3440 P3_R1077_U265 ; P3_R1077_U268
g26527 nand P3_R1077_U8 P3_R1077_U92 ; P3_R1077_U269
g26528 not P3_R1077_U162 ; P3_R1077_U270
g26529 or P3_U3075 P3_U3907 ; P3_R1077_U271
g26530 or P3_U3080 P3_U3445 ; P3_R1077_U272
g26531 or P3_U3074 P3_U3906 ; P3_R1077_U273
g26532 not P3_R1077_U80 ; P3_R1077_U274
g26533 nand P3_U3907 P3_R1077_U274 ; P3_R1077_U275
g26534 nand P3_R1077_U275 P3_R1077_U90 ; P3_R1077_U276
g26535 nand P3_R1077_U80 P3_R1077_U81 ; P3_R1077_U277
g26536 nand P3_R1077_U277 P3_R1077_U276 ; P3_R1077_U278
g26537 nand P3_R1077_U175 P3_R1077_U9 ; P3_R1077_U279
g26538 nand P3_U3074 P3_U3906 ; P3_R1077_U280
g26539 nand P3_R1077_U278 P3_R1077_U279 ; P3_R1077_U281
g26540 or P3_U3443 P3_U3081 ; P3_R1077_U282
g26541 or P3_U3906 P3_U3074 ; P3_R1077_U283
g26542 nand P3_R1077_U162 P3_R1077_U131 ; P3_R1077_U284
g26543 nand P3_R1077_U283 P3_R1077_U281 ; P3_R1077_U285
g26544 not P3_R1077_U159 ; P3_R1077_U286
g26545 or P3_U3905 P3_U3060 ; P3_R1077_U287
g26546 nand P3_R1077_U287 P3_R1077_U159 ; P3_R1077_U288
g26547 nand P3_U3060 P3_U3905 ; P3_R1077_U289
g26548 not P3_R1077_U157 ; P3_R1077_U290
g26549 or P3_U3904 P3_U3065 ; P3_R1077_U291
g26550 nand P3_R1077_U291 P3_R1077_U157 ; P3_R1077_U292
g26551 nand P3_U3065 P3_U3904 ; P3_R1077_U293
g26552 not P3_R1077_U155 ; P3_R1077_U294
g26553 or P3_U3057 P3_U3902 ; P3_R1077_U295
g26554 nand P3_R1077_U176 P3_R1077_U173 ; P3_R1077_U296
g26555 not P3_R1077_U86 ; P3_R1077_U297
g26556 or P3_U3903 P3_U3064 ; P3_R1077_U298
g26557 nand P3_R1077_U155 P3_R1077_U298 P3_R1077_U168 ; P3_R1077_U299
g26558 not P3_R1077_U153 ; P3_R1077_U300
g26559 or P3_U3900 P3_U3052 ; P3_R1077_U301
g26560 nand P3_U3052 P3_U3900 ; P3_R1077_U302
g26561 not P3_R1077_U151 ; P3_R1077_U303
g26562 nand P3_U3899 P3_R1077_U151 ; P3_R1077_U304
g26563 not P3_R1077_U149 ; P3_R1077_U305
g26564 nand P3_R1077_U298 P3_R1077_U155 ; P3_R1077_U306
g26565 not P3_R1077_U89 ; P3_R1077_U307
g26566 or P3_U3902 P3_U3057 ; P3_R1077_U308
g26567 nand P3_R1077_U308 P3_R1077_U89 ; P3_R1077_U309
g26568 nand P3_R1077_U309 P3_R1077_U173 P3_R1077_U154 ; P3_R1077_U310
g26569 nand P3_R1077_U307 P3_R1077_U173 ; P3_R1077_U311
g26570 nand P3_U3901 P3_U3056 ; P3_R1077_U312
g26571 nand P3_R1077_U311 P3_R1077_U312 P3_R1077_U168 ; P3_R1077_U313
g26572 or P3_U3057 P3_U3902 ; P3_R1077_U314
g26573 nand P3_R1077_U282 P3_R1077_U162 ; P3_R1077_U315
g26574 not P3_R1077_U91 ; P3_R1077_U316
g26575 nand P3_R1077_U9 P3_R1077_U91 ; P3_R1077_U317
g26576 nand P3_R1077_U135 P3_R1077_U317 ; P3_R1077_U318
g26577 nand P3_R1077_U317 P3_R1077_U278 ; P3_R1077_U319
g26578 nand P3_R1077_U453 P3_R1077_U319 ; P3_R1077_U320
g26579 or P3_U3445 P3_U3080 ; P3_R1077_U321
g26580 nand P3_R1077_U321 P3_R1077_U91 ; P3_R1077_U322
g26581 nand P3_R1077_U136 P3_R1077_U322 ; P3_R1077_U323
g26582 nand P3_R1077_U316 P3_R1077_U80 ; P3_R1077_U324
g26583 nand P3_U3075 P3_U3907 ; P3_R1077_U325
g26584 nand P3_R1077_U137 P3_R1077_U324 ; P3_R1077_U326
g26585 or P3_U3392 P3_U3077 ; P3_R1077_U327
g26586 not P3_R1077_U161 ; P3_R1077_U328
g26587 or P3_U3080 P3_U3445 ; P3_R1077_U329
g26588 or P3_U3437 P3_U3072 ; P3_R1077_U330
g26589 nand P3_R1077_U330 P3_R1077_U92 ; P3_R1077_U331
g26590 nand P3_R1077_U138 P3_R1077_U331 ; P3_R1077_U332
g26591 nand P3_R1077_U262 P3_R1077_U59 ; P3_R1077_U333
g26592 nand P3_U3440 P3_U3068 ; P3_R1077_U334
g26593 nand P3_R1077_U139 P3_R1077_U333 ; P3_R1077_U335
g26594 or P3_U3072 P3_U3437 ; P3_R1077_U336
g26595 nand P3_R1077_U250 P3_R1077_U167 ; P3_R1077_U337
g26596 not P3_R1077_U93 ; P3_R1077_U338
g26597 or P3_U3425 P3_U3071 ; P3_R1077_U339
g26598 nand P3_R1077_U339 P3_R1077_U93 ; P3_R1077_U340
g26599 nand P3_R1077_U140 P3_R1077_U340 ; P3_R1077_U341
g26600 nand P3_R1077_U338 P3_R1077_U172 ; P3_R1077_U342
g26601 nand P3_U3079 P3_U3428 ; P3_R1077_U343
g26602 nand P3_R1077_U141 P3_R1077_U342 ; P3_R1077_U344
g26603 or P3_U3071 P3_U3425 ; P3_R1077_U345
g26604 or P3_U3416 P3_U3082 ; P3_R1077_U346
g26605 nand P3_R1077_U346 P3_R1077_U40 ; P3_R1077_U347
g26606 nand P3_R1077_U142 P3_R1077_U347 ; P3_R1077_U348
g26607 nand P3_R1077_U206 P3_R1077_U171 ; P3_R1077_U349
g26608 nand P3_U3061 P3_U3419 ; P3_R1077_U350
g26609 nand P3_R1077_U143 P3_R1077_U349 ; P3_R1077_U351
g26610 nand P3_R1077_U207 P3_R1077_U171 ; P3_R1077_U352
g26611 nand P3_R1077_U204 P3_R1077_U61 ; P3_R1077_U353
g26612 nand P3_R1077_U214 P3_R1077_U22 ; P3_R1077_U354
g26613 nand P3_R1077_U228 P3_R1077_U34 ; P3_R1077_U355
g26614 nand P3_R1077_U231 P3_R1077_U180 ; P3_R1077_U356
g26615 nand P3_R1077_U314 P3_R1077_U173 ; P3_R1077_U357
g26616 nand P3_R1077_U298 P3_R1077_U176 ; P3_R1077_U358
g26617 nand P3_R1077_U329 P3_R1077_U80 ; P3_R1077_U359
g26618 nand P3_R1077_U282 P3_R1077_U77 ; P3_R1077_U360
g26619 nand P3_R1077_U336 P3_R1077_U59 ; P3_R1077_U361
g26620 nand P3_R1077_U345 P3_R1077_U172 ; P3_R1077_U362
g26621 nand P3_R1077_U250 P3_R1077_U68 ; P3_R1077_U363
g26622 nand P3_U3899 P3_U3053 ; P3_R1077_U364
g26623 nand P3_R1077_U296 P3_R1077_U168 ; P3_R1077_U365
g26624 nand P3_U3056 P3_R1077_U295 ; P3_R1077_U366
g26625 nand P3_U3901 P3_R1077_U295 ; P3_R1077_U367
g26626 nand P3_R1077_U296 P3_R1077_U168 P3_R1077_U301 ; P3_R1077_U368
g26627 nand P3_R1077_U155 P3_R1077_U168 P3_R1077_U133 ; P3_R1077_U369
g26628 nand P3_R1077_U297 P3_R1077_U301 ; P3_R1077_U370
g26629 nand P3_U3082 P3_R1077_U39 ; P3_R1077_U371
g26630 nand P3_U3416 P3_R1077_U38 ; P3_R1077_U372
g26631 nand P3_R1077_U372 P3_R1077_U371 ; P3_R1077_U373
g26632 nand P3_R1077_U352 P3_R1077_U40 ; P3_R1077_U374
g26633 nand P3_R1077_U373 P3_R1077_U206 ; P3_R1077_U375
g26634 nand P3_U3083 P3_R1077_U36 ; P3_R1077_U376
g26635 nand P3_U3413 P3_R1077_U37 ; P3_R1077_U377
g26636 nand P3_R1077_U377 P3_R1077_U376 ; P3_R1077_U378
g26637 nand P3_R1077_U353 P3_R1077_U144 ; P3_R1077_U379
g26638 nand P3_R1077_U203 P3_R1077_U378 ; P3_R1077_U380
g26639 nand P3_U3069 P3_R1077_U23 ; P3_R1077_U381
g26640 nand P3_U3410 P3_R1077_U21 ; P3_R1077_U382
g26641 nand P3_U3070 P3_R1077_U19 ; P3_R1077_U383
g26642 nand P3_U3407 P3_R1077_U20 ; P3_R1077_U384
g26643 nand P3_R1077_U384 P3_R1077_U383 ; P3_R1077_U385
g26644 nand P3_R1077_U354 P3_R1077_U41 ; P3_R1077_U386
g26645 nand P3_R1077_U385 P3_R1077_U195 ; P3_R1077_U387
g26646 nand P3_U3066 P3_R1077_U35 ; P3_R1077_U388
g26647 nand P3_U3404 P3_R1077_U26 ; P3_R1077_U389
g26648 nand P3_U3059 P3_R1077_U24 ; P3_R1077_U390
g26649 nand P3_U3401 P3_R1077_U25 ; P3_R1077_U391
g26650 nand P3_R1077_U391 P3_R1077_U390 ; P3_R1077_U392
g26651 nand P3_R1077_U355 P3_R1077_U44 ; P3_R1077_U393
g26652 nand P3_R1077_U392 P3_R1077_U221 ; P3_R1077_U394
g26653 nand P3_U3063 P3_R1077_U32 ; P3_R1077_U395
g26654 nand P3_U3398 P3_R1077_U33 ; P3_R1077_U396
g26655 nand P3_R1077_U396 P3_R1077_U395 ; P3_R1077_U397
g26656 nand P3_R1077_U356 P3_R1077_U145 ; P3_R1077_U398
g26657 nand P3_R1077_U230 P3_R1077_U397 ; P3_R1077_U399
g26658 nand P3_U3067 P3_R1077_U27 ; P3_R1077_U400
g26659 nand P3_U3395 P3_R1077_U28 ; P3_R1077_U401
g26660 nand P3_U3054 P3_R1077_U147 ; P3_R1077_U402
g26661 nand P3_U3908 P3_R1077_U146 ; P3_R1077_U403
g26662 nand P3_U3054 P3_R1077_U147 ; P3_R1077_U404
g26663 nand P3_U3908 P3_R1077_U146 ; P3_R1077_U405
g26664 nand P3_R1077_U405 P3_R1077_U404 ; P3_R1077_U406
g26665 nand P3_R1077_U148 P3_R1077_U149 ; P3_R1077_U407
g26666 nand P3_R1077_U305 P3_R1077_U406 ; P3_R1077_U408
g26667 nand P3_U3053 P3_R1077_U88 ; P3_R1077_U409
g26668 nand P3_U3899 P3_R1077_U87 ; P3_R1077_U410
g26669 nand P3_U3053 P3_R1077_U88 ; P3_R1077_U411
g26670 nand P3_U3899 P3_R1077_U87 ; P3_R1077_U412
g26671 nand P3_R1077_U412 P3_R1077_U411 ; P3_R1077_U413
g26672 nand P3_R1077_U150 P3_R1077_U151 ; P3_R1077_U414
g26673 nand P3_R1077_U303 P3_R1077_U413 ; P3_R1077_U415
g26674 nand P3_U3052 P3_R1077_U46 ; P3_R1077_U416
g26675 nand P3_U3900 P3_R1077_U47 ; P3_R1077_U417
g26676 nand P3_U3052 P3_R1077_U46 ; P3_R1077_U418
g26677 nand P3_U3900 P3_R1077_U47 ; P3_R1077_U419
g26678 nand P3_R1077_U419 P3_R1077_U418 ; P3_R1077_U420
g26679 nand P3_R1077_U152 P3_R1077_U153 ; P3_R1077_U421
g26680 nand P3_R1077_U300 P3_R1077_U420 ; P3_R1077_U422
g26681 nand P3_U3056 P3_R1077_U49 ; P3_R1077_U423
g26682 nand P3_U3901 P3_R1077_U48 ; P3_R1077_U424
g26683 nand P3_U3057 P3_R1077_U50 ; P3_R1077_U425
g26684 nand P3_U3902 P3_R1077_U51 ; P3_R1077_U426
g26685 nand P3_R1077_U426 P3_R1077_U425 ; P3_R1077_U427
g26686 nand P3_R1077_U357 P3_R1077_U89 ; P3_R1077_U428
g26687 nand P3_R1077_U427 P3_R1077_U307 ; P3_R1077_U429
g26688 nand P3_U3064 P3_R1077_U52 ; P3_R1077_U430
g26689 nand P3_U3903 P3_R1077_U53 ; P3_R1077_U431
g26690 nand P3_R1077_U431 P3_R1077_U430 ; P3_R1077_U432
g26691 nand P3_R1077_U358 P3_R1077_U155 ; P3_R1077_U433
g26692 nand P3_R1077_U294 P3_R1077_U432 ; P3_R1077_U434
g26693 nand P3_U3065 P3_R1077_U84 ; P3_R1077_U435
g26694 nand P3_U3904 P3_R1077_U85 ; P3_R1077_U436
g26695 nand P3_U3065 P3_R1077_U84 ; P3_R1077_U437
g26696 nand P3_U3904 P3_R1077_U85 ; P3_R1077_U438
g26697 nand P3_R1077_U438 P3_R1077_U437 ; P3_R1077_U439
g26698 nand P3_R1077_U156 P3_R1077_U157 ; P3_R1077_U440
g26699 nand P3_R1077_U290 P3_R1077_U439 ; P3_R1077_U441
g26700 nand P3_U3060 P3_R1077_U82 ; P3_R1077_U442
g26701 nand P3_U3905 P3_R1077_U83 ; P3_R1077_U443
g26702 nand P3_U3060 P3_R1077_U82 ; P3_R1077_U444
g26703 nand P3_U3905 P3_R1077_U83 ; P3_R1077_U445
g26704 nand P3_R1077_U445 P3_R1077_U444 ; P3_R1077_U446
g26705 nand P3_R1077_U158 P3_R1077_U159 ; P3_R1077_U447
g26706 nand P3_R1077_U286 P3_R1077_U446 ; P3_R1077_U448
g26707 nand P3_U3074 P3_R1077_U54 ; P3_R1077_U449
g26708 nand P3_U3906 P3_R1077_U55 ; P3_R1077_U450
g26709 nand P3_U3074 P3_R1077_U54 ; P3_R1077_U451
g26710 nand P3_U3906 P3_R1077_U55 ; P3_R1077_U452
g26711 nand P3_R1077_U452 P3_R1077_U451 ; P3_R1077_U453
g26712 nand P3_U3075 P3_R1077_U81 ; P3_R1077_U454
g26713 nand P3_U3907 P3_R1077_U90 ; P3_R1077_U455
g26714 nand P3_R1077_U182 P3_R1077_U161 ; P3_R1077_U456
g26715 nand P3_R1077_U328 P3_R1077_U31 ; P3_R1077_U457
g26716 nand P3_U3080 P3_R1077_U78 ; P3_R1077_U458
g26717 nand P3_U3445 P3_R1077_U79 ; P3_R1077_U459
g26718 nand P3_R1077_U459 P3_R1077_U458 ; P3_R1077_U460
g26719 nand P3_R1077_U359 P3_R1077_U91 ; P3_R1077_U461
g26720 nand P3_R1077_U460 P3_R1077_U316 ; P3_R1077_U462
g26721 nand P3_U3081 P3_R1077_U75 ; P3_R1077_U463
g26722 nand P3_U3443 P3_R1077_U76 ; P3_R1077_U464
g26723 nand P3_R1077_U464 P3_R1077_U463 ; P3_R1077_U465
g26724 nand P3_R1077_U360 P3_R1077_U162 ; P3_R1077_U466
g26725 nand P3_R1077_U270 P3_R1077_U465 ; P3_R1077_U467
g26726 nand P3_U3068 P3_R1077_U60 ; P3_R1077_U468
g26727 nand P3_U3440 P3_R1077_U58 ; P3_R1077_U469
g26728 nand P3_U3072 P3_R1077_U56 ; P3_R1077_U470
g26729 nand P3_U3437 P3_R1077_U57 ; P3_R1077_U471
g26730 nand P3_R1077_U471 P3_R1077_U470 ; P3_R1077_U472
g26731 nand P3_R1077_U361 P3_R1077_U92 ; P3_R1077_U473
g26732 nand P3_R1077_U472 P3_R1077_U262 ; P3_R1077_U474
g26733 nand P3_U3073 P3_R1077_U73 ; P3_R1077_U475
g26734 nand P3_U3434 P3_R1077_U74 ; P3_R1077_U476
g26735 nand P3_U3073 P3_R1077_U73 ; P3_R1077_U477
g26736 nand P3_U3434 P3_R1077_U74 ; P3_R1077_U478
g26737 nand P3_R1077_U478 P3_R1077_U477 ; P3_R1077_U479
g26738 nand P3_R1077_U163 P3_R1077_U164 ; P3_R1077_U480
g26739 nand P3_R1077_U258 P3_R1077_U479 ; P3_R1077_U481
g26740 nand P3_U3078 P3_R1077_U71 ; P3_R1077_U482
g26741 nand P3_U3431 P3_R1077_U72 ; P3_R1077_U483
g26742 nand P3_U3078 P3_R1077_U71 ; P3_R1077_U484
g26743 nand P3_U3431 P3_R1077_U72 ; P3_R1077_U485
g26744 nand P3_R1077_U485 P3_R1077_U484 ; P3_R1077_U486
g26745 nand P3_R1077_U165 P3_R1077_U166 ; P3_R1077_U487
g26746 nand P3_R1077_U254 P3_R1077_U486 ; P3_R1077_U488
g26747 nand P3_U3079 P3_R1077_U69 ; P3_R1077_U489
g26748 nand P3_U3428 P3_R1077_U70 ; P3_R1077_U490
g26749 nand P3_U3071 P3_R1077_U64 ; P3_R1077_U491
g26750 nand P3_U3425 P3_R1077_U65 ; P3_R1077_U492
g26751 nand P3_R1077_U492 P3_R1077_U491 ; P3_R1077_U493
g26752 nand P3_R1077_U362 P3_R1077_U93 ; P3_R1077_U494
g26753 nand P3_R1077_U493 P3_R1077_U338 ; P3_R1077_U495
g26754 nand P3_U3062 P3_R1077_U66 ; P3_R1077_U496
g26755 nand P3_U3422 P3_R1077_U67 ; P3_R1077_U497
g26756 nand P3_R1077_U497 P3_R1077_U496 ; P3_R1077_U498
g26757 nand P3_R1077_U363 P3_R1077_U167 ; P3_R1077_U499
g26758 nand P3_R1077_U244 P3_R1077_U498 ; P3_R1077_U500
g26759 nand P3_U3061 P3_R1077_U62 ; P3_R1077_U501
g26760 nand P3_U3419 P3_R1077_U63 ; P3_R1077_U502
g26761 nand P3_U3076 P3_R1077_U29 ; P3_R1077_U503
g26762 nand P3_U3387 P3_R1077_U30 ; P3_R1077_U504
g26763 and P3_R1143_U179 P3_R1143_U178 ; P3_R1143_U4
g26764 and P3_R1143_U197 P3_R1143_U196 ; P3_R1143_U5
g26765 and P3_R1143_U237 P3_R1143_U236 ; P3_R1143_U6
g26766 and P3_R1143_U246 P3_R1143_U245 ; P3_R1143_U7
g26767 and P3_R1143_U264 P3_R1143_U263 ; P3_R1143_U8
g26768 and P3_R1143_U272 P3_R1143_U271 ; P3_R1143_U9
g26769 and P3_R1143_U351 P3_R1143_U348 ; P3_R1143_U10
g26770 and P3_R1143_U344 P3_R1143_U341 ; P3_R1143_U11
g26771 and P3_R1143_U335 P3_R1143_U332 ; P3_R1143_U12
g26772 and P3_R1143_U326 P3_R1143_U323 ; P3_R1143_U13
g26773 and P3_R1143_U320 P3_R1143_U318 ; P3_R1143_U14
g26774 and P3_R1143_U313 P3_R1143_U310 ; P3_R1143_U15
g26775 and P3_R1143_U235 P3_R1143_U232 ; P3_R1143_U16
g26776 and P3_R1143_U227 P3_R1143_U224 ; P3_R1143_U17
g26777 and P3_R1143_U213 P3_R1143_U210 ; P3_R1143_U18
g26778 not P3_U3407 ; P3_R1143_U19
g26779 not P3_U3070 ; P3_R1143_U20
g26780 not P3_U3069 ; P3_R1143_U21
g26781 nand P3_U3070 P3_U3407 ; P3_R1143_U22
g26782 not P3_U3410 ; P3_R1143_U23
g26783 not P3_U3401 ; P3_R1143_U24
g26784 not P3_U3059 ; P3_R1143_U25
g26785 not P3_U3066 ; P3_R1143_U26
g26786 not P3_U3395 ; P3_R1143_U27
g26787 not P3_U3067 ; P3_R1143_U28
g26788 not P3_U3387 ; P3_R1143_U29
g26789 not P3_U3076 ; P3_R1143_U30
g26790 nand P3_U3076 P3_U3387 ; P3_R1143_U31
g26791 not P3_U3398 ; P3_R1143_U32
g26792 not P3_U3063 ; P3_R1143_U33
g26793 nand P3_U3059 P3_U3401 ; P3_R1143_U34
g26794 not P3_U3404 ; P3_R1143_U35
g26795 not P3_U3413 ; P3_R1143_U36
g26796 not P3_U3083 ; P3_R1143_U37
g26797 not P3_U3082 ; P3_R1143_U38
g26798 not P3_U3416 ; P3_R1143_U39
g26799 nand P3_R1143_U63 P3_R1143_U205 ; P3_R1143_U40
g26800 nand P3_R1143_U117 P3_R1143_U193 ; P3_R1143_U41
g26801 nand P3_R1143_U182 P3_R1143_U183 ; P3_R1143_U42
g26802 nand P3_U3392 P3_U3077 ; P3_R1143_U43
g26803 nand P3_R1143_U122 P3_R1143_U219 ; P3_R1143_U44
g26804 nand P3_R1143_U216 P3_R1143_U215 ; P3_R1143_U45
g26805 not P3_U3900 ; P3_R1143_U46
g26806 not P3_U3052 ; P3_R1143_U47
g26807 not P3_U3056 ; P3_R1143_U48
g26808 not P3_U3901 ; P3_R1143_U49
g26809 not P3_U3902 ; P3_R1143_U50
g26810 not P3_U3057 ; P3_R1143_U51
g26811 not P3_U3903 ; P3_R1143_U52
g26812 not P3_U3064 ; P3_R1143_U53
g26813 not P3_U3906 ; P3_R1143_U54
g26814 not P3_U3074 ; P3_R1143_U55
g26815 not P3_U3437 ; P3_R1143_U56
g26816 not P3_U3072 ; P3_R1143_U57
g26817 not P3_U3068 ; P3_R1143_U58
g26818 nand P3_U3072 P3_U3437 ; P3_R1143_U59
g26819 not P3_U3440 ; P3_R1143_U60
g26820 not P3_U3419 ; P3_R1143_U61
g26821 not P3_U3061 ; P3_R1143_U62
g26822 nand P3_U3083 P3_U3413 ; P3_R1143_U63
g26823 not P3_U3425 ; P3_R1143_U64
g26824 not P3_U3071 ; P3_R1143_U65
g26825 not P3_U3422 ; P3_R1143_U66
g26826 not P3_U3062 ; P3_R1143_U67
g26827 nand P3_U3062 P3_U3422 ; P3_R1143_U68
g26828 not P3_U3428 ; P3_R1143_U69
g26829 not P3_U3079 ; P3_R1143_U70
g26830 not P3_U3431 ; P3_R1143_U71
g26831 not P3_U3078 ; P3_R1143_U72
g26832 not P3_U3434 ; P3_R1143_U73
g26833 not P3_U3073 ; P3_R1143_U74
g26834 not P3_U3443 ; P3_R1143_U75
g26835 not P3_U3081 ; P3_R1143_U76
g26836 nand P3_U3081 P3_U3443 ; P3_R1143_U77
g26837 not P3_U3445 ; P3_R1143_U78
g26838 not P3_U3080 ; P3_R1143_U79
g26839 nand P3_U3080 P3_U3445 ; P3_R1143_U80
g26840 not P3_U3907 ; P3_R1143_U81
g26841 not P3_U3905 ; P3_R1143_U82
g26842 not P3_U3060 ; P3_R1143_U83
g26843 not P3_U3904 ; P3_R1143_U84
g26844 not P3_U3065 ; P3_R1143_U85
g26845 nand P3_U3901 P3_U3056 ; P3_R1143_U86
g26846 not P3_U3053 ; P3_R1143_U87
g26847 not P3_U3899 ; P3_R1143_U88
g26848 nand P3_R1143_U306 P3_R1143_U176 ; P3_R1143_U89
g26849 not P3_U3075 ; P3_R1143_U90
g26850 nand P3_R1143_U77 P3_R1143_U315 ; P3_R1143_U91
g26851 nand P3_R1143_U261 P3_R1143_U260 ; P3_R1143_U92
g26852 nand P3_R1143_U68 P3_R1143_U337 ; P3_R1143_U93
g26853 nand P3_R1143_U457 P3_R1143_U456 ; P3_R1143_U94
g26854 nand P3_R1143_U504 P3_R1143_U503 ; P3_R1143_U95
g26855 nand P3_R1143_U375 P3_R1143_U374 ; P3_R1143_U96
g26856 nand P3_R1143_U380 P3_R1143_U379 ; P3_R1143_U97
g26857 nand P3_R1143_U387 P3_R1143_U386 ; P3_R1143_U98
g26858 nand P3_R1143_U394 P3_R1143_U393 ; P3_R1143_U99
g26859 nand P3_R1143_U399 P3_R1143_U398 ; P3_R1143_U100
g26860 nand P3_R1143_U408 P3_R1143_U407 ; P3_R1143_U101
g26861 nand P3_R1143_U415 P3_R1143_U414 ; P3_R1143_U102
g26862 nand P3_R1143_U422 P3_R1143_U421 ; P3_R1143_U103
g26863 nand P3_R1143_U429 P3_R1143_U428 ; P3_R1143_U104
g26864 nand P3_R1143_U434 P3_R1143_U433 ; P3_R1143_U105
g26865 nand P3_R1143_U441 P3_R1143_U440 ; P3_R1143_U106
g26866 nand P3_R1143_U448 P3_R1143_U447 ; P3_R1143_U107
g26867 nand P3_R1143_U462 P3_R1143_U461 ; P3_R1143_U108
g26868 nand P3_R1143_U467 P3_R1143_U466 ; P3_R1143_U109
g26869 nand P3_R1143_U474 P3_R1143_U473 ; P3_R1143_U110
g26870 nand P3_R1143_U481 P3_R1143_U480 ; P3_R1143_U111
g26871 nand P3_R1143_U488 P3_R1143_U487 ; P3_R1143_U112
g26872 nand P3_R1143_U495 P3_R1143_U494 ; P3_R1143_U113
g26873 nand P3_R1143_U500 P3_R1143_U499 ; P3_R1143_U114
g26874 and P3_R1143_U189 P3_R1143_U187 ; P3_R1143_U115
g26875 and P3_R1143_U4 P3_R1143_U180 ; P3_R1143_U116
g26876 and P3_R1143_U194 P3_R1143_U192 ; P3_R1143_U117
g26877 and P3_R1143_U201 P3_R1143_U200 ; P3_R1143_U118
g26878 and P3_R1143_U382 P3_R1143_U381 P3_R1143_U22 ; P3_R1143_U119
g26879 and P3_R1143_U212 P3_R1143_U5 ; P3_R1143_U120
g26880 and P3_R1143_U181 P3_R1143_U180 ; P3_R1143_U121
g26881 and P3_R1143_U220 P3_R1143_U218 ; P3_R1143_U122
g26882 and P3_R1143_U389 P3_R1143_U388 P3_R1143_U34 ; P3_R1143_U123
g26883 and P3_R1143_U226 P3_R1143_U4 ; P3_R1143_U124
g26884 and P3_R1143_U234 P3_R1143_U181 ; P3_R1143_U125
g26885 and P3_R1143_U204 P3_R1143_U6 ; P3_R1143_U126
g26886 and P3_R1143_U243 P3_R1143_U239 ; P3_R1143_U127
g26887 and P3_R1143_U250 P3_R1143_U7 ; P3_R1143_U128
g26888 and P3_R1143_U248 P3_R1143_U172 ; P3_R1143_U129
g26889 and P3_R1143_U268 P3_R1143_U267 ; P3_R1143_U130
g26890 and P3_R1143_U9 P3_R1143_U282 P3_R1143_U273 ; P3_R1143_U131
g26891 and P3_R1143_U285 P3_R1143_U280 ; P3_R1143_U132
g26892 and P3_R1143_U301 P3_R1143_U298 ; P3_R1143_U133
g26893 and P3_R1143_U368 P3_R1143_U302 ; P3_R1143_U134
g26894 and P3_R1143_U160 P3_R1143_U278 ; P3_R1143_U135
g26895 and P3_R1143_U455 P3_R1143_U454 P3_R1143_U80 ; P3_R1143_U136
g26896 and P3_R1143_U325 P3_R1143_U9 ; P3_R1143_U137
g26897 and P3_R1143_U469 P3_R1143_U468 P3_R1143_U59 ; P3_R1143_U138
g26898 and P3_R1143_U334 P3_R1143_U8 ; P3_R1143_U139
g26899 and P3_R1143_U490 P3_R1143_U489 P3_R1143_U172 ; P3_R1143_U140
g26900 and P3_R1143_U343 P3_R1143_U7 ; P3_R1143_U141
g26901 and P3_R1143_U502 P3_R1143_U501 P3_R1143_U171 ; P3_R1143_U142
g26902 and P3_R1143_U350 P3_R1143_U6 ; P3_R1143_U143
g26903 nand P3_R1143_U118 P3_R1143_U202 ; P3_R1143_U144
g26904 nand P3_R1143_U217 P3_R1143_U229 ; P3_R1143_U145
g26905 not P3_U3054 ; P3_R1143_U146
g26906 not P3_U3908 ; P3_R1143_U147
g26907 and P3_R1143_U403 P3_R1143_U402 ; P3_R1143_U148
g26908 nand P3_R1143_U304 P3_R1143_U169 P3_R1143_U364 ; P3_R1143_U149
g26909 and P3_R1143_U410 P3_R1143_U409 ; P3_R1143_U150
g26910 nand P3_R1143_U370 P3_R1143_U369 P3_R1143_U134 ; P3_R1143_U151
g26911 and P3_R1143_U417 P3_R1143_U416 ; P3_R1143_U152
g26912 nand P3_R1143_U365 P3_R1143_U299 P3_R1143_U86 ; P3_R1143_U153
g26913 and P3_R1143_U424 P3_R1143_U423 ; P3_R1143_U154
g26914 nand P3_R1143_U293 P3_R1143_U292 ; P3_R1143_U155
g26915 and P3_R1143_U436 P3_R1143_U435 ; P3_R1143_U156
g26916 nand P3_R1143_U289 P3_R1143_U288 ; P3_R1143_U157
g26917 and P3_R1143_U443 P3_R1143_U442 ; P3_R1143_U158
g26918 nand P3_R1143_U132 P3_R1143_U284 ; P3_R1143_U159
g26919 and P3_R1143_U450 P3_R1143_U449 ; P3_R1143_U160
g26920 nand P3_R1143_U43 P3_R1143_U327 ; P3_R1143_U161
g26921 nand P3_R1143_U130 P3_R1143_U269 ; P3_R1143_U162
g26922 and P3_R1143_U476 P3_R1143_U475 ; P3_R1143_U163
g26923 nand P3_R1143_U257 P3_R1143_U256 ; P3_R1143_U164
g26924 and P3_R1143_U483 P3_R1143_U482 ; P3_R1143_U165
g26925 nand P3_R1143_U253 P3_R1143_U252 ; P3_R1143_U166
g26926 nand P3_R1143_U127 P3_R1143_U242 ; P3_R1143_U167
g26927 nand P3_R1143_U367 P3_R1143_U366 ; P3_R1143_U168
g26928 nand P3_U3053 P3_R1143_U151 ; P3_R1143_U169
g26929 not P3_R1143_U34 ; P3_R1143_U170
g26930 nand P3_U3416 P3_U3082 ; P3_R1143_U171
g26931 nand P3_U3071 P3_U3425 ; P3_R1143_U172
g26932 nand P3_U3057 P3_U3902 ; P3_R1143_U173
g26933 not P3_R1143_U68 ; P3_R1143_U174
g26934 not P3_R1143_U77 ; P3_R1143_U175
g26935 nand P3_U3064 P3_U3903 ; P3_R1143_U176
g26936 not P3_R1143_U63 ; P3_R1143_U177
g26937 or P3_U3066 P3_U3404 ; P3_R1143_U178
g26938 or P3_U3059 P3_U3401 ; P3_R1143_U179
g26939 or P3_U3398 P3_U3063 ; P3_R1143_U180
g26940 or P3_U3395 P3_U3067 ; P3_R1143_U181
g26941 not P3_R1143_U31 ; P3_R1143_U182
g26942 or P3_U3392 P3_U3077 ; P3_R1143_U183
g26943 not P3_R1143_U42 ; P3_R1143_U184
g26944 not P3_R1143_U43 ; P3_R1143_U185
g26945 nand P3_R1143_U42 P3_R1143_U43 ; P3_R1143_U186
g26946 nand P3_U3067 P3_U3395 ; P3_R1143_U187
g26947 nand P3_R1143_U186 P3_R1143_U181 ; P3_R1143_U188
g26948 nand P3_U3063 P3_U3398 ; P3_R1143_U189
g26949 nand P3_R1143_U115 P3_R1143_U188 ; P3_R1143_U190
g26950 nand P3_R1143_U35 P3_R1143_U34 ; P3_R1143_U191
g26951 nand P3_U3066 P3_R1143_U191 ; P3_R1143_U192
g26952 nand P3_R1143_U116 P3_R1143_U190 ; P3_R1143_U193
g26953 nand P3_U3404 P3_R1143_U170 ; P3_R1143_U194
g26954 not P3_R1143_U41 ; P3_R1143_U195
g26955 or P3_U3069 P3_U3410 ; P3_R1143_U196
g26956 or P3_U3070 P3_U3407 ; P3_R1143_U197
g26957 not P3_R1143_U22 ; P3_R1143_U198
g26958 nand P3_R1143_U23 P3_R1143_U22 ; P3_R1143_U199
g26959 nand P3_U3069 P3_R1143_U199 ; P3_R1143_U200
g26960 nand P3_U3410 P3_R1143_U198 ; P3_R1143_U201
g26961 nand P3_R1143_U5 P3_R1143_U41 ; P3_R1143_U202
g26962 not P3_R1143_U144 ; P3_R1143_U203
g26963 or P3_U3413 P3_U3083 ; P3_R1143_U204
g26964 nand P3_R1143_U204 P3_R1143_U144 ; P3_R1143_U205
g26965 not P3_R1143_U40 ; P3_R1143_U206
g26966 or P3_U3082 P3_U3416 ; P3_R1143_U207
g26967 or P3_U3407 P3_U3070 ; P3_R1143_U208
g26968 nand P3_R1143_U208 P3_R1143_U41 ; P3_R1143_U209
g26969 nand P3_R1143_U119 P3_R1143_U209 ; P3_R1143_U210
g26970 nand P3_R1143_U195 P3_R1143_U22 ; P3_R1143_U211
g26971 nand P3_U3410 P3_U3069 ; P3_R1143_U212
g26972 nand P3_R1143_U120 P3_R1143_U211 ; P3_R1143_U213
g26973 or P3_U3070 P3_U3407 ; P3_R1143_U214
g26974 nand P3_R1143_U185 P3_R1143_U181 ; P3_R1143_U215
g26975 nand P3_U3067 P3_U3395 ; P3_R1143_U216
g26976 not P3_R1143_U45 ; P3_R1143_U217
g26977 nand P3_R1143_U121 P3_R1143_U184 ; P3_R1143_U218
g26978 nand P3_R1143_U45 P3_R1143_U180 ; P3_R1143_U219
g26979 nand P3_U3063 P3_U3398 ; P3_R1143_U220
g26980 not P3_R1143_U44 ; P3_R1143_U221
g26981 or P3_U3401 P3_U3059 ; P3_R1143_U222
g26982 nand P3_R1143_U222 P3_R1143_U44 ; P3_R1143_U223
g26983 nand P3_R1143_U123 P3_R1143_U223 ; P3_R1143_U224
g26984 nand P3_R1143_U221 P3_R1143_U34 ; P3_R1143_U225
g26985 nand P3_U3404 P3_U3066 ; P3_R1143_U226
g26986 nand P3_R1143_U124 P3_R1143_U225 ; P3_R1143_U227
g26987 or P3_U3059 P3_U3401 ; P3_R1143_U228
g26988 nand P3_R1143_U184 P3_R1143_U181 ; P3_R1143_U229
g26989 not P3_R1143_U145 ; P3_R1143_U230
g26990 nand P3_U3063 P3_U3398 ; P3_R1143_U231
g26991 nand P3_R1143_U401 P3_R1143_U400 P3_R1143_U43 P3_R1143_U42 ; P3_R1143_U232
g26992 nand P3_R1143_U43 P3_R1143_U42 ; P3_R1143_U233
g26993 nand P3_U3067 P3_U3395 ; P3_R1143_U234
g26994 nand P3_R1143_U125 P3_R1143_U233 ; P3_R1143_U235
g26995 or P3_U3082 P3_U3416 ; P3_R1143_U236
g26996 or P3_U3061 P3_U3419 ; P3_R1143_U237
g26997 nand P3_R1143_U177 P3_R1143_U6 ; P3_R1143_U238
g26998 nand P3_U3061 P3_U3419 ; P3_R1143_U239
g26999 nand P3_R1143_U171 P3_R1143_U238 ; P3_R1143_U240
g27000 or P3_U3419 P3_U3061 ; P3_R1143_U241
g27001 nand P3_R1143_U126 P3_R1143_U144 ; P3_R1143_U242
g27002 nand P3_R1143_U241 P3_R1143_U240 ; P3_R1143_U243
g27003 not P3_R1143_U167 ; P3_R1143_U244
g27004 or P3_U3079 P3_U3428 ; P3_R1143_U245
g27005 or P3_U3071 P3_U3425 ; P3_R1143_U246
g27006 nand P3_R1143_U174 P3_R1143_U7 ; P3_R1143_U247
g27007 nand P3_U3079 P3_U3428 ; P3_R1143_U248
g27008 nand P3_R1143_U129 P3_R1143_U247 ; P3_R1143_U249
g27009 or P3_U3422 P3_U3062 ; P3_R1143_U250
g27010 or P3_U3428 P3_U3079 ; P3_R1143_U251
g27011 nand P3_R1143_U128 P3_R1143_U167 ; P3_R1143_U252
g27012 nand P3_R1143_U251 P3_R1143_U249 ; P3_R1143_U253
g27013 not P3_R1143_U166 ; P3_R1143_U254
g27014 or P3_U3431 P3_U3078 ; P3_R1143_U255
g27015 nand P3_R1143_U255 P3_R1143_U166 ; P3_R1143_U256
g27016 nand P3_U3078 P3_U3431 ; P3_R1143_U257
g27017 not P3_R1143_U164 ; P3_R1143_U258
g27018 or P3_U3434 P3_U3073 ; P3_R1143_U259
g27019 nand P3_R1143_U259 P3_R1143_U164 ; P3_R1143_U260
g27020 nand P3_U3073 P3_U3434 ; P3_R1143_U261
g27021 not P3_R1143_U92 ; P3_R1143_U262
g27022 or P3_U3068 P3_U3440 ; P3_R1143_U263
g27023 or P3_U3072 P3_U3437 ; P3_R1143_U264
g27024 not P3_R1143_U59 ; P3_R1143_U265
g27025 nand P3_R1143_U60 P3_R1143_U59 ; P3_R1143_U266
g27026 nand P3_U3068 P3_R1143_U266 ; P3_R1143_U267
g27027 nand P3_U3440 P3_R1143_U265 ; P3_R1143_U268
g27028 nand P3_R1143_U8 P3_R1143_U92 ; P3_R1143_U269
g27029 not P3_R1143_U162 ; P3_R1143_U270
g27030 or P3_U3075 P3_U3907 ; P3_R1143_U271
g27031 or P3_U3080 P3_U3445 ; P3_R1143_U272
g27032 or P3_U3074 P3_U3906 ; P3_R1143_U273
g27033 not P3_R1143_U80 ; P3_R1143_U274
g27034 nand P3_U3907 P3_R1143_U274 ; P3_R1143_U275
g27035 nand P3_R1143_U275 P3_R1143_U90 ; P3_R1143_U276
g27036 nand P3_R1143_U80 P3_R1143_U81 ; P3_R1143_U277
g27037 nand P3_R1143_U277 P3_R1143_U276 ; P3_R1143_U278
g27038 nand P3_R1143_U175 P3_R1143_U9 ; P3_R1143_U279
g27039 nand P3_U3074 P3_U3906 ; P3_R1143_U280
g27040 nand P3_R1143_U278 P3_R1143_U279 ; P3_R1143_U281
g27041 or P3_U3443 P3_U3081 ; P3_R1143_U282
g27042 or P3_U3906 P3_U3074 ; P3_R1143_U283
g27043 nand P3_R1143_U162 P3_R1143_U131 ; P3_R1143_U284
g27044 nand P3_R1143_U283 P3_R1143_U281 ; P3_R1143_U285
g27045 not P3_R1143_U159 ; P3_R1143_U286
g27046 or P3_U3905 P3_U3060 ; P3_R1143_U287
g27047 nand P3_R1143_U287 P3_R1143_U159 ; P3_R1143_U288
g27048 nand P3_U3060 P3_U3905 ; P3_R1143_U289
g27049 not P3_R1143_U157 ; P3_R1143_U290
g27050 or P3_U3904 P3_U3065 ; P3_R1143_U291
g27051 nand P3_R1143_U291 P3_R1143_U157 ; P3_R1143_U292
g27052 nand P3_U3065 P3_U3904 ; P3_R1143_U293
g27053 not P3_R1143_U155 ; P3_R1143_U294
g27054 or P3_U3057 P3_U3902 ; P3_R1143_U295
g27055 nand P3_R1143_U176 P3_R1143_U173 ; P3_R1143_U296
g27056 not P3_R1143_U86 ; P3_R1143_U297
g27057 or P3_U3903 P3_U3064 ; P3_R1143_U298
g27058 nand P3_R1143_U155 P3_R1143_U298 P3_R1143_U168 ; P3_R1143_U299
g27059 not P3_R1143_U153 ; P3_R1143_U300
g27060 or P3_U3900 P3_U3052 ; P3_R1143_U301
g27061 nand P3_U3052 P3_U3900 ; P3_R1143_U302
g27062 not P3_R1143_U151 ; P3_R1143_U303
g27063 nand P3_U3899 P3_R1143_U151 ; P3_R1143_U304
g27064 not P3_R1143_U149 ; P3_R1143_U305
g27065 nand P3_R1143_U298 P3_R1143_U155 ; P3_R1143_U306
g27066 not P3_R1143_U89 ; P3_R1143_U307
g27067 or P3_U3902 P3_U3057 ; P3_R1143_U308
g27068 nand P3_R1143_U308 P3_R1143_U89 ; P3_R1143_U309
g27069 nand P3_R1143_U309 P3_R1143_U173 P3_R1143_U154 ; P3_R1143_U310
g27070 nand P3_R1143_U307 P3_R1143_U173 ; P3_R1143_U311
g27071 nand P3_U3901 P3_U3056 ; P3_R1143_U312
g27072 nand P3_R1143_U311 P3_R1143_U312 P3_R1143_U168 ; P3_R1143_U313
g27073 or P3_U3057 P3_U3902 ; P3_R1143_U314
g27074 nand P3_R1143_U282 P3_R1143_U162 ; P3_R1143_U315
g27075 not P3_R1143_U91 ; P3_R1143_U316
g27076 nand P3_R1143_U9 P3_R1143_U91 ; P3_R1143_U317
g27077 nand P3_R1143_U135 P3_R1143_U317 ; P3_R1143_U318
g27078 nand P3_R1143_U317 P3_R1143_U278 ; P3_R1143_U319
g27079 nand P3_R1143_U453 P3_R1143_U319 ; P3_R1143_U320
g27080 or P3_U3445 P3_U3080 ; P3_R1143_U321
g27081 nand P3_R1143_U321 P3_R1143_U91 ; P3_R1143_U322
g27082 nand P3_R1143_U136 P3_R1143_U322 ; P3_R1143_U323
g27083 nand P3_R1143_U316 P3_R1143_U80 ; P3_R1143_U324
g27084 nand P3_U3075 P3_U3907 ; P3_R1143_U325
g27085 nand P3_R1143_U137 P3_R1143_U324 ; P3_R1143_U326
g27086 or P3_U3392 P3_U3077 ; P3_R1143_U327
g27087 not P3_R1143_U161 ; P3_R1143_U328
g27088 or P3_U3080 P3_U3445 ; P3_R1143_U329
g27089 or P3_U3437 P3_U3072 ; P3_R1143_U330
g27090 nand P3_R1143_U330 P3_R1143_U92 ; P3_R1143_U331
g27091 nand P3_R1143_U138 P3_R1143_U331 ; P3_R1143_U332
g27092 nand P3_R1143_U262 P3_R1143_U59 ; P3_R1143_U333
g27093 nand P3_U3440 P3_U3068 ; P3_R1143_U334
g27094 nand P3_R1143_U139 P3_R1143_U333 ; P3_R1143_U335
g27095 or P3_U3072 P3_U3437 ; P3_R1143_U336
g27096 nand P3_R1143_U250 P3_R1143_U167 ; P3_R1143_U337
g27097 not P3_R1143_U93 ; P3_R1143_U338
g27098 or P3_U3425 P3_U3071 ; P3_R1143_U339
g27099 nand P3_R1143_U339 P3_R1143_U93 ; P3_R1143_U340
g27100 nand P3_R1143_U140 P3_R1143_U340 ; P3_R1143_U341
g27101 nand P3_R1143_U338 P3_R1143_U172 ; P3_R1143_U342
g27102 nand P3_U3079 P3_U3428 ; P3_R1143_U343
g27103 nand P3_R1143_U141 P3_R1143_U342 ; P3_R1143_U344
g27104 or P3_U3071 P3_U3425 ; P3_R1143_U345
g27105 or P3_U3416 P3_U3082 ; P3_R1143_U346
g27106 nand P3_R1143_U346 P3_R1143_U40 ; P3_R1143_U347
g27107 nand P3_R1143_U142 P3_R1143_U347 ; P3_R1143_U348
g27108 nand P3_R1143_U206 P3_R1143_U171 ; P3_R1143_U349
g27109 nand P3_U3061 P3_U3419 ; P3_R1143_U350
g27110 nand P3_R1143_U143 P3_R1143_U349 ; P3_R1143_U351
g27111 nand P3_R1143_U207 P3_R1143_U171 ; P3_R1143_U352
g27112 nand P3_R1143_U204 P3_R1143_U63 ; P3_R1143_U353
g27113 nand P3_R1143_U214 P3_R1143_U22 ; P3_R1143_U354
g27114 nand P3_R1143_U228 P3_R1143_U34 ; P3_R1143_U355
g27115 nand P3_R1143_U231 P3_R1143_U180 ; P3_R1143_U356
g27116 nand P3_R1143_U314 P3_R1143_U173 ; P3_R1143_U357
g27117 nand P3_R1143_U298 P3_R1143_U176 ; P3_R1143_U358
g27118 nand P3_R1143_U329 P3_R1143_U80 ; P3_R1143_U359
g27119 nand P3_R1143_U282 P3_R1143_U77 ; P3_R1143_U360
g27120 nand P3_R1143_U336 P3_R1143_U59 ; P3_R1143_U361
g27121 nand P3_R1143_U345 P3_R1143_U172 ; P3_R1143_U362
g27122 nand P3_R1143_U250 P3_R1143_U68 ; P3_R1143_U363
g27123 nand P3_U3899 P3_U3053 ; P3_R1143_U364
g27124 nand P3_R1143_U296 P3_R1143_U168 ; P3_R1143_U365
g27125 nand P3_U3056 P3_R1143_U295 ; P3_R1143_U366
g27126 nand P3_U3901 P3_R1143_U295 ; P3_R1143_U367
g27127 nand P3_R1143_U296 P3_R1143_U168 P3_R1143_U301 ; P3_R1143_U368
g27128 nand P3_R1143_U155 P3_R1143_U168 P3_R1143_U133 ; P3_R1143_U369
g27129 nand P3_R1143_U297 P3_R1143_U301 ; P3_R1143_U370
g27130 nand P3_U3082 P3_R1143_U39 ; P3_R1143_U371
g27131 nand P3_U3416 P3_R1143_U38 ; P3_R1143_U372
g27132 nand P3_R1143_U372 P3_R1143_U371 ; P3_R1143_U373
g27133 nand P3_R1143_U352 P3_R1143_U40 ; P3_R1143_U374
g27134 nand P3_R1143_U373 P3_R1143_U206 ; P3_R1143_U375
g27135 nand P3_U3083 P3_R1143_U36 ; P3_R1143_U376
g27136 nand P3_U3413 P3_R1143_U37 ; P3_R1143_U377
g27137 nand P3_R1143_U377 P3_R1143_U376 ; P3_R1143_U378
g27138 nand P3_R1143_U353 P3_R1143_U144 ; P3_R1143_U379
g27139 nand P3_R1143_U203 P3_R1143_U378 ; P3_R1143_U380
g27140 nand P3_U3069 P3_R1143_U23 ; P3_R1143_U381
g27141 nand P3_U3410 P3_R1143_U21 ; P3_R1143_U382
g27142 nand P3_U3070 P3_R1143_U19 ; P3_R1143_U383
g27143 nand P3_U3407 P3_R1143_U20 ; P3_R1143_U384
g27144 nand P3_R1143_U384 P3_R1143_U383 ; P3_R1143_U385
g27145 nand P3_R1143_U354 P3_R1143_U41 ; P3_R1143_U386
g27146 nand P3_R1143_U385 P3_R1143_U195 ; P3_R1143_U387
g27147 nand P3_U3066 P3_R1143_U35 ; P3_R1143_U388
g27148 nand P3_U3404 P3_R1143_U26 ; P3_R1143_U389
g27149 nand P3_U3059 P3_R1143_U24 ; P3_R1143_U390
g27150 nand P3_U3401 P3_R1143_U25 ; P3_R1143_U391
g27151 nand P3_R1143_U391 P3_R1143_U390 ; P3_R1143_U392
g27152 nand P3_R1143_U355 P3_R1143_U44 ; P3_R1143_U393
g27153 nand P3_R1143_U392 P3_R1143_U221 ; P3_R1143_U394
g27154 nand P3_U3063 P3_R1143_U32 ; P3_R1143_U395
g27155 nand P3_U3398 P3_R1143_U33 ; P3_R1143_U396
g27156 nand P3_R1143_U396 P3_R1143_U395 ; P3_R1143_U397
g27157 nand P3_R1143_U356 P3_R1143_U145 ; P3_R1143_U398
g27158 nand P3_R1143_U230 P3_R1143_U397 ; P3_R1143_U399
g27159 nand P3_U3067 P3_R1143_U27 ; P3_R1143_U400
g27160 nand P3_U3395 P3_R1143_U28 ; P3_R1143_U401
g27161 nand P3_U3054 P3_R1143_U147 ; P3_R1143_U402
g27162 nand P3_U3908 P3_R1143_U146 ; P3_R1143_U403
g27163 nand P3_U3054 P3_R1143_U147 ; P3_R1143_U404
g27164 nand P3_U3908 P3_R1143_U146 ; P3_R1143_U405
g27165 nand P3_R1143_U405 P3_R1143_U404 ; P3_R1143_U406
g27166 nand P3_R1143_U148 P3_R1143_U149 ; P3_R1143_U407
g27167 nand P3_R1143_U305 P3_R1143_U406 ; P3_R1143_U408
g27168 nand P3_U3053 P3_R1143_U88 ; P3_R1143_U409
g27169 nand P3_U3899 P3_R1143_U87 ; P3_R1143_U410
g27170 nand P3_U3053 P3_R1143_U88 ; P3_R1143_U411
g27171 nand P3_U3899 P3_R1143_U87 ; P3_R1143_U412
g27172 nand P3_R1143_U412 P3_R1143_U411 ; P3_R1143_U413
g27173 nand P3_R1143_U150 P3_R1143_U151 ; P3_R1143_U414
g27174 nand P3_R1143_U303 P3_R1143_U413 ; P3_R1143_U415
g27175 nand P3_U3052 P3_R1143_U46 ; P3_R1143_U416
g27176 nand P3_U3900 P3_R1143_U47 ; P3_R1143_U417
g27177 nand P3_U3052 P3_R1143_U46 ; P3_R1143_U418
g27178 nand P3_U3900 P3_R1143_U47 ; P3_R1143_U419
g27179 nand P3_R1143_U419 P3_R1143_U418 ; P3_R1143_U420
g27180 nand P3_R1143_U152 P3_R1143_U153 ; P3_R1143_U421
g27181 nand P3_R1143_U300 P3_R1143_U420 ; P3_R1143_U422
g27182 nand P3_U3056 P3_R1143_U49 ; P3_R1143_U423
g27183 nand P3_U3901 P3_R1143_U48 ; P3_R1143_U424
g27184 nand P3_U3057 P3_R1143_U50 ; P3_R1143_U425
g27185 nand P3_U3902 P3_R1143_U51 ; P3_R1143_U426
g27186 nand P3_R1143_U426 P3_R1143_U425 ; P3_R1143_U427
g27187 nand P3_R1143_U357 P3_R1143_U89 ; P3_R1143_U428
g27188 nand P3_R1143_U427 P3_R1143_U307 ; P3_R1143_U429
g27189 nand P3_U3064 P3_R1143_U52 ; P3_R1143_U430
g27190 nand P3_U3903 P3_R1143_U53 ; P3_R1143_U431
g27191 nand P3_R1143_U431 P3_R1143_U430 ; P3_R1143_U432
g27192 nand P3_R1143_U358 P3_R1143_U155 ; P3_R1143_U433
g27193 nand P3_R1143_U294 P3_R1143_U432 ; P3_R1143_U434
g27194 nand P3_U3065 P3_R1143_U84 ; P3_R1143_U435
g27195 nand P3_U3904 P3_R1143_U85 ; P3_R1143_U436
g27196 nand P3_U3065 P3_R1143_U84 ; P3_R1143_U437
g27197 nand P3_U3904 P3_R1143_U85 ; P3_R1143_U438
g27198 nand P3_R1143_U438 P3_R1143_U437 ; P3_R1143_U439
g27199 nand P3_R1143_U156 P3_R1143_U157 ; P3_R1143_U440
g27200 nand P3_R1143_U290 P3_R1143_U439 ; P3_R1143_U441
g27201 nand P3_U3060 P3_R1143_U82 ; P3_R1143_U442
g27202 nand P3_U3905 P3_R1143_U83 ; P3_R1143_U443
g27203 nand P3_U3060 P3_R1143_U82 ; P3_R1143_U444
g27204 nand P3_U3905 P3_R1143_U83 ; P3_R1143_U445
g27205 nand P3_R1143_U445 P3_R1143_U444 ; P3_R1143_U446
g27206 nand P3_R1143_U158 P3_R1143_U159 ; P3_R1143_U447
g27207 nand P3_R1143_U286 P3_R1143_U446 ; P3_R1143_U448
g27208 nand P3_U3074 P3_R1143_U54 ; P3_R1143_U449
g27209 nand P3_U3906 P3_R1143_U55 ; P3_R1143_U450
g27210 nand P3_U3074 P3_R1143_U54 ; P3_R1143_U451
g27211 nand P3_U3906 P3_R1143_U55 ; P3_R1143_U452
g27212 nand P3_R1143_U452 P3_R1143_U451 ; P3_R1143_U453
g27213 nand P3_U3075 P3_R1143_U81 ; P3_R1143_U454
g27214 nand P3_U3907 P3_R1143_U90 ; P3_R1143_U455
g27215 nand P3_R1143_U182 P3_R1143_U161 ; P3_R1143_U456
g27216 nand P3_R1143_U328 P3_R1143_U31 ; P3_R1143_U457
g27217 nand P3_U3080 P3_R1143_U78 ; P3_R1143_U458
g27218 nand P3_U3445 P3_R1143_U79 ; P3_R1143_U459
g27219 nand P3_R1143_U459 P3_R1143_U458 ; P3_R1143_U460
g27220 nand P3_R1143_U359 P3_R1143_U91 ; P3_R1143_U461
g27221 nand P3_R1143_U460 P3_R1143_U316 ; P3_R1143_U462
g27222 nand P3_U3081 P3_R1143_U75 ; P3_R1143_U463
g27223 nand P3_U3443 P3_R1143_U76 ; P3_R1143_U464
g27224 nand P3_R1143_U464 P3_R1143_U463 ; P3_R1143_U465
g27225 nand P3_R1143_U360 P3_R1143_U162 ; P3_R1143_U466
g27226 nand P3_R1143_U270 P3_R1143_U465 ; P3_R1143_U467
g27227 nand P3_U3068 P3_R1143_U60 ; P3_R1143_U468
g27228 nand P3_U3440 P3_R1143_U58 ; P3_R1143_U469
g27229 nand P3_U3072 P3_R1143_U56 ; P3_R1143_U470
g27230 nand P3_U3437 P3_R1143_U57 ; P3_R1143_U471
g27231 nand P3_R1143_U471 P3_R1143_U470 ; P3_R1143_U472
g27232 nand P3_R1143_U361 P3_R1143_U92 ; P3_R1143_U473
g27233 nand P3_R1143_U472 P3_R1143_U262 ; P3_R1143_U474
g27234 nand P3_U3073 P3_R1143_U73 ; P3_R1143_U475
g27235 nand P3_U3434 P3_R1143_U74 ; P3_R1143_U476
g27236 nand P3_U3073 P3_R1143_U73 ; P3_R1143_U477
g27237 nand P3_U3434 P3_R1143_U74 ; P3_R1143_U478
g27238 nand P3_R1143_U478 P3_R1143_U477 ; P3_R1143_U479
g27239 nand P3_R1143_U163 P3_R1143_U164 ; P3_R1143_U480
g27240 nand P3_R1143_U258 P3_R1143_U479 ; P3_R1143_U481
g27241 nand P3_U3078 P3_R1143_U71 ; P3_R1143_U482
g27242 nand P3_U3431 P3_R1143_U72 ; P3_R1143_U483
g27243 nand P3_U3078 P3_R1143_U71 ; P3_R1143_U484
g27244 nand P3_U3431 P3_R1143_U72 ; P3_R1143_U485
g27245 nand P3_R1143_U485 P3_R1143_U484 ; P3_R1143_U486
g27246 nand P3_R1143_U165 P3_R1143_U166 ; P3_R1143_U487
g27247 nand P3_R1143_U254 P3_R1143_U486 ; P3_R1143_U488
g27248 nand P3_U3079 P3_R1143_U69 ; P3_R1143_U489
g27249 nand P3_U3428 P3_R1143_U70 ; P3_R1143_U490
g27250 nand P3_U3071 P3_R1143_U64 ; P3_R1143_U491
g27251 nand P3_U3425 P3_R1143_U65 ; P3_R1143_U492
g27252 nand P3_R1143_U492 P3_R1143_U491 ; P3_R1143_U493
g27253 nand P3_R1143_U362 P3_R1143_U93 ; P3_R1143_U494
g27254 nand P3_R1143_U493 P3_R1143_U338 ; P3_R1143_U495
g27255 nand P3_U3062 P3_R1143_U66 ; P3_R1143_U496
g27256 nand P3_U3422 P3_R1143_U67 ; P3_R1143_U497
g27257 nand P3_R1143_U497 P3_R1143_U496 ; P3_R1143_U498
g27258 nand P3_R1143_U363 P3_R1143_U167 ; P3_R1143_U499
g27259 nand P3_R1143_U244 P3_R1143_U498 ; P3_R1143_U500
g27260 nand P3_U3061 P3_R1143_U61 ; P3_R1143_U501
g27261 nand P3_U3419 P3_R1143_U62 ; P3_R1143_U502
g27262 nand P3_U3076 P3_R1143_U29 ; P3_R1143_U503
g27263 nand P3_U3387 P3_R1143_U30 ; P3_R1143_U504
g27264 and P3_R1158_U227 P3_R1158_U226 ; P3_R1158_U4
g27265 and P3_R1158_U238 P3_R1158_U237 ; P3_R1158_U5
g27266 and P3_R1158_U263 P3_R1158_U262 ; P3_R1158_U6
g27267 and P3_R1158_U277 P3_R1158_U276 ; P3_R1158_U7
g27268 and P3_R1158_U289 P3_R1158_U288 ; P3_R1158_U8
g27269 and P3_R1158_U6 P3_R1158_U267 ; P3_R1158_U9
g27270 and P3_R1158_U5 P3_R1158_U235 ; P3_R1158_U10
g27271 and P3_R1158_U9 P3_R1158_U260 ; P3_R1158_U11
g27272 and P3_R1158_U535 P3_R1158_U534 ; P3_R1158_U12
g27273 and P3_R1158_U345 P3_R1158_U342 ; P3_R1158_U13
g27274 and P3_R1158_U336 P3_R1158_U333 ; P3_R1158_U14
g27275 and P3_R1158_U329 P3_R1158_U326 ; P3_R1158_U15
g27276 and P3_R1158_U537 P3_R1158_U536 P3_R1158_U142 ; P3_R1158_U16
g27277 and P3_R1158_U256 P3_R1158_U253 ; P3_R1158_U17
g27278 and P3_R1158_U249 P3_R1158_U246 ; P3_R1158_U18
g27279 nand P3_U3056 P3_R1158_U306 ; P3_R1158_U19
g27280 not P3_U3152 ; P3_R1158_U20
g27281 not P3_U3083 ; P3_R1158_U21
g27282 not P3_U3070 ; P3_R1158_U22
g27283 nand P3_U3070 P3_R1158_U67 ; P3_R1158_U23
g27284 not P3_U3069 ; P3_R1158_U24
g27285 not P3_U3066 ; P3_R1158_U25
g27286 nand P3_U3066 P3_R1158_U69 ; P3_R1158_U26
g27287 not P3_U3067 ; P3_R1158_U27
g27288 nand P3_U3067 P3_R1158_U70 ; P3_R1158_U28
g27289 not P3_U3063 ; P3_R1158_U29
g27290 not P3_U3077 ; P3_R1158_U30
g27291 not P3_U3076 ; P3_R1158_U31
g27292 not P3_U3059 ; P3_R1158_U32
g27293 not P3_U3082 ; P3_R1158_U33
g27294 nand P3_R1158_U359 P3_R1158_U241 P3_R1158_U362 ; P3_R1158_U34
g27295 nand P3_R1158_U379 P3_R1158_U26 ; P3_R1158_U35
g27296 nand P3_R1158_U361 P3_R1158_U224 P3_R1158_U360 ; P3_R1158_U36
g27297 not P3_U3052 ; P3_R1158_U37
g27298 not P3_U3057 ; P3_R1158_U38
g27299 not P3_U3064 ; P3_R1158_U39
g27300 not P3_U3056 ; P3_R1158_U40
g27301 not P3_U3072 ; P3_R1158_U41
g27302 nand P3_U3072 P3_R1158_U79 ; P3_R1158_U42
g27303 not P3_U3068 ; P3_R1158_U43
g27304 not P3_U3078 ; P3_R1158_U44
g27305 not P3_U3071 ; P3_R1158_U45
g27306 not P3_U3062 ; P3_R1158_U46
g27307 nand P3_U3062 P3_R1158_U84 ; P3_R1158_U47
g27308 not P3_U3079 ; P3_R1158_U48
g27309 not P3_U3061 ; P3_R1158_U49
g27310 nand P3_U3061 P3_R1158_U85 ; P3_R1158_U50
g27311 not P3_U3073 ; P3_R1158_U51
g27312 not P3_U3081 ; P3_R1158_U52
g27313 not P3_U3075 ; P3_R1158_U53
g27314 not P3_U3080 ; P3_R1158_U54
g27315 nand P3_U3080 P3_R1158_U88 ; P3_R1158_U55
g27316 not P3_U3074 ; P3_R1158_U56
g27317 not P3_U3060 ; P3_R1158_U57
g27318 not P3_U3065 ; P3_R1158_U58
g27319 nand P3_U3057 P3_R1158_U76 ; P3_R1158_U59
g27320 nand P3_U3064 P3_R1158_U77 ; P3_R1158_U60
g27321 nand P3_R1158_U55 P3_R1158_U322 ; P3_R1158_U61
g27322 nand P3_R1158_U274 P3_R1158_U273 ; P3_R1158_U62
g27323 nand P3_R1158_U365 P3_R1158_U269 ; P3_R1158_U63
g27324 nand P3_R1158_U47 P3_R1158_U338 ; P3_R1158_U64
g27325 nand P3_R1158_U394 P3_R1158_U393 ; P3_R1158_U65
g27326 nand P3_R1158_U426 P3_R1158_U425 ; P3_R1158_U66
g27327 nand P3_R1158_U423 P3_R1158_U422 ; P3_R1158_U67
g27328 nand P3_R1158_U420 P3_R1158_U419 ; P3_R1158_U68
g27329 nand P3_R1158_U417 P3_R1158_U416 ; P3_R1158_U69
g27330 nand P3_R1158_U414 P3_R1158_U413 ; P3_R1158_U70
g27331 nand P3_R1158_U411 P3_R1158_U410 ; P3_R1158_U71
g27332 nand P3_R1158_U405 P3_R1158_U404 ; P3_R1158_U72
g27333 nand P3_R1158_U408 P3_R1158_U407 ; P3_R1158_U73
g27334 nand P3_R1158_U402 P3_R1158_U401 ; P3_R1158_U74
g27335 nand P3_R1158_U466 P3_R1158_U465 ; P3_R1158_U75
g27336 nand P3_R1158_U514 P3_R1158_U513 ; P3_R1158_U76
g27337 nand P3_R1158_U517 P3_R1158_U516 ; P3_R1158_U77
g27338 nand P3_R1158_U511 P3_R1158_U510 ; P3_R1158_U78
g27339 nand P3_R1158_U490 P3_R1158_U489 ; P3_R1158_U79
g27340 nand P3_R1158_U487 P3_R1158_U486 ; P3_R1158_U80
g27341 nand P3_R1158_U481 P3_R1158_U480 ; P3_R1158_U81
g27342 nand P3_R1158_U478 P3_R1158_U477 ; P3_R1158_U82
g27343 nand P3_R1158_U475 P3_R1158_U474 ; P3_R1158_U83
g27344 nand P3_R1158_U472 P3_R1158_U471 ; P3_R1158_U84
g27345 nand P3_R1158_U469 P3_R1158_U468 ; P3_R1158_U85
g27346 nand P3_R1158_U484 P3_R1158_U483 ; P3_R1158_U86
g27347 nand P3_R1158_U493 P3_R1158_U492 ; P3_R1158_U87
g27348 nand P3_R1158_U502 P3_R1158_U501 ; P3_R1158_U88
g27349 nand P3_R1158_U496 P3_R1158_U495 ; P3_R1158_U89
g27350 nand P3_R1158_U499 P3_R1158_U498 ; P3_R1158_U90
g27351 nand P3_R1158_U505 P3_R1158_U504 ; P3_R1158_U91
g27352 nand P3_R1158_U508 P3_R1158_U507 ; P3_R1158_U92
g27353 nand P3_R1158_U523 P3_R1158_U522 ; P3_R1158_U93
g27354 nand P3_R1158_U632 P3_R1158_U631 ; P3_R1158_U94
g27355 nand P3_R1158_U429 P3_R1158_U428 ; P3_R1158_U95
g27356 nand P3_R1158_U436 P3_R1158_U435 ; P3_R1158_U96
g27357 nand P3_R1158_U443 P3_R1158_U442 ; P3_R1158_U97
g27358 nand P3_R1158_U450 P3_R1158_U449 ; P3_R1158_U98
g27359 nand P3_R1158_U457 P3_R1158_U456 ; P3_R1158_U99
g27360 nand P3_R1158_U464 P3_R1158_U463 ; P3_R1158_U100
g27361 nand P3_R1158_U526 P3_R1158_U525 ; P3_R1158_U101
g27362 nand P3_R1158_U533 P3_R1158_U532 ; P3_R1158_U102
g27363 and P3_R1158_U320 P3_R1158_U209 ; P3_R1158_U103
g27364 and P3_R1158_U141 P3_R1158_U12 ; P3_R1158_U104
g27365 nand P3_R1158_U542 P3_R1158_U541 ; P3_R1158_U105
g27366 nand P3_R1158_U547 P3_R1158_U546 ; P3_R1158_U106
g27367 nand P3_R1158_U554 P3_R1158_U553 ; P3_R1158_U107
g27368 nand P3_R1158_U561 P3_R1158_U560 ; P3_R1158_U108
g27369 nand P3_R1158_U568 P3_R1158_U567 ; P3_R1158_U109
g27370 nand P3_R1158_U575 P3_R1158_U574 ; P3_R1158_U110
g27371 nand P3_R1158_U580 P3_R1158_U579 ; P3_R1158_U111
g27372 nand P3_R1158_U587 P3_R1158_U586 ; P3_R1158_U112
g27373 nand P3_R1158_U594 P3_R1158_U593 ; P3_R1158_U113
g27374 nand P3_R1158_U601 P3_R1158_U600 ; P3_R1158_U114
g27375 nand P3_R1158_U608 P3_R1158_U607 ; P3_R1158_U115
g27376 nand P3_R1158_U615 P3_R1158_U614 ; P3_R1158_U116
g27377 nand P3_R1158_U620 P3_R1158_U619 ; P3_R1158_U117
g27378 nand P3_R1158_U627 P3_R1158_U626 ; P3_R1158_U118
g27379 and P3_R1158_U73 P3_U3152 ; P3_R1158_U119
g27380 and P3_R1158_U230 P3_R1158_U229 ; P3_R1158_U120
g27381 and P3_R1158_U242 P3_R1158_U10 ; P3_R1158_U121
g27382 and P3_R1158_U364 P3_R1158_U243 ; P3_R1158_U122
g27383 and P3_R1158_U438 P3_R1158_U437 P3_R1158_U23 ; P3_R1158_U123
g27384 and P3_R1158_U248 P3_R1158_U5 ; P3_R1158_U124
g27385 and P3_R1158_U459 P3_R1158_U458 P3_R1158_U28 ; P3_R1158_U125
g27386 and P3_R1158_U255 P3_R1158_U4 ; P3_R1158_U126
g27387 and P3_R1158_U265 P3_R1158_U213 ; P3_R1158_U127
g27388 and P3_R1158_U270 P3_R1158_U11 ; P3_R1158_U128
g27389 and P3_R1158_U373 P3_R1158_U271 ; P3_R1158_U129
g27390 and P3_R1158_U281 P3_R1158_U280 ; P3_R1158_U130
g27391 and P3_R1158_U293 P3_R1158_U8 ; P3_R1158_U131
g27392 and P3_R1158_U291 P3_R1158_U214 ; P3_R1158_U132
g27393 and P3_R1158_U314 P3_R1158_U376 ; P3_R1158_U133
g27394 and P3_R1158_U316 P3_R1158_U307 ; P3_R1158_U134
g27395 and P3_R1158_U316 P3_R1158_U369 ; P3_R1158_U135
g27396 and P3_R1158_U374 P3_R1158_U315 ; P3_R1158_U136
g27397 nand P3_R1158_U520 P3_R1158_U519 ; P3_R1158_U137
g27398 and P3_R1158_U515 P3_R1158_U38 ; P3_R1158_U138
g27399 and P3_R1158_U320 P3_R1158_U215 ; P3_R1158_U139
g27400 and P3_R1158_U320 P3_R1158_U218 ; P3_R1158_U140
g27401 and P3_R1158_U60 P3_R1158_U59 ; P3_R1158_U141
g27402 and P3_R1158_U391 P3_R1158_U319 P3_R1158_U392 ; P3_R1158_U142
g27403 and P3_R1158_U563 P3_R1158_U562 P3_R1158_U214 ; P3_R1158_U143
g27404 and P3_R1158_U328 P3_R1158_U8 ; P3_R1158_U144
g27405 and P3_R1158_U589 P3_R1158_U588 P3_R1158_U42 ; P3_R1158_U145
g27406 and P3_R1158_U335 P3_R1158_U7 ; P3_R1158_U146
g27407 and P3_R1158_U610 P3_R1158_U609 P3_R1158_U213 ; P3_R1158_U147
g27408 and P3_R1158_U344 P3_R1158_U6 ; P3_R1158_U148
g27409 nand P3_R1158_U629 P3_R1158_U628 ; P3_R1158_U149
g27410 not P3_U3416 ; P3_R1158_U150
g27411 and P3_R1158_U397 P3_R1158_U396 ; P3_R1158_U151
g27412 not P3_U3401 ; P3_R1158_U152
g27413 not P3_U3392 ; P3_R1158_U153
g27414 not P3_U3387 ; P3_R1158_U154
g27415 not P3_U3398 ; P3_R1158_U155
g27416 not P3_U3395 ; P3_R1158_U156
g27417 not P3_U3404 ; P3_R1158_U157
g27418 not P3_U3410 ; P3_R1158_U158
g27419 not P3_U3407 ; P3_R1158_U159
g27420 not P3_U3413 ; P3_R1158_U160
g27421 nand P3_R1158_U122 P3_R1158_U383 ; P3_R1158_U161
g27422 and P3_R1158_U431 P3_R1158_U430 ; P3_R1158_U162
g27423 nand P3_R1158_U363 P3_R1158_U381 ; P3_R1158_U163
g27424 and P3_R1158_U445 P3_R1158_U444 ; P3_R1158_U164
g27425 nand P3_R1158_U233 P3_R1158_U211 P3_R1158_U356 ; P3_R1158_U165
g27426 and P3_R1158_U452 P3_R1158_U451 ; P3_R1158_U166
g27427 nand P3_R1158_U120 P3_R1158_U231 ; P3_R1158_U167
g27428 not P3_U3900 ; P3_R1158_U168
g27429 not P3_U3419 ; P3_R1158_U169
g27430 not P3_U3422 ; P3_R1158_U170
g27431 not P3_U3428 ; P3_R1158_U171
g27432 not P3_U3425 ; P3_R1158_U172
g27433 not P3_U3431 ; P3_R1158_U173
g27434 not P3_U3434 ; P3_R1158_U174
g27435 not P3_U3440 ; P3_R1158_U175
g27436 not P3_U3437 ; P3_R1158_U176
g27437 not P3_U3443 ; P3_R1158_U177
g27438 not P3_U3906 ; P3_R1158_U178
g27439 not P3_U3907 ; P3_R1158_U179
g27440 not P3_U3445 ; P3_R1158_U180
g27441 not P3_U3905 ; P3_R1158_U181
g27442 not P3_U3904 ; P3_R1158_U182
g27443 not P3_U3901 ; P3_R1158_U183
g27444 not P3_U3902 ; P3_R1158_U184
g27445 not P3_U3903 ; P3_R1158_U185
g27446 not P3_U3053 ; P3_R1158_U186
g27447 not P3_U3899 ; P3_R1158_U187
g27448 and P3_R1158_U528 P3_R1158_U527 ; P3_R1158_U188
g27449 nand P3_R1158_U311 P3_R1158_U310 ; P3_R1158_U189
g27450 nand P3_R1158_U309 P3_R1158_U192 ; P3_R1158_U190
g27451 nand P3_R1158_U60 P3_R1158_U190 ; P3_R1158_U191
g27452 nand P3_R1158_U304 P3_R1158_U303 ; P3_R1158_U192
g27453 and P3_R1158_U549 P3_R1158_U548 ; P3_R1158_U193
g27454 nand P3_R1158_U300 P3_R1158_U299 ; P3_R1158_U194
g27455 and P3_R1158_U556 P3_R1158_U555 ; P3_R1158_U195
g27456 nand P3_R1158_U296 P3_R1158_U295 ; P3_R1158_U196
g27457 and P3_R1158_U570 P3_R1158_U569 ; P3_R1158_U197
g27458 nand P3_R1158_U221 P3_R1158_U220 ; P3_R1158_U198
g27459 nand P3_R1158_U286 P3_R1158_U285 ; P3_R1158_U199
g27460 and P3_R1158_U582 P3_R1158_U581 ; P3_R1158_U200
g27461 nand P3_R1158_U130 P3_R1158_U282 ; P3_R1158_U201
g27462 and P3_R1158_U596 P3_R1158_U595 ; P3_R1158_U202
g27463 nand P3_R1158_U129 P3_R1158_U389 ; P3_R1158_U203
g27464 and P3_R1158_U603 P3_R1158_U602 ; P3_R1158_U204
g27465 nand P3_R1158_U372 P3_R1158_U387 ; P3_R1158_U205
g27466 nand P3_R1158_U385 P3_R1158_U50 ; P3_R1158_U206
g27467 and P3_R1158_U622 P3_R1158_U621 ; P3_R1158_U207
g27468 nand P3_R1158_U258 P3_R1158_U210 P3_R1158_U357 ; P3_R1158_U208
g27469 nand P3_R1158_U19 P3_R1158_U367 ; P3_R1158_U209
g27470 nand P3_R1158_U65 P3_R1158_U161 ; P3_R1158_U210
g27471 nand P3_R1158_U74 P3_R1158_U167 ; P3_R1158_U211
g27472 not P3_R1158_U28 ; P3_R1158_U212
g27473 nand P3_U3071 P3_R1158_U82 ; P3_R1158_U213
g27474 nand P3_U3075 P3_R1158_U90 ; P3_R1158_U214
g27475 not P3_R1158_U59 ; P3_R1158_U215
g27476 not P3_R1158_U47 ; P3_R1158_U216
g27477 not P3_R1158_U55 ; P3_R1158_U217
g27478 not P3_R1158_U60 ; P3_R1158_U218
g27479 nand P3_R1158_U409 P3_R1158_U20 ; P3_R1158_U219
g27480 nand P3_U3076 P3_R1158_U219 ; P3_R1158_U220
g27481 nand P3_U3152 P3_R1158_U73 ; P3_R1158_U221
g27482 not P3_R1158_U198 ; P3_R1158_U222
g27483 nand P3_R1158_U406 P3_R1158_U30 ; P3_R1158_U223
g27484 nand P3_U3077 P3_R1158_U72 ; P3_R1158_U224
g27485 not P3_R1158_U36 ; P3_R1158_U225
g27486 nand P3_R1158_U412 P3_R1158_U29 ; P3_R1158_U226
g27487 nand P3_R1158_U415 P3_R1158_U27 ; P3_R1158_U227
g27488 nand P3_R1158_U29 P3_R1158_U28 ; P3_R1158_U228
g27489 nand P3_R1158_U71 P3_R1158_U228 ; P3_R1158_U229
g27490 nand P3_U3063 P3_R1158_U212 ; P3_R1158_U230
g27491 nand P3_R1158_U4 P3_R1158_U36 ; P3_R1158_U231
g27492 not P3_R1158_U167 ; P3_R1158_U232
g27493 nand P3_U3059 P3_R1158_U167 ; P3_R1158_U233
g27494 not P3_R1158_U165 ; P3_R1158_U234
g27495 nand P3_R1158_U418 P3_R1158_U25 ; P3_R1158_U235
g27496 not P3_R1158_U26 ; P3_R1158_U236
g27497 nand P3_R1158_U421 P3_R1158_U24 ; P3_R1158_U237
g27498 nand P3_R1158_U424 P3_R1158_U22 ; P3_R1158_U238
g27499 not P3_R1158_U23 ; P3_R1158_U239
g27500 nand P3_R1158_U24 P3_R1158_U23 ; P3_R1158_U240
g27501 nand P3_U3069 P3_R1158_U239 ; P3_R1158_U241
g27502 nand P3_R1158_U427 P3_R1158_U21 ; P3_R1158_U242
g27503 nand P3_U3083 P3_R1158_U66 ; P3_R1158_U243
g27504 nand P3_R1158_U424 P3_R1158_U22 ; P3_R1158_U244
g27505 nand P3_R1158_U244 P3_R1158_U35 ; P3_R1158_U245
g27506 nand P3_R1158_U123 P3_R1158_U245 ; P3_R1158_U246
g27507 nand P3_R1158_U380 P3_R1158_U23 ; P3_R1158_U247
g27508 nand P3_U3069 P3_R1158_U68 ; P3_R1158_U248
g27509 nand P3_R1158_U124 P3_R1158_U247 ; P3_R1158_U249
g27510 nand P3_R1158_U424 P3_R1158_U22 ; P3_R1158_U250
g27511 nand P3_R1158_U415 P3_R1158_U27 ; P3_R1158_U251
g27512 nand P3_R1158_U251 P3_R1158_U36 ; P3_R1158_U252
g27513 nand P3_R1158_U125 P3_R1158_U252 ; P3_R1158_U253
g27514 nand P3_R1158_U225 P3_R1158_U28 ; P3_R1158_U254
g27515 nand P3_U3063 P3_R1158_U71 ; P3_R1158_U255
g27516 nand P3_R1158_U126 P3_R1158_U254 ; P3_R1158_U256
g27517 nand P3_R1158_U415 P3_R1158_U27 ; P3_R1158_U257
g27518 nand P3_U3082 P3_R1158_U161 ; P3_R1158_U258
g27519 not P3_R1158_U208 ; P3_R1158_U259
g27520 nand P3_R1158_U470 P3_R1158_U49 ; P3_R1158_U260
g27521 not P3_R1158_U50 ; P3_R1158_U261
g27522 nand P3_R1158_U476 P3_R1158_U48 ; P3_R1158_U262
g27523 nand P3_R1158_U479 P3_R1158_U45 ; P3_R1158_U263
g27524 nand P3_R1158_U216 P3_R1158_U6 ; P3_R1158_U264
g27525 nand P3_U3079 P3_R1158_U83 ; P3_R1158_U265
g27526 nand P3_R1158_U127 P3_R1158_U264 ; P3_R1158_U266
g27527 nand P3_R1158_U473 P3_R1158_U46 ; P3_R1158_U267
g27528 nand P3_R1158_U476 P3_R1158_U48 ; P3_R1158_U268
g27529 nand P3_R1158_U268 P3_R1158_U266 ; P3_R1158_U269
g27530 nand P3_R1158_U482 P3_R1158_U44 ; P3_R1158_U270
g27531 nand P3_U3078 P3_R1158_U81 ; P3_R1158_U271
g27532 nand P3_R1158_U485 P3_R1158_U51 ; P3_R1158_U272
g27533 nand P3_R1158_U272 P3_R1158_U203 ; P3_R1158_U273
g27534 nand P3_U3073 P3_R1158_U86 ; P3_R1158_U274
g27535 not P3_R1158_U62 ; P3_R1158_U275
g27536 nand P3_R1158_U488 P3_R1158_U43 ; P3_R1158_U276
g27537 nand P3_R1158_U491 P3_R1158_U41 ; P3_R1158_U277
g27538 not P3_R1158_U42 ; P3_R1158_U278
g27539 nand P3_R1158_U43 P3_R1158_U42 ; P3_R1158_U279
g27540 nand P3_R1158_U80 P3_R1158_U279 ; P3_R1158_U280
g27541 nand P3_U3068 P3_R1158_U278 ; P3_R1158_U281
g27542 nand P3_R1158_U7 P3_R1158_U62 ; P3_R1158_U282
g27543 not P3_R1158_U201 ; P3_R1158_U283
g27544 nand P3_R1158_U494 P3_R1158_U52 ; P3_R1158_U284
g27545 nand P3_R1158_U284 P3_R1158_U201 ; P3_R1158_U285
g27546 nand P3_U3081 P3_R1158_U87 ; P3_R1158_U286
g27547 not P3_R1158_U199 ; P3_R1158_U287
g27548 nand P3_R1158_U497 P3_R1158_U56 ; P3_R1158_U288
g27549 nand P3_R1158_U500 P3_R1158_U53 ; P3_R1158_U289
g27550 nand P3_R1158_U217 P3_R1158_U8 ; P3_R1158_U290
g27551 nand P3_U3074 P3_R1158_U89 ; P3_R1158_U291
g27552 nand P3_R1158_U132 P3_R1158_U290 ; P3_R1158_U292
g27553 nand P3_R1158_U503 P3_R1158_U54 ; P3_R1158_U293
g27554 nand P3_R1158_U497 P3_R1158_U56 ; P3_R1158_U294
g27555 nand P3_R1158_U131 P3_R1158_U199 ; P3_R1158_U295
g27556 nand P3_R1158_U294 P3_R1158_U292 ; P3_R1158_U296
g27557 not P3_R1158_U196 ; P3_R1158_U297
g27558 nand P3_R1158_U506 P3_R1158_U57 ; P3_R1158_U298
g27559 nand P3_R1158_U298 P3_R1158_U196 ; P3_R1158_U299
g27560 nand P3_U3060 P3_R1158_U91 ; P3_R1158_U300
g27561 not P3_R1158_U194 ; P3_R1158_U301
g27562 nand P3_R1158_U509 P3_R1158_U58 ; P3_R1158_U302
g27563 nand P3_R1158_U302 P3_R1158_U194 ; P3_R1158_U303
g27564 nand P3_U3065 P3_R1158_U92 ; P3_R1158_U304
g27565 not P3_R1158_U192 ; P3_R1158_U305
g27566 nand P3_R1158_U515 P3_R1158_U38 ; P3_R1158_U306
g27567 nand P3_R1158_U60 P3_R1158_U59 P3_R1158_U308 ; P3_R1158_U307
g27568 nand P3_U3056 P3_R1158_U78 ; P3_R1158_U308
g27569 nand P3_R1158_U518 P3_R1158_U39 ; P3_R1158_U309
g27570 nand P3_R1158_U369 P3_R1158_U192 ; P3_R1158_U310
g27571 nand P3_R1158_U366 P3_R1158_U307 ; P3_R1158_U311
g27572 not P3_R1158_U189 ; P3_R1158_U312
g27573 nand P3_R1158_U467 P3_R1158_U37 ; P3_R1158_U313
g27574 nand P3_U3052 P3_R1158_U75 ; P3_R1158_U314
g27575 nand P3_U3052 P3_R1158_U75 ; P3_R1158_U315
g27576 nand P3_R1158_U467 P3_R1158_U37 ; P3_R1158_U316
g27577 not P3_R1158_U190 ; P3_R1158_U317
g27578 not P3_R1158_U191 ; P3_R1158_U318
g27579 nand P3_R1158_U138 P3_R1158_U12 ; P3_R1158_U319
g27580 nand P3_U3056 P3_R1158_U78 ; P3_R1158_U320
g27581 nand P3_R1158_U515 P3_R1158_U38 ; P3_R1158_U321
g27582 nand P3_R1158_U293 P3_R1158_U199 ; P3_R1158_U322
g27583 not P3_R1158_U61 ; P3_R1158_U323
g27584 nand P3_R1158_U500 P3_R1158_U53 ; P3_R1158_U324
g27585 nand P3_R1158_U324 P3_R1158_U61 ; P3_R1158_U325
g27586 nand P3_R1158_U143 P3_R1158_U325 ; P3_R1158_U326
g27587 nand P3_R1158_U323 P3_R1158_U214 ; P3_R1158_U327
g27588 nand P3_U3074 P3_R1158_U89 ; P3_R1158_U328
g27589 nand P3_R1158_U144 P3_R1158_U327 ; P3_R1158_U329
g27590 nand P3_R1158_U500 P3_R1158_U53 ; P3_R1158_U330
g27591 nand P3_R1158_U491 P3_R1158_U41 ; P3_R1158_U331
g27592 nand P3_R1158_U331 P3_R1158_U62 ; P3_R1158_U332
g27593 nand P3_R1158_U145 P3_R1158_U332 ; P3_R1158_U333
g27594 nand P3_R1158_U275 P3_R1158_U42 ; P3_R1158_U334
g27595 nand P3_U3068 P3_R1158_U80 ; P3_R1158_U335
g27596 nand P3_R1158_U146 P3_R1158_U334 ; P3_R1158_U336
g27597 nand P3_R1158_U491 P3_R1158_U41 ; P3_R1158_U337
g27598 nand P3_R1158_U267 P3_R1158_U206 ; P3_R1158_U338
g27599 not P3_R1158_U64 ; P3_R1158_U339
g27600 nand P3_R1158_U479 P3_R1158_U45 ; P3_R1158_U340
g27601 nand P3_R1158_U340 P3_R1158_U64 ; P3_R1158_U341
g27602 nand P3_R1158_U147 P3_R1158_U341 ; P3_R1158_U342
g27603 nand P3_R1158_U339 P3_R1158_U213 ; P3_R1158_U343
g27604 nand P3_U3079 P3_R1158_U83 ; P3_R1158_U344
g27605 nand P3_R1158_U148 P3_R1158_U343 ; P3_R1158_U345
g27606 nand P3_R1158_U479 P3_R1158_U45 ; P3_R1158_U346
g27607 nand P3_R1158_U250 P3_R1158_U23 ; P3_R1158_U347
g27608 nand P3_R1158_U257 P3_R1158_U28 ; P3_R1158_U348
g27609 nand P3_R1158_U321 P3_R1158_U59 ; P3_R1158_U349
g27610 nand P3_R1158_U309 P3_R1158_U60 ; P3_R1158_U350
g27611 nand P3_R1158_U330 P3_R1158_U214 ; P3_R1158_U351
g27612 nand P3_R1158_U293 P3_R1158_U55 ; P3_R1158_U352
g27613 nand P3_R1158_U337 P3_R1158_U42 ; P3_R1158_U353
g27614 nand P3_R1158_U346 P3_R1158_U213 ; P3_R1158_U354
g27615 nand P3_R1158_U267 P3_R1158_U47 ; P3_R1158_U355
g27616 nand P3_U3059 P3_R1158_U74 ; P3_R1158_U356
g27617 nand P3_U3082 P3_R1158_U65 ; P3_R1158_U357
g27618 nand P3_R1158_U133 P3_R1158_U310 ; P3_R1158_U358
g27619 nand P3_R1158_U68 P3_R1158_U240 ; P3_R1158_U359
g27620 nand P3_U3076 P3_R1158_U219 P3_R1158_U223 ; P3_R1158_U360
g27621 nand P3_R1158_U119 P3_R1158_U223 ; P3_R1158_U361
g27622 nand P3_R1158_U236 P3_R1158_U5 ; P3_R1158_U362
g27623 not P3_R1158_U34 ; P3_R1158_U363
g27624 nand P3_R1158_U34 P3_R1158_U242 ; P3_R1158_U364
g27625 nand P3_R1158_U261 P3_R1158_U9 ; P3_R1158_U365
g27626 nand P3_R1158_U367 P3_R1158_U308 P3_R1158_U19 ; P3_R1158_U366
g27627 nand P3_R1158_U78 P3_R1158_U306 ; P3_R1158_U367
g27628 not P3_R1158_U19 ; P3_R1158_U368
g27629 nand P3_R1158_U371 P3_R1158_U370 ; P3_R1158_U369
g27630 nand P3_R1158_U309 P3_R1158_U306 P3_R1158_U78 ; P3_R1158_U370
g27631 nand P3_R1158_U368 P3_R1158_U309 ; P3_R1158_U371
g27632 not P3_R1158_U63 ; P3_R1158_U372
g27633 nand P3_R1158_U63 P3_R1158_U270 ; P3_R1158_U373
g27634 nand P3_R1158_U134 P3_R1158_U366 ; P3_R1158_U374
g27635 nand P3_R1158_U135 P3_R1158_U192 ; P3_R1158_U375
g27636 nand P3_R1158_U378 P3_R1158_U377 ; P3_R1158_U376
g27637 nand P3_R1158_U60 P3_R1158_U59 P3_R1158_U308 ; P3_R1158_U377
g27638 nand P3_R1158_U367 P3_R1158_U308 P3_R1158_U19 ; P3_R1158_U378
g27639 nand P3_R1158_U235 P3_R1158_U165 ; P3_R1158_U379
g27640 not P3_R1158_U35 ; P3_R1158_U380
g27641 nand P3_R1158_U10 P3_R1158_U165 ; P3_R1158_U381
g27642 not P3_R1158_U163 ; P3_R1158_U382
g27643 nand P3_R1158_U121 P3_R1158_U165 ; P3_R1158_U383
g27644 not P3_R1158_U161 ; P3_R1158_U384
g27645 nand P3_R1158_U260 P3_R1158_U208 ; P3_R1158_U385
g27646 not P3_R1158_U206 ; P3_R1158_U386
g27647 nand P3_R1158_U11 P3_R1158_U208 ; P3_R1158_U387
g27648 not P3_R1158_U205 ; P3_R1158_U388
g27649 nand P3_R1158_U128 P3_R1158_U208 ; P3_R1158_U389
g27650 not P3_R1158_U203 ; P3_R1158_U390
g27651 nand P3_R1158_U139 P3_R1158_U209 ; P3_R1158_U391
g27652 nand P3_R1158_U140 P3_R1158_U209 ; P3_R1158_U392
g27653 nand P3_U3152 P3_R1158_U150 ; P3_R1158_U393
g27654 nand P3_U3416 P3_R1158_U20 ; P3_R1158_U394
g27655 not P3_R1158_U65 ; P3_R1158_U395
g27656 nand P3_R1158_U395 P3_U3082 ; P3_R1158_U396
g27657 nand P3_R1158_U65 P3_R1158_U33 ; P3_R1158_U397
g27658 nand P3_R1158_U395 P3_U3082 ; P3_R1158_U398
g27659 nand P3_R1158_U65 P3_R1158_U33 ; P3_R1158_U399
g27660 nand P3_R1158_U399 P3_R1158_U398 ; P3_R1158_U400
g27661 nand P3_U3152 P3_R1158_U152 ; P3_R1158_U401
g27662 nand P3_U3401 P3_R1158_U20 ; P3_R1158_U402
g27663 not P3_R1158_U74 ; P3_R1158_U403
g27664 nand P3_U3152 P3_R1158_U153 ; P3_R1158_U404
g27665 nand P3_U3392 P3_R1158_U20 ; P3_R1158_U405
g27666 not P3_R1158_U72 ; P3_R1158_U406
g27667 nand P3_U3152 P3_R1158_U154 ; P3_R1158_U407
g27668 nand P3_U3387 P3_R1158_U20 ; P3_R1158_U408
g27669 not P3_R1158_U73 ; P3_R1158_U409
g27670 nand P3_U3152 P3_R1158_U155 ; P3_R1158_U410
g27671 nand P3_U3398 P3_R1158_U20 ; P3_R1158_U411
g27672 not P3_R1158_U71 ; P3_R1158_U412
g27673 nand P3_U3152 P3_R1158_U156 ; P3_R1158_U413
g27674 nand P3_U3395 P3_R1158_U20 ; P3_R1158_U414
g27675 not P3_R1158_U70 ; P3_R1158_U415
g27676 nand P3_U3152 P3_R1158_U157 ; P3_R1158_U416
g27677 nand P3_U3404 P3_R1158_U20 ; P3_R1158_U417
g27678 not P3_R1158_U69 ; P3_R1158_U418
g27679 nand P3_U3152 P3_R1158_U158 ; P3_R1158_U419
g27680 nand P3_U3410 P3_R1158_U20 ; P3_R1158_U420
g27681 not P3_R1158_U68 ; P3_R1158_U421
g27682 nand P3_U3152 P3_R1158_U159 ; P3_R1158_U422
g27683 nand P3_U3407 P3_R1158_U20 ; P3_R1158_U423
g27684 not P3_R1158_U67 ; P3_R1158_U424
g27685 nand P3_U3152 P3_R1158_U160 ; P3_R1158_U425
g27686 nand P3_U3413 P3_R1158_U20 ; P3_R1158_U426
g27687 not P3_R1158_U66 ; P3_R1158_U427
g27688 nand P3_R1158_U151 P3_R1158_U161 ; P3_R1158_U428
g27689 nand P3_R1158_U384 P3_R1158_U400 ; P3_R1158_U429
g27690 nand P3_R1158_U427 P3_U3083 ; P3_R1158_U430
g27691 nand P3_R1158_U66 P3_R1158_U21 ; P3_R1158_U431
g27692 nand P3_R1158_U427 P3_U3083 ; P3_R1158_U432
g27693 nand P3_R1158_U66 P3_R1158_U21 ; P3_R1158_U433
g27694 nand P3_R1158_U433 P3_R1158_U432 ; P3_R1158_U434
g27695 nand P3_R1158_U162 P3_R1158_U163 ; P3_R1158_U435
g27696 nand P3_R1158_U382 P3_R1158_U434 ; P3_R1158_U436
g27697 nand P3_R1158_U421 P3_U3069 ; P3_R1158_U437
g27698 nand P3_R1158_U68 P3_R1158_U24 ; P3_R1158_U438
g27699 nand P3_R1158_U424 P3_U3070 ; P3_R1158_U439
g27700 nand P3_R1158_U67 P3_R1158_U22 ; P3_R1158_U440
g27701 nand P3_R1158_U440 P3_R1158_U439 ; P3_R1158_U441
g27702 nand P3_R1158_U35 P3_R1158_U347 ; P3_R1158_U442
g27703 nand P3_R1158_U441 P3_R1158_U380 ; P3_R1158_U443
g27704 nand P3_R1158_U418 P3_U3066 ; P3_R1158_U444
g27705 nand P3_R1158_U69 P3_R1158_U25 ; P3_R1158_U445
g27706 nand P3_R1158_U418 P3_U3066 ; P3_R1158_U446
g27707 nand P3_R1158_U69 P3_R1158_U25 ; P3_R1158_U447
g27708 nand P3_R1158_U447 P3_R1158_U446 ; P3_R1158_U448
g27709 nand P3_R1158_U164 P3_R1158_U165 ; P3_R1158_U449
g27710 nand P3_R1158_U234 P3_R1158_U448 ; P3_R1158_U450
g27711 nand P3_R1158_U403 P3_U3059 ; P3_R1158_U451
g27712 nand P3_R1158_U74 P3_R1158_U32 ; P3_R1158_U452
g27713 nand P3_R1158_U403 P3_U3059 ; P3_R1158_U453
g27714 nand P3_R1158_U74 P3_R1158_U32 ; P3_R1158_U454
g27715 nand P3_R1158_U454 P3_R1158_U453 ; P3_R1158_U455
g27716 nand P3_R1158_U166 P3_R1158_U167 ; P3_R1158_U456
g27717 nand P3_R1158_U232 P3_R1158_U455 ; P3_R1158_U457
g27718 nand P3_R1158_U412 P3_U3063 ; P3_R1158_U458
g27719 nand P3_R1158_U71 P3_R1158_U29 ; P3_R1158_U459
g27720 nand P3_R1158_U415 P3_U3067 ; P3_R1158_U460
g27721 nand P3_R1158_U70 P3_R1158_U27 ; P3_R1158_U461
g27722 nand P3_R1158_U461 P3_R1158_U460 ; P3_R1158_U462
g27723 nand P3_R1158_U348 P3_R1158_U36 ; P3_R1158_U463
g27724 nand P3_R1158_U462 P3_R1158_U225 ; P3_R1158_U464
g27725 nand P3_U3152 P3_R1158_U168 ; P3_R1158_U465
g27726 nand P3_U3900 P3_R1158_U20 ; P3_R1158_U466
g27727 not P3_R1158_U75 ; P3_R1158_U467
g27728 nand P3_U3152 P3_R1158_U169 ; P3_R1158_U468
g27729 nand P3_U3419 P3_R1158_U20 ; P3_R1158_U469
g27730 not P3_R1158_U85 ; P3_R1158_U470
g27731 nand P3_U3152 P3_R1158_U170 ; P3_R1158_U471
g27732 nand P3_U3422 P3_R1158_U20 ; P3_R1158_U472
g27733 not P3_R1158_U84 ; P3_R1158_U473
g27734 nand P3_U3152 P3_R1158_U171 ; P3_R1158_U474
g27735 nand P3_U3428 P3_R1158_U20 ; P3_R1158_U475
g27736 not P3_R1158_U83 ; P3_R1158_U476
g27737 nand P3_U3152 P3_R1158_U172 ; P3_R1158_U477
g27738 nand P3_U3425 P3_R1158_U20 ; P3_R1158_U478
g27739 not P3_R1158_U82 ; P3_R1158_U479
g27740 nand P3_U3152 P3_R1158_U173 ; P3_R1158_U480
g27741 nand P3_U3431 P3_R1158_U20 ; P3_R1158_U481
g27742 not P3_R1158_U81 ; P3_R1158_U482
g27743 nand P3_U3152 P3_R1158_U174 ; P3_R1158_U483
g27744 nand P3_U3434 P3_R1158_U20 ; P3_R1158_U484
g27745 not P3_R1158_U86 ; P3_R1158_U485
g27746 nand P3_U3152 P3_R1158_U175 ; P3_R1158_U486
g27747 nand P3_U3440 P3_R1158_U20 ; P3_R1158_U487
g27748 not P3_R1158_U80 ; P3_R1158_U488
g27749 nand P3_U3152 P3_R1158_U176 ; P3_R1158_U489
g27750 nand P3_U3437 P3_R1158_U20 ; P3_R1158_U490
g27751 not P3_R1158_U79 ; P3_R1158_U491
g27752 nand P3_U3152 P3_R1158_U177 ; P3_R1158_U492
g27753 nand P3_U3443 P3_R1158_U20 ; P3_R1158_U493
g27754 not P3_R1158_U87 ; P3_R1158_U494
g27755 nand P3_U3152 P3_R1158_U178 ; P3_R1158_U495
g27756 nand P3_U3906 P3_R1158_U20 ; P3_R1158_U496
g27757 not P3_R1158_U89 ; P3_R1158_U497
g27758 nand P3_U3152 P3_R1158_U179 ; P3_R1158_U498
g27759 nand P3_U3907 P3_R1158_U20 ; P3_R1158_U499
g27760 not P3_R1158_U90 ; P3_R1158_U500
g27761 nand P3_U3152 P3_R1158_U180 ; P3_R1158_U501
g27762 nand P3_U3445 P3_R1158_U20 ; P3_R1158_U502
g27763 not P3_R1158_U88 ; P3_R1158_U503
g27764 nand P3_U3152 P3_R1158_U181 ; P3_R1158_U504
g27765 nand P3_U3905 P3_R1158_U20 ; P3_R1158_U505
g27766 not P3_R1158_U91 ; P3_R1158_U506
g27767 nand P3_U3152 P3_R1158_U182 ; P3_R1158_U507
g27768 nand P3_U3904 P3_R1158_U20 ; P3_R1158_U508
g27769 not P3_R1158_U92 ; P3_R1158_U509
g27770 nand P3_U3152 P3_R1158_U183 ; P3_R1158_U510
g27771 nand P3_U3901 P3_R1158_U20 ; P3_R1158_U511
g27772 not P3_R1158_U78 ; P3_R1158_U512
g27773 nand P3_U3152 P3_R1158_U184 ; P3_R1158_U513
g27774 nand P3_U3902 P3_R1158_U20 ; P3_R1158_U514
g27775 not P3_R1158_U76 ; P3_R1158_U515
g27776 nand P3_U3152 P3_R1158_U185 ; P3_R1158_U516
g27777 nand P3_U3903 P3_R1158_U20 ; P3_R1158_U517
g27778 not P3_R1158_U77 ; P3_R1158_U518
g27779 nand P3_U3152 P3_R1158_U186 ; P3_R1158_U519
g27780 nand P3_U3053 P3_R1158_U20 ; P3_R1158_U520
g27781 not P3_R1158_U137 ; P3_R1158_U521
g27782 nand P3_U3899 P3_R1158_U521 ; P3_R1158_U522
g27783 nand P3_R1158_U137 P3_R1158_U187 ; P3_R1158_U523
g27784 not P3_R1158_U93 ; P3_R1158_U524
g27785 nand P3_R1158_U358 P3_R1158_U313 P3_R1158_U524 ; P3_R1158_U525
g27786 nand P3_R1158_U136 P3_R1158_U375 P3_R1158_U93 ; P3_R1158_U526
g27787 nand P3_R1158_U467 P3_U3052 ; P3_R1158_U527
g27788 nand P3_R1158_U75 P3_R1158_U37 ; P3_R1158_U528
g27789 nand P3_R1158_U467 P3_U3052 ; P3_R1158_U529
g27790 nand P3_R1158_U75 P3_R1158_U37 ; P3_R1158_U530
g27791 nand P3_R1158_U530 P3_R1158_U529 ; P3_R1158_U531
g27792 nand P3_R1158_U188 P3_R1158_U189 ; P3_R1158_U532
g27793 nand P3_R1158_U312 P3_R1158_U531 ; P3_R1158_U533
g27794 nand P3_R1158_U512 P3_U3056 ; P3_R1158_U534
g27795 nand P3_R1158_U78 P3_R1158_U40 ; P3_R1158_U535
g27796 nand P3_R1158_U104 P3_R1158_U190 ; P3_R1158_U536
g27797 nand P3_R1158_U103 P3_R1158_U317 ; P3_R1158_U537
g27798 nand P3_R1158_U515 P3_U3057 ; P3_R1158_U538
g27799 nand P3_R1158_U76 P3_R1158_U38 ; P3_R1158_U539
g27800 nand P3_R1158_U539 P3_R1158_U538 ; P3_R1158_U540
g27801 nand P3_R1158_U349 P3_R1158_U191 ; P3_R1158_U541
g27802 nand P3_R1158_U318 P3_R1158_U540 ; P3_R1158_U542
g27803 nand P3_R1158_U518 P3_U3064 ; P3_R1158_U543
g27804 nand P3_R1158_U77 P3_R1158_U39 ; P3_R1158_U544
g27805 nand P3_R1158_U544 P3_R1158_U543 ; P3_R1158_U545
g27806 nand P3_R1158_U350 P3_R1158_U192 ; P3_R1158_U546
g27807 nand P3_R1158_U305 P3_R1158_U545 ; P3_R1158_U547
g27808 nand P3_R1158_U509 P3_U3065 ; P3_R1158_U548
g27809 nand P3_R1158_U92 P3_R1158_U58 ; P3_R1158_U549
g27810 nand P3_R1158_U509 P3_U3065 ; P3_R1158_U550
g27811 nand P3_R1158_U92 P3_R1158_U58 ; P3_R1158_U551
g27812 nand P3_R1158_U551 P3_R1158_U550 ; P3_R1158_U552
g27813 nand P3_R1158_U193 P3_R1158_U194 ; P3_R1158_U553
g27814 nand P3_R1158_U301 P3_R1158_U552 ; P3_R1158_U554
g27815 nand P3_R1158_U506 P3_U3060 ; P3_R1158_U555
g27816 nand P3_R1158_U91 P3_R1158_U57 ; P3_R1158_U556
g27817 nand P3_R1158_U506 P3_U3060 ; P3_R1158_U557
g27818 nand P3_R1158_U91 P3_R1158_U57 ; P3_R1158_U558
g27819 nand P3_R1158_U558 P3_R1158_U557 ; P3_R1158_U559
g27820 nand P3_R1158_U195 P3_R1158_U196 ; P3_R1158_U560
g27821 nand P3_R1158_U297 P3_R1158_U559 ; P3_R1158_U561
g27822 nand P3_R1158_U497 P3_U3074 ; P3_R1158_U562
g27823 nand P3_R1158_U89 P3_R1158_U56 ; P3_R1158_U563
g27824 nand P3_R1158_U500 P3_U3075 ; P3_R1158_U564
g27825 nand P3_R1158_U90 P3_R1158_U53 ; P3_R1158_U565
g27826 nand P3_R1158_U565 P3_R1158_U564 ; P3_R1158_U566
g27827 nand P3_R1158_U351 P3_R1158_U61 ; P3_R1158_U567
g27828 nand P3_R1158_U566 P3_R1158_U323 ; P3_R1158_U568
g27829 nand P3_R1158_U406 P3_U3077 ; P3_R1158_U569
g27830 nand P3_R1158_U72 P3_R1158_U30 ; P3_R1158_U570
g27831 nand P3_R1158_U406 P3_U3077 ; P3_R1158_U571
g27832 nand P3_R1158_U72 P3_R1158_U30 ; P3_R1158_U572
g27833 nand P3_R1158_U572 P3_R1158_U571 ; P3_R1158_U573
g27834 nand P3_R1158_U197 P3_R1158_U198 ; P3_R1158_U574
g27835 nand P3_R1158_U222 P3_R1158_U573 ; P3_R1158_U575
g27836 nand P3_R1158_U503 P3_U3080 ; P3_R1158_U576
g27837 nand P3_R1158_U88 P3_R1158_U54 ; P3_R1158_U577
g27838 nand P3_R1158_U577 P3_R1158_U576 ; P3_R1158_U578
g27839 nand P3_R1158_U352 P3_R1158_U199 ; P3_R1158_U579
g27840 nand P3_R1158_U287 P3_R1158_U578 ; P3_R1158_U580
g27841 nand P3_R1158_U494 P3_U3081 ; P3_R1158_U581
g27842 nand P3_R1158_U87 P3_R1158_U52 ; P3_R1158_U582
g27843 nand P3_R1158_U494 P3_U3081 ; P3_R1158_U583
g27844 nand P3_R1158_U87 P3_R1158_U52 ; P3_R1158_U584
g27845 nand P3_R1158_U584 P3_R1158_U583 ; P3_R1158_U585
g27846 nand P3_R1158_U200 P3_R1158_U201 ; P3_R1158_U586
g27847 nand P3_R1158_U283 P3_R1158_U585 ; P3_R1158_U587
g27848 nand P3_R1158_U488 P3_U3068 ; P3_R1158_U588
g27849 nand P3_R1158_U80 P3_R1158_U43 ; P3_R1158_U589
g27850 nand P3_R1158_U491 P3_U3072 ; P3_R1158_U590
g27851 nand P3_R1158_U79 P3_R1158_U41 ; P3_R1158_U591
g27852 nand P3_R1158_U591 P3_R1158_U590 ; P3_R1158_U592
g27853 nand P3_R1158_U353 P3_R1158_U62 ; P3_R1158_U593
g27854 nand P3_R1158_U592 P3_R1158_U275 ; P3_R1158_U594
g27855 nand P3_R1158_U485 P3_U3073 ; P3_R1158_U595
g27856 nand P3_R1158_U86 P3_R1158_U51 ; P3_R1158_U596
g27857 nand P3_R1158_U485 P3_U3073 ; P3_R1158_U597
g27858 nand P3_R1158_U86 P3_R1158_U51 ; P3_R1158_U598
g27859 nand P3_R1158_U598 P3_R1158_U597 ; P3_R1158_U599
g27860 nand P3_R1158_U202 P3_R1158_U203 ; P3_R1158_U600
g27861 nand P3_R1158_U390 P3_R1158_U599 ; P3_R1158_U601
g27862 nand P3_R1158_U482 P3_U3078 ; P3_R1158_U602
g27863 nand P3_R1158_U81 P3_R1158_U44 ; P3_R1158_U603
g27864 nand P3_R1158_U482 P3_U3078 ; P3_R1158_U604
g27865 nand P3_R1158_U81 P3_R1158_U44 ; P3_R1158_U605
g27866 nand P3_R1158_U605 P3_R1158_U604 ; P3_R1158_U606
g27867 nand P3_R1158_U204 P3_R1158_U205 ; P3_R1158_U607
g27868 nand P3_R1158_U388 P3_R1158_U606 ; P3_R1158_U608
g27869 nand P3_R1158_U476 P3_U3079 ; P3_R1158_U609
g27870 nand P3_R1158_U83 P3_R1158_U48 ; P3_R1158_U610
g27871 nand P3_R1158_U479 P3_U3071 ; P3_R1158_U611
g27872 nand P3_R1158_U82 P3_R1158_U45 ; P3_R1158_U612
g27873 nand P3_R1158_U612 P3_R1158_U611 ; P3_R1158_U613
g27874 nand P3_R1158_U354 P3_R1158_U64 ; P3_R1158_U614
g27875 nand P3_R1158_U613 P3_R1158_U339 ; P3_R1158_U615
g27876 nand P3_R1158_U473 P3_U3062 ; P3_R1158_U616
g27877 nand P3_R1158_U84 P3_R1158_U46 ; P3_R1158_U617
g27878 nand P3_R1158_U617 P3_R1158_U616 ; P3_R1158_U618
g27879 nand P3_R1158_U206 P3_R1158_U355 ; P3_R1158_U619
g27880 nand P3_R1158_U386 P3_R1158_U618 ; P3_R1158_U620
g27881 nand P3_R1158_U470 P3_U3061 ; P3_R1158_U621
g27882 nand P3_R1158_U85 P3_R1158_U49 ; P3_R1158_U622
g27883 nand P3_R1158_U470 P3_U3061 ; P3_R1158_U623
g27884 nand P3_R1158_U85 P3_R1158_U49 ; P3_R1158_U624
g27885 nand P3_R1158_U624 P3_R1158_U623 ; P3_R1158_U625
g27886 nand P3_R1158_U207 P3_R1158_U208 ; P3_R1158_U626
g27887 nand P3_R1158_U259 P3_R1158_U625 ; P3_R1158_U627
g27888 nand P3_R1158_U73 P3_R1158_U20 ; P3_R1158_U628
g27889 nand P3_R1158_U409 P3_U3152 ; P3_R1158_U629
g27890 not P3_R1158_U149 ; P3_R1158_U630
g27891 nand P3_R1158_U630 P3_U3076 ; P3_R1158_U631
g27892 nand P3_R1158_U149 P3_R1158_U31 ; P3_R1158_U632
g27893 and P3_R1131_U210 P3_R1131_U209 ; P3_R1131_U6
g27894 and P3_R1131_U189 P3_R1131_U245 ; P3_R1131_U7
g27895 and P3_R1131_U247 P3_R1131_U246 ; P3_R1131_U8
g27896 and P3_R1131_U190 P3_R1131_U262 ; P3_R1131_U9
g27897 and P3_R1131_U264 P3_R1131_U263 ; P3_R1131_U10
g27898 and P3_R1131_U191 P3_R1131_U286 ; P3_R1131_U11
g27899 and P3_R1131_U288 P3_R1131_U287 ; P3_R1131_U12
g27900 and P3_R1131_U208 P3_R1131_U194 P3_R1131_U213 ; P3_R1131_U13
g27901 and P3_R1131_U218 P3_R1131_U195 ; P3_R1131_U14
g27902 and P3_R1131_U392 P3_R1131_U391 ; P3_R1131_U15
g27903 nand P3_R1131_U342 P3_R1131_U345 ; P3_R1131_U16
g27904 nand P3_R1131_U331 P3_R1131_U334 ; P3_R1131_U17
g27905 nand P3_R1131_U320 P3_R1131_U323 ; P3_R1131_U18
g27906 nand P3_R1131_U312 P3_R1131_U314 ; P3_R1131_U19
g27907 nand P3_R1131_U162 P3_R1131_U183 P3_R1131_U351 ; P3_R1131_U20
g27908 nand P3_R1131_U241 P3_R1131_U243 ; P3_R1131_U21
g27909 nand P3_R1131_U233 P3_R1131_U236 ; P3_R1131_U22
g27910 nand P3_R1131_U225 P3_R1131_U227 ; P3_R1131_U23
g27911 nand P3_R1131_U172 P3_R1131_U348 ; P3_R1131_U24
g27912 not P3_U3069 ; P3_R1131_U25
g27913 nand P3_U3069 P3_R1131_U39 ; P3_R1131_U26
g27914 not P3_U3083 ; P3_R1131_U27
g27915 not P3_U3413 ; P3_R1131_U28
g27916 not P3_U3395 ; P3_R1131_U29
g27917 not P3_U3387 ; P3_R1131_U30
g27918 not P3_U3077 ; P3_R1131_U31
g27919 not P3_U3398 ; P3_R1131_U32
g27920 not P3_U3067 ; P3_R1131_U33
g27921 nand P3_U3067 P3_R1131_U29 ; P3_R1131_U34
g27922 not P3_U3063 ; P3_R1131_U35
g27923 not P3_U3404 ; P3_R1131_U36
g27924 not P3_U3407 ; P3_R1131_U37
g27925 not P3_U3401 ; P3_R1131_U38
g27926 not P3_U3410 ; P3_R1131_U39
g27927 not P3_U3070 ; P3_R1131_U40
g27928 not P3_U3066 ; P3_R1131_U41
g27929 not P3_U3059 ; P3_R1131_U42
g27930 nand P3_U3059 P3_R1131_U38 ; P3_R1131_U43
g27931 nand P3_R1131_U214 P3_R1131_U212 ; P3_R1131_U44
g27932 not P3_U3416 ; P3_R1131_U45
g27933 not P3_U3082 ; P3_R1131_U46
g27934 nand P3_R1131_U44 P3_R1131_U215 ; P3_R1131_U47
g27935 nand P3_R1131_U43 P3_R1131_U229 ; P3_R1131_U48
g27936 nand P3_R1131_U201 P3_R1131_U185 P3_R1131_U349 ; P3_R1131_U49
g27937 not P3_U3901 ; P3_R1131_U50
g27938 not P3_U3422 ; P3_R1131_U51
g27939 not P3_U3419 ; P3_R1131_U52
g27940 not P3_U3062 ; P3_R1131_U53
g27941 not P3_U3061 ; P3_R1131_U54
g27942 nand P3_U3082 P3_R1131_U45 ; P3_R1131_U55
g27943 not P3_U3425 ; P3_R1131_U56
g27944 not P3_U3071 ; P3_R1131_U57
g27945 not P3_U3428 ; P3_R1131_U58
g27946 not P3_U3079 ; P3_R1131_U59
g27947 not P3_U3437 ; P3_R1131_U60
g27948 not P3_U3434 ; P3_R1131_U61
g27949 not P3_U3431 ; P3_R1131_U62
g27950 not P3_U3072 ; P3_R1131_U63
g27951 not P3_U3073 ; P3_R1131_U64
g27952 not P3_U3078 ; P3_R1131_U65
g27953 nand P3_U3078 P3_R1131_U62 ; P3_R1131_U66
g27954 not P3_U3440 ; P3_R1131_U67
g27955 not P3_U3068 ; P3_R1131_U68
g27956 not P3_U3081 ; P3_R1131_U69
g27957 not P3_U3445 ; P3_R1131_U70
g27958 not P3_U3080 ; P3_R1131_U71
g27959 not P3_U3907 ; P3_R1131_U72
g27960 not P3_U3075 ; P3_R1131_U73
g27961 not P3_U3904 ; P3_R1131_U74
g27962 not P3_U3905 ; P3_R1131_U75
g27963 not P3_U3906 ; P3_R1131_U76
g27964 not P3_U3065 ; P3_R1131_U77
g27965 not P3_U3060 ; P3_R1131_U78
g27966 not P3_U3074 ; P3_R1131_U79
g27967 nand P3_U3074 P3_R1131_U76 ; P3_R1131_U80
g27968 not P3_U3903 ; P3_R1131_U81
g27969 not P3_U3064 ; P3_R1131_U82
g27970 not P3_U3902 ; P3_R1131_U83
g27971 not P3_U3057 ; P3_R1131_U84
g27972 not P3_U3900 ; P3_R1131_U85
g27973 not P3_U3056 ; P3_R1131_U86
g27974 nand P3_U3056 P3_R1131_U50 ; P3_R1131_U87
g27975 not P3_U3052 ; P3_R1131_U88
g27976 not P3_U3899 ; P3_R1131_U89
g27977 not P3_U3053 ; P3_R1131_U90
g27978 nand P3_R1131_U302 P3_R1131_U301 ; P3_R1131_U91
g27979 nand P3_R1131_U80 P3_R1131_U316 ; P3_R1131_U92
g27980 nand P3_R1131_U66 P3_R1131_U327 ; P3_R1131_U93
g27981 nand P3_R1131_U55 P3_R1131_U338 ; P3_R1131_U94
g27982 not P3_U3076 ; P3_R1131_U95
g27983 nand P3_R1131_U402 P3_R1131_U401 ; P3_R1131_U96
g27984 nand P3_R1131_U416 P3_R1131_U415 ; P3_R1131_U97
g27985 nand P3_R1131_U421 P3_R1131_U420 ; P3_R1131_U98
g27986 nand P3_R1131_U437 P3_R1131_U436 ; P3_R1131_U99
g27987 nand P3_R1131_U442 P3_R1131_U441 ; P3_R1131_U100
g27988 nand P3_R1131_U447 P3_R1131_U446 ; P3_R1131_U101
g27989 nand P3_R1131_U452 P3_R1131_U451 ; P3_R1131_U102
g27990 nand P3_R1131_U457 P3_R1131_U456 ; P3_R1131_U103
g27991 nand P3_R1131_U473 P3_R1131_U472 ; P3_R1131_U104
g27992 nand P3_R1131_U478 P3_R1131_U477 ; P3_R1131_U105
g27993 nand P3_R1131_U361 P3_R1131_U360 ; P3_R1131_U106
g27994 nand P3_R1131_U370 P3_R1131_U369 ; P3_R1131_U107
g27995 nand P3_R1131_U377 P3_R1131_U376 ; P3_R1131_U108
g27996 nand P3_R1131_U381 P3_R1131_U380 ; P3_R1131_U109
g27997 nand P3_R1131_U390 P3_R1131_U389 ; P3_R1131_U110
g27998 nand P3_R1131_U411 P3_R1131_U410 ; P3_R1131_U111
g27999 nand P3_R1131_U428 P3_R1131_U427 ; P3_R1131_U112
g28000 nand P3_R1131_U432 P3_R1131_U431 ; P3_R1131_U113
g28001 nand P3_R1131_U464 P3_R1131_U463 ; P3_R1131_U114
g28002 nand P3_R1131_U468 P3_R1131_U467 ; P3_R1131_U115
g28003 nand P3_R1131_U485 P3_R1131_U484 ; P3_R1131_U116
g28004 and P3_R1131_U352 P3_R1131_U193 ; P3_R1131_U117
g28005 and P3_R1131_U205 P3_R1131_U206 ; P3_R1131_U118
g28006 and P3_R1131_U14 P3_R1131_U13 ; P3_R1131_U119
g28007 and P3_R1131_U357 P3_R1131_U354 ; P3_R1131_U120
g28008 and P3_R1131_U363 P3_R1131_U362 P3_R1131_U26 ; P3_R1131_U121
g28009 and P3_R1131_U366 P3_R1131_U195 ; P3_R1131_U122
g28010 and P3_R1131_U235 P3_R1131_U6 ; P3_R1131_U123
g28011 and P3_R1131_U373 P3_R1131_U194 ; P3_R1131_U124
g28012 and P3_R1131_U383 P3_R1131_U382 P3_R1131_U34 ; P3_R1131_U125
g28013 and P3_R1131_U386 P3_R1131_U193 ; P3_R1131_U126
g28014 and P3_R1131_U222 P3_R1131_U7 ; P3_R1131_U127
g28015 and P3_R1131_U267 P3_R1131_U9 ; P3_R1131_U128
g28016 and P3_R1131_U291 P3_R1131_U11 ; P3_R1131_U129
g28017 and P3_R1131_U355 P3_R1131_U192 ; P3_R1131_U130
g28018 and P3_R1131_U306 P3_R1131_U307 ; P3_R1131_U131
g28019 and P3_R1131_U309 P3_R1131_U395 ; P3_R1131_U132
g28020 and P3_R1131_U306 P3_R1131_U307 ; P3_R1131_U133
g28021 and P3_R1131_U15 P3_R1131_U310 ; P3_R1131_U134
g28022 nand P3_R1131_U399 P3_R1131_U398 ; P3_R1131_U135
g28023 and P3_R1131_U404 P3_R1131_U403 P3_R1131_U87 ; P3_R1131_U136
g28024 and P3_R1131_U407 P3_R1131_U192 ; P3_R1131_U137
g28025 nand P3_R1131_U413 P3_R1131_U412 ; P3_R1131_U138
g28026 nand P3_R1131_U418 P3_R1131_U417 ; P3_R1131_U139
g28027 and P3_R1131_U322 P3_R1131_U12 ; P3_R1131_U140
g28028 and P3_R1131_U424 P3_R1131_U191 ; P3_R1131_U141
g28029 nand P3_R1131_U434 P3_R1131_U433 ; P3_R1131_U142
g28030 nand P3_R1131_U439 P3_R1131_U438 ; P3_R1131_U143
g28031 nand P3_R1131_U444 P3_R1131_U443 ; P3_R1131_U144
g28032 nand P3_R1131_U449 P3_R1131_U448 ; P3_R1131_U145
g28033 nand P3_R1131_U454 P3_R1131_U453 ; P3_R1131_U146
g28034 and P3_R1131_U333 P3_R1131_U10 ; P3_R1131_U147
g28035 and P3_R1131_U460 P3_R1131_U190 ; P3_R1131_U148
g28036 nand P3_R1131_U470 P3_R1131_U469 ; P3_R1131_U149
g28037 nand P3_R1131_U475 P3_R1131_U474 ; P3_R1131_U150
g28038 and P3_R1131_U344 P3_R1131_U8 ; P3_R1131_U151
g28039 and P3_R1131_U481 P3_R1131_U189 ; P3_R1131_U152
g28040 and P3_R1131_U359 P3_R1131_U358 ; P3_R1131_U153
g28041 nand P3_R1131_U120 P3_R1131_U356 ; P3_R1131_U154
g28042 and P3_R1131_U368 P3_R1131_U367 ; P3_R1131_U155
g28043 and P3_R1131_U375 P3_R1131_U374 ; P3_R1131_U156
g28044 and P3_R1131_U379 P3_R1131_U378 ; P3_R1131_U157
g28045 nand P3_R1131_U118 P3_R1131_U203 ; P3_R1131_U158
g28046 and P3_R1131_U388 P3_R1131_U387 ; P3_R1131_U159
g28047 not P3_U3908 ; P3_R1131_U160
g28048 not P3_U3054 ; P3_R1131_U161
g28049 and P3_R1131_U397 P3_R1131_U396 ; P3_R1131_U162
g28050 nand P3_R1131_U131 P3_R1131_U304 ; P3_R1131_U163
g28051 and P3_R1131_U409 P3_R1131_U408 ; P3_R1131_U164
g28052 nand P3_R1131_U298 P3_R1131_U297 ; P3_R1131_U165
g28053 nand P3_R1131_U294 P3_R1131_U293 ; P3_R1131_U166
g28054 and P3_R1131_U426 P3_R1131_U425 ; P3_R1131_U167
g28055 and P3_R1131_U430 P3_R1131_U429 ; P3_R1131_U168
g28056 nand P3_R1131_U284 P3_R1131_U283 ; P3_R1131_U169
g28057 nand P3_R1131_U280 P3_R1131_U279 ; P3_R1131_U170
g28058 not P3_U3392 ; P3_R1131_U171
g28059 nand P3_U3387 P3_R1131_U95 ; P3_R1131_U172
g28060 nand P3_R1131_U276 P3_R1131_U184 P3_R1131_U350 ; P3_R1131_U173
g28061 not P3_U3443 ; P3_R1131_U174
g28062 nand P3_R1131_U274 P3_R1131_U273 ; P3_R1131_U175
g28063 nand P3_R1131_U270 P3_R1131_U269 ; P3_R1131_U176
g28064 and P3_R1131_U462 P3_R1131_U461 ; P3_R1131_U177
g28065 and P3_R1131_U466 P3_R1131_U465 ; P3_R1131_U178
g28066 nand P3_R1131_U260 P3_R1131_U259 ; P3_R1131_U179
g28067 nand P3_R1131_U256 P3_R1131_U255 ; P3_R1131_U180
g28068 nand P3_R1131_U252 P3_R1131_U251 ; P3_R1131_U181
g28069 and P3_R1131_U483 P3_R1131_U482 ; P3_R1131_U182
g28070 nand P3_R1131_U132 P3_R1131_U163 ; P3_R1131_U183
g28071 nand P3_R1131_U175 P3_R1131_U174 ; P3_R1131_U184
g28072 nand P3_R1131_U172 P3_R1131_U171 ; P3_R1131_U185
g28073 not P3_R1131_U87 ; P3_R1131_U186
g28074 not P3_R1131_U34 ; P3_R1131_U187
g28075 not P3_R1131_U26 ; P3_R1131_U188
g28076 nand P3_U3419 P3_R1131_U54 ; P3_R1131_U189
g28077 nand P3_U3434 P3_R1131_U64 ; P3_R1131_U190
g28078 nand P3_U3905 P3_R1131_U78 ; P3_R1131_U191
g28079 nand P3_U3901 P3_R1131_U86 ; P3_R1131_U192
g28080 nand P3_U3395 P3_R1131_U33 ; P3_R1131_U193
g28081 nand P3_U3404 P3_R1131_U41 ; P3_R1131_U194
g28082 nand P3_U3410 P3_R1131_U25 ; P3_R1131_U195
g28083 not P3_R1131_U66 ; P3_R1131_U196
g28084 not P3_R1131_U80 ; P3_R1131_U197
g28085 not P3_R1131_U43 ; P3_R1131_U198
g28086 not P3_R1131_U55 ; P3_R1131_U199
g28087 not P3_R1131_U172 ; P3_R1131_U200
g28088 nand P3_U3077 P3_R1131_U172 ; P3_R1131_U201
g28089 not P3_R1131_U49 ; P3_R1131_U202
g28090 nand P3_R1131_U117 P3_R1131_U49 ; P3_R1131_U203
g28091 nand P3_R1131_U35 P3_R1131_U34 ; P3_R1131_U204
g28092 nand P3_R1131_U204 P3_R1131_U32 ; P3_R1131_U205
g28093 nand P3_U3063 P3_R1131_U187 ; P3_R1131_U206
g28094 not P3_R1131_U158 ; P3_R1131_U207
g28095 nand P3_U3407 P3_R1131_U40 ; P3_R1131_U208
g28096 nand P3_U3070 P3_R1131_U37 ; P3_R1131_U209
g28097 nand P3_U3066 P3_R1131_U36 ; P3_R1131_U210
g28098 nand P3_R1131_U198 P3_R1131_U194 ; P3_R1131_U211
g28099 nand P3_R1131_U6 P3_R1131_U211 ; P3_R1131_U212
g28100 nand P3_U3401 P3_R1131_U42 ; P3_R1131_U213
g28101 nand P3_U3407 P3_R1131_U40 ; P3_R1131_U214
g28102 nand P3_R1131_U13 P3_R1131_U158 ; P3_R1131_U215
g28103 not P3_R1131_U44 ; P3_R1131_U216
g28104 not P3_R1131_U47 ; P3_R1131_U217
g28105 nand P3_U3413 P3_R1131_U27 ; P3_R1131_U218
g28106 nand P3_R1131_U27 P3_R1131_U26 ; P3_R1131_U219
g28107 nand P3_U3083 P3_R1131_U188 ; P3_R1131_U220
g28108 not P3_R1131_U154 ; P3_R1131_U221
g28109 nand P3_U3416 P3_R1131_U46 ; P3_R1131_U222
g28110 nand P3_R1131_U222 P3_R1131_U55 ; P3_R1131_U223
g28111 nand P3_R1131_U217 P3_R1131_U26 ; P3_R1131_U224
g28112 nand P3_R1131_U122 P3_R1131_U224 ; P3_R1131_U225
g28113 nand P3_R1131_U47 P3_R1131_U195 ; P3_R1131_U226
g28114 nand P3_R1131_U121 P3_R1131_U226 ; P3_R1131_U227
g28115 nand P3_R1131_U26 P3_R1131_U195 ; P3_R1131_U228
g28116 nand P3_R1131_U213 P3_R1131_U158 ; P3_R1131_U229
g28117 not P3_R1131_U48 ; P3_R1131_U230
g28118 nand P3_U3066 P3_R1131_U36 ; P3_R1131_U231
g28119 nand P3_R1131_U230 P3_R1131_U231 ; P3_R1131_U232
g28120 nand P3_R1131_U124 P3_R1131_U232 ; P3_R1131_U233
g28121 nand P3_R1131_U48 P3_R1131_U194 ; P3_R1131_U234
g28122 nand P3_U3407 P3_R1131_U40 ; P3_R1131_U235
g28123 nand P3_R1131_U123 P3_R1131_U234 ; P3_R1131_U236
g28124 nand P3_U3066 P3_R1131_U36 ; P3_R1131_U237
g28125 nand P3_R1131_U194 P3_R1131_U237 ; P3_R1131_U238
g28126 nand P3_R1131_U213 P3_R1131_U43 ; P3_R1131_U239
g28127 nand P3_R1131_U202 P3_R1131_U34 ; P3_R1131_U240
g28128 nand P3_R1131_U126 P3_R1131_U240 ; P3_R1131_U241
g28129 nand P3_R1131_U49 P3_R1131_U193 ; P3_R1131_U242
g28130 nand P3_R1131_U125 P3_R1131_U242 ; P3_R1131_U243
g28131 nand P3_R1131_U193 P3_R1131_U34 ; P3_R1131_U244
g28132 nand P3_U3422 P3_R1131_U53 ; P3_R1131_U245
g28133 nand P3_U3062 P3_R1131_U51 ; P3_R1131_U246
g28134 nand P3_U3061 P3_R1131_U52 ; P3_R1131_U247
g28135 nand P3_R1131_U199 P3_R1131_U7 ; P3_R1131_U248
g28136 nand P3_R1131_U8 P3_R1131_U248 ; P3_R1131_U249
g28137 nand P3_U3422 P3_R1131_U53 ; P3_R1131_U250
g28138 nand P3_R1131_U127 P3_R1131_U154 ; P3_R1131_U251
g28139 nand P3_R1131_U250 P3_R1131_U249 ; P3_R1131_U252
g28140 not P3_R1131_U181 ; P3_R1131_U253
g28141 nand P3_U3425 P3_R1131_U57 ; P3_R1131_U254
g28142 nand P3_R1131_U254 P3_R1131_U181 ; P3_R1131_U255
g28143 nand P3_U3071 P3_R1131_U56 ; P3_R1131_U256
g28144 not P3_R1131_U180 ; P3_R1131_U257
g28145 nand P3_U3428 P3_R1131_U59 ; P3_R1131_U258
g28146 nand P3_R1131_U258 P3_R1131_U180 ; P3_R1131_U259
g28147 nand P3_U3079 P3_R1131_U58 ; P3_R1131_U260
g28148 not P3_R1131_U179 ; P3_R1131_U261
g28149 nand P3_U3437 P3_R1131_U63 ; P3_R1131_U262
g28150 nand P3_U3072 P3_R1131_U60 ; P3_R1131_U263
g28151 nand P3_U3073 P3_R1131_U61 ; P3_R1131_U264
g28152 nand P3_R1131_U196 P3_R1131_U9 ; P3_R1131_U265
g28153 nand P3_R1131_U10 P3_R1131_U265 ; P3_R1131_U266
g28154 nand P3_U3431 P3_R1131_U65 ; P3_R1131_U267
g28155 nand P3_U3437 P3_R1131_U63 ; P3_R1131_U268
g28156 nand P3_R1131_U128 P3_R1131_U179 ; P3_R1131_U269
g28157 nand P3_R1131_U268 P3_R1131_U266 ; P3_R1131_U270
g28158 not P3_R1131_U176 ; P3_R1131_U271
g28159 nand P3_U3440 P3_R1131_U68 ; P3_R1131_U272
g28160 nand P3_R1131_U272 P3_R1131_U176 ; P3_R1131_U273
g28161 nand P3_U3068 P3_R1131_U67 ; P3_R1131_U274
g28162 not P3_R1131_U175 ; P3_R1131_U275
g28163 nand P3_U3081 P3_R1131_U175 ; P3_R1131_U276
g28164 not P3_R1131_U173 ; P3_R1131_U277
g28165 nand P3_U3445 P3_R1131_U71 ; P3_R1131_U278
g28166 nand P3_R1131_U278 P3_R1131_U173 ; P3_R1131_U279
g28167 nand P3_U3080 P3_R1131_U70 ; P3_R1131_U280
g28168 not P3_R1131_U170 ; P3_R1131_U281
g28169 nand P3_U3907 P3_R1131_U73 ; P3_R1131_U282
g28170 nand P3_R1131_U282 P3_R1131_U170 ; P3_R1131_U283
g28171 nand P3_U3075 P3_R1131_U72 ; P3_R1131_U284
g28172 not P3_R1131_U169 ; P3_R1131_U285
g28173 nand P3_U3904 P3_R1131_U77 ; P3_R1131_U286
g28174 nand P3_U3065 P3_R1131_U74 ; P3_R1131_U287
g28175 nand P3_U3060 P3_R1131_U75 ; P3_R1131_U288
g28176 nand P3_R1131_U197 P3_R1131_U11 ; P3_R1131_U289
g28177 nand P3_R1131_U12 P3_R1131_U289 ; P3_R1131_U290
g28178 nand P3_U3906 P3_R1131_U79 ; P3_R1131_U291
g28179 nand P3_U3904 P3_R1131_U77 ; P3_R1131_U292
g28180 nand P3_R1131_U129 P3_R1131_U169 ; P3_R1131_U293
g28181 nand P3_R1131_U292 P3_R1131_U290 ; P3_R1131_U294
g28182 not P3_R1131_U166 ; P3_R1131_U295
g28183 nand P3_U3903 P3_R1131_U82 ; P3_R1131_U296
g28184 nand P3_R1131_U296 P3_R1131_U166 ; P3_R1131_U297
g28185 nand P3_U3064 P3_R1131_U81 ; P3_R1131_U298
g28186 not P3_R1131_U165 ; P3_R1131_U299
g28187 nand P3_U3902 P3_R1131_U84 ; P3_R1131_U300
g28188 nand P3_R1131_U300 P3_R1131_U165 ; P3_R1131_U301
g28189 nand P3_U3057 P3_R1131_U83 ; P3_R1131_U302
g28190 not P3_R1131_U91 ; P3_R1131_U303
g28191 nand P3_R1131_U130 P3_R1131_U91 ; P3_R1131_U304
g28192 nand P3_R1131_U88 P3_R1131_U87 ; P3_R1131_U305
g28193 nand P3_R1131_U305 P3_R1131_U85 ; P3_R1131_U306
g28194 nand P3_U3052 P3_R1131_U186 ; P3_R1131_U307
g28195 not P3_R1131_U163 ; P3_R1131_U308
g28196 nand P3_U3899 P3_R1131_U90 ; P3_R1131_U309
g28197 nand P3_U3053 P3_R1131_U89 ; P3_R1131_U310
g28198 nand P3_R1131_U303 P3_R1131_U87 ; P3_R1131_U311
g28199 nand P3_R1131_U137 P3_R1131_U311 ; P3_R1131_U312
g28200 nand P3_R1131_U91 P3_R1131_U192 ; P3_R1131_U313
g28201 nand P3_R1131_U136 P3_R1131_U313 ; P3_R1131_U314
g28202 nand P3_R1131_U192 P3_R1131_U87 ; P3_R1131_U315
g28203 nand P3_R1131_U291 P3_R1131_U169 ; P3_R1131_U316
g28204 not P3_R1131_U92 ; P3_R1131_U317
g28205 nand P3_U3060 P3_R1131_U75 ; P3_R1131_U318
g28206 nand P3_R1131_U317 P3_R1131_U318 ; P3_R1131_U319
g28207 nand P3_R1131_U141 P3_R1131_U319 ; P3_R1131_U320
g28208 nand P3_R1131_U92 P3_R1131_U191 ; P3_R1131_U321
g28209 nand P3_U3904 P3_R1131_U77 ; P3_R1131_U322
g28210 nand P3_R1131_U140 P3_R1131_U321 ; P3_R1131_U323
g28211 nand P3_U3060 P3_R1131_U75 ; P3_R1131_U324
g28212 nand P3_R1131_U191 P3_R1131_U324 ; P3_R1131_U325
g28213 nand P3_R1131_U291 P3_R1131_U80 ; P3_R1131_U326
g28214 nand P3_R1131_U267 P3_R1131_U179 ; P3_R1131_U327
g28215 not P3_R1131_U93 ; P3_R1131_U328
g28216 nand P3_U3073 P3_R1131_U61 ; P3_R1131_U329
g28217 nand P3_R1131_U328 P3_R1131_U329 ; P3_R1131_U330
g28218 nand P3_R1131_U148 P3_R1131_U330 ; P3_R1131_U331
g28219 nand P3_R1131_U93 P3_R1131_U190 ; P3_R1131_U332
g28220 nand P3_U3437 P3_R1131_U63 ; P3_R1131_U333
g28221 nand P3_R1131_U147 P3_R1131_U332 ; P3_R1131_U334
g28222 nand P3_U3073 P3_R1131_U61 ; P3_R1131_U335
g28223 nand P3_R1131_U190 P3_R1131_U335 ; P3_R1131_U336
g28224 nand P3_R1131_U267 P3_R1131_U66 ; P3_R1131_U337
g28225 nand P3_R1131_U222 P3_R1131_U154 ; P3_R1131_U338
g28226 not P3_R1131_U94 ; P3_R1131_U339
g28227 nand P3_U3061 P3_R1131_U52 ; P3_R1131_U340
g28228 nand P3_R1131_U339 P3_R1131_U340 ; P3_R1131_U341
g28229 nand P3_R1131_U152 P3_R1131_U341 ; P3_R1131_U342
g28230 nand P3_R1131_U94 P3_R1131_U189 ; P3_R1131_U343
g28231 nand P3_U3422 P3_R1131_U53 ; P3_R1131_U344
g28232 nand P3_R1131_U151 P3_R1131_U343 ; P3_R1131_U345
g28233 nand P3_U3061 P3_R1131_U52 ; P3_R1131_U346
g28234 nand P3_R1131_U189 P3_R1131_U346 ; P3_R1131_U347
g28235 nand P3_U3076 P3_R1131_U30 ; P3_R1131_U348
g28236 nand P3_U3077 P3_R1131_U171 ; P3_R1131_U349
g28237 nand P3_U3081 P3_R1131_U174 ; P3_R1131_U350
g28238 nand P3_R1131_U133 P3_R1131_U304 P3_R1131_U134 ; P3_R1131_U351
g28239 nand P3_U3398 P3_R1131_U35 ; P3_R1131_U352
g28240 nand P3_U3413 P3_R1131_U220 ; P3_R1131_U353
g28241 nand P3_R1131_U353 P3_R1131_U219 ; P3_R1131_U354
g28242 nand P3_U3900 P3_R1131_U88 ; P3_R1131_U355
g28243 nand P3_R1131_U119 P3_R1131_U158 ; P3_R1131_U356
g28244 nand P3_R1131_U216 P3_R1131_U14 ; P3_R1131_U357
g28245 nand P3_U3416 P3_R1131_U46 ; P3_R1131_U358
g28246 nand P3_U3082 P3_R1131_U45 ; P3_R1131_U359
g28247 nand P3_R1131_U223 P3_R1131_U154 ; P3_R1131_U360
g28248 nand P3_R1131_U221 P3_R1131_U153 ; P3_R1131_U361
g28249 nand P3_U3413 P3_R1131_U27 ; P3_R1131_U362
g28250 nand P3_U3083 P3_R1131_U28 ; P3_R1131_U363
g28251 nand P3_U3413 P3_R1131_U27 ; P3_R1131_U364
g28252 nand P3_U3083 P3_R1131_U28 ; P3_R1131_U365
g28253 nand P3_R1131_U365 P3_R1131_U364 ; P3_R1131_U366
g28254 nand P3_U3410 P3_R1131_U25 ; P3_R1131_U367
g28255 nand P3_U3069 P3_R1131_U39 ; P3_R1131_U368
g28256 nand P3_R1131_U228 P3_R1131_U47 ; P3_R1131_U369
g28257 nand P3_R1131_U155 P3_R1131_U217 ; P3_R1131_U370
g28258 nand P3_U3407 P3_R1131_U40 ; P3_R1131_U371
g28259 nand P3_U3070 P3_R1131_U37 ; P3_R1131_U372
g28260 nand P3_R1131_U372 P3_R1131_U371 ; P3_R1131_U373
g28261 nand P3_U3404 P3_R1131_U41 ; P3_R1131_U374
g28262 nand P3_U3066 P3_R1131_U36 ; P3_R1131_U375
g28263 nand P3_R1131_U238 P3_R1131_U48 ; P3_R1131_U376
g28264 nand P3_R1131_U156 P3_R1131_U230 ; P3_R1131_U377
g28265 nand P3_U3401 P3_R1131_U42 ; P3_R1131_U378
g28266 nand P3_U3059 P3_R1131_U38 ; P3_R1131_U379
g28267 nand P3_R1131_U239 P3_R1131_U158 ; P3_R1131_U380
g28268 nand P3_R1131_U207 P3_R1131_U157 ; P3_R1131_U381
g28269 nand P3_U3398 P3_R1131_U35 ; P3_R1131_U382
g28270 nand P3_U3063 P3_R1131_U32 ; P3_R1131_U383
g28271 nand P3_U3398 P3_R1131_U35 ; P3_R1131_U384
g28272 nand P3_U3063 P3_R1131_U32 ; P3_R1131_U385
g28273 nand P3_R1131_U385 P3_R1131_U384 ; P3_R1131_U386
g28274 nand P3_U3395 P3_R1131_U33 ; P3_R1131_U387
g28275 nand P3_U3067 P3_R1131_U29 ; P3_R1131_U388
g28276 nand P3_R1131_U244 P3_R1131_U49 ; P3_R1131_U389
g28277 nand P3_R1131_U159 P3_R1131_U202 ; P3_R1131_U390
g28278 nand P3_U3908 P3_R1131_U161 ; P3_R1131_U391
g28279 nand P3_U3054 P3_R1131_U160 ; P3_R1131_U392
g28280 nand P3_U3908 P3_R1131_U161 ; P3_R1131_U393
g28281 nand P3_U3054 P3_R1131_U160 ; P3_R1131_U394
g28282 nand P3_R1131_U394 P3_R1131_U393 ; P3_R1131_U395
g28283 nand P3_U3053 P3_R1131_U395 P3_R1131_U89 ; P3_R1131_U396
g28284 nand P3_R1131_U15 P3_R1131_U90 P3_U3899 ; P3_R1131_U397
g28285 nand P3_U3899 P3_R1131_U90 ; P3_R1131_U398
g28286 nand P3_U3053 P3_R1131_U89 ; P3_R1131_U399
g28287 not P3_R1131_U135 ; P3_R1131_U400
g28288 nand P3_R1131_U308 P3_R1131_U400 ; P3_R1131_U401
g28289 nand P3_R1131_U135 P3_R1131_U163 ; P3_R1131_U402
g28290 nand P3_U3900 P3_R1131_U88 ; P3_R1131_U403
g28291 nand P3_U3052 P3_R1131_U85 ; P3_R1131_U404
g28292 nand P3_U3900 P3_R1131_U88 ; P3_R1131_U405
g28293 nand P3_U3052 P3_R1131_U85 ; P3_R1131_U406
g28294 nand P3_R1131_U406 P3_R1131_U405 ; P3_R1131_U407
g28295 nand P3_U3901 P3_R1131_U86 ; P3_R1131_U408
g28296 nand P3_U3056 P3_R1131_U50 ; P3_R1131_U409
g28297 nand P3_R1131_U315 P3_R1131_U91 ; P3_R1131_U410
g28298 nand P3_R1131_U164 P3_R1131_U303 ; P3_R1131_U411
g28299 nand P3_U3902 P3_R1131_U84 ; P3_R1131_U412
g28300 nand P3_U3057 P3_R1131_U83 ; P3_R1131_U413
g28301 not P3_R1131_U138 ; P3_R1131_U414
g28302 nand P3_R1131_U299 P3_R1131_U414 ; P3_R1131_U415
g28303 nand P3_R1131_U138 P3_R1131_U165 ; P3_R1131_U416
g28304 nand P3_U3903 P3_R1131_U82 ; P3_R1131_U417
g28305 nand P3_U3064 P3_R1131_U81 ; P3_R1131_U418
g28306 not P3_R1131_U139 ; P3_R1131_U419
g28307 nand P3_R1131_U295 P3_R1131_U419 ; P3_R1131_U420
g28308 nand P3_R1131_U139 P3_R1131_U166 ; P3_R1131_U421
g28309 nand P3_U3904 P3_R1131_U77 ; P3_R1131_U422
g28310 nand P3_U3065 P3_R1131_U74 ; P3_R1131_U423
g28311 nand P3_R1131_U423 P3_R1131_U422 ; P3_R1131_U424
g28312 nand P3_U3905 P3_R1131_U78 ; P3_R1131_U425
g28313 nand P3_U3060 P3_R1131_U75 ; P3_R1131_U426
g28314 nand P3_R1131_U325 P3_R1131_U92 ; P3_R1131_U427
g28315 nand P3_R1131_U167 P3_R1131_U317 ; P3_R1131_U428
g28316 nand P3_U3906 P3_R1131_U79 ; P3_R1131_U429
g28317 nand P3_U3074 P3_R1131_U76 ; P3_R1131_U430
g28318 nand P3_R1131_U326 P3_R1131_U169 ; P3_R1131_U431
g28319 nand P3_R1131_U285 P3_R1131_U168 ; P3_R1131_U432
g28320 nand P3_U3907 P3_R1131_U73 ; P3_R1131_U433
g28321 nand P3_U3075 P3_R1131_U72 ; P3_R1131_U434
g28322 not P3_R1131_U142 ; P3_R1131_U435
g28323 nand P3_R1131_U281 P3_R1131_U435 ; P3_R1131_U436
g28324 nand P3_R1131_U142 P3_R1131_U170 ; P3_R1131_U437
g28325 nand P3_U3392 P3_R1131_U31 ; P3_R1131_U438
g28326 nand P3_U3077 P3_R1131_U171 ; P3_R1131_U439
g28327 not P3_R1131_U143 ; P3_R1131_U440
g28328 nand P3_R1131_U200 P3_R1131_U440 ; P3_R1131_U441
g28329 nand P3_R1131_U143 P3_R1131_U172 ; P3_R1131_U442
g28330 nand P3_U3445 P3_R1131_U71 ; P3_R1131_U443
g28331 nand P3_U3080 P3_R1131_U70 ; P3_R1131_U444
g28332 not P3_R1131_U144 ; P3_R1131_U445
g28333 nand P3_R1131_U277 P3_R1131_U445 ; P3_R1131_U446
g28334 nand P3_R1131_U144 P3_R1131_U173 ; P3_R1131_U447
g28335 nand P3_U3443 P3_R1131_U69 ; P3_R1131_U448
g28336 nand P3_U3081 P3_R1131_U174 ; P3_R1131_U449
g28337 not P3_R1131_U145 ; P3_R1131_U450
g28338 nand P3_R1131_U275 P3_R1131_U450 ; P3_R1131_U451
g28339 nand P3_R1131_U145 P3_R1131_U175 ; P3_R1131_U452
g28340 nand P3_U3440 P3_R1131_U68 ; P3_R1131_U453
g28341 nand P3_U3068 P3_R1131_U67 ; P3_R1131_U454
g28342 not P3_R1131_U146 ; P3_R1131_U455
g28343 nand P3_R1131_U271 P3_R1131_U455 ; P3_R1131_U456
g28344 nand P3_R1131_U146 P3_R1131_U176 ; P3_R1131_U457
g28345 nand P3_U3437 P3_R1131_U63 ; P3_R1131_U458
g28346 nand P3_U3072 P3_R1131_U60 ; P3_R1131_U459
g28347 nand P3_R1131_U459 P3_R1131_U458 ; P3_R1131_U460
g28348 nand P3_U3434 P3_R1131_U64 ; P3_R1131_U461
g28349 nand P3_U3073 P3_R1131_U61 ; P3_R1131_U462
g28350 nand P3_R1131_U336 P3_R1131_U93 ; P3_R1131_U463
g28351 nand P3_R1131_U177 P3_R1131_U328 ; P3_R1131_U464
g28352 nand P3_U3431 P3_R1131_U65 ; P3_R1131_U465
g28353 nand P3_U3078 P3_R1131_U62 ; P3_R1131_U466
g28354 nand P3_R1131_U337 P3_R1131_U179 ; P3_R1131_U467
g28355 nand P3_R1131_U261 P3_R1131_U178 ; P3_R1131_U468
g28356 nand P3_U3428 P3_R1131_U59 ; P3_R1131_U469
g28357 nand P3_U3079 P3_R1131_U58 ; P3_R1131_U470
g28358 not P3_R1131_U149 ; P3_R1131_U471
g28359 nand P3_R1131_U257 P3_R1131_U471 ; P3_R1131_U472
g28360 nand P3_R1131_U149 P3_R1131_U180 ; P3_R1131_U473
g28361 nand P3_U3425 P3_R1131_U57 ; P3_R1131_U474
g28362 nand P3_U3071 P3_R1131_U56 ; P3_R1131_U475
g28363 not P3_R1131_U150 ; P3_R1131_U476
g28364 nand P3_R1131_U253 P3_R1131_U476 ; P3_R1131_U477
g28365 nand P3_R1131_U150 P3_R1131_U181 ; P3_R1131_U478
g28366 nand P3_U3422 P3_R1131_U53 ; P3_R1131_U479
g28367 nand P3_U3062 P3_R1131_U51 ; P3_R1131_U480
g28368 nand P3_R1131_U480 P3_R1131_U479 ; P3_R1131_U481
g28369 nand P3_U3419 P3_R1131_U54 ; P3_R1131_U482
g28370 nand P3_U3061 P3_R1131_U52 ; P3_R1131_U483
g28371 nand P3_R1131_U347 P3_R1131_U94 ; P3_R1131_U484
g28372 nand P3_R1131_U182 P3_R1131_U339 ; P3_R1131_U485
g28373 and P3_R1054_U102 P3_R1054_U118 ; P3_R1054_U6
g28374 and P3_R1054_U120 P3_R1054_U119 ; P3_R1054_U7
g28375 and P3_R1054_U99 P3_R1054_U157 ; P3_R1054_U8
g28376 and P3_R1054_U159 P3_R1054_U158 ; P3_R1054_U9
g28377 and P3_R1054_U100 P3_R1054_U174 ; P3_R1054_U10
g28378 and P3_R1054_U176 P3_R1054_U175 ; P3_R1054_U11
g28379 nand P3_R1054_U207 P3_R1054_U210 ; P3_R1054_U12
g28380 nand P3_R1054_U196 P3_R1054_U199 ; P3_R1054_U13
g28381 nand P3_R1054_U153 P3_R1054_U155 ; P3_R1054_U14
g28382 nand P3_R1054_U145 P3_R1054_U148 ; P3_R1054_U15
g28383 nand P3_R1054_U137 P3_R1054_U139 ; P3_R1054_U16
g28384 nand P3_R1054_U21 P3_R1054_U213 ; P3_R1054_U17
g28385 not P3_U3409 ; P3_R1054_U18
g28386 not P3_U3394 ; P3_R1054_U19
g28387 not P3_U3386 ; P3_R1054_U20
g28388 nand P3_U3386 P3_R1054_U65 ; P3_R1054_U21
g28389 not P3_U3573 ; P3_R1054_U22
g28390 not P3_U3397 ; P3_R1054_U23
g28391 not P3_U3562 ; P3_R1054_U24
g28392 nand P3_U3562 P3_R1054_U19 ; P3_R1054_U25
g28393 not P3_U3561 ; P3_R1054_U26
g28394 not P3_U3406 ; P3_R1054_U27
g28395 not P3_U3403 ; P3_R1054_U28
g28396 not P3_U3400 ; P3_R1054_U29
g28397 not P3_U3558 ; P3_R1054_U30
g28398 not P3_U3559 ; P3_R1054_U31
g28399 not P3_U3560 ; P3_R1054_U32
g28400 nand P3_U3560 P3_R1054_U29 ; P3_R1054_U33
g28401 not P3_U3412 ; P3_R1054_U34
g28402 not P3_U3557 ; P3_R1054_U35
g28403 nand P3_U3557 P3_R1054_U18 ; P3_R1054_U36
g28404 not P3_U3556 ; P3_R1054_U37
g28405 not P3_U3415 ; P3_R1054_U38
g28406 not P3_U3555 ; P3_R1054_U39
g28407 nand P3_R1054_U126 P3_R1054_U125 ; P3_R1054_U40
g28408 nand P3_R1054_U33 P3_R1054_U141 ; P3_R1054_U41
g28409 nand P3_R1054_U110 P3_R1054_U109 ; P3_R1054_U42
g28410 not P3_U3421 ; P3_R1054_U43
g28411 not P3_U3418 ; P3_R1054_U44
g28412 not P3_U3571 ; P3_R1054_U45
g28413 not P3_U3572 ; P3_R1054_U46
g28414 nand P3_U3555 P3_R1054_U38 ; P3_R1054_U47
g28415 not P3_U3424 ; P3_R1054_U48
g28416 not P3_U3570 ; P3_R1054_U49
g28417 not P3_U3427 ; P3_R1054_U50
g28418 not P3_U3569 ; P3_R1054_U51
g28419 not P3_U3436 ; P3_R1054_U52
g28420 not P3_U3433 ; P3_R1054_U53
g28421 not P3_U3430 ; P3_R1054_U54
g28422 not P3_U3566 ; P3_R1054_U55
g28423 not P3_U3567 ; P3_R1054_U56
g28424 not P3_U3568 ; P3_R1054_U57
g28425 nand P3_U3568 P3_R1054_U54 ; P3_R1054_U58
g28426 not P3_U3439 ; P3_R1054_U59
g28427 not P3_U3565 ; P3_R1054_U60
g28428 nand P3_R1054_U186 P3_R1054_U185 ; P3_R1054_U61
g28429 not P3_U3564 ; P3_R1054_U62
g28430 nand P3_R1054_U58 P3_R1054_U192 ; P3_R1054_U63
g28431 nand P3_R1054_U47 P3_R1054_U203 ; P3_R1054_U64
g28432 not P3_U3574 ; P3_R1054_U65
g28433 nand P3_R1054_U251 P3_R1054_U250 ; P3_R1054_U66
g28434 nand P3_R1054_U256 P3_R1054_U255 ; P3_R1054_U67
g28435 nand P3_R1054_U261 P3_R1054_U260 ; P3_R1054_U68
g28436 nand P3_R1054_U266 P3_R1054_U265 ; P3_R1054_U69
g28437 nand P3_R1054_U282 P3_R1054_U281 ; P3_R1054_U70
g28438 nand P3_R1054_U287 P3_R1054_U286 ; P3_R1054_U71
g28439 nand P3_R1054_U217 P3_R1054_U216 ; P3_R1054_U72
g28440 nand P3_R1054_U226 P3_R1054_U225 ; P3_R1054_U73
g28441 nand P3_R1054_U233 P3_R1054_U232 ; P3_R1054_U74
g28442 nand P3_R1054_U237 P3_R1054_U236 ; P3_R1054_U75
g28443 nand P3_R1054_U246 P3_R1054_U245 ; P3_R1054_U76
g28444 nand P3_R1054_U273 P3_R1054_U272 ; P3_R1054_U77
g28445 nand P3_R1054_U277 P3_R1054_U276 ; P3_R1054_U78
g28446 nand P3_R1054_U294 P3_R1054_U293 ; P3_R1054_U79
g28447 nand P3_R1054_U248 P3_R1054_U247 ; P3_R1054_U80
g28448 nand P3_R1054_U253 P3_R1054_U252 ; P3_R1054_U81
g28449 nand P3_R1054_U258 P3_R1054_U257 ; P3_R1054_U82
g28450 nand P3_R1054_U263 P3_R1054_U262 ; P3_R1054_U83
g28451 nand P3_R1054_U279 P3_R1054_U278 ; P3_R1054_U84
g28452 nand P3_R1054_U284 P3_R1054_U283 ; P3_R1054_U85
g28453 nand P3_R1054_U131 P3_R1054_U132 P3_R1054_U129 ; P3_R1054_U86
g28454 nand P3_R1054_U115 P3_R1054_U116 P3_R1054_U113 ; P3_R1054_U87
g28455 not P3_U3391 ; P3_R1054_U88
g28456 not P3_U3379 ; P3_R1054_U89
g28457 not P3_U3563 ; P3_R1054_U90
g28458 nand P3_R1054_U190 P3_R1054_U189 ; P3_R1054_U91
g28459 not P3_U3442 ; P3_R1054_U92
g28460 nand P3_R1054_U182 P3_R1054_U181 ; P3_R1054_U93
g28461 nand P3_R1054_U172 P3_R1054_U171 ; P3_R1054_U94
g28462 nand P3_R1054_U168 P3_R1054_U167 ; P3_R1054_U95
g28463 nand P3_R1054_U164 P3_R1054_U163 ; P3_R1054_U96
g28464 not P3_R1054_U25 ; P3_R1054_U97
g28465 not P3_R1054_U36 ; P3_R1054_U98
g28466 nand P3_U3418 P3_R1054_U46 ; P3_R1054_U99
g28467 nand P3_U3433 P3_R1054_U56 ; P3_R1054_U100
g28468 nand P3_U3394 P3_R1054_U24 ; P3_R1054_U101
g28469 nand P3_U3403 P3_R1054_U31 ; P3_R1054_U102
g28470 nand P3_U3409 P3_R1054_U35 ; P3_R1054_U103
g28471 not P3_R1054_U58 ; P3_R1054_U104
g28472 not P3_R1054_U33 ; P3_R1054_U105
g28473 not P3_R1054_U47 ; P3_R1054_U106
g28474 not P3_R1054_U21 ; P3_R1054_U107
g28475 nand P3_R1054_U107 P3_R1054_U22 ; P3_R1054_U108
g28476 nand P3_R1054_U108 P3_R1054_U88 ; P3_R1054_U109
g28477 nand P3_U3573 P3_R1054_U21 ; P3_R1054_U110
g28478 not P3_R1054_U42 ; P3_R1054_U111
g28479 nand P3_U3397 P3_R1054_U26 ; P3_R1054_U112
g28480 nand P3_R1054_U112 P3_R1054_U101 P3_R1054_U42 ; P3_R1054_U113
g28481 nand P3_R1054_U26 P3_R1054_U25 ; P3_R1054_U114
g28482 nand P3_R1054_U114 P3_R1054_U23 ; P3_R1054_U115
g28483 nand P3_U3561 P3_R1054_U97 ; P3_R1054_U116
g28484 not P3_R1054_U87 ; P3_R1054_U117
g28485 nand P3_U3406 P3_R1054_U30 ; P3_R1054_U118
g28486 nand P3_U3558 P3_R1054_U27 ; P3_R1054_U119
g28487 nand P3_U3559 P3_R1054_U28 ; P3_R1054_U120
g28488 nand P3_R1054_U105 P3_R1054_U6 ; P3_R1054_U121
g28489 nand P3_R1054_U7 P3_R1054_U121 ; P3_R1054_U122
g28490 nand P3_U3400 P3_R1054_U32 ; P3_R1054_U123
g28491 nand P3_U3406 P3_R1054_U30 ; P3_R1054_U124
g28492 nand P3_R1054_U123 P3_R1054_U6 P3_R1054_U87 ; P3_R1054_U125
g28493 nand P3_R1054_U124 P3_R1054_U122 ; P3_R1054_U126
g28494 not P3_R1054_U40 ; P3_R1054_U127
g28495 nand P3_U3412 P3_R1054_U37 ; P3_R1054_U128
g28496 nand P3_R1054_U128 P3_R1054_U103 P3_R1054_U40 ; P3_R1054_U129
g28497 nand P3_R1054_U37 P3_R1054_U36 ; P3_R1054_U130
g28498 nand P3_R1054_U130 P3_R1054_U34 ; P3_R1054_U131
g28499 nand P3_U3556 P3_R1054_U98 ; P3_R1054_U132
g28500 not P3_R1054_U86 ; P3_R1054_U133
g28501 nand P3_U3415 P3_R1054_U39 ; P3_R1054_U134
g28502 nand P3_R1054_U134 P3_R1054_U47 ; P3_R1054_U135
g28503 nand P3_R1054_U127 P3_R1054_U36 ; P3_R1054_U136
g28504 nand P3_R1054_U222 P3_R1054_U103 P3_R1054_U136 ; P3_R1054_U137
g28505 nand P3_R1054_U40 P3_R1054_U103 ; P3_R1054_U138
g28506 nand P3_R1054_U219 P3_R1054_U218 P3_R1054_U36 P3_R1054_U138 ; P3_R1054_U139
g28507 nand P3_R1054_U36 P3_R1054_U103 ; P3_R1054_U140
g28508 nand P3_R1054_U123 P3_R1054_U87 ; P3_R1054_U141
g28509 not P3_R1054_U41 ; P3_R1054_U142
g28510 nand P3_U3559 P3_R1054_U28 ; P3_R1054_U143
g28511 nand P3_R1054_U142 P3_R1054_U143 ; P3_R1054_U144
g28512 nand P3_R1054_U229 P3_R1054_U102 P3_R1054_U144 ; P3_R1054_U145
g28513 nand P3_R1054_U41 P3_R1054_U102 ; P3_R1054_U146
g28514 nand P3_U3406 P3_R1054_U30 ; P3_R1054_U147
g28515 nand P3_R1054_U147 P3_R1054_U7 P3_R1054_U146 ; P3_R1054_U148
g28516 nand P3_U3559 P3_R1054_U28 ; P3_R1054_U149
g28517 nand P3_R1054_U102 P3_R1054_U149 ; P3_R1054_U150
g28518 nand P3_R1054_U123 P3_R1054_U33 ; P3_R1054_U151
g28519 nand P3_R1054_U111 P3_R1054_U25 ; P3_R1054_U152
g28520 nand P3_R1054_U242 P3_R1054_U101 P3_R1054_U152 ; P3_R1054_U153
g28521 nand P3_R1054_U42 P3_R1054_U101 ; P3_R1054_U154
g28522 nand P3_R1054_U239 P3_R1054_U238 P3_R1054_U25 P3_R1054_U154 ; P3_R1054_U155
g28523 nand P3_R1054_U25 P3_R1054_U101 ; P3_R1054_U156
g28524 nand P3_U3421 P3_R1054_U45 ; P3_R1054_U157
g28525 nand P3_U3571 P3_R1054_U43 ; P3_R1054_U158
g28526 nand P3_U3572 P3_R1054_U44 ; P3_R1054_U159
g28527 nand P3_R1054_U106 P3_R1054_U8 ; P3_R1054_U160
g28528 nand P3_R1054_U9 P3_R1054_U160 ; P3_R1054_U161
g28529 nand P3_U3421 P3_R1054_U45 ; P3_R1054_U162
g28530 nand P3_R1054_U134 P3_R1054_U8 P3_R1054_U86 ; P3_R1054_U163
g28531 nand P3_R1054_U162 P3_R1054_U161 ; P3_R1054_U164
g28532 not P3_R1054_U96 ; P3_R1054_U165
g28533 nand P3_U3424 P3_R1054_U49 ; P3_R1054_U166
g28534 nand P3_R1054_U166 P3_R1054_U96 ; P3_R1054_U167
g28535 nand P3_U3570 P3_R1054_U48 ; P3_R1054_U168
g28536 not P3_R1054_U95 ; P3_R1054_U169
g28537 nand P3_U3427 P3_R1054_U51 ; P3_R1054_U170
g28538 nand P3_R1054_U170 P3_R1054_U95 ; P3_R1054_U171
g28539 nand P3_U3569 P3_R1054_U50 ; P3_R1054_U172
g28540 not P3_R1054_U94 ; P3_R1054_U173
g28541 nand P3_U3436 P3_R1054_U55 ; P3_R1054_U174
g28542 nand P3_U3566 P3_R1054_U52 ; P3_R1054_U175
g28543 nand P3_U3567 P3_R1054_U53 ; P3_R1054_U176
g28544 nand P3_R1054_U104 P3_R1054_U10 ; P3_R1054_U177
g28545 nand P3_R1054_U11 P3_R1054_U177 ; P3_R1054_U178
g28546 nand P3_U3430 P3_R1054_U57 ; P3_R1054_U179
g28547 nand P3_U3436 P3_R1054_U55 ; P3_R1054_U180
g28548 nand P3_R1054_U179 P3_R1054_U10 P3_R1054_U94 ; P3_R1054_U181
g28549 nand P3_R1054_U180 P3_R1054_U178 ; P3_R1054_U182
g28550 not P3_R1054_U93 ; P3_R1054_U183
g28551 nand P3_U3439 P3_R1054_U60 ; P3_R1054_U184
g28552 nand P3_R1054_U184 P3_R1054_U93 ; P3_R1054_U185
g28553 nand P3_U3565 P3_R1054_U59 ; P3_R1054_U186
g28554 not P3_R1054_U61 ; P3_R1054_U187
g28555 nand P3_R1054_U187 P3_R1054_U62 ; P3_R1054_U188
g28556 nand P3_R1054_U188 P3_R1054_U92 ; P3_R1054_U189
g28557 nand P3_U3564 P3_R1054_U61 ; P3_R1054_U190
g28558 not P3_R1054_U91 ; P3_R1054_U191
g28559 nand P3_R1054_U179 P3_R1054_U94 ; P3_R1054_U192
g28560 not P3_R1054_U63 ; P3_R1054_U193
g28561 nand P3_U3567 P3_R1054_U53 ; P3_R1054_U194
g28562 nand P3_R1054_U193 P3_R1054_U194 ; P3_R1054_U195
g28563 nand P3_R1054_U269 P3_R1054_U100 P3_R1054_U195 ; P3_R1054_U196
g28564 nand P3_R1054_U63 P3_R1054_U100 ; P3_R1054_U197
g28565 nand P3_U3436 P3_R1054_U55 ; P3_R1054_U198
g28566 nand P3_R1054_U198 P3_R1054_U11 P3_R1054_U197 ; P3_R1054_U199
g28567 nand P3_U3567 P3_R1054_U53 ; P3_R1054_U200
g28568 nand P3_R1054_U100 P3_R1054_U200 ; P3_R1054_U201
g28569 nand P3_R1054_U179 P3_R1054_U58 ; P3_R1054_U202
g28570 nand P3_R1054_U134 P3_R1054_U86 ; P3_R1054_U203
g28571 not P3_R1054_U64 ; P3_R1054_U204
g28572 nand P3_U3572 P3_R1054_U44 ; P3_R1054_U205
g28573 nand P3_R1054_U204 P3_R1054_U205 ; P3_R1054_U206
g28574 nand P3_R1054_U290 P3_R1054_U99 P3_R1054_U206 ; P3_R1054_U207
g28575 nand P3_R1054_U64 P3_R1054_U99 ; P3_R1054_U208
g28576 nand P3_U3421 P3_R1054_U45 ; P3_R1054_U209
g28577 nand P3_R1054_U209 P3_R1054_U9 P3_R1054_U208 ; P3_R1054_U210
g28578 nand P3_U3572 P3_R1054_U44 ; P3_R1054_U211
g28579 nand P3_R1054_U99 P3_R1054_U211 ; P3_R1054_U212
g28580 nand P3_U3574 P3_R1054_U20 ; P3_R1054_U213
g28581 nand P3_U3415 P3_R1054_U39 ; P3_R1054_U214
g28582 nand P3_U3555 P3_R1054_U38 ; P3_R1054_U215
g28583 nand P3_R1054_U135 P3_R1054_U86 ; P3_R1054_U216
g28584 nand P3_R1054_U215 P3_R1054_U214 P3_R1054_U133 ; P3_R1054_U217
g28585 nand P3_U3412 P3_R1054_U37 ; P3_R1054_U218
g28586 nand P3_U3556 P3_R1054_U34 ; P3_R1054_U219
g28587 nand P3_U3412 P3_R1054_U37 ; P3_R1054_U220
g28588 nand P3_U3556 P3_R1054_U34 ; P3_R1054_U221
g28589 nand P3_R1054_U221 P3_R1054_U220 ; P3_R1054_U222
g28590 nand P3_U3409 P3_R1054_U35 ; P3_R1054_U223
g28591 nand P3_U3557 P3_R1054_U18 ; P3_R1054_U224
g28592 nand P3_R1054_U140 P3_R1054_U40 ; P3_R1054_U225
g28593 nand P3_R1054_U224 P3_R1054_U223 P3_R1054_U127 ; P3_R1054_U226
g28594 nand P3_U3406 P3_R1054_U30 ; P3_R1054_U227
g28595 nand P3_U3558 P3_R1054_U27 ; P3_R1054_U228
g28596 nand P3_R1054_U228 P3_R1054_U227 ; P3_R1054_U229
g28597 nand P3_U3403 P3_R1054_U31 ; P3_R1054_U230
g28598 nand P3_U3559 P3_R1054_U28 ; P3_R1054_U231
g28599 nand P3_R1054_U150 P3_R1054_U41 ; P3_R1054_U232
g28600 nand P3_R1054_U231 P3_R1054_U230 P3_R1054_U142 ; P3_R1054_U233
g28601 nand P3_U3400 P3_R1054_U32 ; P3_R1054_U234
g28602 nand P3_U3560 P3_R1054_U29 ; P3_R1054_U235
g28603 nand P3_R1054_U151 P3_R1054_U87 ; P3_R1054_U236
g28604 nand P3_R1054_U235 P3_R1054_U234 P3_R1054_U117 ; P3_R1054_U237
g28605 nand P3_U3397 P3_R1054_U26 ; P3_R1054_U238
g28606 nand P3_U3561 P3_R1054_U23 ; P3_R1054_U239
g28607 nand P3_U3397 P3_R1054_U26 ; P3_R1054_U240
g28608 nand P3_U3561 P3_R1054_U23 ; P3_R1054_U241
g28609 nand P3_R1054_U241 P3_R1054_U240 ; P3_R1054_U242
g28610 nand P3_U3394 P3_R1054_U24 ; P3_R1054_U243
g28611 nand P3_U3562 P3_R1054_U19 ; P3_R1054_U244
g28612 nand P3_R1054_U156 P3_R1054_U42 ; P3_R1054_U245
g28613 nand P3_R1054_U244 P3_R1054_U243 P3_R1054_U111 ; P3_R1054_U246
g28614 nand P3_U3391 P3_R1054_U22 ; P3_R1054_U247
g28615 nand P3_U3573 P3_R1054_U88 ; P3_R1054_U248
g28616 not P3_R1054_U80 ; P3_R1054_U249
g28617 nand P3_R1054_U249 P3_R1054_U107 ; P3_R1054_U250
g28618 nand P3_R1054_U80 P3_R1054_U21 ; P3_R1054_U251
g28619 nand P3_U3379 P3_R1054_U90 ; P3_R1054_U252
g28620 nand P3_U3563 P3_R1054_U89 ; P3_R1054_U253
g28621 not P3_R1054_U81 ; P3_R1054_U254
g28622 nand P3_R1054_U191 P3_R1054_U254 ; P3_R1054_U255
g28623 nand P3_R1054_U81 P3_R1054_U91 ; P3_R1054_U256
g28624 nand P3_U3442 P3_R1054_U62 ; P3_R1054_U257
g28625 nand P3_U3564 P3_R1054_U92 ; P3_R1054_U258
g28626 not P3_R1054_U82 ; P3_R1054_U259
g28627 nand P3_R1054_U259 P3_R1054_U187 ; P3_R1054_U260
g28628 nand P3_R1054_U82 P3_R1054_U61 ; P3_R1054_U261
g28629 nand P3_U3439 P3_R1054_U60 ; P3_R1054_U262
g28630 nand P3_U3565 P3_R1054_U59 ; P3_R1054_U263
g28631 not P3_R1054_U83 ; P3_R1054_U264
g28632 nand P3_R1054_U183 P3_R1054_U264 ; P3_R1054_U265
g28633 nand P3_R1054_U83 P3_R1054_U93 ; P3_R1054_U266
g28634 nand P3_U3436 P3_R1054_U55 ; P3_R1054_U267
g28635 nand P3_U3566 P3_R1054_U52 ; P3_R1054_U268
g28636 nand P3_R1054_U268 P3_R1054_U267 ; P3_R1054_U269
g28637 nand P3_U3433 P3_R1054_U56 ; P3_R1054_U270
g28638 nand P3_U3567 P3_R1054_U53 ; P3_R1054_U271
g28639 nand P3_R1054_U201 P3_R1054_U63 ; P3_R1054_U272
g28640 nand P3_R1054_U271 P3_R1054_U270 P3_R1054_U193 ; P3_R1054_U273
g28641 nand P3_U3430 P3_R1054_U57 ; P3_R1054_U274
g28642 nand P3_U3568 P3_R1054_U54 ; P3_R1054_U275
g28643 nand P3_R1054_U202 P3_R1054_U94 ; P3_R1054_U276
g28644 nand P3_R1054_U275 P3_R1054_U274 P3_R1054_U173 ; P3_R1054_U277
g28645 nand P3_U3427 P3_R1054_U51 ; P3_R1054_U278
g28646 nand P3_U3569 P3_R1054_U50 ; P3_R1054_U279
g28647 not P3_R1054_U84 ; P3_R1054_U280
g28648 nand P3_R1054_U169 P3_R1054_U280 ; P3_R1054_U281
g28649 nand P3_R1054_U84 P3_R1054_U95 ; P3_R1054_U282
g28650 nand P3_U3424 P3_R1054_U49 ; P3_R1054_U283
g28651 nand P3_U3570 P3_R1054_U48 ; P3_R1054_U284
g28652 not P3_R1054_U85 ; P3_R1054_U285
g28653 nand P3_R1054_U165 P3_R1054_U285 ; P3_R1054_U286
g28654 nand P3_R1054_U85 P3_R1054_U96 ; P3_R1054_U287
g28655 nand P3_U3421 P3_R1054_U45 ; P3_R1054_U288
g28656 nand P3_U3571 P3_R1054_U43 ; P3_R1054_U289
g28657 nand P3_R1054_U289 P3_R1054_U288 ; P3_R1054_U290
g28658 nand P3_U3418 P3_R1054_U46 ; P3_R1054_U291
g28659 nand P3_U3572 P3_R1054_U44 ; P3_R1054_U292
g28660 nand P3_R1054_U212 P3_R1054_U64 ; P3_R1054_U293
g28661 nand P3_R1054_U292 P3_R1054_U291 P3_R1054_U204 ; P3_R1054_U294
g28662 and P3_R1161_U179 P3_R1161_U178 ; P3_R1161_U4
g28663 and P3_R1161_U197 P3_R1161_U196 ; P3_R1161_U5
g28664 and P3_R1161_U237 P3_R1161_U236 ; P3_R1161_U6
g28665 and P3_R1161_U246 P3_R1161_U245 ; P3_R1161_U7
g28666 and P3_R1161_U264 P3_R1161_U263 ; P3_R1161_U8
g28667 and P3_R1161_U272 P3_R1161_U271 ; P3_R1161_U9
g28668 and P3_R1161_U351 P3_R1161_U348 ; P3_R1161_U10
g28669 and P3_R1161_U344 P3_R1161_U341 ; P3_R1161_U11
g28670 and P3_R1161_U335 P3_R1161_U332 ; P3_R1161_U12
g28671 and P3_R1161_U326 P3_R1161_U323 ; P3_R1161_U13
g28672 and P3_R1161_U320 P3_R1161_U318 ; P3_R1161_U14
g28673 and P3_R1161_U313 P3_R1161_U310 ; P3_R1161_U15
g28674 and P3_R1161_U235 P3_R1161_U232 ; P3_R1161_U16
g28675 and P3_R1161_U227 P3_R1161_U224 ; P3_R1161_U17
g28676 and P3_R1161_U213 P3_R1161_U210 ; P3_R1161_U18
g28677 not P3_U3407 ; P3_R1161_U19
g28678 not P3_U3070 ; P3_R1161_U20
g28679 not P3_U3069 ; P3_R1161_U21
g28680 nand P3_U3070 P3_U3407 ; P3_R1161_U22
g28681 not P3_U3410 ; P3_R1161_U23
g28682 not P3_U3401 ; P3_R1161_U24
g28683 not P3_U3059 ; P3_R1161_U25
g28684 not P3_U3066 ; P3_R1161_U26
g28685 not P3_U3395 ; P3_R1161_U27
g28686 not P3_U3067 ; P3_R1161_U28
g28687 not P3_U3387 ; P3_R1161_U29
g28688 not P3_U3076 ; P3_R1161_U30
g28689 nand P3_U3076 P3_U3387 ; P3_R1161_U31
g28690 not P3_U3398 ; P3_R1161_U32
g28691 not P3_U3063 ; P3_R1161_U33
g28692 nand P3_U3059 P3_U3401 ; P3_R1161_U34
g28693 not P3_U3404 ; P3_R1161_U35
g28694 not P3_U3413 ; P3_R1161_U36
g28695 not P3_U3083 ; P3_R1161_U37
g28696 not P3_U3082 ; P3_R1161_U38
g28697 not P3_U3416 ; P3_R1161_U39
g28698 nand P3_R1161_U63 P3_R1161_U205 ; P3_R1161_U40
g28699 nand P3_R1161_U117 P3_R1161_U193 ; P3_R1161_U41
g28700 nand P3_R1161_U182 P3_R1161_U183 ; P3_R1161_U42
g28701 nand P3_U3392 P3_U3077 ; P3_R1161_U43
g28702 nand P3_R1161_U122 P3_R1161_U219 ; P3_R1161_U44
g28703 nand P3_R1161_U216 P3_R1161_U215 ; P3_R1161_U45
g28704 not P3_U3900 ; P3_R1161_U46
g28705 not P3_U3052 ; P3_R1161_U47
g28706 not P3_U3056 ; P3_R1161_U48
g28707 not P3_U3901 ; P3_R1161_U49
g28708 not P3_U3902 ; P3_R1161_U50
g28709 not P3_U3057 ; P3_R1161_U51
g28710 not P3_U3903 ; P3_R1161_U52
g28711 not P3_U3064 ; P3_R1161_U53
g28712 not P3_U3906 ; P3_R1161_U54
g28713 not P3_U3074 ; P3_R1161_U55
g28714 not P3_U3437 ; P3_R1161_U56
g28715 not P3_U3072 ; P3_R1161_U57
g28716 not P3_U3068 ; P3_R1161_U58
g28717 nand P3_U3072 P3_U3437 ; P3_R1161_U59
g28718 not P3_U3440 ; P3_R1161_U60
g28719 not P3_U3419 ; P3_R1161_U61
g28720 not P3_U3061 ; P3_R1161_U62
g28721 nand P3_U3083 P3_U3413 ; P3_R1161_U63
g28722 not P3_U3425 ; P3_R1161_U64
g28723 not P3_U3071 ; P3_R1161_U65
g28724 not P3_U3422 ; P3_R1161_U66
g28725 not P3_U3062 ; P3_R1161_U67
g28726 nand P3_U3062 P3_U3422 ; P3_R1161_U68
g28727 not P3_U3428 ; P3_R1161_U69
g28728 not P3_U3079 ; P3_R1161_U70
g28729 not P3_U3431 ; P3_R1161_U71
g28730 not P3_U3078 ; P3_R1161_U72
g28731 not P3_U3434 ; P3_R1161_U73
g28732 not P3_U3073 ; P3_R1161_U74
g28733 not P3_U3443 ; P3_R1161_U75
g28734 not P3_U3081 ; P3_R1161_U76
g28735 nand P3_U3081 P3_U3443 ; P3_R1161_U77
g28736 not P3_U3445 ; P3_R1161_U78
g28737 not P3_U3080 ; P3_R1161_U79
g28738 nand P3_U3080 P3_U3445 ; P3_R1161_U80
g28739 not P3_U3907 ; P3_R1161_U81
g28740 not P3_U3905 ; P3_R1161_U82
g28741 not P3_U3060 ; P3_R1161_U83
g28742 not P3_U3904 ; P3_R1161_U84
g28743 not P3_U3065 ; P3_R1161_U85
g28744 nand P3_U3901 P3_U3056 ; P3_R1161_U86
g28745 not P3_U3053 ; P3_R1161_U87
g28746 not P3_U3899 ; P3_R1161_U88
g28747 nand P3_R1161_U306 P3_R1161_U176 ; P3_R1161_U89
g28748 not P3_U3075 ; P3_R1161_U90
g28749 nand P3_R1161_U77 P3_R1161_U315 ; P3_R1161_U91
g28750 nand P3_R1161_U261 P3_R1161_U260 ; P3_R1161_U92
g28751 nand P3_R1161_U68 P3_R1161_U337 ; P3_R1161_U93
g28752 nand P3_R1161_U457 P3_R1161_U456 ; P3_R1161_U94
g28753 nand P3_R1161_U504 P3_R1161_U503 ; P3_R1161_U95
g28754 nand P3_R1161_U375 P3_R1161_U374 ; P3_R1161_U96
g28755 nand P3_R1161_U380 P3_R1161_U379 ; P3_R1161_U97
g28756 nand P3_R1161_U387 P3_R1161_U386 ; P3_R1161_U98
g28757 nand P3_R1161_U394 P3_R1161_U393 ; P3_R1161_U99
g28758 nand P3_R1161_U399 P3_R1161_U398 ; P3_R1161_U100
g28759 nand P3_R1161_U408 P3_R1161_U407 ; P3_R1161_U101
g28760 nand P3_R1161_U415 P3_R1161_U414 ; P3_R1161_U102
g28761 nand P3_R1161_U422 P3_R1161_U421 ; P3_R1161_U103
g28762 nand P3_R1161_U429 P3_R1161_U428 ; P3_R1161_U104
g28763 nand P3_R1161_U434 P3_R1161_U433 ; P3_R1161_U105
g28764 nand P3_R1161_U441 P3_R1161_U440 ; P3_R1161_U106
g28765 nand P3_R1161_U448 P3_R1161_U447 ; P3_R1161_U107
g28766 nand P3_R1161_U462 P3_R1161_U461 ; P3_R1161_U108
g28767 nand P3_R1161_U467 P3_R1161_U466 ; P3_R1161_U109
g28768 nand P3_R1161_U474 P3_R1161_U473 ; P3_R1161_U110
g28769 nand P3_R1161_U481 P3_R1161_U480 ; P3_R1161_U111
g28770 nand P3_R1161_U488 P3_R1161_U487 ; P3_R1161_U112
g28771 nand P3_R1161_U495 P3_R1161_U494 ; P3_R1161_U113
g28772 nand P3_R1161_U500 P3_R1161_U499 ; P3_R1161_U114
g28773 and P3_R1161_U189 P3_R1161_U187 ; P3_R1161_U115
g28774 and P3_R1161_U4 P3_R1161_U180 ; P3_R1161_U116
g28775 and P3_R1161_U194 P3_R1161_U192 ; P3_R1161_U117
g28776 and P3_R1161_U201 P3_R1161_U200 ; P3_R1161_U118
g28777 and P3_R1161_U382 P3_R1161_U381 P3_R1161_U22 ; P3_R1161_U119
g28778 and P3_R1161_U212 P3_R1161_U5 ; P3_R1161_U120
g28779 and P3_R1161_U181 P3_R1161_U180 ; P3_R1161_U121
g28780 and P3_R1161_U220 P3_R1161_U218 ; P3_R1161_U122
g28781 and P3_R1161_U389 P3_R1161_U388 P3_R1161_U34 ; P3_R1161_U123
g28782 and P3_R1161_U226 P3_R1161_U4 ; P3_R1161_U124
g28783 and P3_R1161_U234 P3_R1161_U181 ; P3_R1161_U125
g28784 and P3_R1161_U204 P3_R1161_U6 ; P3_R1161_U126
g28785 and P3_R1161_U243 P3_R1161_U239 ; P3_R1161_U127
g28786 and P3_R1161_U250 P3_R1161_U7 ; P3_R1161_U128
g28787 and P3_R1161_U248 P3_R1161_U172 ; P3_R1161_U129
g28788 and P3_R1161_U268 P3_R1161_U267 ; P3_R1161_U130
g28789 and P3_R1161_U9 P3_R1161_U282 P3_R1161_U273 ; P3_R1161_U131
g28790 and P3_R1161_U285 P3_R1161_U280 ; P3_R1161_U132
g28791 and P3_R1161_U301 P3_R1161_U298 ; P3_R1161_U133
g28792 and P3_R1161_U368 P3_R1161_U302 ; P3_R1161_U134
g28793 and P3_R1161_U160 P3_R1161_U278 ; P3_R1161_U135
g28794 and P3_R1161_U455 P3_R1161_U454 P3_R1161_U80 ; P3_R1161_U136
g28795 and P3_R1161_U325 P3_R1161_U9 ; P3_R1161_U137
g28796 and P3_R1161_U469 P3_R1161_U468 P3_R1161_U59 ; P3_R1161_U138
g28797 and P3_R1161_U334 P3_R1161_U8 ; P3_R1161_U139
g28798 and P3_R1161_U490 P3_R1161_U489 P3_R1161_U172 ; P3_R1161_U140
g28799 and P3_R1161_U343 P3_R1161_U7 ; P3_R1161_U141
g28800 and P3_R1161_U502 P3_R1161_U501 P3_R1161_U171 ; P3_R1161_U142
g28801 and P3_R1161_U350 P3_R1161_U6 ; P3_R1161_U143
g28802 nand P3_R1161_U118 P3_R1161_U202 ; P3_R1161_U144
g28803 nand P3_R1161_U217 P3_R1161_U229 ; P3_R1161_U145
g28804 not P3_U3054 ; P3_R1161_U146
g28805 not P3_U3908 ; P3_R1161_U147
g28806 and P3_R1161_U403 P3_R1161_U402 ; P3_R1161_U148
g28807 nand P3_R1161_U304 P3_R1161_U169 P3_R1161_U364 ; P3_R1161_U149
g28808 and P3_R1161_U410 P3_R1161_U409 ; P3_R1161_U150
g28809 nand P3_R1161_U370 P3_R1161_U369 P3_R1161_U134 ; P3_R1161_U151
g28810 and P3_R1161_U417 P3_R1161_U416 ; P3_R1161_U152
g28811 nand P3_R1161_U365 P3_R1161_U299 P3_R1161_U86 ; P3_R1161_U153
g28812 and P3_R1161_U424 P3_R1161_U423 ; P3_R1161_U154
g28813 nand P3_R1161_U293 P3_R1161_U292 ; P3_R1161_U155
g28814 and P3_R1161_U436 P3_R1161_U435 ; P3_R1161_U156
g28815 nand P3_R1161_U289 P3_R1161_U288 ; P3_R1161_U157
g28816 and P3_R1161_U443 P3_R1161_U442 ; P3_R1161_U158
g28817 nand P3_R1161_U132 P3_R1161_U284 ; P3_R1161_U159
g28818 and P3_R1161_U450 P3_R1161_U449 ; P3_R1161_U160
g28819 nand P3_R1161_U43 P3_R1161_U327 ; P3_R1161_U161
g28820 nand P3_R1161_U130 P3_R1161_U269 ; P3_R1161_U162
g28821 and P3_R1161_U476 P3_R1161_U475 ; P3_R1161_U163
g28822 nand P3_R1161_U257 P3_R1161_U256 ; P3_R1161_U164
g28823 and P3_R1161_U483 P3_R1161_U482 ; P3_R1161_U165
g28824 nand P3_R1161_U253 P3_R1161_U252 ; P3_R1161_U166
g28825 nand P3_R1161_U127 P3_R1161_U242 ; P3_R1161_U167
g28826 nand P3_R1161_U367 P3_R1161_U366 ; P3_R1161_U168
g28827 nand P3_U3053 P3_R1161_U151 ; P3_R1161_U169
g28828 not P3_R1161_U34 ; P3_R1161_U170
g28829 nand P3_U3416 P3_U3082 ; P3_R1161_U171
g28830 nand P3_U3071 P3_U3425 ; P3_R1161_U172
g28831 nand P3_U3057 P3_U3902 ; P3_R1161_U173
g28832 not P3_R1161_U68 ; P3_R1161_U174
g28833 not P3_R1161_U77 ; P3_R1161_U175
g28834 nand P3_U3064 P3_U3903 ; P3_R1161_U176
g28835 not P3_R1161_U63 ; P3_R1161_U177
g28836 or P3_U3066 P3_U3404 ; P3_R1161_U178
g28837 or P3_U3059 P3_U3401 ; P3_R1161_U179
g28838 or P3_U3398 P3_U3063 ; P3_R1161_U180
g28839 or P3_U3395 P3_U3067 ; P3_R1161_U181
g28840 not P3_R1161_U31 ; P3_R1161_U182
g28841 or P3_U3392 P3_U3077 ; P3_R1161_U183
g28842 not P3_R1161_U42 ; P3_R1161_U184
g28843 not P3_R1161_U43 ; P3_R1161_U185
g28844 nand P3_R1161_U42 P3_R1161_U43 ; P3_R1161_U186
g28845 nand P3_U3067 P3_U3395 ; P3_R1161_U187
g28846 nand P3_R1161_U186 P3_R1161_U181 ; P3_R1161_U188
g28847 nand P3_U3063 P3_U3398 ; P3_R1161_U189
g28848 nand P3_R1161_U115 P3_R1161_U188 ; P3_R1161_U190
g28849 nand P3_R1161_U35 P3_R1161_U34 ; P3_R1161_U191
g28850 nand P3_U3066 P3_R1161_U191 ; P3_R1161_U192
g28851 nand P3_R1161_U116 P3_R1161_U190 ; P3_R1161_U193
g28852 nand P3_U3404 P3_R1161_U170 ; P3_R1161_U194
g28853 not P3_R1161_U41 ; P3_R1161_U195
g28854 or P3_U3069 P3_U3410 ; P3_R1161_U196
g28855 or P3_U3070 P3_U3407 ; P3_R1161_U197
g28856 not P3_R1161_U22 ; P3_R1161_U198
g28857 nand P3_R1161_U23 P3_R1161_U22 ; P3_R1161_U199
g28858 nand P3_U3069 P3_R1161_U199 ; P3_R1161_U200
g28859 nand P3_U3410 P3_R1161_U198 ; P3_R1161_U201
g28860 nand P3_R1161_U5 P3_R1161_U41 ; P3_R1161_U202
g28861 not P3_R1161_U144 ; P3_R1161_U203
g28862 or P3_U3413 P3_U3083 ; P3_R1161_U204
g28863 nand P3_R1161_U204 P3_R1161_U144 ; P3_R1161_U205
g28864 not P3_R1161_U40 ; P3_R1161_U206
g28865 or P3_U3082 P3_U3416 ; P3_R1161_U207
g28866 or P3_U3407 P3_U3070 ; P3_R1161_U208
g28867 nand P3_R1161_U208 P3_R1161_U41 ; P3_R1161_U209
g28868 nand P3_R1161_U119 P3_R1161_U209 ; P3_R1161_U210
g28869 nand P3_R1161_U195 P3_R1161_U22 ; P3_R1161_U211
g28870 nand P3_U3410 P3_U3069 ; P3_R1161_U212
g28871 nand P3_R1161_U120 P3_R1161_U211 ; P3_R1161_U213
g28872 or P3_U3070 P3_U3407 ; P3_R1161_U214
g28873 nand P3_R1161_U185 P3_R1161_U181 ; P3_R1161_U215
g28874 nand P3_U3067 P3_U3395 ; P3_R1161_U216
g28875 not P3_R1161_U45 ; P3_R1161_U217
g28876 nand P3_R1161_U121 P3_R1161_U184 ; P3_R1161_U218
g28877 nand P3_R1161_U45 P3_R1161_U180 ; P3_R1161_U219
g28878 nand P3_U3063 P3_U3398 ; P3_R1161_U220
g28879 not P3_R1161_U44 ; P3_R1161_U221
g28880 or P3_U3401 P3_U3059 ; P3_R1161_U222
g28881 nand P3_R1161_U222 P3_R1161_U44 ; P3_R1161_U223
g28882 nand P3_R1161_U123 P3_R1161_U223 ; P3_R1161_U224
g28883 nand P3_R1161_U221 P3_R1161_U34 ; P3_R1161_U225
g28884 nand P3_U3404 P3_U3066 ; P3_R1161_U226
g28885 nand P3_R1161_U124 P3_R1161_U225 ; P3_R1161_U227
g28886 or P3_U3059 P3_U3401 ; P3_R1161_U228
g28887 nand P3_R1161_U184 P3_R1161_U181 ; P3_R1161_U229
g28888 not P3_R1161_U145 ; P3_R1161_U230
g28889 nand P3_U3063 P3_U3398 ; P3_R1161_U231
g28890 nand P3_R1161_U401 P3_R1161_U400 P3_R1161_U43 P3_R1161_U42 ; P3_R1161_U232
g28891 nand P3_R1161_U43 P3_R1161_U42 ; P3_R1161_U233
g28892 nand P3_U3067 P3_U3395 ; P3_R1161_U234
g28893 nand P3_R1161_U125 P3_R1161_U233 ; P3_R1161_U235
g28894 or P3_U3082 P3_U3416 ; P3_R1161_U236
g28895 or P3_U3061 P3_U3419 ; P3_R1161_U237
g28896 nand P3_R1161_U177 P3_R1161_U6 ; P3_R1161_U238
g28897 nand P3_U3061 P3_U3419 ; P3_R1161_U239
g28898 nand P3_R1161_U171 P3_R1161_U238 ; P3_R1161_U240
g28899 or P3_U3419 P3_U3061 ; P3_R1161_U241
g28900 nand P3_R1161_U126 P3_R1161_U144 ; P3_R1161_U242
g28901 nand P3_R1161_U241 P3_R1161_U240 ; P3_R1161_U243
g28902 not P3_R1161_U167 ; P3_R1161_U244
g28903 or P3_U3079 P3_U3428 ; P3_R1161_U245
g28904 or P3_U3071 P3_U3425 ; P3_R1161_U246
g28905 nand P3_R1161_U174 P3_R1161_U7 ; P3_R1161_U247
g28906 nand P3_U3079 P3_U3428 ; P3_R1161_U248
g28907 nand P3_R1161_U129 P3_R1161_U247 ; P3_R1161_U249
g28908 or P3_U3422 P3_U3062 ; P3_R1161_U250
g28909 or P3_U3428 P3_U3079 ; P3_R1161_U251
g28910 nand P3_R1161_U128 P3_R1161_U167 ; P3_R1161_U252
g28911 nand P3_R1161_U251 P3_R1161_U249 ; P3_R1161_U253
g28912 not P3_R1161_U166 ; P3_R1161_U254
g28913 or P3_U3431 P3_U3078 ; P3_R1161_U255
g28914 nand P3_R1161_U255 P3_R1161_U166 ; P3_R1161_U256
g28915 nand P3_U3078 P3_U3431 ; P3_R1161_U257
g28916 not P3_R1161_U164 ; P3_R1161_U258
g28917 or P3_U3434 P3_U3073 ; P3_R1161_U259
g28918 nand P3_R1161_U259 P3_R1161_U164 ; P3_R1161_U260
g28919 nand P3_U3073 P3_U3434 ; P3_R1161_U261
g28920 not P3_R1161_U92 ; P3_R1161_U262
g28921 or P3_U3068 P3_U3440 ; P3_R1161_U263
g28922 or P3_U3072 P3_U3437 ; P3_R1161_U264
g28923 not P3_R1161_U59 ; P3_R1161_U265
g28924 nand P3_R1161_U60 P3_R1161_U59 ; P3_R1161_U266
g28925 nand P3_U3068 P3_R1161_U266 ; P3_R1161_U267
g28926 nand P3_U3440 P3_R1161_U265 ; P3_R1161_U268
g28927 nand P3_R1161_U8 P3_R1161_U92 ; P3_R1161_U269
g28928 not P3_R1161_U162 ; P3_R1161_U270
g28929 or P3_U3075 P3_U3907 ; P3_R1161_U271
g28930 or P3_U3080 P3_U3445 ; P3_R1161_U272
g28931 or P3_U3074 P3_U3906 ; P3_R1161_U273
g28932 not P3_R1161_U80 ; P3_R1161_U274
g28933 nand P3_U3907 P3_R1161_U274 ; P3_R1161_U275
g28934 nand P3_R1161_U275 P3_R1161_U90 ; P3_R1161_U276
g28935 nand P3_R1161_U80 P3_R1161_U81 ; P3_R1161_U277
g28936 nand P3_R1161_U277 P3_R1161_U276 ; P3_R1161_U278
g28937 nand P3_R1161_U175 P3_R1161_U9 ; P3_R1161_U279
g28938 nand P3_U3074 P3_U3906 ; P3_R1161_U280
g28939 nand P3_R1161_U278 P3_R1161_U279 ; P3_R1161_U281
g28940 or P3_U3443 P3_U3081 ; P3_R1161_U282
g28941 or P3_U3906 P3_U3074 ; P3_R1161_U283
g28942 nand P3_R1161_U162 P3_R1161_U131 ; P3_R1161_U284
g28943 nand P3_R1161_U283 P3_R1161_U281 ; P3_R1161_U285
g28944 not P3_R1161_U159 ; P3_R1161_U286
g28945 or P3_U3905 P3_U3060 ; P3_R1161_U287
g28946 nand P3_R1161_U287 P3_R1161_U159 ; P3_R1161_U288
g28947 nand P3_U3060 P3_U3905 ; P3_R1161_U289
g28948 not P3_R1161_U157 ; P3_R1161_U290
g28949 or P3_U3904 P3_U3065 ; P3_R1161_U291
g28950 nand P3_R1161_U291 P3_R1161_U157 ; P3_R1161_U292
g28951 nand P3_U3065 P3_U3904 ; P3_R1161_U293
g28952 not P3_R1161_U155 ; P3_R1161_U294
g28953 or P3_U3057 P3_U3902 ; P3_R1161_U295
g28954 nand P3_R1161_U176 P3_R1161_U173 ; P3_R1161_U296
g28955 not P3_R1161_U86 ; P3_R1161_U297
g28956 or P3_U3903 P3_U3064 ; P3_R1161_U298
g28957 nand P3_R1161_U155 P3_R1161_U298 P3_R1161_U168 ; P3_R1161_U299
g28958 not P3_R1161_U153 ; P3_R1161_U300
g28959 or P3_U3900 P3_U3052 ; P3_R1161_U301
g28960 nand P3_U3052 P3_U3900 ; P3_R1161_U302
g28961 not P3_R1161_U151 ; P3_R1161_U303
g28962 nand P3_U3899 P3_R1161_U151 ; P3_R1161_U304
g28963 not P3_R1161_U149 ; P3_R1161_U305
g28964 nand P3_R1161_U298 P3_R1161_U155 ; P3_R1161_U306
g28965 not P3_R1161_U89 ; P3_R1161_U307
g28966 or P3_U3902 P3_U3057 ; P3_R1161_U308
g28967 nand P3_R1161_U308 P3_R1161_U89 ; P3_R1161_U309
g28968 nand P3_R1161_U309 P3_R1161_U173 P3_R1161_U154 ; P3_R1161_U310
g28969 nand P3_R1161_U307 P3_R1161_U173 ; P3_R1161_U311
g28970 nand P3_U3901 P3_U3056 ; P3_R1161_U312
g28971 nand P3_R1161_U311 P3_R1161_U312 P3_R1161_U168 ; P3_R1161_U313
g28972 or P3_U3057 P3_U3902 ; P3_R1161_U314
g28973 nand P3_R1161_U282 P3_R1161_U162 ; P3_R1161_U315
g28974 not P3_R1161_U91 ; P3_R1161_U316
g28975 nand P3_R1161_U9 P3_R1161_U91 ; P3_R1161_U317
g28976 nand P3_R1161_U135 P3_R1161_U317 ; P3_R1161_U318
g28977 nand P3_R1161_U317 P3_R1161_U278 ; P3_R1161_U319
g28978 nand P3_R1161_U453 P3_R1161_U319 ; P3_R1161_U320
g28979 or P3_U3445 P3_U3080 ; P3_R1161_U321
g28980 nand P3_R1161_U321 P3_R1161_U91 ; P3_R1161_U322
g28981 nand P3_R1161_U136 P3_R1161_U322 ; P3_R1161_U323
g28982 nand P3_R1161_U316 P3_R1161_U80 ; P3_R1161_U324
g28983 nand P3_U3075 P3_U3907 ; P3_R1161_U325
g28984 nand P3_R1161_U137 P3_R1161_U324 ; P3_R1161_U326
g28985 or P3_U3392 P3_U3077 ; P3_R1161_U327
g28986 not P3_R1161_U161 ; P3_R1161_U328
g28987 or P3_U3080 P3_U3445 ; P3_R1161_U329
g28988 or P3_U3437 P3_U3072 ; P3_R1161_U330
g28989 nand P3_R1161_U330 P3_R1161_U92 ; P3_R1161_U331
g28990 nand P3_R1161_U138 P3_R1161_U331 ; P3_R1161_U332
g28991 nand P3_R1161_U262 P3_R1161_U59 ; P3_R1161_U333
g28992 nand P3_U3440 P3_U3068 ; P3_R1161_U334
g28993 nand P3_R1161_U139 P3_R1161_U333 ; P3_R1161_U335
g28994 or P3_U3072 P3_U3437 ; P3_R1161_U336
g28995 nand P3_R1161_U250 P3_R1161_U167 ; P3_R1161_U337
g28996 not P3_R1161_U93 ; P3_R1161_U338
g28997 or P3_U3425 P3_U3071 ; P3_R1161_U339
g28998 nand P3_R1161_U339 P3_R1161_U93 ; P3_R1161_U340
g28999 nand P3_R1161_U140 P3_R1161_U340 ; P3_R1161_U341
g29000 nand P3_R1161_U338 P3_R1161_U172 ; P3_R1161_U342
g29001 nand P3_U3079 P3_U3428 ; P3_R1161_U343
g29002 nand P3_R1161_U141 P3_R1161_U342 ; P3_R1161_U344
g29003 or P3_U3071 P3_U3425 ; P3_R1161_U345
g29004 or P3_U3416 P3_U3082 ; P3_R1161_U346
g29005 nand P3_R1161_U346 P3_R1161_U40 ; P3_R1161_U347
g29006 nand P3_R1161_U142 P3_R1161_U347 ; P3_R1161_U348
g29007 nand P3_R1161_U206 P3_R1161_U171 ; P3_R1161_U349
g29008 nand P3_U3061 P3_U3419 ; P3_R1161_U350
g29009 nand P3_R1161_U143 P3_R1161_U349 ; P3_R1161_U351
g29010 nand P3_R1161_U207 P3_R1161_U171 ; P3_R1161_U352
g29011 nand P3_R1161_U204 P3_R1161_U63 ; P3_R1161_U353
g29012 nand P3_R1161_U214 P3_R1161_U22 ; P3_R1161_U354
g29013 nand P3_R1161_U228 P3_R1161_U34 ; P3_R1161_U355
g29014 nand P3_R1161_U231 P3_R1161_U180 ; P3_R1161_U356
g29015 nand P3_R1161_U314 P3_R1161_U173 ; P3_R1161_U357
g29016 nand P3_R1161_U298 P3_R1161_U176 ; P3_R1161_U358
g29017 nand P3_R1161_U329 P3_R1161_U80 ; P3_R1161_U359
g29018 nand P3_R1161_U282 P3_R1161_U77 ; P3_R1161_U360
g29019 nand P3_R1161_U336 P3_R1161_U59 ; P3_R1161_U361
g29020 nand P3_R1161_U345 P3_R1161_U172 ; P3_R1161_U362
g29021 nand P3_R1161_U250 P3_R1161_U68 ; P3_R1161_U363
g29022 nand P3_U3899 P3_U3053 ; P3_R1161_U364
g29023 nand P3_R1161_U296 P3_R1161_U168 ; P3_R1161_U365
g29024 nand P3_U3056 P3_R1161_U295 ; P3_R1161_U366
g29025 nand P3_U3901 P3_R1161_U295 ; P3_R1161_U367
g29026 nand P3_R1161_U296 P3_R1161_U168 P3_R1161_U301 ; P3_R1161_U368
g29027 nand P3_R1161_U155 P3_R1161_U168 P3_R1161_U133 ; P3_R1161_U369
g29028 nand P3_R1161_U297 P3_R1161_U301 ; P3_R1161_U370
g29029 nand P3_U3082 P3_R1161_U39 ; P3_R1161_U371
g29030 nand P3_U3416 P3_R1161_U38 ; P3_R1161_U372
g29031 nand P3_R1161_U372 P3_R1161_U371 ; P3_R1161_U373
g29032 nand P3_R1161_U352 P3_R1161_U40 ; P3_R1161_U374
g29033 nand P3_R1161_U373 P3_R1161_U206 ; P3_R1161_U375
g29034 nand P3_U3083 P3_R1161_U36 ; P3_R1161_U376
g29035 nand P3_U3413 P3_R1161_U37 ; P3_R1161_U377
g29036 nand P3_R1161_U377 P3_R1161_U376 ; P3_R1161_U378
g29037 nand P3_R1161_U353 P3_R1161_U144 ; P3_R1161_U379
g29038 nand P3_R1161_U203 P3_R1161_U378 ; P3_R1161_U380
g29039 nand P3_U3069 P3_R1161_U23 ; P3_R1161_U381
g29040 nand P3_U3410 P3_R1161_U21 ; P3_R1161_U382
g29041 nand P3_U3070 P3_R1161_U19 ; P3_R1161_U383
g29042 nand P3_U3407 P3_R1161_U20 ; P3_R1161_U384
g29043 nand P3_R1161_U384 P3_R1161_U383 ; P3_R1161_U385
g29044 nand P3_R1161_U354 P3_R1161_U41 ; P3_R1161_U386
g29045 nand P3_R1161_U385 P3_R1161_U195 ; P3_R1161_U387
g29046 nand P3_U3066 P3_R1161_U35 ; P3_R1161_U388
g29047 nand P3_U3404 P3_R1161_U26 ; P3_R1161_U389
g29048 nand P3_U3059 P3_R1161_U24 ; P3_R1161_U390
g29049 nand P3_U3401 P3_R1161_U25 ; P3_R1161_U391
g29050 nand P3_R1161_U391 P3_R1161_U390 ; P3_R1161_U392
g29051 nand P3_R1161_U355 P3_R1161_U44 ; P3_R1161_U393
g29052 nand P3_R1161_U392 P3_R1161_U221 ; P3_R1161_U394
g29053 nand P3_U3063 P3_R1161_U32 ; P3_R1161_U395
g29054 nand P3_U3398 P3_R1161_U33 ; P3_R1161_U396
g29055 nand P3_R1161_U396 P3_R1161_U395 ; P3_R1161_U397
g29056 nand P3_R1161_U356 P3_R1161_U145 ; P3_R1161_U398
g29057 nand P3_R1161_U230 P3_R1161_U397 ; P3_R1161_U399
g29058 nand P3_U3067 P3_R1161_U27 ; P3_R1161_U400
g29059 nand P3_U3395 P3_R1161_U28 ; P3_R1161_U401
g29060 nand P3_U3054 P3_R1161_U147 ; P3_R1161_U402
g29061 nand P3_U3908 P3_R1161_U146 ; P3_R1161_U403
g29062 nand P3_U3054 P3_R1161_U147 ; P3_R1161_U404
g29063 nand P3_U3908 P3_R1161_U146 ; P3_R1161_U405
g29064 nand P3_R1161_U405 P3_R1161_U404 ; P3_R1161_U406
g29065 nand P3_R1161_U148 P3_R1161_U149 ; P3_R1161_U407
g29066 nand P3_R1161_U305 P3_R1161_U406 ; P3_R1161_U408
g29067 nand P3_U3053 P3_R1161_U88 ; P3_R1161_U409
g29068 nand P3_U3899 P3_R1161_U87 ; P3_R1161_U410
g29069 nand P3_U3053 P3_R1161_U88 ; P3_R1161_U411
g29070 nand P3_U3899 P3_R1161_U87 ; P3_R1161_U412
g29071 nand P3_R1161_U412 P3_R1161_U411 ; P3_R1161_U413
g29072 nand P3_R1161_U150 P3_R1161_U151 ; P3_R1161_U414
g29073 nand P3_R1161_U303 P3_R1161_U413 ; P3_R1161_U415
g29074 nand P3_U3052 P3_R1161_U46 ; P3_R1161_U416
g29075 nand P3_U3900 P3_R1161_U47 ; P3_R1161_U417
g29076 nand P3_U3052 P3_R1161_U46 ; P3_R1161_U418
g29077 nand P3_U3900 P3_R1161_U47 ; P3_R1161_U419
g29078 nand P3_R1161_U419 P3_R1161_U418 ; P3_R1161_U420
g29079 nand P3_R1161_U152 P3_R1161_U153 ; P3_R1161_U421
g29080 nand P3_R1161_U300 P3_R1161_U420 ; P3_R1161_U422
g29081 nand P3_U3056 P3_R1161_U49 ; P3_R1161_U423
g29082 nand P3_U3901 P3_R1161_U48 ; P3_R1161_U424
g29083 nand P3_U3057 P3_R1161_U50 ; P3_R1161_U425
g29084 nand P3_U3902 P3_R1161_U51 ; P3_R1161_U426
g29085 nand P3_R1161_U426 P3_R1161_U425 ; P3_R1161_U427
g29086 nand P3_R1161_U357 P3_R1161_U89 ; P3_R1161_U428
g29087 nand P3_R1161_U427 P3_R1161_U307 ; P3_R1161_U429
g29088 nand P3_U3064 P3_R1161_U52 ; P3_R1161_U430
g29089 nand P3_U3903 P3_R1161_U53 ; P3_R1161_U431
g29090 nand P3_R1161_U431 P3_R1161_U430 ; P3_R1161_U432
g29091 nand P3_R1161_U358 P3_R1161_U155 ; P3_R1161_U433
g29092 nand P3_R1161_U294 P3_R1161_U432 ; P3_R1161_U434
g29093 nand P3_U3065 P3_R1161_U84 ; P3_R1161_U435
g29094 nand P3_U3904 P3_R1161_U85 ; P3_R1161_U436
g29095 nand P3_U3065 P3_R1161_U84 ; P3_R1161_U437
g29096 nand P3_U3904 P3_R1161_U85 ; P3_R1161_U438
g29097 nand P3_R1161_U438 P3_R1161_U437 ; P3_R1161_U439
g29098 nand P3_R1161_U156 P3_R1161_U157 ; P3_R1161_U440
g29099 nand P3_R1161_U290 P3_R1161_U439 ; P3_R1161_U441
g29100 nand P3_U3060 P3_R1161_U82 ; P3_R1161_U442
g29101 nand P3_U3905 P3_R1161_U83 ; P3_R1161_U443
g29102 nand P3_U3060 P3_R1161_U82 ; P3_R1161_U444
g29103 nand P3_U3905 P3_R1161_U83 ; P3_R1161_U445
g29104 nand P3_R1161_U445 P3_R1161_U444 ; P3_R1161_U446
g29105 nand P3_R1161_U158 P3_R1161_U159 ; P3_R1161_U447
g29106 nand P3_R1161_U286 P3_R1161_U446 ; P3_R1161_U448
g29107 nand P3_U3074 P3_R1161_U54 ; P3_R1161_U449
g29108 nand P3_U3906 P3_R1161_U55 ; P3_R1161_U450
g29109 nand P3_U3074 P3_R1161_U54 ; P3_R1161_U451
g29110 nand P3_U3906 P3_R1161_U55 ; P3_R1161_U452
g29111 nand P3_R1161_U452 P3_R1161_U451 ; P3_R1161_U453
g29112 nand P3_U3075 P3_R1161_U81 ; P3_R1161_U454
g29113 nand P3_U3907 P3_R1161_U90 ; P3_R1161_U455
g29114 nand P3_R1161_U182 P3_R1161_U161 ; P3_R1161_U456
g29115 nand P3_R1161_U328 P3_R1161_U31 ; P3_R1161_U457
g29116 nand P3_U3080 P3_R1161_U78 ; P3_R1161_U458
g29117 nand P3_U3445 P3_R1161_U79 ; P3_R1161_U459
g29118 nand P3_R1161_U459 P3_R1161_U458 ; P3_R1161_U460
g29119 nand P3_R1161_U359 P3_R1161_U91 ; P3_R1161_U461
g29120 nand P3_R1161_U460 P3_R1161_U316 ; P3_R1161_U462
g29121 nand P3_U3081 P3_R1161_U75 ; P3_R1161_U463
g29122 nand P3_U3443 P3_R1161_U76 ; P3_R1161_U464
g29123 nand P3_R1161_U464 P3_R1161_U463 ; P3_R1161_U465
g29124 nand P3_R1161_U360 P3_R1161_U162 ; P3_R1161_U466
g29125 nand P3_R1161_U270 P3_R1161_U465 ; P3_R1161_U467
g29126 nand P3_U3068 P3_R1161_U60 ; P3_R1161_U468
g29127 nand P3_U3440 P3_R1161_U58 ; P3_R1161_U469
g29128 nand P3_U3072 P3_R1161_U56 ; P3_R1161_U470
g29129 nand P3_U3437 P3_R1161_U57 ; P3_R1161_U471
g29130 nand P3_R1161_U471 P3_R1161_U470 ; P3_R1161_U472
g29131 nand P3_R1161_U361 P3_R1161_U92 ; P3_R1161_U473
g29132 nand P3_R1161_U472 P3_R1161_U262 ; P3_R1161_U474
g29133 nand P3_U3073 P3_R1161_U73 ; P3_R1161_U475
g29134 nand P3_U3434 P3_R1161_U74 ; P3_R1161_U476
g29135 nand P3_U3073 P3_R1161_U73 ; P3_R1161_U477
g29136 nand P3_U3434 P3_R1161_U74 ; P3_R1161_U478
g29137 nand P3_R1161_U478 P3_R1161_U477 ; P3_R1161_U479
g29138 nand P3_R1161_U163 P3_R1161_U164 ; P3_R1161_U480
g29139 nand P3_R1161_U258 P3_R1161_U479 ; P3_R1161_U481
g29140 nand P3_U3078 P3_R1161_U71 ; P3_R1161_U482
g29141 nand P3_U3431 P3_R1161_U72 ; P3_R1161_U483
g29142 nand P3_U3078 P3_R1161_U71 ; P3_R1161_U484
g29143 nand P3_U3431 P3_R1161_U72 ; P3_R1161_U485
g29144 nand P3_R1161_U485 P3_R1161_U484 ; P3_R1161_U486
g29145 nand P3_R1161_U165 P3_R1161_U166 ; P3_R1161_U487
g29146 nand P3_R1161_U254 P3_R1161_U486 ; P3_R1161_U488
g29147 nand P3_U3079 P3_R1161_U69 ; P3_R1161_U489
g29148 nand P3_U3428 P3_R1161_U70 ; P3_R1161_U490
g29149 nand P3_U3071 P3_R1161_U64 ; P3_R1161_U491
g29150 nand P3_U3425 P3_R1161_U65 ; P3_R1161_U492
g29151 nand P3_R1161_U492 P3_R1161_U491 ; P3_R1161_U493
g29152 nand P3_R1161_U362 P3_R1161_U93 ; P3_R1161_U494
g29153 nand P3_R1161_U493 P3_R1161_U338 ; P3_R1161_U495
g29154 nand P3_U3062 P3_R1161_U66 ; P3_R1161_U496
g29155 nand P3_U3422 P3_R1161_U67 ; P3_R1161_U497
g29156 nand P3_R1161_U497 P3_R1161_U496 ; P3_R1161_U498
g29157 nand P3_R1161_U363 P3_R1161_U167 ; P3_R1161_U499
g29158 nand P3_R1161_U244 P3_R1161_U498 ; P3_R1161_U500
g29159 nand P3_U3061 P3_R1161_U61 ; P3_R1161_U501
g29160 nand P3_U3419 P3_R1161_U62 ; P3_R1161_U502
g29161 nand P3_U3076 P3_R1161_U29 ; P3_R1161_U503
g29162 nand P3_U3387 P3_R1161_U30 ; P3_R1161_U504
