i DATAI_31_
i DATAI_30_
i DATAI_29_
i DATAI_28_
i DATAI_27_
i DATAI_26_
i DATAI_25_
i DATAI_24_
i DATAI_23_
i DATAI_22_
i DATAI_21_
i DATAI_20_
i DATAI_19_
i DATAI_18_
i DATAI_17_
i DATAI_16_
i DATAI_15_
i DATAI_14_
i DATAI_13_
i DATAI_12_
i DATAI_11_
i DATAI_10_
i DATAI_9_
i DATAI_8_
i DATAI_7_
i DATAI_6_
i DATAI_5_
i DATAI_4_
i DATAI_3_
i DATAI_2_
i DATAI_1_
i DATAI_0_
i MEMORYFETCH_REG_SCAN_IN
i NA_N
i BS16_N
i READY_N
i HOLD
i READREQUEST_REG_SCAN_IN
i ADS_N_REG_SCAN_IN
i CODEFETCH_REG_SCAN_IN
i M_IO_N_REG_SCAN_IN
i D_C_N_REG_SCAN_IN
i REQUESTPENDING_REG_SCAN_IN
i STATEBS16_REG_SCAN_IN
i MORE_REG_SCAN_IN
i FLUSH_REG_SCAN_IN
i W_R_N_REG_SCAN_IN
i BYTEENABLE_REG_0__SCAN_IN
i BYTEENABLE_REG_1__SCAN_IN
i BYTEENABLE_REG_2__SCAN_IN
i BYTEENABLE_REG_3__SCAN_IN
i REIP_REG_31__SCAN_IN
i REIP_REG_30__SCAN_IN
i REIP_REG_29__SCAN_IN
i REIP_REG_28__SCAN_IN
i REIP_REG_27__SCAN_IN
i REIP_REG_26__SCAN_IN
i REIP_REG_25__SCAN_IN
i REIP_REG_24__SCAN_IN
i REIP_REG_23__SCAN_IN
i REIP_REG_22__SCAN_IN
i REIP_REG_21__SCAN_IN
i REIP_REG_20__SCAN_IN
i REIP_REG_19__SCAN_IN
i REIP_REG_18__SCAN_IN
i REIP_REG_17__SCAN_IN
i REIP_REG_16__SCAN_IN
i BE_N_REG_3__SCAN_IN
i BE_N_REG_2__SCAN_IN
i BE_N_REG_1__SCAN_IN
i BE_N_REG_0__SCAN_IN
i ADDRESS_REG_29__SCAN_IN
i ADDRESS_REG_28__SCAN_IN
i ADDRESS_REG_27__SCAN_IN
i ADDRESS_REG_26__SCAN_IN
i ADDRESS_REG_25__SCAN_IN
i ADDRESS_REG_24__SCAN_IN
i ADDRESS_REG_23__SCAN_IN
i ADDRESS_REG_22__SCAN_IN
i ADDRESS_REG_21__SCAN_IN
i ADDRESS_REG_20__SCAN_IN
i ADDRESS_REG_19__SCAN_IN
i ADDRESS_REG_18__SCAN_IN
i ADDRESS_REG_17__SCAN_IN
i ADDRESS_REG_16__SCAN_IN
i ADDRESS_REG_15__SCAN_IN
i ADDRESS_REG_14__SCAN_IN
i ADDRESS_REG_13__SCAN_IN
i ADDRESS_REG_12__SCAN_IN
i ADDRESS_REG_11__SCAN_IN
i ADDRESS_REG_10__SCAN_IN
i ADDRESS_REG_9__SCAN_IN
i ADDRESS_REG_8__SCAN_IN
i ADDRESS_REG_7__SCAN_IN
i ADDRESS_REG_6__SCAN_IN
i ADDRESS_REG_5__SCAN_IN
i ADDRESS_REG_4__SCAN_IN
i ADDRESS_REG_3__SCAN_IN
i ADDRESS_REG_2__SCAN_IN
i ADDRESS_REG_1__SCAN_IN
i ADDRESS_REG_0__SCAN_IN
i STATE_REG_2__SCAN_IN
i STATE_REG_1__SCAN_IN
i STATE_REG_0__SCAN_IN
i DATAWIDTH_REG_0__SCAN_IN
i DATAWIDTH_REG_1__SCAN_IN
i DATAWIDTH_REG_2__SCAN_IN
i DATAWIDTH_REG_3__SCAN_IN
i DATAWIDTH_REG_4__SCAN_IN
i DATAWIDTH_REG_5__SCAN_IN
i DATAWIDTH_REG_6__SCAN_IN
i DATAWIDTH_REG_7__SCAN_IN
i DATAWIDTH_REG_8__SCAN_IN
i DATAWIDTH_REG_9__SCAN_IN
i DATAWIDTH_REG_10__SCAN_IN
i DATAWIDTH_REG_11__SCAN_IN
i DATAWIDTH_REG_12__SCAN_IN
i DATAWIDTH_REG_13__SCAN_IN
i DATAWIDTH_REG_14__SCAN_IN
i DATAWIDTH_REG_15__SCAN_IN
i DATAWIDTH_REG_16__SCAN_IN
i DATAWIDTH_REG_17__SCAN_IN
i DATAWIDTH_REG_18__SCAN_IN
i DATAWIDTH_REG_19__SCAN_IN
i DATAWIDTH_REG_20__SCAN_IN
i DATAWIDTH_REG_21__SCAN_IN
i DATAWIDTH_REG_22__SCAN_IN
i DATAWIDTH_REG_23__SCAN_IN
i DATAWIDTH_REG_24__SCAN_IN
i DATAWIDTH_REG_25__SCAN_IN
i DATAWIDTH_REG_26__SCAN_IN
i DATAWIDTH_REG_27__SCAN_IN
i DATAWIDTH_REG_28__SCAN_IN
i DATAWIDTH_REG_29__SCAN_IN
i DATAWIDTH_REG_30__SCAN_IN
i DATAWIDTH_REG_31__SCAN_IN
i STATE2_REG_3__SCAN_IN
i STATE2_REG_2__SCAN_IN
i STATE2_REG_1__SCAN_IN
i STATE2_REG_0__SCAN_IN
i INSTQUEUE_REG_15__7__SCAN_IN
i INSTQUEUE_REG_15__6__SCAN_IN
i INSTQUEUE_REG_15__5__SCAN_IN
i INSTQUEUE_REG_15__4__SCAN_IN
i INSTQUEUE_REG_15__3__SCAN_IN
i INSTQUEUE_REG_15__2__SCAN_IN
i INSTQUEUE_REG_15__1__SCAN_IN
i INSTQUEUE_REG_15__0__SCAN_IN
i INSTQUEUE_REG_14__7__SCAN_IN
i INSTQUEUE_REG_14__6__SCAN_IN
i INSTQUEUE_REG_14__5__SCAN_IN
i INSTQUEUE_REG_14__4__SCAN_IN
i INSTQUEUE_REG_14__3__SCAN_IN
i INSTQUEUE_REG_14__2__SCAN_IN
i INSTQUEUE_REG_14__1__SCAN_IN
i INSTQUEUE_REG_14__0__SCAN_IN
i INSTQUEUE_REG_13__7__SCAN_IN
i INSTQUEUE_REG_13__6__SCAN_IN
i INSTQUEUE_REG_13__5__SCAN_IN
i INSTQUEUE_REG_13__4__SCAN_IN
i INSTQUEUE_REG_13__3__SCAN_IN
i INSTQUEUE_REG_13__2__SCAN_IN
i INSTQUEUE_REG_13__1__SCAN_IN
i INSTQUEUE_REG_13__0__SCAN_IN
i INSTQUEUE_REG_12__7__SCAN_IN
i INSTQUEUE_REG_12__6__SCAN_IN
i INSTQUEUE_REG_12__5__SCAN_IN
i INSTQUEUE_REG_12__4__SCAN_IN
i INSTQUEUE_REG_12__3__SCAN_IN
i INSTQUEUE_REG_12__2__SCAN_IN
i INSTQUEUE_REG_12__1__SCAN_IN
i INSTQUEUE_REG_12__0__SCAN_IN
i INSTQUEUE_REG_11__7__SCAN_IN
i INSTQUEUE_REG_11__6__SCAN_IN
i INSTQUEUE_REG_11__5__SCAN_IN
i INSTQUEUE_REG_11__4__SCAN_IN
i INSTQUEUE_REG_11__3__SCAN_IN
i INSTQUEUE_REG_11__2__SCAN_IN
i INSTQUEUE_REG_11__1__SCAN_IN
i INSTQUEUE_REG_11__0__SCAN_IN
i INSTQUEUE_REG_10__7__SCAN_IN
i INSTQUEUE_REG_10__6__SCAN_IN
i INSTQUEUE_REG_10__5__SCAN_IN
i INSTQUEUE_REG_10__4__SCAN_IN
i INSTQUEUE_REG_10__3__SCAN_IN
i INSTQUEUE_REG_10__2__SCAN_IN
i INSTQUEUE_REG_10__1__SCAN_IN
i INSTQUEUE_REG_10__0__SCAN_IN
i INSTQUEUE_REG_9__7__SCAN_IN
i INSTQUEUE_REG_9__6__SCAN_IN
i INSTQUEUE_REG_9__5__SCAN_IN
i INSTQUEUE_REG_9__4__SCAN_IN
i INSTQUEUE_REG_9__3__SCAN_IN
i INSTQUEUE_REG_9__2__SCAN_IN
i INSTQUEUE_REG_9__1__SCAN_IN
i INSTQUEUE_REG_9__0__SCAN_IN
i INSTQUEUE_REG_8__7__SCAN_IN
i INSTQUEUE_REG_8__6__SCAN_IN
i INSTQUEUE_REG_8__5__SCAN_IN
i INSTQUEUE_REG_8__4__SCAN_IN
i INSTQUEUE_REG_8__3__SCAN_IN
i INSTQUEUE_REG_8__2__SCAN_IN
i INSTQUEUE_REG_8__1__SCAN_IN
i INSTQUEUE_REG_8__0__SCAN_IN
i INSTQUEUE_REG_7__7__SCAN_IN
i INSTQUEUE_REG_7__6__SCAN_IN
i INSTQUEUE_REG_7__5__SCAN_IN
i INSTQUEUE_REG_7__4__SCAN_IN
i INSTQUEUE_REG_7__3__SCAN_IN
i INSTQUEUE_REG_7__2__SCAN_IN
i INSTQUEUE_REG_7__1__SCAN_IN
i INSTQUEUE_REG_7__0__SCAN_IN
i INSTQUEUE_REG_6__7__SCAN_IN
i INSTQUEUE_REG_6__6__SCAN_IN
i INSTQUEUE_REG_6__5__SCAN_IN
i INSTQUEUE_REG_6__4__SCAN_IN
i INSTQUEUE_REG_6__3__SCAN_IN
i INSTQUEUE_REG_6__2__SCAN_IN
i INSTQUEUE_REG_6__1__SCAN_IN
i INSTQUEUE_REG_6__0__SCAN_IN
i INSTQUEUE_REG_5__7__SCAN_IN
i INSTQUEUE_REG_5__6__SCAN_IN
i INSTQUEUE_REG_5__5__SCAN_IN
i INSTQUEUE_REG_5__4__SCAN_IN
i INSTQUEUE_REG_5__3__SCAN_IN
i INSTQUEUE_REG_5__2__SCAN_IN
i INSTQUEUE_REG_5__1__SCAN_IN
i INSTQUEUE_REG_5__0__SCAN_IN
i INSTQUEUE_REG_4__7__SCAN_IN
i INSTQUEUE_REG_4__6__SCAN_IN
i INSTQUEUE_REG_4__5__SCAN_IN
i INSTQUEUE_REG_4__4__SCAN_IN
i INSTQUEUE_REG_4__3__SCAN_IN
i INSTQUEUE_REG_4__2__SCAN_IN
i INSTQUEUE_REG_4__1__SCAN_IN
i INSTQUEUE_REG_4__0__SCAN_IN
i INSTQUEUE_REG_3__7__SCAN_IN
i INSTQUEUE_REG_3__6__SCAN_IN
i INSTQUEUE_REG_3__5__SCAN_IN
i INSTQUEUE_REG_3__4__SCAN_IN
i INSTQUEUE_REG_3__3__SCAN_IN
i INSTQUEUE_REG_3__2__SCAN_IN
i INSTQUEUE_REG_3__1__SCAN_IN
i INSTQUEUE_REG_3__0__SCAN_IN
i INSTQUEUE_REG_2__7__SCAN_IN
i INSTQUEUE_REG_2__6__SCAN_IN
i INSTQUEUE_REG_2__5__SCAN_IN
i INSTQUEUE_REG_2__4__SCAN_IN
i INSTQUEUE_REG_2__3__SCAN_IN
i INSTQUEUE_REG_2__2__SCAN_IN
i INSTQUEUE_REG_2__1__SCAN_IN
i INSTQUEUE_REG_2__0__SCAN_IN
i INSTQUEUE_REG_1__7__SCAN_IN
i INSTQUEUE_REG_1__6__SCAN_IN
i INSTQUEUE_REG_1__5__SCAN_IN
i INSTQUEUE_REG_1__4__SCAN_IN
i INSTQUEUE_REG_1__3__SCAN_IN
i INSTQUEUE_REG_1__2__SCAN_IN
i INSTQUEUE_REG_1__1__SCAN_IN
i INSTQUEUE_REG_1__0__SCAN_IN
i INSTQUEUE_REG_0__7__SCAN_IN
i INSTQUEUE_REG_0__6__SCAN_IN
i INSTQUEUE_REG_0__5__SCAN_IN
i INSTQUEUE_REG_0__4__SCAN_IN
i INSTQUEUE_REG_0__3__SCAN_IN
i INSTQUEUE_REG_0__2__SCAN_IN
i INSTQUEUE_REG_0__1__SCAN_IN
i INSTQUEUE_REG_0__0__SCAN_IN
i INSTQUEUERD_ADDR_REG_4__SCAN_IN
i INSTQUEUERD_ADDR_REG_3__SCAN_IN
i INSTQUEUERD_ADDR_REG_2__SCAN_IN
i INSTQUEUERD_ADDR_REG_1__SCAN_IN
i INSTQUEUERD_ADDR_REG_0__SCAN_IN
i INSTQUEUEWR_ADDR_REG_4__SCAN_IN
i INSTQUEUEWR_ADDR_REG_3__SCAN_IN
i INSTQUEUEWR_ADDR_REG_2__SCAN_IN
i INSTQUEUEWR_ADDR_REG_1__SCAN_IN
i INSTQUEUEWR_ADDR_REG_0__SCAN_IN
i INSTADDRPOINTER_REG_0__SCAN_IN
i INSTADDRPOINTER_REG_1__SCAN_IN
i INSTADDRPOINTER_REG_2__SCAN_IN
i INSTADDRPOINTER_REG_3__SCAN_IN
i INSTADDRPOINTER_REG_4__SCAN_IN
i INSTADDRPOINTER_REG_5__SCAN_IN
i INSTADDRPOINTER_REG_6__SCAN_IN
i INSTADDRPOINTER_REG_7__SCAN_IN
i INSTADDRPOINTER_REG_8__SCAN_IN
i INSTADDRPOINTER_REG_9__SCAN_IN
i INSTADDRPOINTER_REG_10__SCAN_IN
i INSTADDRPOINTER_REG_11__SCAN_IN
i INSTADDRPOINTER_REG_12__SCAN_IN
i INSTADDRPOINTER_REG_13__SCAN_IN
i INSTADDRPOINTER_REG_14__SCAN_IN
i INSTADDRPOINTER_REG_15__SCAN_IN
i INSTADDRPOINTER_REG_16__SCAN_IN
i INSTADDRPOINTER_REG_17__SCAN_IN
i INSTADDRPOINTER_REG_18__SCAN_IN
i INSTADDRPOINTER_REG_19__SCAN_IN
i INSTADDRPOINTER_REG_20__SCAN_IN
i INSTADDRPOINTER_REG_21__SCAN_IN
i INSTADDRPOINTER_REG_22__SCAN_IN
i INSTADDRPOINTER_REG_23__SCAN_IN
i INSTADDRPOINTER_REG_24__SCAN_IN
i INSTADDRPOINTER_REG_25__SCAN_IN
i INSTADDRPOINTER_REG_26__SCAN_IN
i INSTADDRPOINTER_REG_27__SCAN_IN
i INSTADDRPOINTER_REG_28__SCAN_IN
i INSTADDRPOINTER_REG_29__SCAN_IN
i INSTADDRPOINTER_REG_30__SCAN_IN
i INSTADDRPOINTER_REG_31__SCAN_IN
i PHYADDRPOINTER_REG_0__SCAN_IN
i PHYADDRPOINTER_REG_1__SCAN_IN
i PHYADDRPOINTER_REG_2__SCAN_IN
i PHYADDRPOINTER_REG_3__SCAN_IN
i PHYADDRPOINTER_REG_4__SCAN_IN
i PHYADDRPOINTER_REG_5__SCAN_IN
i PHYADDRPOINTER_REG_6__SCAN_IN
i PHYADDRPOINTER_REG_7__SCAN_IN
i PHYADDRPOINTER_REG_8__SCAN_IN
i PHYADDRPOINTER_REG_9__SCAN_IN
i PHYADDRPOINTER_REG_10__SCAN_IN
i PHYADDRPOINTER_REG_11__SCAN_IN
i PHYADDRPOINTER_REG_12__SCAN_IN
i PHYADDRPOINTER_REG_13__SCAN_IN
i PHYADDRPOINTER_REG_14__SCAN_IN
i PHYADDRPOINTER_REG_15__SCAN_IN
i PHYADDRPOINTER_REG_16__SCAN_IN
i PHYADDRPOINTER_REG_17__SCAN_IN
i PHYADDRPOINTER_REG_18__SCAN_IN
i PHYADDRPOINTER_REG_19__SCAN_IN
i PHYADDRPOINTER_REG_20__SCAN_IN
i PHYADDRPOINTER_REG_21__SCAN_IN
i PHYADDRPOINTER_REG_22__SCAN_IN
i PHYADDRPOINTER_REG_23__SCAN_IN
i PHYADDRPOINTER_REG_24__SCAN_IN
i PHYADDRPOINTER_REG_25__SCAN_IN
i PHYADDRPOINTER_REG_26__SCAN_IN
i PHYADDRPOINTER_REG_27__SCAN_IN
i PHYADDRPOINTER_REG_28__SCAN_IN
i PHYADDRPOINTER_REG_29__SCAN_IN
i PHYADDRPOINTER_REG_30__SCAN_IN
i PHYADDRPOINTER_REG_31__SCAN_IN
i LWORD_REG_15__SCAN_IN
i LWORD_REG_14__SCAN_IN
i LWORD_REG_13__SCAN_IN
i LWORD_REG_12__SCAN_IN
i LWORD_REG_11__SCAN_IN
i LWORD_REG_10__SCAN_IN
i LWORD_REG_9__SCAN_IN
i LWORD_REG_8__SCAN_IN
i LWORD_REG_7__SCAN_IN
i LWORD_REG_6__SCAN_IN
i LWORD_REG_5__SCAN_IN
i LWORD_REG_4__SCAN_IN
i LWORD_REG_3__SCAN_IN
i LWORD_REG_2__SCAN_IN
i LWORD_REG_1__SCAN_IN
i LWORD_REG_0__SCAN_IN
i UWORD_REG_14__SCAN_IN
i UWORD_REG_13__SCAN_IN
i UWORD_REG_12__SCAN_IN
i UWORD_REG_11__SCAN_IN
i UWORD_REG_10__SCAN_IN
i UWORD_REG_9__SCAN_IN
i UWORD_REG_8__SCAN_IN
i UWORD_REG_7__SCAN_IN
i UWORD_REG_6__SCAN_IN
i UWORD_REG_5__SCAN_IN
i UWORD_REG_4__SCAN_IN
i UWORD_REG_3__SCAN_IN
i UWORD_REG_2__SCAN_IN
i UWORD_REG_1__SCAN_IN
i UWORD_REG_0__SCAN_IN
i DATAO_REG_0__SCAN_IN
i DATAO_REG_1__SCAN_IN
i DATAO_REG_2__SCAN_IN
i DATAO_REG_3__SCAN_IN
i DATAO_REG_4__SCAN_IN
i DATAO_REG_5__SCAN_IN
i DATAO_REG_6__SCAN_IN
i DATAO_REG_7__SCAN_IN
i DATAO_REG_8__SCAN_IN
i DATAO_REG_9__SCAN_IN
i DATAO_REG_10__SCAN_IN
i DATAO_REG_11__SCAN_IN
i DATAO_REG_12__SCAN_IN
i DATAO_REG_13__SCAN_IN
i DATAO_REG_14__SCAN_IN
i DATAO_REG_15__SCAN_IN
i DATAO_REG_16__SCAN_IN
i DATAO_REG_17__SCAN_IN
i DATAO_REG_18__SCAN_IN
i DATAO_REG_19__SCAN_IN
i DATAO_REG_20__SCAN_IN
i DATAO_REG_21__SCAN_IN
i DATAO_REG_22__SCAN_IN
i DATAO_REG_23__SCAN_IN
i DATAO_REG_24__SCAN_IN
i DATAO_REG_25__SCAN_IN
i DATAO_REG_26__SCAN_IN
i DATAO_REG_27__SCAN_IN
i DATAO_REG_28__SCAN_IN
i DATAO_REG_29__SCAN_IN
i DATAO_REG_30__SCAN_IN
i DATAO_REG_31__SCAN_IN
i EAX_REG_0__SCAN_IN
i EAX_REG_1__SCAN_IN
i EAX_REG_2__SCAN_IN
i EAX_REG_3__SCAN_IN
i EAX_REG_4__SCAN_IN
i EAX_REG_5__SCAN_IN
i EAX_REG_6__SCAN_IN
i EAX_REG_7__SCAN_IN
i EAX_REG_8__SCAN_IN
i EAX_REG_9__SCAN_IN
i EAX_REG_10__SCAN_IN
i EAX_REG_11__SCAN_IN
i EAX_REG_12__SCAN_IN
i EAX_REG_13__SCAN_IN
i EAX_REG_14__SCAN_IN
i EAX_REG_15__SCAN_IN
i EAX_REG_16__SCAN_IN
i EAX_REG_17__SCAN_IN
i EAX_REG_18__SCAN_IN
i EAX_REG_19__SCAN_IN
i EAX_REG_20__SCAN_IN
i EAX_REG_21__SCAN_IN
i EAX_REG_22__SCAN_IN
i EAX_REG_23__SCAN_IN
i EAX_REG_24__SCAN_IN
i EAX_REG_25__SCAN_IN
i EAX_REG_26__SCAN_IN
i EAX_REG_27__SCAN_IN
i EAX_REG_28__SCAN_IN
i EAX_REG_29__SCAN_IN
i EAX_REG_30__SCAN_IN
i EAX_REG_31__SCAN_IN
i EBX_REG_0__SCAN_IN
i EBX_REG_1__SCAN_IN
i EBX_REG_2__SCAN_IN
i EBX_REG_3__SCAN_IN
i EBX_REG_4__SCAN_IN
i EBX_REG_5__SCAN_IN
i EBX_REG_6__SCAN_IN
i EBX_REG_7__SCAN_IN
i EBX_REG_8__SCAN_IN
i EBX_REG_9__SCAN_IN
i EBX_REG_10__SCAN_IN
i EBX_REG_11__SCAN_IN
i EBX_REG_12__SCAN_IN
i EBX_REG_13__SCAN_IN
i EBX_REG_14__SCAN_IN
i EBX_REG_15__SCAN_IN
i EBX_REG_16__SCAN_IN
i EBX_REG_17__SCAN_IN
i EBX_REG_18__SCAN_IN
i EBX_REG_19__SCAN_IN
i EBX_REG_20__SCAN_IN
i EBX_REG_21__SCAN_IN
i EBX_REG_22__SCAN_IN
i EBX_REG_23__SCAN_IN
i EBX_REG_24__SCAN_IN
i EBX_REG_25__SCAN_IN
i EBX_REG_26__SCAN_IN
i EBX_REG_27__SCAN_IN
i EBX_REG_28__SCAN_IN
i EBX_REG_29__SCAN_IN
i EBX_REG_30__SCAN_IN
i EBX_REG_31__SCAN_IN
i REIP_REG_0__SCAN_IN
i REIP_REG_1__SCAN_IN
i REIP_REG_2__SCAN_IN
i REIP_REG_3__SCAN_IN
i REIP_REG_4__SCAN_IN
i REIP_REG_5__SCAN_IN
i REIP_REG_6__SCAN_IN
i REIP_REG_7__SCAN_IN
i REIP_REG_8__SCAN_IN
i REIP_REG_9__SCAN_IN
i REIP_REG_10__SCAN_IN
i REIP_REG_11__SCAN_IN
i REIP_REG_12__SCAN_IN
i REIP_REG_13__SCAN_IN
i REIP_REG_14__SCAN_IN
i REIP_REG_15__SCAN_IN
o BE_N_REG_3__SCAN_IN
o BE_N_REG_2__SCAN_IN
o BE_N_REG_1__SCAN_IN
o BE_N_REG_0__SCAN_IN
o ADDRESS_REG_29__SCAN_IN
o ADDRESS_REG_28__SCAN_IN
o ADDRESS_REG_27__SCAN_IN
o ADDRESS_REG_26__SCAN_IN
o ADDRESS_REG_25__SCAN_IN
o ADDRESS_REG_24__SCAN_IN
o ADDRESS_REG_23__SCAN_IN
o ADDRESS_REG_22__SCAN_IN
o ADDRESS_REG_21__SCAN_IN
o ADDRESS_REG_20__SCAN_IN
o ADDRESS_REG_19__SCAN_IN
o ADDRESS_REG_18__SCAN_IN
o ADDRESS_REG_17__SCAN_IN
o ADDRESS_REG_16__SCAN_IN
o ADDRESS_REG_15__SCAN_IN
o ADDRESS_REG_14__SCAN_IN
o ADDRESS_REG_13__SCAN_IN
o ADDRESS_REG_12__SCAN_IN
o ADDRESS_REG_11__SCAN_IN
o ADDRESS_REG_10__SCAN_IN
o ADDRESS_REG_9__SCAN_IN
o ADDRESS_REG_8__SCAN_IN
o ADDRESS_REG_7__SCAN_IN
o ADDRESS_REG_6__SCAN_IN
o ADDRESS_REG_5__SCAN_IN
o ADDRESS_REG_4__SCAN_IN
o ADDRESS_REG_3__SCAN_IN
o ADDRESS_REG_2__SCAN_IN
o ADDRESS_REG_1__SCAN_IN
o ADDRESS_REG_0__SCAN_IN
o W_R_N_REG_SCAN_IN
o D_C_N_REG_SCAN_IN
o M_IO_N_REG_SCAN_IN
o ADS_N_REG_SCAN_IN
o DATAO_REG_31__SCAN_IN
o DATAO_REG_30__SCAN_IN
o DATAO_REG_29__SCAN_IN
o DATAO_REG_28__SCAN_IN
o DATAO_REG_27__SCAN_IN
o DATAO_REG_26__SCAN_IN
o DATAO_REG_25__SCAN_IN
o DATAO_REG_24__SCAN_IN
o DATAO_REG_23__SCAN_IN
o DATAO_REG_22__SCAN_IN
o DATAO_REG_21__SCAN_IN
o DATAO_REG_20__SCAN_IN
o DATAO_REG_19__SCAN_IN
o DATAO_REG_18__SCAN_IN
o DATAO_REG_17__SCAN_IN
o DATAO_REG_16__SCAN_IN
o DATAO_REG_15__SCAN_IN
o DATAO_REG_14__SCAN_IN
o DATAO_REG_13__SCAN_IN
o DATAO_REG_12__SCAN_IN
o DATAO_REG_11__SCAN_IN
o DATAO_REG_10__SCAN_IN
o DATAO_REG_9__SCAN_IN
o DATAO_REG_8__SCAN_IN
o DATAO_REG_7__SCAN_IN
o DATAO_REG_6__SCAN_IN
o DATAO_REG_5__SCAN_IN
o DATAO_REG_4__SCAN_IN
o DATAO_REG_3__SCAN_IN
o DATAO_REG_2__SCAN_IN
o DATAO_REG_1__SCAN_IN
o DATAO_REG_0__SCAN_IN
o U3445
o U3446
o U3447
o U3448
o U3213
o U3212
o U3211
o U3210
o U3209
o U3208
o U3207
o U3206
o U3205
o U3204
o U3203
o U3202
o U3201
o U3200
o U3199
o U3198
o U3197
o U3196
o U3195
o U3194
o U3193
o U3192
o U3191
o U3190
o U3189
o U3188
o U3187
o U3186
o U3185
o U3184
o U3183
o U3182
o U3181
o U3451
o U3452
o U3180
o U3179
o U3178
o U3177
o U3176
o U3175
o U3174
o U3173
o U3172
o U3171
o U3170
o U3169
o U3168
o U3167
o U3166
o U3165
o U3164
o U3163
o U3162
o U3161
o U3160
o U3159
o U3158
o U3157
o U3156
o U3155
o U3154
o U3153
o U3152
o U3151
o U3453
o U3150
o U3149
o U3148
o U3147
o U3146
o U3145
o U3144
o U3143
o U3142
o U3141
o U3140
o U3139
o U3138
o U3137
o U3136
o U3135
o U3134
o U3133
o U3132
o U3131
o U3130
o U3129
o U3128
o U3127
o U3126
o U3125
o U3124
o U3123
o U3122
o U3121
o U3120
o U3119
o U3118
o U3117
o U3116
o U3115
o U3114
o U3113
o U3112
o U3111
o U3110
o U3109
o U3108
o U3107
o U3106
o U3105
o U3104
o U3103
o U3102
o U3101
o U3100
o U3099
o U3098
o U3097
o U3096
o U3095
o U3094
o U3093
o U3092
o U3091
o U3090
o U3089
o U3088
o U3087
o U3086
o U3085
o U3084
o U3083
o U3082
o U3081
o U3080
o U3079
o U3078
o U3077
o U3076
o U3075
o U3074
o U3073
o U3072
o U3071
o U3070
o U3069
o U3068
o U3067
o U3066
o U3065
o U3064
o U3063
o U3062
o U3061
o U3060
o U3059
o U3058
o U3057
o U3056
o U3055
o U3054
o U3053
o U3052
o U3051
o U3050
o U3049
o U3048
o U3047
o U3046
o U3045
o U3044
o U3043
o U3042
o U3041
o U3040
o U3039
o U3038
o U3037
o U3036
o U3035
o U3034
o U3033
o U3032
o U3031
o U3030
o U3029
o U3028
o U3027
o U3026
o U3025
o U3024
o U3023
o U3022
o U3021
o U3020
o U3455
o U3456
o U3459
o U3460
o U3461
o U3019
o U3462
o U3463
o U3464
o U3465
o U3018
o U3017
o U3016
o U3015
o U3014
o U3013
o U3012
o U3011
o U3010
o U3009
o U3008
o U3007
o U3006
o U3005
o U3004
o U3003
o U3002
o U3001
o U3000
o U2999
o U2998
o U2997
o U2996
o U2995
o U2994
o U2993
o U2992
o U2991
o U2990
o U2989
o U2988
o U2987
o U2986
o U2985
o U2984
o U2983
o U2982
o U2981
o U2980
o U2979
o U2978
o U2977
o U2976
o U2975
o U2974
o U2973
o U2972
o U2971
o U2970
o U2969
o U2968
o U2967
o U2966
o U2965
o U2964
o U2963
o U2962
o U2961
o U2960
o U2959
o U2958
o U2957
o U2956
o U2955
o U2954
o U2953
o U2952
o U2951
o U2950
o U2949
o U2948
o U2947
o U2946
o U2945
o U2944
o U2943
o U2942
o U2941
o U2940
o U2939
o U2938
o U2937
o U2936
o U2935
o U2934
o U2933
o U2932
o U2931
o U2930
o U2929
o U2928
o U2927
o U2926
o U2925
o U2924
o U2923
o U2922
o U2921
o U2920
o U2919
o U2918
o U2917
o U2916
o U2915
o U2914
o U2913
o U2912
o U2911
o U2910
o U2909
o U2908
o U2907
o U2906
o U2905
o U2904
o U2903
o U2902
o U2901
o U2900
o U2899
o U2898
o U2897
o U2896
o U2895
o U2894
o U2893
o U2892
o U2891
o U2890
o U2889
o U2888
o U2887
o U2886
o U2885
o U2884
o U2883
o U2882
o U2881
o U2880
o U2879
o U2878
o U2877
o U2876
o U2875
o U2874
o U2873
o U2872
o U2871
o U2870
o U2869
o U2868
o U2867
o U2866
o U2865
o U2864
o U2863
o U2862
o U2861
o U2860
o U2859
o U2858
o U2857
o U2856
o U2855
o U2854
o U2853
o U2852
o U2851
o U2850
o U2849
o U2848
o U2847
o U2846
o U2845
o U2844
o U2843
o U2842
o U2841
o U2840
o U2839
o U2838
o U2837
o U2836
o U2835
o U2834
o U2833
o U2832
o U2831
o U2830
o U2829
o U2828
o U2827
o U2826
o U2825
o U2824
o U2823
o U2822
o U2821
o U2820
o U2819
o U2818
o U2817
o U2816
o U2815
o U2814
o U2813
o U2812
o U2811
o U2810
o U2809
o U2808
o U2807
o U2806
o U2805
o U2804
o U2803
o U2802
o U2801
o U2800
o U2799
o U2798
o U2797
o U2796
o U2795
o U3468
o U2794
o U3469
o U3470
o U2793
o U3471
o U2792
o U3472
o U2791
o U3473
o U2790
o U2789
o U3474
o U2788
g1 nor STATE2_REG_2__SCAN_IN STATEBS16_REG_SCAN_IN ; U2352
g2 and U4219 STATE2_REG_2__SCAN_IN ; U2353
g3 and U4253 U4465 ; U2354
g4 and U3221 U2450 ; U2355
g5 and R2238_U6 U4180 ; U2356
g6 and U5947 U3853 R2167_U17 ; U2357
g7 and U2388 U4212 ; U2358
g8 and U3418 STATE2_REG_2__SCAN_IN ; U2359
g9 and U3401 STATE2_REG_2__SCAN_IN ; U2360
g10 and U4212 STATE2_REG_3__SCAN_IN ; U2361
g11 and U2359 U4196 ; U2362
g12 and U2359 U4198 ; U2363
g13 and U3852 U3403 ; U2364
g14 and U4249 U3403 ; U2365
g15 and U3418 U3417 STATE2_REG_1__SCAN_IN ; U2366
g16 and U3418 R2337_U58 STATE2_REG_1__SCAN_IN ; U2367
g17 and U4223 STATE2_REG_0__SCAN_IN ; U2368
g18 and U2362 U4485 ; U2369
g19 and U3401 U3250 ; U2370
g20 and U4210 U4437 ; U2371
g21 and U3403 STATE2_REG_0__SCAN_IN ; U2372
g22 and U3418 STATE2_REG_3__SCAN_IN ; U2373
g23 and U2360 U4202 ; U2374
g24 and U2360 U4204 ; U2375
g25 and U5786 U3403 ; U2376
g26 and U3750 U3401 ; U2377
g27 and U2360 U5557 ; U2378
g28 and U2363 U3267 ; U2379
g29 and U2360 U7596 ; U2380
g30 and U2357 U3258 ; U2381
g31 and U2357 U4465 ; U2382
g32 and U4210 U3378 ; U2383
g33 and U3404 STATE2_REG_0__SCAN_IN ; U2384
g34 and U3404 U3281 ; U2385
g35 and U4211 U3410 ; U2386
g36 and U3872 U4211 ; U2387
g37 and U4197 STATEBS16_REG_SCAN_IN ; U2388
g38 and U2452 U7482 ; U2389
g39 and DATAI_0_ U4212 ; U2390
g40 and DATAI_1_ U4212 ; U2391
g41 and DATAI_2_ U4212 ; U2392
g42 and DATAI_3_ U4212 ; U2393
g43 and DATAI_4_ U4212 ; U2394
g44 and DATAI_5_ U4212 ; U2395
g45 and DATAI_6_ U4212 ; U2396
g46 and DATAI_7_ U4212 ; U2397
g47 and DATAI_24_ U2358 ; U2398
g48 and DATAI_16_ U2358 ; U2399
g49 and DATAI_25_ U2358 ; U2400
g50 and DATAI_17_ U2358 ; U2401
g51 and DATAI_26_ U2358 ; U2402
g52 and DATAI_18_ U2358 ; U2403
g53 and DATAI_27_ U2358 ; U2404
g54 and DATAI_19_ U2358 ; U2405
g55 and DATAI_28_ U2358 ; U2406
g56 and DATAI_20_ U2358 ; U2407
g57 and DATAI_29_ U2358 ; U2408
g58 and DATAI_21_ U2358 ; U2409
g59 and DATAI_30_ U2358 ; U2410
g60 and DATAI_22_ U2358 ; U2411
g61 and DATAI_31_ U2358 ; U2412
g62 and DATAI_23_ U2358 ; U2413
g63 and U2361 U3258 ; U2414
g64 and U2361 U3378 ; U2415
g65 and U2361 U3264 ; U2416
g66 and U2361 U3271 ; U2417
g67 and U2361 U3270 ; U2418
g68 and U2361 U3265 ; U2419
g69 and U2361 U4161 ; U2420
g70 and U2361 U4159 ; U2421
g71 and U4211 U5449 ; U2422
g72 and U4211 U4219 ; U2423
g73 and U2384 U3271 ; U2424
g74 and U2368 U2448 ; U2425
g75 and U3877 U3418 ; U2426
g76 nor STATE2_REG_3__SCAN_IN STATE2_REG_1__SCAN_IN ; U2427
g77 and STATE2_REG_2__SCAN_IN STATE2_REG_1__SCAN_IN ; U2428
g78 and U6354 U3418 ; U2429
g79 and U3374 STATE2_REG_1__SCAN_IN ; U2430
g80 and U4187 U7482 ; U2431
g81 and U3442 U3347 ; U2432
g82 and U4528 U3442 ; U2433
g83 and U7684 U3347 ; U2434
g84 and U4528 U7684 ; U2435
g85 and U3222 U3288 ; U2436
g86 and U4531 U3288 ; U2437
g87 and R2182_U42 R2182_U25 ; U2438
g88 and R2182_U42 U3303 ; U2439
g89 and R2182_U25 U3304 ; U2440
g90 nor R2182_U42 R2182_U25 ; U2441
g91 and R2182_U33 R2182_U34 ; U2442
g92 and R2182_U33 U3305 ; U2443
g93 and R2182_U34 U3306 ; U2444
g94 nor R2182_U33 R2182_U34 ; U2445
g95 and U3458 STATE2_REG_1__SCAN_IN ; U2446
g96 and U3565 U2452 ; U2447
g97 and R2167_U17 U3271 ; U2448
g98 and U4482 U3258 ; U2449
g99 and U4388 STATE2_REG_0__SCAN_IN ; U2450
g100 and U4239 STATE2_REG_0__SCAN_IN ; U2451
g101 and U4388 U3264 U3378 U4161 ; U2452
g102 and INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2453
g103 and U3253 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U2454
g104 and U3253 INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U2455
g105 and U3252 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2456
g106 and U3252 INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2457
g107 and U3495 U4366 ; U2458
g108 and U3251 INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2459
g109 and U3251 U3253 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U2460
g110 and U3494 U3493 ; U2461
g111 and U3251 U3252 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2462
g112 and U3492 U3491 ; U2463
g113 and U4368 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U2464
g114 and U3490 U3489 ; U2465
g115 and U3488 U3487 ; U2466
g116 and U3257 U4366 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U2467
g117 and U3486 U3485 ; U2468
g118 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U2469
g119 and U3253 U2469 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U2470
g120 and U3252 U2469 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2471
g121 and U4368 U3257 ; U2472
g122 and U7668 U7667 U3393 ; U2473
g123 and R2144_U49 U3299 ; U2474
g124 and U3441 U3345 ; U2475
g125 and R2144_U8 R2144_U49 ; U2476
g126 and U4516 U2476 ; U2477
g127 and INSTQUEUEWR_ADDR_REG_3__SCAN_IN INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U2478
g128 and U3290 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U2479
g129 and U3302 U4536 ; U2480
g130 and U4512 U2476 ; U2481
g131 and U3314 U4594 ; U2482
g132 and U4513 U2476 ; U2483
g133 and U3321 U4653 ; U2484
g134 and U4514 R2144_U43 ; U2485
g135 nor R2144_U43 R2144_U50 ; U2486
g136 and U2486 U2476 ; U2487
g137 nor INSTQUEUEWR_ADDR_REG_1__SCAN_IN INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; U2488
g138 and U3325 U4710 ; U2489
g139 and U7681 U3345 ; U2490
g140 and U4517 U4516 ; U2491
g141 and U3330 U4768 ; U2492
g142 and U4517 U4512 ; U2493
g143 and U3334 U4825 ; U2494
g144 and U4517 U4513 ; U2495
g145 and U3337 U4883 ; U2496
g146 and U4517 U2486 ; U2497
g147 and U3341 U4940 ; U2498
g148 and U4519 U3441 ; U2499
g149 and U3346 U3344 ; U2500
g150 and U4512 U2474 ; U2501
g151 and U3351 U5053 ; U2502
g152 and U4513 U2474 ; U2503
g153 and U3354 U5111 ; U2504
g154 and U2486 U2474 ; U2505
g155 and U3358 U5168 ; U2506
g156 and U4519 U7681 ; U2507
g157 nor R2144_U49 R2144_U8 ; U2508
g158 and U2508 U4516 ; U2509
g159 nor INSTQUEUEWR_ADDR_REG_3__SCAN_IN INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U2510
g160 and U3361 U5226 ; U2511
g161 and U2508 U4512 ; U2512
g162 and U3365 U5283 ; U2513
g163 and U2508 U4513 ; U2514
g164 and U3368 U5341 ; U2515
g165 and U2508 U2486 ; U2516
g166 and U3372 U5398 ; U2517
g167 and U7688 U7687 U5456 ; U2518
g168 and U3732 U5487 ; U2519
g169 and U4207 U3433 ; U2520
g170 and U3389 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2521
g171 and U5471 U5499 ; U2522
g172 and U2522 U2521 ; U2523
g173 and U3253 U3389 ; U2524
g174 and U2522 U2524 ; U2525
g175 and U5507 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U2526
g176 and U2522 U2526 ; U2527
g177 and U5507 U3253 ; U2528
g178 and U2522 U2528 ; U2529
g179 and U5471 U3388 ; U2530
g180 and U2530 U2521 ; U2531
g181 and U2530 U2524 ; U2532
g182 and U2530 U2526 ; U2533
g183 and U2530 U2528 ; U2534
g184 and U5499 U3425 ; U2535
g185 and U2535 U2521 ; U2536
g186 and U2535 U2524 ; U2537
g187 and U2535 U2526 ; U2538
g188 and U2535 U2528 ; U2539
g189 and U3425 U3388 ; U2540
g190 and U2521 U2540 ; U2541
g191 and U2524 U2540 ; U2542
g192 and U2526 U2540 ; U2543
g193 and U2528 U2540 ; U2544
g194 and U5468 U7708 ; U2545
g195 and U2545 U2454 ; U2546
g196 and U2545 U3486 ; U2547
g197 and U2545 U4366 ; U2548
g198 and U2545 U2456 ; U2549
g199 and U5468 U3443 ; U2550
g200 and U2550 U2454 ; U2551
g201 and U2550 U3486 ; U2552
g202 and U2550 U4366 ; U2553
g203 and U2550 U2456 ; U2554
g204 and U7708 U3429 ; U2555
g205 and U2555 U2454 ; U2556
g206 and U2555 U3486 ; U2557
g207 and U2555 U4366 ; U2558
g208 and U2555 U2456 ; U2559
g209 and U3443 U3429 ; U2560
g210 and U2560 U2454 ; U2561
g211 and U2560 U3486 ; U2562
g212 and U2560 U4366 ; U2563
g213 and U2560 U2456 ; U2564
g214 and U7053 U4367 ; U2565
g215 and U7053 U2460 ; U2566
g216 and U7053 U2462 ; U2567
g217 and U7053 U4368 ; U2568
g218 and U7053 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U2569
g219 and U2569 U3486 ; U2570
g220 and U2569 U2454 ; U2571
g221 and U2569 U2456 ; U2572
g222 and U2569 U4366 ; U2573
g223 and U4367 U3432 ; U2574
g224 and U2460 U3432 ; U2575
g225 and U2462 U3432 ; U2576
g226 and U4368 U3432 ; U2577
g227 and U3432 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U2578
g228 and U2578 U3486 ; U2579
g229 and U2578 U2454 ; U2580
g230 and U2578 U2456 ; U2581
g231 and U2578 U4366 ; U2582
g232 and U7778 U4172 ; U2583
g233 and U2583 U2524 ; U2584
g234 and U2583 U2521 ; U2585
g235 and U2583 U2528 ; U2586
g236 and U2583 U2526 ; U2587
g237 and U7778 U3439 ; U2588
g238 and U2588 U2524 ; U2589
g239 and U2588 U2521 ; U2590
g240 and U2588 U2528 ; U2591
g241 and U2588 U2526 ; U2592
g242 and U4172 U3444 ; U2593
g243 and U2593 U2524 ; U2594
g244 and U2593 U2521 ; U2595
g245 and U2593 U2528 ; U2596
g246 and U2593 U2526 ; U2597
g247 and U3444 U3439 ; U2598
g248 and U2598 U2524 ; U2599
g249 and U2598 U2521 ; U2600
g250 and U2598 U2528 ; U2601
g251 and U2598 U2526 ; U2602
g252 and U3376 STATE2_REG_0__SCAN_IN ; U2603
g253 and U2379 EBX_REG_31__SCAN_IN ; U2604
g254 and U3521 U2607 U3520 U3519 U3518 ; U2605
g255 and U7492 U3414 ; U2606
g256 and U7660 U7659 ; U2607
g257 and U7775 U7774 ; U2608
g258 nand U6744 U3993 ; U2609
g259 nand U6741 U3992 ; U2610
g260 nand U6738 U3991 ; U2611
g261 nand U6735 U3990 ; U2612
g262 nand U6844 U4014 ; U2613
g263 nand U6841 U6842 U6843 ; U2614
g264 nand U6838 U6839 U6840 ; U2615
g265 nand U6835 U6836 U6837 ; U2616
g266 nand U6832 U6833 U6834 ; U2617
g267 nand U6829 U6830 U6831 ; U2618
g268 and R2144_U145 U6734 ; U2620
g269 and R2144_U145 U6734 ; U2621
g270 and R2144_U145 U6734 ; U2622
g271 and R2144_U145 U6734 ; U2623
g272 and R2144_U145 U6734 ; U2624
g273 and R2144_U145 U6734 ; U2625
g274 and R2144_U145 U6734 ; U2626
g275 and R2144_U145 U6734 ; U2627
g276 and R2144_U145 U6734 ; U2628
g277 and R2144_U145 U6734 ; U2629
g278 and R2144_U145 U6734 ; U2630
g279 and R2144_U145 U6734 ; U2631
g280 and R2144_U145 U6734 ; U2632
g281 and R2144_U145 U6734 ; U2633
g282 and R2144_U11 U6734 ; U2634
g283 and R2144_U37 U6734 ; U2635
g284 and R2144_U38 U6734 ; U2636
g285 and R2144_U39 U6734 ; U2637
g286 and R2144_U40 U6734 ; U2638
g287 and R2144_U41 U6734 ; U2639
g288 and R2144_U42 U6734 ; U2640
g289 and R2144_U30 U6734 ; U2641
g290 and R2144_U80 U6734 ; U2642
g291 and R2144_U10 U6734 ; U2643
g292 and R2144_U9 U6734 ; U2644
g293 and R2144_U45 U6734 ; U2645
g294 and R2144_U47 U6734 ; U2646
g295 and R2144_U8 U6734 ; U2647
g296 nand U3427 U6857 ; U2648
g297 and R2144_U50 U6734 ; U2649
g298 and U6858 STATE2_REG_2__SCAN_IN ; U2650
g299 nand U6757 U6756 U6758 ; U2651
g300 nand U6759 U3997 ; U2652
g301 nand U6768 U3999 ; U2653
g302 nand U6772 U4000 ; U2654
g303 nand U6776 U4001 ; U2655
g304 nand U6780 U4002 ; U2656
g305 nand U6784 U4003 ; U2657
g306 nand U6788 U4004 ; U2658
g307 nand U6792 U4005 ; U2659
g308 nand U6796 U4006 ; U2660
g309 nand U6800 U4007 ; U2661
g310 nand U6804 U4008 ; U2662
g311 nand U6813 U4010 ; U2663
g312 nand U6817 U4011 ; U2664
g313 nand U6821 U4012 ; U2665
g314 nand U6825 U4013 ; U2666
g315 nand U6747 U3994 ; U2667
g316 nand U6755 U6754 U3996 U6751 ; U2668
g317 nand U6767 U6766 U3998 U6763 ; U2669
g318 nand U6812 U6811 U4009 U6808 ; U2670
g319 nand U6851 U6850 U4015 U6847 ; U2671
g320 nand U6854 U6852 U6853 U6856 U6855 ; U2672
g321 nand U7446 U7445 ; U2673
g322 nand U7448 U7447 ; U2674
g323 nand U4156 U7451 ; U2675
g324 nand U4157 U7454 ; U2676
g325 nand U7782 U7781 U7455 ; U2677
g326 nand U7444 U3271 ; U2678
g327 nand U7393 U7392 ; U2679
g328 nand U7395 U7394 ; U2680
g329 nand U7399 U7398 ; U2681
g330 nand U7401 U7400 ; U2682
g331 nand U7403 U7402 ; U2683
g332 nand U7405 U7404 ; U2684
g333 nand U7407 U7406 ; U2685
g334 nand U7409 U7408 ; U2686
g335 nand U7411 U7410 ; U2687
g336 nand U7413 U7412 ; U2688
g337 nand U7415 U7414 ; U2689
g338 nand U7417 U7416 ; U2690
g339 nand U7421 U7420 ; U2691
g340 nand U7423 U7422 ; U2692
g341 nand U7425 U7424 ; U2693
g342 nand U7427 U7426 ; U2694
g343 nand U7429 U7428 ; U2695
g344 nand U7431 U7430 ; U2696
g345 nand U7433 U7432 ; U2697
g346 nand U7435 U7434 ; U2698
g347 nand U7437 U7436 ; U2699
g348 nand U7439 U7438 ; U2700
g349 nand U7381 U7380 ; U2701
g350 nand U7383 U7382 ; U2702
g351 nand U7385 U7384 ; U2703
g352 nand U7387 U7386 ; U2704
g353 nand U7389 U7388 ; U2705
g354 nand U7391 U7390 ; U2706
g355 nand U7397 U7396 ; U2707
g356 nand U7419 U7418 ; U2708
g357 nand U7441 U7440 ; U2709
g358 nand U7443 U7442 ; U2710
g359 nand U7365 U7364 ; U2711
g360 nand U7367 U7366 ; U2712
g361 nand U4153 U4227 ; U2713
g362 nand U7374 U7373 U4154 U3421 ; U2714
g363 nand U4227 U4155 ; U2715
g364 nand U7353 U7352 ; U2716
g365 nand U7355 U7354 ; U2717
g366 nand U4149 U7356 ; U2718
g367 nand U4150 U7358 ; U2719
g368 nand U4151 U7360 ; U2720
g369 nand U4152 U7362 ; U2721
g370 nand U4147 U4180 ; U2722
g371 and U7224 U7071 ; U2723
g372 and U7241 U7071 ; U2724
g373 and U7258 U7071 ; U2725
g374 and U7608 U7071 ; U2726
g375 and U7290 U7071 ; U2727
g376 and U7307 U7071 ; U2728
g377 and U7324 U7071 ; U2729
g378 and U7341 U7071 ; U2730
g379 nand U2606 U7342 ; U2731
g380 and U7071 U7070 ; U2732
g381 and U7102 U7071 ; U2733
g382 and U7119 U7071 ; U2734
g383 and U7606 U7071 ; U2735
g384 and U7151 U7071 ; U2736
g385 and U7168 U7071 ; U2737
g386 and U7185 U7071 ; U2738
g387 and U7202 U7071 ; U2739
g388 and U7051 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; U2740
g389 nand U4066 U7084 ; U2741
g390 and U7480 U7479 ; U2742
g391 and U7494 U7458 ; U2743
g392 and U7467 U7466 ; U2744
g393 nand U7036 U7035 ; U2745
g394 nand U7038 U7037 ; U2746
g395 nand U7040 U7039 ; U2747
g396 nand U7604 U7041 ; U2748
g397 nand U7043 U7042 ; U2749
g398 nand U7045 U7044 ; U2750
g399 nand U4049 U7046 ; U2751
g400 nand U4050 U7048 U7049 ; U2752
g401 and U6945 U6897 ; U2753
g402 and U6962 U6897 ; U2754
g403 and U6979 U6897 ; U2755
g404 and U7603 U6897 ; U2756
g405 and U7011 U6897 ; U2757
g406 and U7028 U6897 ; U2758
g407 and U6897 U6896 ; U2759
g408 and U6914 U6897 ; U2760
g409 nand U6916 U6915 ; U2761
g410 nand U6918 U6917 ; U2762
g411 nand U6920 U6919 ; U2763
g412 nand U6922 U6921 ; U2764
g413 nand U6924 U6923 U6925 ; U2765
g414 nand U6927 U6926 U6928 ; U2766
g415 nand U7031 U7029 U7030 ; U2767
g416 nand U7034 U7032 U7033 ; U2768
g417 and R2144_U145 U4147 ; U2769
g418 and U4147 R2144_U145 ; U2770
g419 and U4147 R2144_U11 ; U2771
g420 and U4147 R2144_U37 ; U2772
g421 and U4147 R2144_U38 ; U2773
g422 and U4147 R2144_U39 ; U2774
g423 and U4147 R2144_U40 ; U2775
g424 and U4147 R2144_U41 ; U2776
g425 and U4147 R2144_U42 ; U2777
g426 and U4147 R2144_U30 ; U2778
g427 nand U6860 U6859 ; U2779
g428 nand U6862 U6861 ; U2780
g429 nand U6864 U6863 ; U2781
g430 nand U6866 U6865 ; U2782
g431 nand U6868 U6867 ; U2783
g432 nand U6870 U6869 ; U2784
g433 nand U6872 U6873 U6871 ; U2785
g434 nand U4016 U6875 U6874 ; U2786
g435 nand U6878 U6879 U6877 ; U2787
g436 nand U6605 U3419 U7486 ; U2788
g437 nand U7638 U6601 ; U2789
g438 nand U6600 U6599 ; U2790
g439 nand U7757 U7756 U4231 ; U2791
g440 nand U7753 U7752 U4231 ; U2792
g441 nand U6589 U4236 ; U2793
g442 nand U7745 U7744 U4228 ; U2794
g443 nand U7735 U7734 U4228 ; U2795
g444 nand U6581 U3936 U3937 U6579 U6583 ; U2796
g445 nand U6574 U3934 U3935 U6572 U6576 ; U2797
g446 nand U6567 U3932 U3933 U6565 U6569 ; U2798
g447 nand U6560 U3930 U3931 U6558 U6562 ; U2799
g448 nand U6553 U3928 U3929 U6551 U6555 ; U2800
g449 nand U6546 U3926 U3927 U6544 U6548 ; U2801
g450 nand U6539 U3924 U3925 U6537 U6541 ; U2802
g451 nand U6532 U3922 U3923 U6530 U6534 ; U2803
g452 nand U6525 U3920 U3921 U6523 U6527 ; U2804
g453 nand U6518 U3918 U3919 U6516 U6520 ; U2805
g454 nand U6511 U3916 U3917 U6509 U6513 ; U2806
g455 nand U6504 U3914 U3915 U6502 U6506 ; U2807
g456 nand U3912 U6497 U3913 U6495 U6499 ; U2808
g457 nand U3910 U6490 U3911 U6488 U6492 ; U2809
g458 nand U3908 U6483 U3909 U6481 U6485 ; U2810
g459 nand U6476 U6475 U3907 U3906 U6478 ; U2811
g460 nand U6469 U6468 U3905 U3904 U6471 ; U2812
g461 nand U3903 U6462 U3902 U6461 U6464 ; U2813
g462 nand U3901 U6455 U3900 U6454 U6457 ; U2814
g463 nand U3899 U6448 U3898 U6447 U6450 ; U2815
g464 nand U3897 U6441 U3896 U6440 U6443 ; U2816
g465 nand U3895 U6434 U3894 U6433 U6436 ; U2817
g466 nand U3893 U6427 U3892 U6426 U6429 ; U2818
g467 nand U3891 U6420 U3890 U6419 U6422 ; U2819
g468 nand U3889 U6413 U3888 U6412 U6415 ; U2820
g469 nand U3887 U6406 U3886 U6405 U6408 ; U2821
g470 nand U3884 U6397 U6398 U3885 ; U2822
g471 nand U3882 U6389 U3883 U6391 U6390 ; U2823
g472 nand U6381 U6380 U6382 U3881 ; U2824
g473 nand U6373 U6372 U6374 U3880 ; U2825
g474 nand U6365 U6364 U6366 U3879 ; U2826
g475 nand U6357 U6356 U6358 U3878 ; U2827
g476 nand U6347 U6346 ; U2828
g477 nand U6344 U6345 U6343 ; U2829
g478 nand U6341 U6342 U6340 ; U2830
g479 nand U6338 U6339 U6337 ; U2831
g480 nand U6335 U6336 U6334 ; U2832
g481 nand U6332 U6333 U6331 ; U2833
g482 nand U6329 U6330 U6328 ; U2834
g483 nand U6326 U6327 U6325 ; U2835
g484 nand U6323 U6324 U6322 ; U2836
g485 nand U6320 U6321 U6319 ; U2837
g486 nand U6317 U6318 U6316 ; U2838
g487 nand U6314 U6315 U6313 ; U2839
g488 nand U6311 U6312 U6310 ; U2840
g489 nand U6308 U6309 U6307 ; U2841
g490 nand U6305 U6306 U6304 ; U2842
g491 nand U6302 U6303 U6301 ; U2843
g492 nand U6299 U6300 U6298 ; U2844
g493 nand U6296 U6297 U6295 ; U2845
g494 nand U6293 U6294 U6292 ; U2846
g495 nand U6290 U6291 U6289 ; U2847
g496 nand U6287 U6288 U6286 ; U2848
g497 nand U6284 U6285 U6283 ; U2849
g498 nand U6281 U6282 U6280 ; U2850
g499 nand U6278 U6279 U6277 ; U2851
g500 nand U6275 U6276 U6274 ; U2852
g501 nand U6272 U6273 U6271 ; U2853
g502 nand U6269 U6270 U6268 ; U2854
g503 nand U6266 U6267 U6265 ; U2855
g504 nand U6263 U6264 U6262 ; U2856
g505 nand U6260 U6261 U6259 ; U2857
g506 nand U6257 U6258 U6256 ; U2858
g507 nand U6254 U6253 U6255 ; U2859
g508 nand U4164 U6250 ; U2860
g509 nand U6247 U6246 U6249 U6248 ; U2861
g510 nand U6243 U6242 U6245 U6244 ; U2862
g511 nand U6239 U6238 U6241 U6240 ; U2863
g512 nand U6235 U6234 U6237 U6236 ; U2864
g513 nand U6231 U6230 U6233 U6232 ; U2865
g514 nand U6227 U6226 U6229 U6228 ; U2866
g515 nand U6223 U6222 U6225 U6224 ; U2867
g516 nand U6219 U6218 U6221 U6220 ; U2868
g517 nand U6215 U6214 U6217 U6216 ; U2869
g518 nand U6211 U6210 U6213 U6212 ; U2870
g519 nand U6207 U6206 U6209 U6208 ; U2871
g520 nand U6203 U6202 U6205 U6204 ; U2872
g521 nand U6199 U6198 U6201 U6200 ; U2873
g522 nand U6195 U6194 U6197 U6196 ; U2874
g523 nand U6191 U6190 U6193 U6192 ; U2875
g524 nand U6189 U6187 U6188 ; U2876
g525 nand U6186 U6184 U6185 ; U2877
g526 nand U6183 U6181 U6182 ; U2878
g527 nand U6180 U6178 U6179 ; U2879
g528 nand U6177 U6175 U6176 ; U2880
g529 nand U6174 U6172 U6173 ; U2881
g530 nand U6171 U6169 U6170 ; U2882
g531 nand U6168 U6166 U6167 ; U2883
g532 nand U6165 U6163 U6164 ; U2884
g533 nand U6162 U6160 U6161 ; U2885
g534 nand U6159 U6157 U6158 ; U2886
g535 nand U6156 U6154 U6155 ; U2887
g536 nand U6153 U6151 U6152 ; U2888
g537 nand U6150 U6148 U6149 ; U2889
g538 nand U6146 U6145 U6147 ; U2890
g539 nand U6143 U6142 U6144 ; U2891
g540 and U6043 DATAO_REG_31__SCAN_IN ; U2892
g541 nand U3870 U6134 ; U2893
g542 nand U3869 U6131 ; U2894
g543 nand U3868 U6128 ; U2895
g544 nand U3867 U6125 ; U2896
g545 nand U3866 U6122 ; U2897
g546 nand U3865 U6119 ; U2898
g547 nand U3864 U6116 ; U2899
g548 nand U3863 U6113 ; U2900
g549 nand U3862 U6110 ; U2901
g550 nand U3861 U6107 ; U2902
g551 nand U3860 U6104 ; U2903
g552 nand U3859 U6101 ; U2904
g553 nand U3858 U6098 ; U2905
g554 nand U3857 U6095 ; U2906
g555 nand U3856 U6092 ; U2907
g556 nand U6090 U6089 U6091 ; U2908
g557 nand U6087 U6086 U6088 ; U2909
g558 nand U6084 U6083 U6085 ; U2910
g559 nand U6081 U6080 U6082 ; U2911
g560 nand U6078 U6077 U6079 ; U2912
g561 nand U6075 U6074 U6076 ; U2913
g562 nand U6072 U6071 U6073 ; U2914
g563 nand U6069 U6068 U6070 ; U2915
g564 nand U6066 U6065 U6067 ; U2916
g565 nand U6063 U6062 U6064 ; U2917
g566 nand U6060 U6059 U6061 ; U2918
g567 nand U6057 U6056 U6058 ; U2919
g568 nand U6054 U6053 U6055 ; U2920
g569 nand U6051 U6050 U6052 ; U2921
g570 nand U6048 U6047 U6049 ; U2922
g571 nand U6045 U6044 U6046 ; U2923
g572 nand U7528 U7530 ; U2924
g573 nand U7527 U7532 ; U2925
g574 nand U7526 U7534 ; U2926
g575 nand U7525 U7536 ; U2927
g576 nand U7524 U7538 ; U2928
g577 nand U7523 U7540 ; U2929
g578 nand U7522 U7542 ; U2930
g579 nand U7521 U7544 ; U2931
g580 nand U7520 U7546 ; U2932
g581 nand U7519 U7548 ; U2933
g582 nand U7518 U7550 ; U2934
g583 nand U7517 U7552 ; U2935
g584 nand U7516 U7554 ; U2936
g585 nand U7515 U7556 ; U2937
g586 nand U7514 U7558 ; U2938
g587 nand U7513 U7560 ; U2939
g588 nand U7512 U7562 ; U2940
g589 nand U7511 U7564 ; U2941
g590 nand U7510 U7566 ; U2942
g591 nand U7509 U7568 ; U2943
g592 nand U7508 U7570 ; U2944
g593 nand U7507 U7572 ; U2945
g594 nand U7506 U7574 ; U2946
g595 nand U7505 U7576 ; U2947
g596 nand U7504 U7578 ; U2948
g597 nand U7503 U7580 ; U2949
g598 nand U7502 U7582 ; U2950
g599 nand U7501 U7584 ; U2951
g600 nand U7500 U7586 ; U2952
g601 nand U7499 U7588 ; U2953
g602 nand U7498 U7590 ; U2954
g603 nand U5944 U5942 U5946 U5943 U5945 ; U2955
g604 nand U5939 U5937 U5941 U5938 U5940 ; U2956
g605 nand U5934 U5932 U5936 U5933 U5935 ; U2957
g606 nand U5929 U5927 U5931 U5928 U5930 ; U2958
g607 nand U5924 U5922 U5926 U5923 U5925 ; U2959
g608 nand U5919 U5917 U5921 U5918 U5920 ; U2960
g609 nand U5914 U5912 U5916 U5913 U5915 ; U2961
g610 nand U5909 U5907 U5911 U5908 U5910 ; U2962
g611 nand U5904 U5902 U5906 U5903 U5905 ; U2963
g612 nand U5899 U5897 U5901 U5898 U5900 ; U2964
g613 nand U5894 U5892 U5896 U5893 U5895 ; U2965
g614 nand U5889 U5887 U5891 U5888 U5890 ; U2966
g615 nand U5884 U5882 U5886 U5883 U5885 ; U2967
g616 nand U5879 U5877 U5881 U5878 U5880 ; U2968
g617 nand U5874 U5872 U5876 U5873 U5875 ; U2969
g618 nand U5869 U5867 U5871 U5868 U5870 ; U2970
g619 nand U5864 U5862 U5866 U5863 U5865 ; U2971
g620 nand U5859 U5857 U5861 U5858 U5860 ; U2972
g621 nand U5854 U5852 U5856 U5853 U5855 ; U2973
g622 nand U5849 U5847 U5851 U5848 U5850 ; U2974
g623 nand U5844 U5842 U5846 U5843 U5845 ; U2975
g624 nand U5839 U5837 U5841 U5838 U5840 ; U2976
g625 nand U5834 U5832 U5836 U5833 U5835 ; U2977
g626 nand U5829 U5827 U5831 U5828 U5830 ; U2978
g627 nand U5824 U5822 U5823 U5826 U5825 ; U2979
g628 nand U5819 U5817 U5818 U5821 U5820 ; U2980
g629 nand U5814 U5812 U5813 U5816 U5815 ; U2981
g630 nand U5809 U5807 U5808 U5811 U5810 ; U2982
g631 nand U5804 U5802 U5803 U5806 U5805 ; U2983
g632 nand U5799 U5797 U5798 U5801 U5800 ; U2984
g633 nand U5793 U5792 U5794 U5796 U5795 ; U2985
g634 nand U5788 U5787 U5789 U5791 U5790 ; U2986
g635 nand U3849 U3847 U5775 U5777 ; U2987
g636 nand U3846 U3844 U5768 U5770 ; U2988
g637 nand U3843 U3841 U5761 U5763 ; U2989
g638 nand U3840 U3838 U5754 U5756 ; U2990
g639 nand U3837 U3835 U5747 U5749 ; U2991
g640 nand U3834 U3832 U5740 U5742 ; U2992
g641 nand U3831 U3829 U5733 U5735 ; U2993
g642 nand U3828 U3826 U5726 U5728 ; U2994
g643 nand U3825 U3823 U5719 U5721 ; U2995
g644 nand U3822 U3820 U5712 U5714 ; U2996
g645 nand U3819 U3817 U5705 U5707 ; U2997
g646 nand U3816 U3814 U5698 U5700 ; U2998
g647 nand U3813 U3811 U5691 U5693 ; U2999
g648 nand U3810 U3808 U5684 U5686 ; U3000
g649 nand U3807 U3805 U5677 U5679 ; U3001
g650 nand U3804 U3802 U5670 U5672 ; U3002
g651 nand U3801 U3799 U5663 U5665 ; U3003
g652 nand U3798 U3796 U5656 U5658 ; U3004
g653 nand U3795 U3793 U5649 U5651 ; U3005
g654 nand U3790 U3792 U5644 ; U3006
g655 nand U3787 U3789 U5637 ; U3007
g656 nand U3784 U3786 U5630 ; U3008
g657 nand U3781 U3783 U5623 ; U3009
g658 nand U3778 U3780 U5616 ; U3010
g659 nand U3775 U3777 U5609 ; U3011
g660 nand U3772 U3774 U5602 ; U3012
g661 nand U3769 U3771 U5595 ; U3013
g662 nand U3766 U3768 U5588 ; U3014
g663 nand U3763 U3764 ; U3015
g664 nand U3760 U3759 U3762 ; U3016
g665 nand U3756 U3755 U3758 ; U3017
g666 nand U3752 U3751 U3754 ; U3018
g667 and U5525 INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; U3019
g668 nand U5448 U5447 U3718 ; U3020
g669 nand U5443 U5442 U3717 ; U3021
g670 nand U5438 U5437 U3716 ; U3022
g671 nand U5433 U5432 U3715 ; U3023
g672 nand U7600 U5428 U3714 ; U3024
g673 nand U5424 U5423 U3713 ; U3025
g674 nand U5419 U5418 U3712 ; U3026
g675 nand U5414 U5413 U3711 ; U3027
g676 nand U5392 U5391 U3709 ; U3028
g677 nand U5387 U5386 U3708 ; U3029
g678 nand U5382 U5381 U3707 ; U3030
g679 nand U5377 U5376 U3706 ; U3031
g680 nand U5372 U5371 U3705 ; U3032
g681 nand U5367 U5366 U3704 ; U3033
g682 nand U5362 U5361 U3703 ; U3034
g683 nand U5357 U5356 U3702 ; U3035
g684 nand U5334 U5333 U3700 ; U3036
g685 nand U5329 U5328 U3699 ; U3037
g686 nand U5324 U5323 U3698 ; U3038
g687 nand U5319 U5318 U3697 ; U3039
g688 nand U5314 U5313 U3696 ; U3040
g689 nand U5309 U5308 U3695 ; U3041
g690 nand U5304 U5303 U3694 ; U3042
g691 nand U5299 U5298 U3693 ; U3043
g692 nand U5277 U5276 U3691 ; U3044
g693 nand U5272 U5271 U3690 ; U3045
g694 nand U5267 U5266 U3689 ; U3046
g695 nand U5262 U5261 U3688 ; U3047
g696 nand U5257 U5256 U3687 ; U3048
g697 nand U5252 U5251 U3686 ; U3049
g698 nand U5247 U5246 U3685 ; U3050
g699 nand U5242 U5241 U3684 ; U3051
g700 nand U5219 U5218 U3682 ; U3052
g701 nand U5214 U5213 U3681 ; U3053
g702 nand U5209 U5208 U3680 ; U3054
g703 nand U5204 U5203 U3679 ; U3055
g704 nand U5199 U5198 U3678 ; U3056
g705 nand U5194 U5193 U3677 ; U3057
g706 nand U5189 U5188 U3676 ; U3058
g707 nand U5184 U5183 U3675 ; U3059
g708 nand U5162 U5161 U3673 ; U3060
g709 nand U5157 U5156 U3672 ; U3061
g710 nand U5152 U5151 U3671 ; U3062
g711 nand U5147 U5146 U3670 ; U3063
g712 nand U5142 U5141 U3669 ; U3064
g713 nand U5137 U5136 U3668 ; U3065
g714 nand U5132 U5131 U3667 ; U3066
g715 nand U5127 U5126 U3666 ; U3067
g716 nand U5104 U5103 U3664 ; U3068
g717 nand U5099 U5098 U3663 ; U3069
g718 nand U5094 U5093 U3662 ; U3070
g719 nand U5089 U5088 U3661 ; U3071
g720 nand U5084 U5083 U3660 ; U3072
g721 nand U5079 U5078 U3659 ; U3073
g722 nand U5074 U5073 U3658 ; U3074
g723 nand U5069 U5068 U3657 ; U3075
g724 nand U5047 U5046 U3655 ; U3076
g725 nand U5042 U5041 U3654 ; U3077
g726 nand U5037 U5036 U3653 ; U3078
g727 nand U5032 U5031 U3652 ; U3079
g728 nand U5027 U5026 U3651 ; U3080
g729 nand U5022 U5021 U3650 ; U3081
g730 nand U5017 U5016 U3649 ; U3082
g731 nand U5012 U5011 U3648 ; U3083
g732 nand U4991 U4990 U3646 ; U3084
g733 nand U4986 U4985 U3645 ; U3085
g734 nand U4981 U4980 U3644 ; U3086
g735 nand U4976 U4975 U3643 ; U3087
g736 nand U4971 U4970 U3642 ; U3088
g737 nand U4966 U4965 U3641 ; U3089
g738 nand U4961 U4960 U3640 ; U3090
g739 nand U4956 U4955 U3639 ; U3091
g740 nand U4934 U4933 U3637 ; U3092
g741 nand U4929 U4928 U3636 ; U3093
g742 nand U4924 U4923 U3635 ; U3094
g743 nand U4919 U4918 U3634 ; U3095
g744 nand U4914 U4913 U3633 ; U3096
g745 nand U4909 U4908 U3632 ; U3097
g746 nand U4904 U4903 U3631 ; U3098
g747 nand U4899 U4898 U3630 ; U3099
g748 nand U4876 U4875 U3628 ; U3100
g749 nand U4871 U4870 U3627 ; U3101
g750 nand U4866 U4865 U3626 ; U3102
g751 nand U4861 U4860 U3625 ; U3103
g752 nand U4856 U4855 U3624 ; U3104
g753 nand U4851 U4850 U3623 ; U3105
g754 nand U4846 U4845 U3622 ; U3106
g755 nand U4841 U4840 U3621 ; U3107
g756 nand U4819 U4818 U3619 ; U3108
g757 nand U4814 U4813 U3618 ; U3109
g758 nand U4809 U4808 U3617 ; U3110
g759 nand U4804 U4803 U3616 ; U3111
g760 nand U4799 U4798 U3615 ; U3112
g761 nand U4794 U4793 U3614 ; U3113
g762 nand U4789 U4788 U3613 ; U3114
g763 nand U4784 U4783 U3612 ; U3115
g764 nand U4761 U4760 U3610 ; U3116
g765 nand U4756 U4755 U3609 ; U3117
g766 nand U4751 U4750 U3608 ; U3118
g767 nand U4746 U4745 U3607 ; U3119
g768 nand U4741 U4740 U3606 ; U3120
g769 nand U4736 U4735 U3605 ; U3121
g770 nand U4731 U4730 U3604 ; U3122
g771 nand U4726 U4725 U3603 ; U3123
g772 nand U4704 U4703 U3601 ; U3124
g773 nand U4699 U4698 U3600 ; U3125
g774 nand U4694 U4693 U3599 ; U3126
g775 nand U4689 U4688 U3598 ; U3127
g776 nand U4684 U4683 U3597 ; U3128
g777 nand U4679 U4678 U3596 ; U3129
g778 nand U4674 U4673 U3595 ; U3130
g779 nand U4669 U4668 U3594 ; U3131
g780 nand U4645 U4644 U3592 ; U3132
g781 nand U4640 U4639 U3591 ; U3133
g782 nand U4635 U4634 U3590 ; U3134
g783 nand U4630 U4629 U3589 ; U3135
g784 nand U4625 U4624 U3588 ; U3136
g785 nand U4620 U4619 U3587 ; U3137
g786 nand U4615 U4614 U3586 ; U3138
g787 nand U4610 U4609 U3585 ; U3139
g788 nand U4587 U4586 U3583 ; U3140
g789 nand U4582 U4581 U3582 ; U3141
g790 nand U4577 U4576 U3581 ; U3142
g791 nand U4572 U4571 U3580 ; U3143
g792 nand U4567 U4566 U3579 ; U3144
g793 nand U4562 U4561 U3578 ; U3145
g794 nand U4557 U4556 U3577 ; U3146
g795 nand U4552 U4551 U3576 ; U3147
g796 nand U7678 U7677 U3574 ; U3148
g797 nand U4508 U4507 U4506 U4232 ; U3149
g798 nand U3570 U4504 ; U3150
g799 and U7638 DATAWIDTH_REG_31__SCAN_IN ; U3151
g800 and U7638 DATAWIDTH_REG_30__SCAN_IN ; U3152
g801 and U7638 DATAWIDTH_REG_29__SCAN_IN ; U3153
g802 and U7638 DATAWIDTH_REG_28__SCAN_IN ; U3154
g803 and U7638 DATAWIDTH_REG_27__SCAN_IN ; U3155
g804 and U7638 DATAWIDTH_REG_26__SCAN_IN ; U3156
g805 and U7638 DATAWIDTH_REG_25__SCAN_IN ; U3157
g806 and U7638 DATAWIDTH_REG_24__SCAN_IN ; U3158
g807 and U7638 DATAWIDTH_REG_23__SCAN_IN ; U3159
g808 and U7638 DATAWIDTH_REG_22__SCAN_IN ; U3160
g809 and U7638 DATAWIDTH_REG_21__SCAN_IN ; U3161
g810 and U7638 DATAWIDTH_REG_20__SCAN_IN ; U3162
g811 and U7638 DATAWIDTH_REG_19__SCAN_IN ; U3163
g812 and U7638 DATAWIDTH_REG_18__SCAN_IN ; U3164
g813 and U7638 DATAWIDTH_REG_17__SCAN_IN ; U3165
g814 and U7638 DATAWIDTH_REG_16__SCAN_IN ; U3166
g815 and U7638 DATAWIDTH_REG_15__SCAN_IN ; U3167
g816 and U7638 DATAWIDTH_REG_14__SCAN_IN ; U3168
g817 and U7638 DATAWIDTH_REG_13__SCAN_IN ; U3169
g818 and U7638 DATAWIDTH_REG_12__SCAN_IN ; U3170
g819 and U7638 DATAWIDTH_REG_11__SCAN_IN ; U3171
g820 and U7638 DATAWIDTH_REG_10__SCAN_IN ; U3172
g821 and U7638 DATAWIDTH_REG_9__SCAN_IN ; U3173
g822 and U7638 DATAWIDTH_REG_8__SCAN_IN ; U3174
g823 and U7638 DATAWIDTH_REG_7__SCAN_IN ; U3175
g824 and U7638 DATAWIDTH_REG_6__SCAN_IN ; U3176
g825 and U7638 DATAWIDTH_REG_5__SCAN_IN ; U3177
g826 and U7638 DATAWIDTH_REG_4__SCAN_IN ; U3178
g827 and U7638 DATAWIDTH_REG_3__SCAN_IN ; U3179
g828 and U7638 DATAWIDTH_REG_2__SCAN_IN ; U3180
g829 nand U7635 U7634 U4363 ; U3181
g830 nand U7633 U7632 U3483 ; U3182
g831 nand U3482 U4357 ; U3183
g832 nand U4343 U4342 U4344 ; U3184
g833 nand U4340 U4339 U4341 ; U3185
g834 nand U4337 U4336 U4338 ; U3186
g835 nand U4334 U4333 U4335 ; U3187
g836 nand U4331 U4330 U4332 ; U3188
g837 nand U4328 U4327 U4329 ; U3189
g838 nand U4325 U4324 U4326 ; U3190
g839 nand U4322 U4321 U4323 ; U3191
g840 nand U4319 U4318 U4320 ; U3192
g841 nand U4316 U4315 U4317 ; U3193
g842 nand U4313 U4312 U4314 ; U3194
g843 nand U4310 U4309 U4311 ; U3195
g844 nand U4307 U4306 U4308 ; U3196
g845 nand U4304 U4303 U4305 ; U3197
g846 nand U4301 U4300 U4302 ; U3198
g847 nand U4298 U4297 U4299 ; U3199
g848 nand U4295 U4294 U4296 ; U3200
g849 nand U4292 U4291 U4293 ; U3201
g850 nand U4289 U4288 U4290 ; U3202
g851 nand U4286 U4285 U4287 ; U3203
g852 nand U4283 U4282 U4284 ; U3204
g853 nand U4280 U4279 U4281 ; U3205
g854 nand U4277 U4276 U4278 ; U3206
g855 nand U4274 U4273 U4275 ; U3207
g856 nand U4271 U4270 U4272 ; U3208
g857 nand U4268 U4267 U4269 ; U3209
g858 nand U4265 U4264 U4266 ; U3210
g859 nand U4262 U4261 U4263 ; U3211
g860 nand U4259 U4258 U4260 ; U3212
g861 nand U4256 U4255 U4257 ; U3213
g862 nand U3989 U3988 U3987 U3986 ; U3214
g863 nand U3985 U3984 U3983 U3982 ; U3215
g864 nand U3981 U3980 U3979 U3978 ; U3216
g865 nand U3977 U3976 U3975 U3974 ; U3217
g866 nand U3973 U3972 U3971 U3970 ; U3218
g867 nand U3969 U3968 U3967 U3966 ; U3219
g868 nand U3965 U3964 U3963 U3962 ; U3220
g869 nand U3961 U3960 U3959 U3958 ; U3221
g870 nand U3316 U3310 ; U3222
g871 nand U2432 U3222 ; U3223
g872 nand U2432 U4531 ; U3224
g873 nand U2434 U3222 ; U3225
g874 nand U2434 U4531 ; U3226
g875 nand U2433 U3222 ; U3227
g876 nand U2433 U4531 ; U3228
g877 nand U2435 U3222 ; U3229
g878 nand U2435 U4531 ; U3230
g879 nand U3378 U3381 U5451 ; U3231
g880 nand U7074 U5452 ; U3232
g881 nand U7780 U7779 U4146 U4144 ; U3233
g882 not REQUESTPENDING_REG_SCAN_IN ; U3234
g883 not STATE_REG_1__SCAN_IN ; U3235
g884 nand U3245 STATE_REG_1__SCAN_IN ; U3236
g885 nand U4209 U3238 ; U3237
g886 not STATE_REG_2__SCAN_IN ; U3238
g887 nand U4209 STATE_REG_2__SCAN_IN ; U3239
g888 not REIP_REG_1__SCAN_IN ; U3240
g889 nand U3238 STATE_REG_1__SCAN_IN ; U3241
g890 or STATE_REG_2__SCAN_IN STATE_REG_1__SCAN_IN ; U3242
g891 not HOLD ; U3243
g892 not READY_N ; U3244
g893 not STATE_REG_0__SCAN_IN ; U3245
g894 nand U3247 STATE_REG_0__SCAN_IN ; U3246
g895 nand U3243 REQUESTPENDING_REG_SCAN_IN ; U3247
g896 or HOLD REQUESTPENDING_REG_SCAN_IN ; U3248
g897 not STATE2_REG_1__SCAN_IN ; U3249
g898 not STATE2_REG_2__SCAN_IN ; U3250
g899 not INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3251
g900 not INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3252
g901 not INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3253
g902 nand U3257 INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3254
g903 or INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3255
g904 or INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3256
g905 not INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3257
g906 nand U3555 U3554 U3553 U3552 ; U3258
g907 nand U4484 U3245 ; U3259
g908 not R2167_U17 ; U3260
g909 nand U3257 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3261
g910 nand INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3262
g911 nand U3507 U3506 U3505 U3504 ; U3263
g912 nand U3527 U4158 U3526 U3525 U3524 ; U3264
g913 nand U3545 U3544 U3543 U3542 ; U3265
g914 nand U3547 U3546 ; U3266
g915 or READY_N STATEBS16_REG_SCAN_IN ; U3267
g916 nand R2167_U17 U4485 ; U3268
g917 nand U4465 U3271 ; U3269
g918 nand U3499 U3498 U3497 U3496 ; U3270
g919 nand U3551 U3550 U3549 U3548 ; U3271
g920 nand U2473 U4489 ; U3272
g921 nand U2389 U3270 ; U3273
g922 nand U4482 U4465 ; U3274
g923 nand U4237 U2447 ; U3275
g924 nand U4448 U3378 U4161 U3265 ; U3276
g925 nand U3258 U3270 ; U3277
g926 nand U4178 U3271 ; U3278
g927 nand U4244 U2431 ; U3279
g928 nand U4166 U4497 U7614 U4213 LT_563_U6 ; U3280
g929 not STATE2_REG_0__SCAN_IN ; U3281
g930 nand U7592 STATE2_REG_0__SCAN_IN ; U3282
g931 not STATE2_REG_3__SCAN_IN ; U3283
g932 nand U3249 STATE2_REG_2__SCAN_IN ; U3284
g933 or STATE2_REG_2__SCAN_IN STATE2_REG_1__SCAN_IN ; U3285
g934 nand R2167_U17 STATE2_REG_3__SCAN_IN ; U3286
g935 nand U4535 U3281 ; U3287
g936 not INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; U3288
g937 not INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; U3289
g938 not INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; U3290
g939 not INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U3291
g940 nand INSTQUEUEWR_ADDR_REG_1__SCAN_IN INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; U3292
g941 nand U4521 U2478 ; U3293
g942 or STATE2_REG_3__SCAN_IN STATE2_REG_2__SCAN_IN ; U3294
g943 not STATEBS16_REG_SCAN_IN ; U3295
g944 not R2144_U43 ; U3296
g945 not R2144_U50 ; U3297
g946 not R2144_U49 ; U3298
g947 not R2144_U8 ; U3299
g948 nand R2144_U50 R2144_U43 ; U3300
g949 nand U3319 U3296 ; U3301
g950 nand U4515 U2475 ; U3302
g951 not R2182_U25 ; U3303
g952 not R2182_U42 ; U3304
g953 not R2182_U34 ; U3305
g954 not R2182_U33 ; U3306
g955 nand U4197 U3295 ; U3307
g956 nand U3293 U4523 ; U3308
g957 nand U3293 U4532 ; U3309
g958 nand U3288 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; U3310
g959 nand U4530 U2478 ; U3311
g960 nand R2144_U50 U3296 ; U3312
g961 nand R2144_U43 U3319 ; U3313
g962 nand U4588 U2475 ; U3314
g963 nand U3311 U4591 ; U3315
g964 nand U3289 INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; U3316
g965 nand U4529 U2478 ; U3317
g966 nand R2144_U43 U3297 ; U3318
g967 nand U3312 U3318 ; U3319
g968 nand U4514 U3296 ; U3320
g969 nand U4646 U2475 ; U3321
g970 nand U3317 U4649 ; U3322
g971 nand U3317 U4651 ; U3323
g972 nand U2488 U2478 ; U3324
g973 nand U2485 U2475 ; U3325
g974 nand U3324 U4707 ; U3326
g975 nand U3291 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; U3327
g976 nand U4526 U4521 ; U3328
g977 nand R2144_U8 U3298 ; U3329
g978 nand U2490 U4515 ; U3330
g979 nand U3328 U4764 ; U3331
g980 nand U3328 U4766 ; U3332
g981 nand U4526 U4530 ; U3333
g982 nand U2490 U4588 ; U3334
g983 nand U3333 U4822 ; U3335
g984 nand U4526 U4529 ; U3336
g985 nand U2490 U4646 ; U3337
g986 nand U3336 U4879 ; U3338
g987 nand U3336 U4881 ; U3339
g988 nand U4526 U2488 ; U3340
g989 nand U2490 U2485 ; U3341
g990 nand U3340 U4937 ; U3342
g991 nand U2479 U4521 ; U3343
g992 nand U2474 U4516 ; U3344
g993 nand U3329 U4518 U3344 ; U3345
g994 nand U2499 U4515 ; U3346
g995 nand U3327 U4527 U3343 ; U3347
g996 nand U3343 U4993 ; U3348
g997 nand U3343 U4995 ; U3349
g998 nand U4530 U2479 ; U3350
g999 nand U2499 U4588 ; U3351
g1000 nand U3350 U5050 ; U3352
g1001 nand U4529 U2479 ; U3353
g1002 nand U2499 U4646 ; U3354
g1003 nand U3353 U5107 ; U3355
g1004 nand U3353 U5109 ; U3356
g1005 nand U2488 U2479 ; U3357
g1006 nand U2499 U2485 ; U3358
g1007 nand U3357 U5165 ; U3359
g1008 nand U2510 U4521 ; U3360
g1009 nand U2507 U4515 ; U3361
g1010 nand U3360 U5222 ; U3362
g1011 nand U3360 U5224 ; U3363
g1012 nand U2510 U4530 ; U3364
g1013 nand U2507 U4588 ; U3365
g1014 nand U3364 U5280 ; U3366
g1015 nand U2510 U4529 ; U3367
g1016 nand U2507 U4646 ; U3368
g1017 nand U3367 U5337 ; U3369
g1018 nand U3367 U5339 ; U3370
g1019 nand U2510 U2488 ; U3371
g1020 nand U2507 U2485 ; U3372
g1021 nand U3371 U5395 ; U3373
g1022 not FLUSH_REG_SCAN_IN ; U3374
g1023 not GTE_485_U6 ; U3375
g1024 nand U3271 U3265 ; U3376
g1025 nand U3271 U3258 ; U3377
g1026 nand U3503 U3502 U3501 U3500 ; U3378
g1027 nand U5478 U5477 U7616 ; U3379
g1028 nand U4387 U3271 ; U3380
g1029 nand U2605 U3264 ; U3381
g1030 nand U4387 U7482 U4482 ; U3382
g1031 nand U3729 U4235 ; U3383
g1032 nand U7482 U4465 U2605 U4482 U4387 ; U3384
g1033 nand U2605 U4448 U4159 U4437 U4388 ; U3385
g1034 nand U4187 U4465 U4222 ; U3386
g1035 nand U2449 U2447 ; U3387
g1036 nand U3431 U5498 ; U3388
g1037 nand U3256 U3262 ; U3389
g1038 not LT_589_U6 ; U3390
g1039 nand U4230 U3287 U5524 ; U3391
g1040 nand U3265 U3271 STATE2_REG_0__SCAN_IN ; U3392
g1041 nand U3258 U3260 ; U3393
g1042 nand U3264 U3378 ; U3394
g1043 nand U2427 U3281 ; U3395
g1044 nand U4448 U3378 ; U3396
g1045 nand U4241 U3265 ; U3397
g1046 nand U4178 U2452 ; U3398
g1047 nand U3258 STATE2_REG_2__SCAN_IN ; U3399
g1048 not REIP_REG_0__SCAN_IN ; U3400
g1049 nand U3744 U5550 ; U3401
g1050 nand U4388 U4161 ; U3402
g1051 nand U3851 U4236 ; U3403
g1052 nand U6042 U6041 ; U3404
g1053 nand U4482 STATE2_REG_0__SCAN_IN ; U3405
g1054 nand U4387 U7482 ; U3406
g1055 nand U4194 U4465 ; U3407
g1056 nand U4182 U2431 ; U3408
g1057 nand U4198 STATE2_REG_0__SCAN_IN ; U3409
g1058 nand U4491 U3378 ; U3410
g1059 nand U4223 U6141 ; U3411
g1060 nand U4204 STATE2_REG_0__SCAN_IN ; U3412
g1061 nand U4223 U6252 ; U3413
g1062 nand U4237 U3874 U2452 STATE2_REG_0__SCAN_IN ; U3414
g1063 nand U3854 U2447 ; U3415
g1064 not EBX_REG_31__SCAN_IN ; U3416
g1065 not R2337_U58 ; U3417
g1066 nand U4216 U3875 ; U3418
g1067 nand U4197 U3249 ; U3419
g1068 nand U3950 U3946 U3943 U3940 ; U3420
g1069 nand U4194 U3258 ; U3421
g1070 not CODEFETCH_REG_SCAN_IN ; U3422
g1071 not READREQUEST_REG_SCAN_IN ; U3423
g1072 nand U2447 U4486 ; U3424
g1073 nand U3254 U5470 ; U3425
g1074 nand U4437 STATE2_REG_2__SCAN_IN ; U3426
g1075 nand U3250 STATEBS16_REG_SCAN_IN ; U3427
g1076 not U3221 ; U3428
g1077 nand U5467 U5466 ; U3429
g1078 nand U2450 U3428 ; U3430
g1079 nand U3251 INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3431
g1080 nand U3261 U7052 ; U3432
g1081 nand U4185 U4222 ; U3433
g1082 nand U4219 U4388 U4238 ; U3434
g1083 nand U4219 U3265 U4238 ; U3435
g1084 nand U4465 U4484 ; U3436
g1085 nand U4062 U7081 U4063 U4065 ; U3437
g1086 nand U4242 U4254 ; U3438
g1087 nand U4171 U3255 ; U3439
g1088 nand U2605 STATE2_REG_0__SCAN_IN ; U3440
g1089 nand U7680 U7679 ; U3441
g1090 nand U7683 U7682 ; U3442
g1091 nand U7707 U7706 ; U3443
g1092 nand U7777 U7776 ; U3444
g1093 nand U7622 U7621 ; U3445
g1094 nand U7624 U7623 ; U3446
g1095 nand U7626 U7625 ; U3447
g1096 nand U7628 U7627 ; U3448
g1097 nand U7637 U7636 ; U3449
g1098 and U3242 U4167 ; U3450
g1099 nand U7640 U7639 ; U3451
g1100 nand U7642 U7641 ; U3452
g1101 nand U7674 U7673 ; U3453
g1102 and U2427 U4203 R2182_U24 ; U3454
g1103 nand U7690 U7689 ; U3455
g1104 nand U7697 U7696 ; U3456
g1105 nand U7699 U7698 ; U3457
g1106 nand U7702 U7701 ; U3458
g1107 nand U7710 U7709 ; U3459
g1108 nand U7712 U7711 ; U3460
g1109 nand U7716 U7715 ; U3461
g1110 nand U7718 U7717 ; U3462
g1111 nand U7723 U7722 ; U3463
g1112 nand U7725 U7724 ; U3464
g1113 nand U7727 U7726 ; U3465
g1114 and R2358_U91 U4437 ; U3466
g1115 nor DATAWIDTH_REG_1__SCAN_IN REIP_REG_1__SCAN_IN ; U3467
g1116 nand U7743 U7742 ; U3468
g1117 nand U7747 U7746 ; U3469
g1118 nand U7749 U7748 ; U3470
g1119 nand U7751 U7750 ; U3471
g1120 nand U7755 U7754 ; U3472
g1121 nand U7759 U7758 ; U3473
g1122 nand U7761 U7760 ; U3474
g1123 and R2182_U24 U4203 ; U3475
g1124 nand U7763 U7762 ; U3476
g1125 nand U7765 U7764 ; U3477
g1126 nand U7767 U7766 ; U3478
g1127 nand U7769 U7768 ; U3479
g1128 nand U7771 U7770 ; U3480
g1129 and READY_N STATE_REG_1__SCAN_IN ; U3481
g1130 and U4356 U3239 ; U3482
g1131 and U4358 U3237 ; U3483
g1132 and STATE_REG_0__SCAN_IN REQUESTPENDING_REG_SCAN_IN ; U3484
g1133 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3485
g1134 and INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3486
g1135 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3487
g1136 and INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3488
g1137 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3489
g1138 and INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3490
g1139 nor INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3491
g1140 and INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3492
g1141 nor INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3493
g1142 and INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3494
g1143 and INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3495
g1144 and U4374 U4373 U4372 U4371 ; U3496
g1145 and U4378 U4377 U4376 U4375 ; U3497
g1146 and U4382 U4381 U4380 U4379 ; U3498
g1147 and U4386 U4385 U4384 U4383 ; U3499
g1148 and U4424 U4423 U4422 U4421 ; U3500
g1149 and U4428 U4427 U4426 U4425 ; U3501
g1150 and U4432 U4431 U4430 U4429 ; U3502
g1151 and U4436 U4435 U4434 U4433 ; U3503
g1152 and U4407 U4406 U4405 U4404 ; U3504
g1153 and U4411 U4410 U4409 U4408 ; U3505
g1154 and U4415 U4414 U4413 U4412 ; U3506
g1155 and U4419 U4418 U4417 U4416 ; U3507
g1156 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3508
g1157 and INSTQUEUE_REG_5__5__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3509
g1158 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3510
g1159 and INSTQUEUE_REG_6__5__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3511
g1160 and INSTQUEUE_REG_8__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3512
g1161 nor INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3513
g1162 and INSTQUEUE_REG_10__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3514
g1163 and INSTQUEUE_REG_12__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3515
g1164 nor INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3516
g1165 and INSTQUEUE_REG_9__5__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3517
g1166 and U4392 U4391 U4390 U4389 ; U3518
g1167 and U4396 U4395 U4394 U4393 ; U3519
g1168 and U4400 U4399 U4398 U4397 ; U3520
g1169 and U4402 U4401 ; U3521
g1170 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3522
g1171 and INSTQUEUE_REG_3__6__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3523
g1172 and U4441 U4440 U4439 U4438 ; U3524
g1173 and U4443 U4442 U4444 ; U3525
g1174 and U4446 U4445 U4447 ; U3526
g1175 and U7666 U7665 U7664 U7663 ; U3527
g1176 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3528
g1177 and INSTQUEUE_REG_1__4__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3529
g1178 nor INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3530
g1179 and INSTQUEUE_REG_4__4__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3531
g1180 nor INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3532
g1181 and INSTQUEUE_REG_12__4__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3533
g1182 and INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3534
g1183 and INSTQUEUE_REG_13__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3535
g1184 nor INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U3536
g1185 and INSTQUEUE_REG_6__4__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U3537
g1186 and INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3538
g1187 and INSTQUEUE_REG_14__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3539
g1188 nor INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U3540
g1189 and INSTQUEUE_REG_9__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U3541
g1190 and U7646 U7645 U7644 U7643 ; U3542
g1191 and U7650 U7649 U7648 U7647 ; U3543
g1192 and U7654 U7653 U7652 U7651 ; U3544
g1193 and U7658 U7657 U7656 U7655 ; U3545
g1194 and U3378 U3270 U7482 ; U3546
g1195 and U4448 U2605 U4388 ; U3547
g1196 and U4469 U4468 U4467 U4466 ; U3548
g1197 and U4473 U4472 U4471 U4470 ; U3549
g1198 and U4477 U4476 U4475 U4474 ; U3550
g1199 and U4481 U4480 U4479 U4478 ; U3551
g1200 and U4452 U4451 U4450 U4449 ; U3552
g1201 and U4456 U4455 U4454 U4453 ; U3553
g1202 and U4460 U4459 U4458 U4457 ; U3554
g1203 and U4464 U4463 U4462 U4461 ; U3555
g1204 and U4365 U4196 ; U3556
g1205 and U4407 U4406 U4405 U4404 ; U3557
g1206 and U4411 U4410 U4409 U4408 ; U3558
g1207 and U4415 U4414 U4413 U4412 ; U3559
g1208 and U4419 U4418 U4417 U4416 ; U3560
g1209 and U4392 U4391 U4390 U4389 ; U3561
g1210 and U4396 U4395 U4394 U4393 ; U3562
g1211 and U4400 U4399 U4398 U4397 ; U3563
g1212 and U4402 U4401 ; U3564
g1213 and U4387 U4159 ; U3565
g1214 and U4237 U3270 ; U3566
g1215 and U3271 U3270 U4388 U7482 ; U3567
g1216 and U4205 U3387 ; U3568
g1217 and U7591 STATE2_REG_2__SCAN_IN ; U3569
g1218 and U4503 U3284 ; U3570
g1219 and U2427 U3244 ; U3571
g1220 and STATE2_REG_3__SCAN_IN STATE2_REG_0__SCAN_IN ; U3572
g1221 and U4234 U4229 ; U3573
g1222 and U3573 U4511 ; U3574
g1223 and U4540 U4541 U4212 ; U3575
g1224 and U4549 U4548 U4550 ; U3576
g1225 and U4554 U4553 U4555 ; U3577
g1226 and U4559 U4558 U4560 ; U3578
g1227 and U4564 U4563 U4565 ; U3579
g1228 and U4569 U4568 U4570 ; U3580
g1229 and U4574 U4573 U4575 ; U3581
g1230 and U4579 U4578 U4580 ; U3582
g1231 and U4584 U4583 U4585 ; U3583
g1232 and U4598 U4599 U4212 ; U3584
g1233 and U4607 U4606 U4608 ; U3585
g1234 and U4612 U4611 U4613 ; U3586
g1235 and U4617 U4616 U4618 ; U3587
g1236 and U4622 U4621 U4623 ; U3588
g1237 and U4627 U4626 U4628 ; U3589
g1238 and U4632 U4631 U4633 ; U3590
g1239 and U4637 U4636 U4638 ; U3591
g1240 and U4642 U4641 U4643 ; U3592
g1241 and U4657 U4658 U4212 ; U3593
g1242 and U4666 U4665 U4667 ; U3594
g1243 and U4671 U4670 U4672 ; U3595
g1244 and U4676 U4675 U4677 ; U3596
g1245 and U4681 U4680 U4682 ; U3597
g1246 and U4686 U4685 U4687 ; U3598
g1247 and U4691 U4690 U4692 ; U3599
g1248 and U4696 U4695 U4697 ; U3600
g1249 and U4701 U4700 U4702 ; U3601
g1250 and U4714 U4715 U4212 ; U3602
g1251 and U4723 U4722 U4724 ; U3603
g1252 and U4728 U4727 U4729 ; U3604
g1253 and U4733 U4732 U4734 ; U3605
g1254 and U4738 U4737 U4739 ; U3606
g1255 and U4743 U4742 U4744 ; U3607
g1256 and U4748 U4747 U4749 ; U3608
g1257 and U4753 U4752 U4754 ; U3609
g1258 and U4758 U4757 U4759 ; U3610
g1259 and U4772 U4773 U4212 ; U3611
g1260 and U4781 U4780 U4782 ; U3612
g1261 and U4786 U4785 U4787 ; U3613
g1262 and U4791 U4790 U4792 ; U3614
g1263 and U4796 U4795 U4797 ; U3615
g1264 and U4801 U4800 U4802 ; U3616
g1265 and U4806 U4805 U4807 ; U3617
g1266 and U4811 U4810 U4812 ; U3618
g1267 and U4816 U4815 U4817 ; U3619
g1268 and U4829 U4830 U4212 ; U3620
g1269 and U4838 U4837 U4839 ; U3621
g1270 and U4843 U4842 U4844 ; U3622
g1271 and U4848 U4847 U4849 ; U3623
g1272 and U4853 U4852 U4854 ; U3624
g1273 and U4858 U4857 U4859 ; U3625
g1274 and U4863 U4862 U4864 ; U3626
g1275 and U4868 U4867 U4869 ; U3627
g1276 and U4873 U4872 U4874 ; U3628
g1277 and U4887 U4888 U4212 ; U3629
g1278 and U4896 U4895 U4897 ; U3630
g1279 and U4901 U4900 U4902 ; U3631
g1280 and U4906 U4905 U4907 ; U3632
g1281 and U4911 U4910 U4912 ; U3633
g1282 and U4916 U4915 U4917 ; U3634
g1283 and U4921 U4920 U4922 ; U3635
g1284 and U4926 U4925 U4927 ; U3636
g1285 and U4931 U4930 U4932 ; U3637
g1286 and U4944 U4945 U4212 ; U3638
g1287 and U4953 U4952 U4954 ; U3639
g1288 and U4958 U4957 U4959 ; U3640
g1289 and U4963 U4962 U4964 ; U3641
g1290 and U4968 U4967 U4969 ; U3642
g1291 and U4973 U4972 U4974 ; U3643
g1292 and U4978 U4977 U4979 ; U3644
g1293 and U4983 U4982 U4984 ; U3645
g1294 and U4988 U4987 U4989 ; U3646
g1295 and U5000 U5001 U4212 ; U3647
g1296 and U5009 U5008 U5010 ; U3648
g1297 and U5014 U5013 U5015 ; U3649
g1298 and U5019 U5018 U5020 ; U3650
g1299 and U5024 U5023 U5025 ; U3651
g1300 and U5029 U5028 U5030 ; U3652
g1301 and U5034 U5033 U5035 ; U3653
g1302 and U5039 U5038 U5040 ; U3654
g1303 and U5044 U5043 U5045 ; U3655
g1304 and U5057 U5058 U4212 ; U3656
g1305 and U5066 U5065 U5067 ; U3657
g1306 and U5071 U5070 U5072 ; U3658
g1307 and U5076 U5075 U5077 ; U3659
g1308 and U5081 U5080 U5082 ; U3660
g1309 and U5086 U5085 U5087 ; U3661
g1310 and U5091 U5090 U5092 ; U3662
g1311 and U5096 U5095 U5097 ; U3663
g1312 and U5101 U5100 U5102 ; U3664
g1313 and U5115 U5116 U4212 ; U3665
g1314 and U5124 U5123 U5125 ; U3666
g1315 and U5129 U5128 U5130 ; U3667
g1316 and U5134 U5133 U5135 ; U3668
g1317 and U5139 U5138 U5140 ; U3669
g1318 and U5144 U5143 U5145 ; U3670
g1319 and U5149 U5148 U5150 ; U3671
g1320 and U5154 U5153 U5155 ; U3672
g1321 and U5159 U5158 U5160 ; U3673
g1322 and U5172 U5173 U4212 ; U3674
g1323 and U5181 U5180 U5182 ; U3675
g1324 and U5186 U5185 U5187 ; U3676
g1325 and U5191 U5190 U5192 ; U3677
g1326 and U5196 U5195 U5197 ; U3678
g1327 and U5201 U5200 U5202 ; U3679
g1328 and U5206 U5205 U5207 ; U3680
g1329 and U5211 U5210 U5212 ; U3681
g1330 and U5216 U5215 U5217 ; U3682
g1331 and U5230 U5231 U4212 ; U3683
g1332 and U5239 U5238 U5240 ; U3684
g1333 and U5244 U5243 U5245 ; U3685
g1334 and U5249 U5248 U5250 ; U3686
g1335 and U5254 U5253 U5255 ; U3687
g1336 and U5259 U5258 U5260 ; U3688
g1337 and U5264 U5263 U5265 ; U3689
g1338 and U5269 U5268 U5270 ; U3690
g1339 and U5274 U5273 U5275 ; U3691
g1340 and U5287 U5288 U4212 ; U3692
g1341 and U5296 U5295 U5297 ; U3693
g1342 and U5301 U5300 U5302 ; U3694
g1343 and U5306 U5305 U5307 ; U3695
g1344 and U5311 U5310 U5312 ; U3696
g1345 and U5316 U5315 U5317 ; U3697
g1346 and U5321 U5320 U5322 ; U3698
g1347 and U5326 U5325 U5327 ; U3699
g1348 and U5331 U5330 U5332 ; U3700
g1349 and U5345 U5346 U4212 ; U3701
g1350 and U5354 U5353 U5355 ; U3702
g1351 and U5359 U5358 U5360 ; U3703
g1352 and U5364 U5363 U5365 ; U3704
g1353 and U5369 U5368 U5370 ; U3705
g1354 and U5374 U5373 U5375 ; U3706
g1355 and U5379 U5378 U5380 ; U3707
g1356 and U5384 U5383 U5385 ; U3708
g1357 and U5389 U5388 U5390 ; U3709
g1358 and U5402 U5403 U4212 ; U3710
g1359 and U5411 U5410 U5412 ; U3711
g1360 and U5416 U5415 U5417 ; U3712
g1361 and U5421 U5420 U5422 ; U3713
g1362 and U5426 U5425 U5427 ; U3714
g1363 and U5430 U5429 U5431 ; U3715
g1364 and U5435 U5434 U5436 ; U3716
g1365 and U5440 U5439 U5441 ; U3717
g1366 and U5445 U5444 U5446 ; U3718
g1367 and STATE2_REG_0__SCAN_IN FLUSH_REG_SCAN_IN ; U3719
g1368 and U4482 U4387 ; U3720
g1369 and U4485 U3244 ; U3721
g1370 and U4198 U3244 ; U3722
g1371 and U7484 U4205 ; U3723
g1372 and U5459 U5460 ; U3724
g1373 and U3724 U5458 ; U3725
g1374 and U3725 U2518 ; U3726
g1375 and U5463 U4230 ; U3727
g1376 and U5474 U5473 ; U3728
g1377 and U4437 U4388 ; U3729
g1378 and U5484 U3380 ; U3730
g1379 and U5486 U5485 ; U3731
g1380 and U5488 U7615 U3730 U3731 ; U3732
g1381 and U4251 U3384 ; U3733
g1382 and U3398 U3275 U3733 U2520 U3266 ; U3734
g1383 and U3736 U5490 ; U3735
g1384 and U5493 U5492 ; U3736
g1385 and U7705 U7704 U5501 ; U3737
g1386 and U5512 U5510 ; U3738
g1387 and U5531 U5532 ; U3739
g1388 and U5535 U5536 ; U3740
g1389 and U5540 U5541 ; U3741
g1390 and U5546 U3244 ; U3742
g1391 and U3271 U3394 ; U3743
g1392 and U5551 U5549 ; U3744
g1393 and U3385 U3386 U5555 ; U3745
g1394 and U2520 U5556 U3745 ; U3746
g1395 and U4174 U3271 ; U3747
g1396 and U3275 U4205 U3435 ; U3748
g1397 and U5554 U7495 ; U3749
g1398 and U7496 STATE2_REG_2__SCAN_IN ; U3750
g1399 and U5559 U5558 ; U3751
g1400 and U5561 U5560 ; U3752
g1401 and U5563 U5564 ; U3753
g1402 and U3753 U5562 ; U3754
g1403 and U5566 U5565 ; U3755
g1404 and U5568 U5567 ; U3756
g1405 and U5570 U5571 ; U3757
g1406 and U3757 U5569 ; U3758
g1407 and U5573 U5572 ; U3759
g1408 and U5575 U5574 ; U3760
g1409 and U5577 U5578 ; U3761
g1410 and U3761 U5576 ; U3762
g1411 and U5580 U5579 U5582 ; U3763
g1412 and U3765 U5583 U5581 ; U3764
g1413 and U5584 U5585 ; U3765
g1414 and U5587 U5586 U5589 ; U3766
g1415 and U5591 U5592 ; U3767
g1416 and U3767 U5590 ; U3768
g1417 and U5594 U5593 U5596 ; U3769
g1418 and U5598 U5599 ; U3770
g1419 and U3770 U5597 ; U3771
g1420 and U5601 U5600 U5603 ; U3772
g1421 and U5605 U5606 ; U3773
g1422 and U3773 U5604 ; U3774
g1423 and U5608 U5607 U5610 ; U3775
g1424 and U5612 U5613 ; U3776
g1425 and U3776 U5611 ; U3777
g1426 and U5615 U5614 U5617 ; U3778
g1427 and U5619 U5620 ; U3779
g1428 and U3779 U5618 ; U3780
g1429 and U5622 U5621 U5624 ; U3781
g1430 and U5626 U5627 ; U3782
g1431 and U3782 U5625 ; U3783
g1432 and U5629 U5628 U5631 ; U3784
g1433 and U5633 U5634 ; U3785
g1434 and U3785 U5632 ; U3786
g1435 and U5636 U5635 U5638 ; U3787
g1436 and U5640 U5641 ; U3788
g1437 and U3788 U5639 ; U3789
g1438 and U5643 U5642 U5645 ; U3790
g1439 and U5647 U5648 ; U3791
g1440 and U3791 U5646 ; U3792
g1441 and U5650 U5652 ; U3793
g1442 and U5654 U5655 ; U3794
g1443 and U3794 U5653 ; U3795
g1444 and U5657 U5659 ; U3796
g1445 and U5661 U5662 ; U3797
g1446 and U3797 U5660 ; U3798
g1447 and U5664 U5666 ; U3799
g1448 and U5668 U5669 ; U3800
g1449 and U3800 U5667 ; U3801
g1450 and U5671 U5673 ; U3802
g1451 and U5675 U5676 ; U3803
g1452 and U3803 U5674 ; U3804
g1453 and U5678 U5680 ; U3805
g1454 and U5682 U5683 ; U3806
g1455 and U3806 U5681 ; U3807
g1456 and U5685 U5687 ; U3808
g1457 and U5689 U5690 ; U3809
g1458 and U3809 U5688 ; U3810
g1459 and U5692 U5694 ; U3811
g1460 and U5696 U5697 ; U3812
g1461 and U3812 U5695 ; U3813
g1462 and U5699 U5701 ; U3814
g1463 and U5703 U5704 ; U3815
g1464 and U3815 U5702 ; U3816
g1465 and U5706 U5708 ; U3817
g1466 and U5710 U5711 ; U3818
g1467 and U3818 U5709 ; U3819
g1468 and U5713 U5715 ; U3820
g1469 and U5717 U5718 ; U3821
g1470 and U3821 U5716 ; U3822
g1471 and U5720 U5722 ; U3823
g1472 and U5724 U5725 ; U3824
g1473 and U3824 U5723 ; U3825
g1474 and U5727 U5729 ; U3826
g1475 and U5731 U5732 ; U3827
g1476 and U3827 U5730 ; U3828
g1477 and U5734 U5736 ; U3829
g1478 and U5738 U5739 ; U3830
g1479 and U3830 U5737 ; U3831
g1480 and U5741 U5743 ; U3832
g1481 and U5745 U5746 ; U3833
g1482 and U3833 U5744 ; U3834
g1483 and U5748 U5750 ; U3835
g1484 and U5752 U5753 ; U3836
g1485 and U3836 U5751 ; U3837
g1486 and U5755 U5757 ; U3838
g1487 and U5759 U5760 ; U3839
g1488 and U3839 U5758 ; U3840
g1489 and U5762 U5764 ; U3841
g1490 and U5766 U5767 ; U3842
g1491 and U3842 U5765 ; U3843
g1492 and U5769 U5771 ; U3844
g1493 and U5773 U5774 ; U3845
g1494 and U3845 U5772 ; U3846
g1495 and U5776 U5778 ; U3847
g1496 and U5780 U5781 ; U3848
g1497 and U3848 U5779 ; U3849
g1498 and U3270 U3249 U7482 ; U3850
g1499 and U5782 U3395 ; U3851
g1500 and STATE2_REG_1__SCAN_IN STATEBS16_REG_SCAN_IN ; U3852
g1501 and U2368 U3271 ; U3853
g1502 and U2449 STATE2_REG_0__SCAN_IN ; U3854
g1503 and U4196 U2368 ; U3855
g1504 and U6093 U6094 ; U3856
g1505 and U6096 U6097 ; U3857
g1506 and U6099 U6100 ; U3858
g1507 and U6102 U6103 ; U3859
g1508 and U6105 U6106 ; U3860
g1509 and U6108 U6109 ; U3861
g1510 and U6111 U6112 ; U3862
g1511 and U6114 U6115 ; U3863
g1512 and U6117 U6118 ; U3864
g1513 and U6120 U6121 ; U3865
g1514 and U6123 U6124 ; U3866
g1515 and U6126 U6127 ; U3867
g1516 and U6129 U6130 ; U3868
g1517 and U6132 U6133 ; U3869
g1518 and U6135 U6136 ; U3870
g1519 and U6139 U6138 ; U3871
g1520 and U2605 U3378 ; U3872
g1521 and U3258 U7482 STATE2_REG_0__SCAN_IN ; U3873
g1522 and U4387 U4159 ; U3874
g1523 and U4229 U4232 U6350 ; U3875
g1524 nor READY_N STATEBS16_REG_SCAN_IN ; U3876
g1525 and U4482 U4174 ; U3877
g1526 and U6361 U6360 U6363 U6362 U6359 ; U3878
g1527 and U6369 U6368 U6371 U6370 U6367 ; U3879
g1528 and U6377 U6376 U6379 U6378 U6375 ; U3880
g1529 and U6385 U6384 U6387 U6386 U6383 ; U3881
g1530 and U6388 U4215 ; U3882
g1531 and U6393 U6392 U6395 U6394 ; U3883
g1532 and U6396 U4215 ; U3884
g1533 and U6401 U6400 U6403 U6402 U6399 ; U3885
g1534 and U6404 U4215 ; U3886
g1535 and U6410 U6407 U6409 ; U3887
g1536 and U6411 U4215 ; U3888
g1537 and U6417 U6414 U6416 ; U3889
g1538 and U6418 U4215 ; U3890
g1539 and U6424 U6421 U6423 ; U3891
g1540 and U6425 U4215 ; U3892
g1541 and U6431 U6428 U6430 ; U3893
g1542 and U6432 U4215 ; U3894
g1543 and U6438 U6435 U6437 ; U3895
g1544 and U6439 U4215 ; U3896
g1545 and U6445 U6442 U6444 ; U3897
g1546 and U6446 U4215 ; U3898
g1547 and U6452 U6449 U6451 ; U3899
g1548 and U6453 U4215 ; U3900
g1549 and U6459 U6456 U6458 ; U3901
g1550 and U6460 U4215 ; U3902
g1551 and U6466 U6463 U6465 ; U3903
g1552 and U6467 U4215 ; U3904
g1553 and U6473 U6470 U6472 ; U3905
g1554 and U6474 U4215 ; U3906
g1555 and U6480 U6477 U6479 ; U3907
g1556 and U4215 U6482 ; U3908
g1557 and U6487 U6484 U6486 ; U3909
g1558 and U4215 U6489 ; U3910
g1559 and U6494 U6491 U6493 ; U3911
g1560 and U4215 U6496 ; U3912
g1561 and U6501 U6498 U6500 ; U3913
g1562 and U6505 U6503 ; U3914
g1563 and U6507 U6508 ; U3915
g1564 and U6512 U6510 ; U3916
g1565 and U6514 U6515 ; U3917
g1566 and U6519 U6517 ; U3918
g1567 and U6521 U6522 ; U3919
g1568 and U6526 U6524 ; U3920
g1569 and U6528 U6529 ; U3921
g1570 and U6533 U6531 ; U3922
g1571 and U6535 U6536 ; U3923
g1572 and U6540 U6538 ; U3924
g1573 and U6542 U6543 ; U3925
g1574 and U6547 U6545 ; U3926
g1575 and U6549 U6550 ; U3927
g1576 and U6554 U6552 ; U3928
g1577 and U6556 U6557 ; U3929
g1578 and U6561 U6559 ; U3930
g1579 and U6563 U6564 ; U3931
g1580 and U6568 U6566 ; U3932
g1581 and U6570 U6571 ; U3933
g1582 and U6575 U6573 ; U3934
g1583 and U6577 U6578 ; U3935
g1584 and U6582 U6580 ; U3936
g1585 and U6584 U6585 ; U3937
g1586 nor DATAWIDTH_REG_2__SCAN_IN DATAWIDTH_REG_3__SCAN_IN DATAWIDTH_REG_4__SCAN_IN DATAWIDTH_REG_5__SCAN_IN ; U3938
g1587 nor DATAWIDTH_REG_6__SCAN_IN DATAWIDTH_REG_7__SCAN_IN DATAWIDTH_REG_8__SCAN_IN DATAWIDTH_REG_9__SCAN_IN ; U3939
g1588 and U3939 U3938 ; U3940
g1589 nor DATAWIDTH_REG_10__SCAN_IN DATAWIDTH_REG_11__SCAN_IN DATAWIDTH_REG_12__SCAN_IN DATAWIDTH_REG_13__SCAN_IN ; U3941
g1590 nor DATAWIDTH_REG_14__SCAN_IN DATAWIDTH_REG_15__SCAN_IN DATAWIDTH_REG_16__SCAN_IN DATAWIDTH_REG_17__SCAN_IN ; U3942
g1591 and U3942 U3941 ; U3943
g1592 nor DATAWIDTH_REG_18__SCAN_IN DATAWIDTH_REG_19__SCAN_IN DATAWIDTH_REG_20__SCAN_IN DATAWIDTH_REG_21__SCAN_IN ; U3944
g1593 nor DATAWIDTH_REG_22__SCAN_IN DATAWIDTH_REG_23__SCAN_IN DATAWIDTH_REG_24__SCAN_IN DATAWIDTH_REG_25__SCAN_IN ; U3945
g1594 and U3945 U3944 ; U3946
g1595 nor DATAWIDTH_REG_26__SCAN_IN DATAWIDTH_REG_27__SCAN_IN ; U3947
g1596 nor DATAWIDTH_REG_28__SCAN_IN DATAWIDTH_REG_29__SCAN_IN ; U3948
g1597 nor DATAWIDTH_REG_30__SCAN_IN DATAWIDTH_REG_31__SCAN_IN ; U3949
g1598 and U3949 U6586 U3948 U3947 ; U3950
g1599 nor DATAWIDTH_REG_0__SCAN_IN DATAWIDTH_REG_1__SCAN_IN REIP_REG_0__SCAN_IN ; U3951
g1600 and U3244 STATE2_REG_2__SCAN_IN ; U3952
g1601 and U6596 U3285 ; U3953
g1602 nor READY_N STATE2_REG_0__SCAN_IN ; U3954
g1603 and U3294 U3395 U6590 ; U3955
g1604 and U3274 STATE2_REG_2__SCAN_IN ; U3956
g1605 and U4223 U4194 ; U3957
g1606 and U6609 U6608 U6607 U6606 ; U3958
g1607 and U6613 U6612 U6611 U6610 ; U3959
g1608 and U6617 U6616 U6615 U6614 ; U3960
g1609 and U6621 U6620 U6619 U6618 ; U3961
g1610 and U6625 U6624 U6623 U6622 ; U3962
g1611 and U6629 U6628 U6627 U6626 ; U3963
g1612 and U6633 U6632 U6631 U6630 ; U3964
g1613 and U6637 U6636 U6635 U6634 ; U3965
g1614 and U6641 U6640 U6639 U6638 ; U3966
g1615 and U6645 U6644 U6643 U6642 ; U3967
g1616 and U6649 U6648 U6647 U6646 ; U3968
g1617 and U6653 U6652 U6651 U6650 ; U3969
g1618 and U6657 U6656 U6655 U6654 ; U3970
g1619 and U6661 U6660 U6659 U6658 ; U3971
g1620 and U6665 U6664 U6663 U6662 ; U3972
g1621 and U7601 U6668 U6667 U6666 ; U3973
g1622 and U6672 U6671 U6670 U6669 ; U3974
g1623 and U6676 U6675 U6674 U6673 ; U3975
g1624 and U6680 U6679 U6678 U6677 ; U3976
g1625 and U6684 U6683 U6682 U6681 ; U3977
g1626 and U6688 U6687 U6686 U6685 ; U3978
g1627 and U6692 U6691 U6690 U6689 ; U3979
g1628 and U6696 U6695 U6694 U6693 ; U3980
g1629 and U6700 U6699 U6698 U6697 ; U3981
g1630 and U6704 U6703 U6702 U6701 ; U3982
g1631 and U6708 U6707 U6706 U6705 ; U3983
g1632 and U6712 U6711 U6710 U6709 ; U3984
g1633 and U6716 U6715 U6714 U6713 ; U3985
g1634 and U6720 U6719 U6718 U6717 ; U3986
g1635 and U6724 U6723 U6722 U6721 ; U3987
g1636 and U6728 U6727 U6726 U6725 ; U3988
g1637 and U6732 U6731 U6730 U6729 ; U3989
g1638 and U6737 U6736 ; U3990
g1639 and U6740 U6739 ; U3991
g1640 and U6743 U6742 ; U3992
g1641 and U6746 U6745 ; U3993
g1642 and U6748 U3995 ; U3994
g1643 and U6750 U6749 ; U3995
g1644 and U6752 U6753 ; U3996
g1645 and U6760 U6761 U6762 ; U3997
g1646 and U6764 U6765 ; U3998
g1647 and U6769 U6770 U6771 ; U3999
g1648 and U6773 U6774 U6775 ; U4000
g1649 and U6777 U6778 U6779 ; U4001
g1650 and U6781 U6782 U6783 ; U4002
g1651 and U6785 U6786 U6787 ; U4003
g1652 and U6789 U6790 U6791 ; U4004
g1653 and U6793 U6794 U6795 ; U4005
g1654 and U6797 U6798 U6799 ; U4006
g1655 and U6801 U6802 U6803 ; U4007
g1656 and U6805 U6806 U6807 ; U4008
g1657 and U6809 U6810 ; U4009
g1658 and U6814 U6815 U6816 ; U4010
g1659 and U6818 U6819 U6820 ; U4011
g1660 and U6822 U6823 U6824 ; U4012
g1661 and U6826 U6827 U6828 ; U4013
g1662 and U6846 U6845 ; U4014
g1663 and U6848 U6849 ; U4015
g1664 and U7482 U6876 U3270 ; U4016
g1665 and U6883 U6882 U6881 U6880 ; U4017
g1666 and U6887 U6886 U6885 U6884 ; U4018
g1667 and U6891 U6890 U6889 U6888 ; U4019
g1668 and U6895 U6894 U6893 U6892 ; U4020
g1669 and U6901 U6900 U6899 U6898 ; U4021
g1670 and U6905 U6904 U6903 U6902 ; U4022
g1671 and U6909 U6908 U6907 U6906 ; U4023
g1672 and U6913 U6912 U6911 U6910 ; U4024
g1673 and U6932 U6931 U6930 U6929 ; U4025
g1674 and U6936 U6935 U6934 U6933 ; U4026
g1675 and U6940 U6939 U6938 U6937 ; U4027
g1676 and U6944 U6943 U6942 U6941 ; U4028
g1677 and U6949 U6948 U6947 U6946 ; U4029
g1678 and U6953 U6952 U6951 U6950 ; U4030
g1679 and U6957 U6956 U6955 U6954 ; U4031
g1680 and U6961 U6960 U6959 U6958 ; U4032
g1681 and U6966 U6965 U6964 U6963 ; U4033
g1682 and U6970 U6969 U6968 U6967 ; U4034
g1683 and U6974 U6973 U6972 U6971 ; U4035
g1684 and U6978 U6977 U6976 U6975 ; U4036
g1685 and U6983 U6982 U6981 U6980 ; U4037
g1686 and U6987 U6986 U6985 U6984 ; U4038
g1687 and U6991 U6990 U6989 U6988 ; U4039
g1688 and U7602 U6994 U6993 U6992 ; U4040
g1689 and U6998 U6997 U6996 U6995 ; U4041
g1690 and U7002 U7001 U7000 U6999 ; U4042
g1691 and U7006 U7005 U7004 U7003 ; U4043
g1692 and U7010 U7009 U7008 U7007 ; U4044
g1693 and U7015 U7014 U7013 U7012 ; U4045
g1694 and U7019 U7018 U7017 U7016 ; U4046
g1695 and U7023 U7022 U7021 U7020 ; U4047
g1696 and U7027 U7026 U7025 U7024 ; U4048
g1697 and U7047 U3430 ; U4049
g1698 and U7050 STATE2_REG_0__SCAN_IN ; U4050
g1699 and U7057 U7056 U7055 U7054 ; U4051
g1700 and U7061 U7060 U7059 U7058 ; U4052
g1701 and U7065 U7064 U7063 U7062 ; U4053
g1702 and U7069 U7068 U7067 U7066 ; U4054
g1703 and U4244 STATE2_REG_0__SCAN_IN ; U4055
g1704 and U4393 U4392 U4391 U4389 ; U4056
g1705 and U4395 U4394 U4396 ; U4057
g1706 and U4400 U4399 U4398 U4397 ; U4058
g1707 and U4402 U4401 ; U4059
g1708 and U4388 U3378 ; U4060
g1709 and U3271 STATE2_REG_0__SCAN_IN ; U4061
g1710 and U7078 U7077 ; U4062
g1711 and U7460 U3421 U7461 ; U4063
g1712 and U7463 U7464 U7462 ; U4064
g1713 and U2606 U7465 U4064 ; U4065
g1714 and U7085 U7083 ; U4066
g1715 and U7089 U7088 U7087 U7086 ; U4067
g1716 and U7093 U7092 U7091 U7090 ; U4068
g1717 and U7097 U7096 U7095 U7094 ; U4069
g1718 and U7101 U7100 U7099 U7098 ; U4070
g1719 and U7106 U7105 U7104 U7103 ; U4071
g1720 and U7110 U7109 U7108 U7107 ; U4072
g1721 and U7114 U7113 U7112 U7111 ; U4073
g1722 and U7118 U7117 U7116 U7115 ; U4074
g1723 and U7123 U7122 U7121 U7120 ; U4075
g1724 and U7127 U7126 U7125 U7124 ; U4076
g1725 and U7131 U7130 U7129 U7128 ; U4077
g1726 and U7133 U7132 ; U4078
g1727 and U7605 U7134 U4078 ; U4079
g1728 and U7138 U7137 U7136 U7135 ; U4080
g1729 and U7142 U7141 U7140 U7139 ; U4081
g1730 and U7146 U7145 U7144 U7143 ; U4082
g1731 and U7150 U7149 U7148 U7147 ; U4083
g1732 and U7155 U7154 U7153 U7152 ; U4084
g1733 and U7159 U7158 U7157 U7156 ; U4085
g1734 and U7163 U7162 U7161 U7160 ; U4086
g1735 and U7167 U7166 U7165 U7164 ; U4087
g1736 and U7172 U7171 U7170 U7169 ; U4088
g1737 and U7176 U7175 U7174 U7173 ; U4089
g1738 and U7180 U7179 U7178 U7177 ; U4090
g1739 and U7184 U7183 U7182 U7181 ; U4091
g1740 and U7189 U7188 U7187 U7186 ; U4092
g1741 and U7193 U7192 U7191 U7190 ; U4093
g1742 and U7197 U7196 U7195 U7194 ; U4094
g1743 and U7201 U7200 U7199 U7198 ; U4095
g1744 and U7203 U3251 ; U4096
g1745 and U7204 U7203 ; U4097
g1746 and U7205 U3252 ; U4098
g1747 and U7077 U3414 ; U4099
g1748 and U7206 U7205 ; U4100
g1749 and U4100 U7460 U7461 ; U4101
g1750 and U7078 U3421 U4099 U4101 ; U4102
g1751 and U7474 U7468 U7464 U7462 ; U4103
g1752 and U7493 U7477 U7476 U7475 ; U4104
g1753 and U7078 U7077 ; U4105
g1754 and U7460 U3421 U7461 ; U4106
g1755 and U7463 U7464 U7462 ; U4107
g1756 and U2608 U7465 U2606 U4107 ; U4108
g1757 and U7211 U7210 U7209 U7208 ; U4109
g1758 and U7215 U7214 U7213 U7212 ; U4110
g1759 and U7219 U7218 U7217 U7216 ; U4111
g1760 and U7223 U7222 U7221 U7220 ; U4112
g1761 and U7228 U7227 U7226 U7225 ; U4113
g1762 and U7232 U7231 U7230 U7229 ; U4114
g1763 and U7236 U7235 U7234 U7233 ; U4115
g1764 and U7240 U7239 U7238 U7237 ; U4116
g1765 and U7245 U7244 U7243 U7242 ; U4117
g1766 and U7249 U7248 U7247 U7246 ; U4118
g1767 and U7253 U7252 U7251 U7250 ; U4119
g1768 and U7257 U7256 U7255 U7254 ; U4120
g1769 and U7262 U7261 U7260 U7259 ; U4121
g1770 and U7266 U7265 U7264 U7263 ; U4122
g1771 and U7270 U7269 U7268 U7267 ; U4123
g1772 and U7607 U7273 U7272 U7271 ; U4124
g1773 and U7277 U7276 U7275 U7274 ; U4125
g1774 and U7281 U7280 U7279 U7278 ; U4126
g1775 and U7285 U7284 U7283 U7282 ; U4127
g1776 and U7289 U7288 U7287 U7286 ; U4128
g1777 and U7294 U7293 U7292 U7291 ; U4129
g1778 and U7298 U7297 U7296 U7295 ; U4130
g1779 and U7302 U7301 U7300 U7299 ; U4131
g1780 and U7306 U7305 U7304 U7303 ; U4132
g1781 and U7311 U7310 U7309 U7308 ; U4133
g1782 and U7315 U7314 U7313 U7312 ; U4134
g1783 and U7319 U7318 U7317 U7316 ; U4135
g1784 and U7323 U7322 U7321 U7320 ; U4136
g1785 and U7328 U7327 U7326 U7325 ; U4137
g1786 and U7332 U7331 U7330 U7329 ; U4138
g1787 and U7336 U7335 U7334 U7333 ; U4139
g1788 and U7340 U7339 U7338 U7337 ; U4140
g1789 and U3271 U3406 ; U4141
g1790 and U3270 U3378 ; U4142
g1791 and U7345 U7346 U4251 ; U4143
g1792 and U4143 U7347 ; U4144
g1793 and U2427 STATE2_REG_0__SCAN_IN ; U4145
g1794 and U4145 U7348 ; U4146
g1795 and U3258 U4161 ; U4147
g1796 and U4161 STATE2_REG_0__SCAN_IN ; U4148
g1797 and U7357 STATE2_REG_0__SCAN_IN ; U4149
g1798 and U7359 U2603 ; U4150
g1799 and U7361 STATE2_REG_0__SCAN_IN ; U4151
g1800 and U7363 U2603 ; U4152
g1801 and U7370 U7371 ; U4153
g1802 and U3440 U7372 ; U4154
g1803 and U7377 U7376 U7375 ; U4155
g1804 and U7450 U7449 ; U4156
g1805 and U7453 U7452 ; U4157
g1806 and U7662 U7661 ; U4158
g1807 nand U3560 U3559 U3558 U3557 ; U4159
g1808 nand U3727 U5462 ; U4160
g1809 nand U3564 U2607 U3563 U3562 U3561 ; U4161
g1810 not INSTADDRPOINTER_REG_31__SCAN_IN ; U4162
g1811 and U7714 U7713 ; U4163
g1812 and U7733 U7732 ; U4164
g1813 nand U2368 U3272 ; U4165
g1814 nand U4496 U3378 ; U4166
g1815 not BS16_N ; U4167
g1816 nand U3955 U4216 ; U4168
g1817 nand U4216 U3419 ; U4169
g1818 nand U7686 U7685 U3726 ; U4170
g1819 nand U3256 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U4171
g1820 not U3439 ; U4172
g1821 nand HOLD U3244 ; U4173
g1822 not U3399 ; U4174
g1823 not U3427 ; U4175
g1824 not U3426 ; U4176
g1825 not U3380 ; U4177
g1826 not U3277 ; U4178
g1827 not U3436 ; U4179
g1828 not U3392 ; U4180
g1829 not U3421 ; U4181
g1830 not U3407 ; U4182
g1831 nand U4253 U3258 ; U4183
g1832 nand U4448 U2605 ; U4184
g1833 not U3383 ; U4185
g1834 not U3412 ; U4186
g1835 not U3276 ; U4187
g1836 not U3408 ; U4188
g1837 not U3409 ; U4189
g1838 not U3415 ; U4190
g1839 not U3395 ; U4191
g1840 not U3414 ; U4192
g1841 nand U3873 U4177 U4185 ; U4193
g1842 not U3405 ; U4194
g1843 not U3430 ; U4195
g1844 not U3269 ; U4196
g1845 not U3294 ; U4197
g1846 not U3377 ; U4198
g1847 not U3433 ; U4199
g1848 not U3434 ; U4200
g1849 not U3435 ; U4201
g1850 not U3387 ; U4202
g1851 not U3275 ; U4203
g1852 not U3279 ; U4204
g1853 nand U3566 U2431 ; U4205
g1854 not U3386 ; U4206
g1855 nand U4437 U3258 ; U4207
g1856 not U3420 ; U4208
g1857 not U3236 ; U4209
g1858 not U3413 ; U4210
g1859 not U3411 ; U4211
g1860 not U3287 ; U4212
g1861 not LT_563_1260_U6 ; U4213
g1862 not U3307 ; U4214
g1863 nand U4243 U3418 ; U4215
g1864 nand U4223 U7488 ; U4216
g1865 nand U2362 U3259 ; U4217
g1866 nand U2363 U4365 ; U4218
g1867 not U3394 ; U4219
g1868 not U3239 ; U4220
g1869 not U3237 ; U4221
g1870 not U3382 ; U4222
g1871 not U3284 ; U4223
g1872 not U3385 ; U4224
g1873 not U4166 ; U4225
g1874 not U3344 ; U4226
g1875 nand U4465 U7369 ; U4227
g1876 nand U3951 U4208 ; U4228
g1877 nand U3572 U4249 ; U4229
g1878 nand U3719 U2428 ; U4230
g1879 nand U4352 U3245 ; U4231
g1880 nand U3281 U2352 STATE2_REG_1__SCAN_IN ; U4232
g1881 nand U2428 U3390 ; U4233
g1882 nand READY_N U3250 STATE2_REG_0__SCAN_IN ; U4234
g1883 not U3381 ; U4235
g1884 nand U2451 U2353 U3850 U2448 ; U4236
g1885 not U3274 ; U4237
g1886 not U3384 ; U4238
g1887 not U3402 ; U4239
g1888 not U3286 ; U4240
g1889 not U3396 ; U4241
g1890 not U3406 ; U4242
g1891 not U3419 ; U4243
g1892 not U3278 ; U4244
g1893 not U3376 ; U4245
g1894 not U3241 ; U4246
g1895 not U3268 ; U4247
g1896 not U3393 ; U4248
g1897 not U3285 ; U4249
g1898 not U3273 ; U4250
g1899 nand U4224 U4387 ; U4251
g1900 not U3398 ; U4252
g1901 not U3440 ; U4253
g1902 not U3397 ; U4254
g1903 nand U4221 REIP_REG_31__SCAN_IN ; U4255
g1904 nand U4220 REIP_REG_30__SCAN_IN ; U4256
g1905 nand U3236 ADDRESS_REG_29__SCAN_IN ; U4257
g1906 nand U4221 REIP_REG_30__SCAN_IN ; U4258
g1907 nand U4220 REIP_REG_29__SCAN_IN ; U4259
g1908 nand U3236 ADDRESS_REG_28__SCAN_IN ; U4260
g1909 nand U4221 REIP_REG_29__SCAN_IN ; U4261
g1910 nand U4220 REIP_REG_28__SCAN_IN ; U4262
g1911 nand U3236 ADDRESS_REG_27__SCAN_IN ; U4263
g1912 nand U4221 REIP_REG_28__SCAN_IN ; U4264
g1913 nand U4220 REIP_REG_27__SCAN_IN ; U4265
g1914 nand U3236 ADDRESS_REG_26__SCAN_IN ; U4266
g1915 nand U4221 REIP_REG_27__SCAN_IN ; U4267
g1916 nand U4220 REIP_REG_26__SCAN_IN ; U4268
g1917 nand U3236 ADDRESS_REG_25__SCAN_IN ; U4269
g1918 nand U4221 REIP_REG_26__SCAN_IN ; U4270
g1919 nand U4220 REIP_REG_25__SCAN_IN ; U4271
g1920 nand U3236 ADDRESS_REG_24__SCAN_IN ; U4272
g1921 nand U4221 REIP_REG_25__SCAN_IN ; U4273
g1922 nand U4220 REIP_REG_24__SCAN_IN ; U4274
g1923 nand U3236 ADDRESS_REG_23__SCAN_IN ; U4275
g1924 nand U4221 REIP_REG_24__SCAN_IN ; U4276
g1925 nand U4220 REIP_REG_23__SCAN_IN ; U4277
g1926 nand U3236 ADDRESS_REG_22__SCAN_IN ; U4278
g1927 nand U4221 REIP_REG_23__SCAN_IN ; U4279
g1928 nand U4220 REIP_REG_22__SCAN_IN ; U4280
g1929 nand U3236 ADDRESS_REG_21__SCAN_IN ; U4281
g1930 nand U4221 REIP_REG_22__SCAN_IN ; U4282
g1931 nand U4220 REIP_REG_21__SCAN_IN ; U4283
g1932 nand U3236 ADDRESS_REG_20__SCAN_IN ; U4284
g1933 nand U4221 REIP_REG_21__SCAN_IN ; U4285
g1934 nand U4220 REIP_REG_20__SCAN_IN ; U4286
g1935 nand U3236 ADDRESS_REG_19__SCAN_IN ; U4287
g1936 nand U4221 REIP_REG_20__SCAN_IN ; U4288
g1937 nand U4220 REIP_REG_19__SCAN_IN ; U4289
g1938 nand U3236 ADDRESS_REG_18__SCAN_IN ; U4290
g1939 nand U4221 REIP_REG_19__SCAN_IN ; U4291
g1940 nand U4220 REIP_REG_18__SCAN_IN ; U4292
g1941 nand U3236 ADDRESS_REG_17__SCAN_IN ; U4293
g1942 nand U4221 REIP_REG_18__SCAN_IN ; U4294
g1943 nand U4220 REIP_REG_17__SCAN_IN ; U4295
g1944 nand U3236 ADDRESS_REG_16__SCAN_IN ; U4296
g1945 nand U4221 REIP_REG_17__SCAN_IN ; U4297
g1946 nand U4220 REIP_REG_16__SCAN_IN ; U4298
g1947 nand U3236 ADDRESS_REG_15__SCAN_IN ; U4299
g1948 nand U4221 REIP_REG_16__SCAN_IN ; U4300
g1949 nand U4220 REIP_REG_15__SCAN_IN ; U4301
g1950 nand U3236 ADDRESS_REG_14__SCAN_IN ; U4302
g1951 nand U4221 REIP_REG_15__SCAN_IN ; U4303
g1952 nand U4220 REIP_REG_14__SCAN_IN ; U4304
g1953 nand U3236 ADDRESS_REG_13__SCAN_IN ; U4305
g1954 nand U4221 REIP_REG_14__SCAN_IN ; U4306
g1955 nand U4220 REIP_REG_13__SCAN_IN ; U4307
g1956 nand U3236 ADDRESS_REG_12__SCAN_IN ; U4308
g1957 nand U4221 REIP_REG_13__SCAN_IN ; U4309
g1958 nand U4220 REIP_REG_12__SCAN_IN ; U4310
g1959 nand U3236 ADDRESS_REG_11__SCAN_IN ; U4311
g1960 nand U4221 REIP_REG_12__SCAN_IN ; U4312
g1961 nand U4220 REIP_REG_11__SCAN_IN ; U4313
g1962 nand U3236 ADDRESS_REG_10__SCAN_IN ; U4314
g1963 nand U4221 REIP_REG_11__SCAN_IN ; U4315
g1964 nand U4220 REIP_REG_10__SCAN_IN ; U4316
g1965 nand U3236 ADDRESS_REG_9__SCAN_IN ; U4317
g1966 nand U4221 REIP_REG_10__SCAN_IN ; U4318
g1967 nand U4220 REIP_REG_9__SCAN_IN ; U4319
g1968 nand U3236 ADDRESS_REG_8__SCAN_IN ; U4320
g1969 nand U4221 REIP_REG_9__SCAN_IN ; U4321
g1970 nand U4220 REIP_REG_8__SCAN_IN ; U4322
g1971 nand U3236 ADDRESS_REG_7__SCAN_IN ; U4323
g1972 nand U4221 REIP_REG_8__SCAN_IN ; U4324
g1973 nand U4220 REIP_REG_7__SCAN_IN ; U4325
g1974 nand U3236 ADDRESS_REG_6__SCAN_IN ; U4326
g1975 nand U4221 REIP_REG_7__SCAN_IN ; U4327
g1976 nand U4220 REIP_REG_6__SCAN_IN ; U4328
g1977 nand U3236 ADDRESS_REG_5__SCAN_IN ; U4329
g1978 nand U4221 REIP_REG_6__SCAN_IN ; U4330
g1979 nand U4220 REIP_REG_5__SCAN_IN ; U4331
g1980 nand U3236 ADDRESS_REG_4__SCAN_IN ; U4332
g1981 nand U4221 REIP_REG_5__SCAN_IN ; U4333
g1982 nand U4220 REIP_REG_4__SCAN_IN ; U4334
g1983 nand U3236 ADDRESS_REG_3__SCAN_IN ; U4335
g1984 nand U4221 REIP_REG_4__SCAN_IN ; U4336
g1985 nand U4220 REIP_REG_3__SCAN_IN ; U4337
g1986 nand U3236 ADDRESS_REG_2__SCAN_IN ; U4338
g1987 nand U4221 REIP_REG_3__SCAN_IN ; U4339
g1988 nand U4220 REIP_REG_2__SCAN_IN ; U4340
g1989 nand U3236 ADDRESS_REG_1__SCAN_IN ; U4341
g1990 nand U4221 REIP_REG_2__SCAN_IN ; U4342
g1991 nand U4220 REIP_REG_1__SCAN_IN ; U4343
g1992 nand U3236 ADDRESS_REG_0__SCAN_IN ; U4344
g1993 not U3247 ; U4345
g1994 nand U4345 U3244 ; U4346
g1995 nand NA_N U4246 ; U4347
g1996 not U3248 ; U4348
g1997 nand U4348 U3244 ; U4349
g1998 or NA_N STATE_REG_0__SCAN_IN ; U4350
g1999 nand U7610 U4350 U7611 ; U4351
g2000 not U3242 ; U4352
g2001 nand HOLD U3234 U4352 ; U4353
g2002 nand U3481 U3248 ; U4354
g2003 nand U4354 U4353 ; U4355
g2004 nand U4347 U4355 STATE_REG_0__SCAN_IN ; U4356
g2005 nand U4351 STATE_REG_2__SCAN_IN ; U4357
g2006 nand READY_N U4209 ; U4358
g2007 nand U3484 U7613 ; U4359
g2008 nand U3247 STATE_REG_2__SCAN_IN ; U4360
g2009 nand NA_N U3245 ; U4361
g2010 nand U4361 U4360 ; U4362
g2011 nand U4362 U3235 ; U4363
g2012 nand U4167 U3242 ; U4364
g2013 not U3267 ; U4365
g2014 not U3256 ; U4366
g2015 not U3431 ; U4367
g2016 not U3255 ; U4368
g2017 not U3261 ; U4369
g2018 not U3254 ; U4370
g2019 nand U4370 INSTQUEUE_REG_7__3__SCAN_IN ; U4371
g2020 nand U2472 INSTQUEUE_REG_0__3__SCAN_IN ; U4372
g2021 nand U2471 INSTQUEUE_REG_1__3__SCAN_IN ; U4373
g2022 nand U2470 INSTQUEUE_REG_2__3__SCAN_IN ; U4374
g2023 nand U2468 INSTQUEUE_REG_3__3__SCAN_IN ; U4375
g2024 nand U2467 INSTQUEUE_REG_4__3__SCAN_IN ; U4376
g2025 nand U2466 INSTQUEUE_REG_5__3__SCAN_IN ; U4377
g2026 nand U2465 INSTQUEUE_REG_6__3__SCAN_IN ; U4378
g2027 nand U2464 INSTQUEUE_REG_8__3__SCAN_IN ; U4379
g2028 nand U2463 INSTQUEUE_REG_9__3__SCAN_IN ; U4380
g2029 nand U2461 INSTQUEUE_REG_10__3__SCAN_IN ; U4381
g2030 nand U2459 INSTQUEUE_REG_11__3__SCAN_IN ; U4382
g2031 nand U2458 INSTQUEUE_REG_12__3__SCAN_IN ; U4383
g2032 nand U2457 INSTQUEUE_REG_13__3__SCAN_IN ; U4384
g2033 nand U2455 INSTQUEUE_REG_14__3__SCAN_IN ; U4385
g2034 nand U2453 INSTQUEUE_REG_15__3__SCAN_IN ; U4386
g2035 not U3270 ; U4387
g2036 not U3265 ; U4388
g2037 nand U3257 INSTQUEUE_REG_7__5__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U4389
g2038 nand U3257 U4368 INSTQUEUE_REG_0__5__SCAN_IN ; U4390
g2039 nand U2469 U3252 INSTQUEUE_REG_1__5__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U4391
g2040 nand U2469 U3253 INSTQUEUE_REG_2__5__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U4392
g2041 nand U4366 U3257 INSTQUEUE_REG_4__5__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U4393
g2042 nand U3508 U3509 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U4394
g2043 nand U3510 U3511 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U4395
g2044 nand U3512 U4368 ; U4396
g2045 nand U3513 U3514 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U4397
g2046 nand U3251 INSTQUEUE_REG_11__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U4398
g2047 nand U4366 U3515 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U4399
g2048 nand U3252 INSTQUEUE_REG_13__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U4400
g2049 nand U3253 INSTQUEUE_REG_14__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U4401
g2050 nand INSTQUEUE_REG_15__5__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U4402
g2051 not U4161 ; U4403
g2052 nand U4370 INSTQUEUE_REG_7__2__SCAN_IN ; U4404
g2053 nand U2472 INSTQUEUE_REG_0__2__SCAN_IN ; U4405
g2054 nand U2471 INSTQUEUE_REG_1__2__SCAN_IN ; U4406
g2055 nand U2470 INSTQUEUE_REG_2__2__SCAN_IN ; U4407
g2056 nand U2468 INSTQUEUE_REG_3__2__SCAN_IN ; U4408
g2057 nand U2467 INSTQUEUE_REG_4__2__SCAN_IN ; U4409
g2058 nand U2466 INSTQUEUE_REG_5__2__SCAN_IN ; U4410
g2059 nand U2465 INSTQUEUE_REG_6__2__SCAN_IN ; U4411
g2060 nand U2464 INSTQUEUE_REG_8__2__SCAN_IN ; U4412
g2061 nand U2463 INSTQUEUE_REG_9__2__SCAN_IN ; U4413
g2062 nand U2461 INSTQUEUE_REG_10__2__SCAN_IN ; U4414
g2063 nand U2459 INSTQUEUE_REG_11__2__SCAN_IN ; U4415
g2064 nand U2458 INSTQUEUE_REG_12__2__SCAN_IN ; U4416
g2065 nand U2457 INSTQUEUE_REG_13__2__SCAN_IN ; U4417
g2066 nand U2455 INSTQUEUE_REG_14__2__SCAN_IN ; U4418
g2067 nand U2453 INSTQUEUE_REG_15__2__SCAN_IN ; U4419
g2068 not U4159 ; U4420
g2069 nand U4370 INSTQUEUE_REG_7__7__SCAN_IN ; U4421
g2070 nand U2472 INSTQUEUE_REG_0__7__SCAN_IN ; U4422
g2071 nand U2471 INSTQUEUE_REG_1__7__SCAN_IN ; U4423
g2072 nand U2470 INSTQUEUE_REG_2__7__SCAN_IN ; U4424
g2073 nand U2468 INSTQUEUE_REG_3__7__SCAN_IN ; U4425
g2074 nand U2467 INSTQUEUE_REG_4__7__SCAN_IN ; U4426
g2075 nand U2466 INSTQUEUE_REG_5__7__SCAN_IN ; U4427
g2076 nand U2465 INSTQUEUE_REG_6__7__SCAN_IN ; U4428
g2077 nand U2464 INSTQUEUE_REG_8__7__SCAN_IN ; U4429
g2078 nand U2463 INSTQUEUE_REG_9__7__SCAN_IN ; U4430
g2079 nand U2461 INSTQUEUE_REG_10__7__SCAN_IN ; U4431
g2080 nand U2459 INSTQUEUE_REG_11__7__SCAN_IN ; U4432
g2081 nand U2458 INSTQUEUE_REG_12__7__SCAN_IN ; U4433
g2082 nand U2457 INSTQUEUE_REG_13__7__SCAN_IN ; U4434
g2083 nand U2455 INSTQUEUE_REG_14__7__SCAN_IN ; U4435
g2084 nand U2453 INSTQUEUE_REG_15__7__SCAN_IN ; U4436
g2085 not U3378 ; U4437
g2086 nand U3486 U4369 INSTQUEUE_REG_7__6__SCAN_IN ; U4438
g2087 nand U2469 U2456 INSTQUEUE_REG_1__6__SCAN_IN ; U4439
g2088 nand U2469 U2454 INSTQUEUE_REG_2__6__SCAN_IN ; U4440
g2089 nand U4366 U4369 INSTQUEUE_REG_4__6__SCAN_IN ; U4441
g2090 nand U2456 U4369 INSTQUEUE_REG_5__6__SCAN_IN ; U4442
g2091 nand U2454 U4369 INSTQUEUE_REG_6__6__SCAN_IN ; U4443
g2092 nand U4366 U3495 INSTQUEUE_REG_12__6__SCAN_IN ; U4444
g2093 nand U3495 U2456 INSTQUEUE_REG_13__6__SCAN_IN ; U4445
g2094 nand U3495 U2454 INSTQUEUE_REG_14__6__SCAN_IN ; U4446
g2095 nand U3495 U3486 INSTQUEUE_REG_15__6__SCAN_IN ; U4447
g2096 not U3264 ; U4448
g2097 nand U4370 INSTQUEUE_REG_7__1__SCAN_IN ; U4449
g2098 nand U2472 INSTQUEUE_REG_0__1__SCAN_IN ; U4450
g2099 nand U2471 INSTQUEUE_REG_1__1__SCAN_IN ; U4451
g2100 nand U2470 INSTQUEUE_REG_2__1__SCAN_IN ; U4452
g2101 nand U2468 INSTQUEUE_REG_3__1__SCAN_IN ; U4453
g2102 nand U2467 INSTQUEUE_REG_4__1__SCAN_IN ; U4454
g2103 nand U2466 INSTQUEUE_REG_5__1__SCAN_IN ; U4455
g2104 nand U2465 INSTQUEUE_REG_6__1__SCAN_IN ; U4456
g2105 nand U2464 INSTQUEUE_REG_8__1__SCAN_IN ; U4457
g2106 nand U2463 INSTQUEUE_REG_9__1__SCAN_IN ; U4458
g2107 nand U2461 INSTQUEUE_REG_10__1__SCAN_IN ; U4459
g2108 nand U2459 INSTQUEUE_REG_11__1__SCAN_IN ; U4460
g2109 nand U2458 INSTQUEUE_REG_12__1__SCAN_IN ; U4461
g2110 nand U2457 INSTQUEUE_REG_13__1__SCAN_IN ; U4462
g2111 nand U2455 INSTQUEUE_REG_14__1__SCAN_IN ; U4463
g2112 nand U2453 INSTQUEUE_REG_15__1__SCAN_IN ; U4464
g2113 not U3258 ; U4465
g2114 nand U4370 INSTQUEUE_REG_7__0__SCAN_IN ; U4466
g2115 nand U2472 INSTQUEUE_REG_0__0__SCAN_IN ; U4467
g2116 nand U2471 INSTQUEUE_REG_1__0__SCAN_IN ; U4468
g2117 nand U2470 INSTQUEUE_REG_2__0__SCAN_IN ; U4469
g2118 nand U2468 INSTQUEUE_REG_3__0__SCAN_IN ; U4470
g2119 nand U2467 INSTQUEUE_REG_4__0__SCAN_IN ; U4471
g2120 nand U2466 INSTQUEUE_REG_5__0__SCAN_IN ; U4472
g2121 nand U2465 INSTQUEUE_REG_6__0__SCAN_IN ; U4473
g2122 nand U2464 INSTQUEUE_REG_8__0__SCAN_IN ; U4474
g2123 nand U2463 INSTQUEUE_REG_9__0__SCAN_IN ; U4475
g2124 nand U2461 INSTQUEUE_REG_10__0__SCAN_IN ; U4476
g2125 nand U2459 INSTQUEUE_REG_11__0__SCAN_IN ; U4477
g2126 nand U2458 INSTQUEUE_REG_12__0__SCAN_IN ; U4478
g2127 nand U2457 INSTQUEUE_REG_13__0__SCAN_IN ; U4479
g2128 nand U2455 INSTQUEUE_REG_14__0__SCAN_IN ; U4480
g2129 nand U2453 INSTQUEUE_REG_15__0__SCAN_IN ; U4481
g2130 not U3271 ; U4482
g2131 nand U3235 STATE_REG_2__SCAN_IN ; U4483
g2132 nand U3241 U4483 ; U4484
g2133 not U3259 ; U4485
g2134 nand U4465 U3375 ; U4486
g2135 not U3424 ; U4487
g2136 nand U3259 U3377 U3274 ; U4488
g2137 nand U4488 U3244 ; U4489
g2138 not U3272 ; U4490
g2139 nand U4448 U4161 ; U4491
g2140 nand U4184 U3273 ; U4492
g2141 nand U4492 U3567 ; U4493
g2142 nand U3568 U4493 ; U4494
g2143 nand U4203 U3375 ; U4495
g2144 nand U7670 U7669 U4495 ; U4496
g2145 nand U2448 U4250 ; U4497
g2146 or FLUSH_REG_SCAN_IN MORE_REG_SCAN_IN ; U4498
g2147 not U3280 ; U4499
g2148 nand U4499 U3249 ; U4500
g2149 nand READY_N STATE2_REG_1__SCAN_IN ; U4501
g2150 not U3282 ; U4502
g2151 nand U7676 U7675 STATE2_REG_1__SCAN_IN ; U4503
g2152 nand U3282 STATE2_REG_2__SCAN_IN ; U4504
g2153 nand U7592 U4234 ; U4505
g2154 nand U3571 U4502 ; U4506
g2155 nand U4505 STATE2_REG_1__SCAN_IN ; U4507
g2156 nand U2368 U7592 ; U4508
g2157 nand U4240 U4249 ; U4509
g2158 nand U7592 U4233 ; U4510
g2159 nand U2368 U3280 ; U4511
g2160 not U3312 ; U4512
g2161 not U3318 ; U4513
g2162 not U3319 ; U4514
g2163 not U3301 ; U4515
g2164 not U3300 ; U4516
g2165 not U3329 ; U4517
g2166 nand R2144_U8 U3300 ; U4518
g2167 not U3345 ; U4519
g2168 not U3302 ; U4520
g2169 not U3292 ; U4521
g2170 not U3293 ; U4522
g2171 nand U2438 U2442 ; U4523
g2172 not U3308 ; U4524
g2173 not U3343 ; U4525
g2174 not U3327 ; U4526
g2175 nand U3292 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; U4527
g2176 not U3347 ; U4528
g2177 not U3316 ; U4529
g2178 not U3310 ; U4530
g2179 not U3222 ; U4531
g2180 nand U2432 U2436 ; U4532
g2181 not U3309 ; U4533
g2182 nand U3250 STATE2_REG_1__SCAN_IN ; U4534
g2183 nand U4534 U3284 U3286 ; U4535
g2184 nand U4516 U2476 ; U4536
g2185 nand U2480 U2358 ; U4537
g2186 nand U3307 U4537 ; U4538
g2187 nand U4524 U4538 ; U4539
g2188 nand U3293 STATE2_REG_3__SCAN_IN ; U4540
g2189 nand U4533 STATE2_REG_2__SCAN_IN ; U4541
g2190 nand U4539 U3575 ; U4542
g2191 nand U2480 U2388 ; U4543
g2192 nand U3307 U4543 ; U4544
g2193 nand U4544 U3308 ; U4545
g2194 nand U3309 STATE2_REG_2__SCAN_IN ; U4546
g2195 nand U4546 U4545 ; U4547
g2196 nand U2415 U4522 ; U4548
g2197 nand U2413 U2477 ; U4549
g2198 nand U2412 U4520 ; U4550
g2199 nand U2397 U4547 ; U4551
g2200 nand U4542 INSTQUEUE_REG_15__7__SCAN_IN ; U4552
g2201 nand U2416 U4522 ; U4553
g2202 nand U2411 U2477 ; U4554
g2203 nand U2410 U4520 ; U4555
g2204 nand U2396 U4547 ; U4556
g2205 nand U4542 INSTQUEUE_REG_15__6__SCAN_IN ; U4557
g2206 nand U2420 U4522 ; U4558
g2207 nand U2409 U2477 ; U4559
g2208 nand U2408 U4520 ; U4560
g2209 nand U2395 U4547 ; U4561
g2210 nand U4542 INSTQUEUE_REG_15__5__SCAN_IN ; U4562
g2211 nand U2419 U4522 ; U4563
g2212 nand U2407 U2477 ; U4564
g2213 nand U2406 U4520 ; U4565
g2214 nand U2394 U4547 ; U4566
g2215 nand U4542 INSTQUEUE_REG_15__4__SCAN_IN ; U4567
g2216 nand U2418 U4522 ; U4568
g2217 nand U2405 U2477 ; U4569
g2218 nand U2404 U4520 ; U4570
g2219 nand U2393 U4547 ; U4571
g2220 nand U4542 INSTQUEUE_REG_15__3__SCAN_IN ; U4572
g2221 nand U2421 U4522 ; U4573
g2222 nand U2403 U2477 ; U4574
g2223 nand U2402 U4520 ; U4575
g2224 nand U2392 U4547 ; U4576
g2225 nand U4542 INSTQUEUE_REG_15__2__SCAN_IN ; U4577
g2226 nand U2414 U4522 ; U4578
g2227 nand U2401 U2477 ; U4579
g2228 nand U2400 U4520 ; U4580
g2229 nand U2391 U4547 ; U4581
g2230 nand U4542 INSTQUEUE_REG_15__1__SCAN_IN ; U4582
g2231 nand U2417 U4522 ; U4583
g2232 nand U2399 U2477 ; U4584
g2233 nand U2398 U4520 ; U4585
g2234 nand U2390 U4547 ; U4586
g2235 nand U4542 INSTQUEUE_REG_15__0__SCAN_IN ; U4587
g2236 not U3313 ; U4588
g2237 not U3314 ; U4589
g2238 not U3311 ; U4590
g2239 nand U2443 U2438 ; U4591
g2240 not U3315 ; U4592
g2241 not U3223 ; U4593
g2242 nand U4512 U2476 ; U4594
g2243 nand U2482 U2358 ; U4595
g2244 nand U3307 U4595 ; U4596
g2245 nand U4592 U4596 ; U4597
g2246 nand U3311 STATE2_REG_3__SCAN_IN ; U4598
g2247 nand U3223 STATE2_REG_2__SCAN_IN ; U4599
g2248 nand U4597 U3584 ; U4600
g2249 nand U2482 U2388 ; U4601
g2250 nand U3307 U4601 ; U4602
g2251 nand U4602 U3315 ; U4603
g2252 nand U4593 STATE2_REG_2__SCAN_IN ; U4604
g2253 nand U4604 U4603 ; U4605
g2254 nand U4590 U2415 ; U4606
g2255 nand U2481 U2413 ; U4607
g2256 nand U4589 U2412 ; U4608
g2257 nand U2397 U4605 ; U4609
g2258 nand U4600 INSTQUEUE_REG_14__7__SCAN_IN ; U4610
g2259 nand U4590 U2416 ; U4611
g2260 nand U2481 U2411 ; U4612
g2261 nand U4589 U2410 ; U4613
g2262 nand U2396 U4605 ; U4614
g2263 nand U4600 INSTQUEUE_REG_14__6__SCAN_IN ; U4615
g2264 nand U4590 U2420 ; U4616
g2265 nand U2481 U2409 ; U4617
g2266 nand U4589 U2408 ; U4618
g2267 nand U2395 U4605 ; U4619
g2268 nand U4600 INSTQUEUE_REG_14__5__SCAN_IN ; U4620
g2269 nand U4590 U2419 ; U4621
g2270 nand U2481 U2407 ; U4622
g2271 nand U4589 U2406 ; U4623
g2272 nand U2394 U4605 ; U4624
g2273 nand U4600 INSTQUEUE_REG_14__4__SCAN_IN ; U4625
g2274 nand U4590 U2418 ; U4626
g2275 nand U2481 U2405 ; U4627
g2276 nand U4589 U2404 ; U4628
g2277 nand U2393 U4605 ; U4629
g2278 nand U4600 INSTQUEUE_REG_14__3__SCAN_IN ; U4630
g2279 nand U4590 U2421 ; U4631
g2280 nand U2481 U2403 ; U4632
g2281 nand U4589 U2402 ; U4633
g2282 nand U2392 U4605 ; U4634
g2283 nand U4600 INSTQUEUE_REG_14__2__SCAN_IN ; U4635
g2284 nand U4590 U2414 ; U4636
g2285 nand U2481 U2401 ; U4637
g2286 nand U4589 U2400 ; U4638
g2287 nand U2391 U4605 ; U4639
g2288 nand U4600 INSTQUEUE_REG_14__1__SCAN_IN ; U4640
g2289 nand U4590 U2417 ; U4641
g2290 nand U2481 U2399 ; U4642
g2291 nand U4589 U2398 ; U4643
g2292 nand U2390 U4605 ; U4644
g2293 nand U4600 INSTQUEUE_REG_14__0__SCAN_IN ; U4645
g2294 not U3320 ; U4646
g2295 not U3321 ; U4647
g2296 not U3317 ; U4648
g2297 nand U2444 U2438 ; U4649
g2298 not U3322 ; U4650
g2299 nand U2437 U2432 ; U4651
g2300 not U3323 ; U4652
g2301 nand U4513 U2476 ; U4653
g2302 nand U2484 U2358 ; U4654
g2303 nand U3307 U4654 ; U4655
g2304 nand U4650 U4655 ; U4656
g2305 nand U3317 STATE2_REG_3__SCAN_IN ; U4657
g2306 nand U4652 STATE2_REG_2__SCAN_IN ; U4658
g2307 nand U4656 U3593 ; U4659
g2308 nand U2484 U2388 ; U4660
g2309 nand U3307 U4660 ; U4661
g2310 nand U4661 U3322 ; U4662
g2311 nand U3323 STATE2_REG_2__SCAN_IN ; U4663
g2312 nand U4663 U4662 ; U4664
g2313 nand U4648 U2415 ; U4665
g2314 nand U2483 U2413 ; U4666
g2315 nand U4647 U2412 ; U4667
g2316 nand U2397 U4664 ; U4668
g2317 nand U4659 INSTQUEUE_REG_13__7__SCAN_IN ; U4669
g2318 nand U4648 U2416 ; U4670
g2319 nand U2483 U2411 ; U4671
g2320 nand U4647 U2410 ; U4672
g2321 nand U2396 U4664 ; U4673
g2322 nand U4659 INSTQUEUE_REG_13__6__SCAN_IN ; U4674
g2323 nand U4648 U2420 ; U4675
g2324 nand U2483 U2409 ; U4676
g2325 nand U4647 U2408 ; U4677
g2326 nand U2395 U4664 ; U4678
g2327 nand U4659 INSTQUEUE_REG_13__5__SCAN_IN ; U4679
g2328 nand U4648 U2419 ; U4680
g2329 nand U2483 U2407 ; U4681
g2330 nand U4647 U2406 ; U4682
g2331 nand U2394 U4664 ; U4683
g2332 nand U4659 INSTQUEUE_REG_13__4__SCAN_IN ; U4684
g2333 nand U4648 U2418 ; U4685
g2334 nand U2483 U2405 ; U4686
g2335 nand U4647 U2404 ; U4687
g2336 nand U2393 U4664 ; U4688
g2337 nand U4659 INSTQUEUE_REG_13__3__SCAN_IN ; U4689
g2338 nand U4648 U2421 ; U4690
g2339 nand U2483 U2403 ; U4691
g2340 nand U4647 U2402 ; U4692
g2341 nand U2392 U4664 ; U4693
g2342 nand U4659 INSTQUEUE_REG_13__2__SCAN_IN ; U4694
g2343 nand U4648 U2414 ; U4695
g2344 nand U2483 U2401 ; U4696
g2345 nand U4647 U2400 ; U4697
g2346 nand U2391 U4664 ; U4698
g2347 nand U4659 INSTQUEUE_REG_13__1__SCAN_IN ; U4699
g2348 nand U4648 U2417 ; U4700
g2349 nand U2483 U2399 ; U4701
g2350 nand U4647 U2398 ; U4702
g2351 nand U2390 U4664 ; U4703
g2352 nand U4659 INSTQUEUE_REG_13__0__SCAN_IN ; U4704
g2353 not U3325 ; U4705
g2354 not U3324 ; U4706
g2355 nand U2445 U2438 ; U4707
g2356 not U3326 ; U4708
g2357 not U3224 ; U4709
g2358 nand U2486 U2476 ; U4710
g2359 nand U2489 U2358 ; U4711
g2360 nand U3307 U4711 ; U4712
g2361 nand U4708 U4712 ; U4713
g2362 nand U3324 STATE2_REG_3__SCAN_IN ; U4714
g2363 nand U3224 STATE2_REG_2__SCAN_IN ; U4715
g2364 nand U4713 U3602 ; U4716
g2365 nand U2489 U2388 ; U4717
g2366 nand U3307 U4717 ; U4718
g2367 nand U4718 U3326 ; U4719
g2368 nand U4709 STATE2_REG_2__SCAN_IN ; U4720
g2369 nand U4720 U4719 ; U4721
g2370 nand U4706 U2415 ; U4722
g2371 nand U2487 U2413 ; U4723
g2372 nand U4705 U2412 ; U4724
g2373 nand U2397 U4721 ; U4725
g2374 nand U4716 INSTQUEUE_REG_12__7__SCAN_IN ; U4726
g2375 nand U4706 U2416 ; U4727
g2376 nand U2487 U2411 ; U4728
g2377 nand U4705 U2410 ; U4729
g2378 nand U2396 U4721 ; U4730
g2379 nand U4716 INSTQUEUE_REG_12__6__SCAN_IN ; U4731
g2380 nand U4706 U2420 ; U4732
g2381 nand U2487 U2409 ; U4733
g2382 nand U4705 U2408 ; U4734
g2383 nand U2395 U4721 ; U4735
g2384 nand U4716 INSTQUEUE_REG_12__5__SCAN_IN ; U4736
g2385 nand U4706 U2419 ; U4737
g2386 nand U2487 U2407 ; U4738
g2387 nand U4705 U2406 ; U4739
g2388 nand U2394 U4721 ; U4740
g2389 nand U4716 INSTQUEUE_REG_12__4__SCAN_IN ; U4741
g2390 nand U4706 U2418 ; U4742
g2391 nand U2487 U2405 ; U4743
g2392 nand U4705 U2404 ; U4744
g2393 nand U2393 U4721 ; U4745
g2394 nand U4716 INSTQUEUE_REG_12__3__SCAN_IN ; U4746
g2395 nand U4706 U2421 ; U4747
g2396 nand U2487 U2403 ; U4748
g2397 nand U4705 U2402 ; U4749
g2398 nand U2392 U4721 ; U4750
g2399 nand U4716 INSTQUEUE_REG_12__2__SCAN_IN ; U4751
g2400 nand U4706 U2414 ; U4752
g2401 nand U2487 U2401 ; U4753
g2402 nand U4705 U2400 ; U4754
g2403 nand U2391 U4721 ; U4755
g2404 nand U4716 INSTQUEUE_REG_12__1__SCAN_IN ; U4756
g2405 nand U4706 U2417 ; U4757
g2406 nand U2487 U2399 ; U4758
g2407 nand U4705 U2398 ; U4759
g2408 nand U2390 U4721 ; U4760
g2409 nand U4716 INSTQUEUE_REG_12__0__SCAN_IN ; U4761
g2410 not U3330 ; U4762
g2411 not U3328 ; U4763
g2412 nand U2440 U2442 ; U4764
g2413 not U3331 ; U4765
g2414 nand U2434 U2436 ; U4766
g2415 not U3332 ; U4767
g2416 nand U4517 U4516 ; U4768
g2417 nand U2492 U2358 ; U4769
g2418 nand U3307 U4769 ; U4770
g2419 nand U4765 U4770 ; U4771
g2420 nand U3328 STATE2_REG_3__SCAN_IN ; U4772
g2421 nand U4767 STATE2_REG_2__SCAN_IN ; U4773
g2422 nand U4771 U3611 ; U4774
g2423 nand U2492 U2388 ; U4775
g2424 nand U3307 U4775 ; U4776
g2425 nand U4776 U3331 ; U4777
g2426 nand U3332 STATE2_REG_2__SCAN_IN ; U4778
g2427 nand U4778 U4777 ; U4779
g2428 nand U4763 U2415 ; U4780
g2429 nand U2491 U2413 ; U4781
g2430 nand U4762 U2412 ; U4782
g2431 nand U2397 U4779 ; U4783
g2432 nand U4774 INSTQUEUE_REG_11__7__SCAN_IN ; U4784
g2433 nand U4763 U2416 ; U4785
g2434 nand U2491 U2411 ; U4786
g2435 nand U4762 U2410 ; U4787
g2436 nand U2396 U4779 ; U4788
g2437 nand U4774 INSTQUEUE_REG_11__6__SCAN_IN ; U4789
g2438 nand U4763 U2420 ; U4790
g2439 nand U2491 U2409 ; U4791
g2440 nand U4762 U2408 ; U4792
g2441 nand U2395 U4779 ; U4793
g2442 nand U4774 INSTQUEUE_REG_11__5__SCAN_IN ; U4794
g2443 nand U4763 U2419 ; U4795
g2444 nand U2491 U2407 ; U4796
g2445 nand U4762 U2406 ; U4797
g2446 nand U2394 U4779 ; U4798
g2447 nand U4774 INSTQUEUE_REG_11__4__SCAN_IN ; U4799
g2448 nand U4763 U2418 ; U4800
g2449 nand U2491 U2405 ; U4801
g2450 nand U4762 U2404 ; U4802
g2451 nand U2393 U4779 ; U4803
g2452 nand U4774 INSTQUEUE_REG_11__3__SCAN_IN ; U4804
g2453 nand U4763 U2421 ; U4805
g2454 nand U2491 U2403 ; U4806
g2455 nand U4762 U2402 ; U4807
g2456 nand U2392 U4779 ; U4808
g2457 nand U4774 INSTQUEUE_REG_11__2__SCAN_IN ; U4809
g2458 nand U4763 U2414 ; U4810
g2459 nand U2491 U2401 ; U4811
g2460 nand U4762 U2400 ; U4812
g2461 nand U2391 U4779 ; U4813
g2462 nand U4774 INSTQUEUE_REG_11__1__SCAN_IN ; U4814
g2463 nand U4763 U2417 ; U4815
g2464 nand U2491 U2399 ; U4816
g2465 nand U4762 U2398 ; U4817
g2466 nand U2390 U4779 ; U4818
g2467 nand U4774 INSTQUEUE_REG_11__0__SCAN_IN ; U4819
g2468 not U3334 ; U4820
g2469 not U3333 ; U4821
g2470 nand U2440 U2443 ; U4822
g2471 not U3335 ; U4823
g2472 not U3225 ; U4824
g2473 nand U4517 U4512 ; U4825
g2474 nand U2494 U2358 ; U4826
g2475 nand U3307 U4826 ; U4827
g2476 nand U4823 U4827 ; U4828
g2477 nand U3333 STATE2_REG_3__SCAN_IN ; U4829
g2478 nand U3225 STATE2_REG_2__SCAN_IN ; U4830
g2479 nand U4828 U3620 ; U4831
g2480 nand U2494 U2388 ; U4832
g2481 nand U3307 U4832 ; U4833
g2482 nand U4833 U3335 ; U4834
g2483 nand U4824 STATE2_REG_2__SCAN_IN ; U4835
g2484 nand U4835 U4834 ; U4836
g2485 nand U4821 U2415 ; U4837
g2486 nand U2493 U2413 ; U4838
g2487 nand U4820 U2412 ; U4839
g2488 nand U2397 U4836 ; U4840
g2489 nand U4831 INSTQUEUE_REG_10__7__SCAN_IN ; U4841
g2490 nand U4821 U2416 ; U4842
g2491 nand U2493 U2411 ; U4843
g2492 nand U4820 U2410 ; U4844
g2493 nand U2396 U4836 ; U4845
g2494 nand U4831 INSTQUEUE_REG_10__6__SCAN_IN ; U4846
g2495 nand U4821 U2420 ; U4847
g2496 nand U2493 U2409 ; U4848
g2497 nand U4820 U2408 ; U4849
g2498 nand U2395 U4836 ; U4850
g2499 nand U4831 INSTQUEUE_REG_10__5__SCAN_IN ; U4851
g2500 nand U4821 U2419 ; U4852
g2501 nand U2493 U2407 ; U4853
g2502 nand U4820 U2406 ; U4854
g2503 nand U2394 U4836 ; U4855
g2504 nand U4831 INSTQUEUE_REG_10__4__SCAN_IN ; U4856
g2505 nand U4821 U2418 ; U4857
g2506 nand U2493 U2405 ; U4858
g2507 nand U4820 U2404 ; U4859
g2508 nand U2393 U4836 ; U4860
g2509 nand U4831 INSTQUEUE_REG_10__3__SCAN_IN ; U4861
g2510 nand U4821 U2421 ; U4862
g2511 nand U2493 U2403 ; U4863
g2512 nand U4820 U2402 ; U4864
g2513 nand U2392 U4836 ; U4865
g2514 nand U4831 INSTQUEUE_REG_10__2__SCAN_IN ; U4866
g2515 nand U4821 U2414 ; U4867
g2516 nand U2493 U2401 ; U4868
g2517 nand U4820 U2400 ; U4869
g2518 nand U2391 U4836 ; U4870
g2519 nand U4831 INSTQUEUE_REG_10__1__SCAN_IN ; U4871
g2520 nand U4821 U2417 ; U4872
g2521 nand U2493 U2399 ; U4873
g2522 nand U4820 U2398 ; U4874
g2523 nand U2390 U4836 ; U4875
g2524 nand U4831 INSTQUEUE_REG_10__0__SCAN_IN ; U4876
g2525 not U3337 ; U4877
g2526 not U3336 ; U4878
g2527 nand U2440 U2444 ; U4879
g2528 not U3338 ; U4880
g2529 nand U2434 U2437 ; U4881
g2530 not U3339 ; U4882
g2531 nand U4517 U4513 ; U4883
g2532 nand U2496 U2358 ; U4884
g2533 nand U3307 U4884 ; U4885
g2534 nand U4880 U4885 ; U4886
g2535 nand U3336 STATE2_REG_3__SCAN_IN ; U4887
g2536 nand U4882 STATE2_REG_2__SCAN_IN ; U4888
g2537 nand U4886 U3629 ; U4889
g2538 nand U2496 U2388 ; U4890
g2539 nand U3307 U4890 ; U4891
g2540 nand U4891 U3338 ; U4892
g2541 nand U3339 STATE2_REG_2__SCAN_IN ; U4893
g2542 nand U4893 U4892 ; U4894
g2543 nand U4878 U2415 ; U4895
g2544 nand U2495 U2413 ; U4896
g2545 nand U4877 U2412 ; U4897
g2546 nand U2397 U4894 ; U4898
g2547 nand U4889 INSTQUEUE_REG_9__7__SCAN_IN ; U4899
g2548 nand U4878 U2416 ; U4900
g2549 nand U2495 U2411 ; U4901
g2550 nand U4877 U2410 ; U4902
g2551 nand U2396 U4894 ; U4903
g2552 nand U4889 INSTQUEUE_REG_9__6__SCAN_IN ; U4904
g2553 nand U4878 U2420 ; U4905
g2554 nand U2495 U2409 ; U4906
g2555 nand U4877 U2408 ; U4907
g2556 nand U2395 U4894 ; U4908
g2557 nand U4889 INSTQUEUE_REG_9__5__SCAN_IN ; U4909
g2558 nand U4878 U2419 ; U4910
g2559 nand U2495 U2407 ; U4911
g2560 nand U4877 U2406 ; U4912
g2561 nand U2394 U4894 ; U4913
g2562 nand U4889 INSTQUEUE_REG_9__4__SCAN_IN ; U4914
g2563 nand U4878 U2418 ; U4915
g2564 nand U2495 U2405 ; U4916
g2565 nand U4877 U2404 ; U4917
g2566 nand U2393 U4894 ; U4918
g2567 nand U4889 INSTQUEUE_REG_9__3__SCAN_IN ; U4919
g2568 nand U4878 U2421 ; U4920
g2569 nand U2495 U2403 ; U4921
g2570 nand U4877 U2402 ; U4922
g2571 nand U2392 U4894 ; U4923
g2572 nand U4889 INSTQUEUE_REG_9__2__SCAN_IN ; U4924
g2573 nand U4878 U2414 ; U4925
g2574 nand U2495 U2401 ; U4926
g2575 nand U4877 U2400 ; U4927
g2576 nand U2391 U4894 ; U4928
g2577 nand U4889 INSTQUEUE_REG_9__1__SCAN_IN ; U4929
g2578 nand U4878 U2417 ; U4930
g2579 nand U2495 U2399 ; U4931
g2580 nand U4877 U2398 ; U4932
g2581 nand U2390 U4894 ; U4933
g2582 nand U4889 INSTQUEUE_REG_9__0__SCAN_IN ; U4934
g2583 not U3341 ; U4935
g2584 not U3340 ; U4936
g2585 nand U2440 U2445 ; U4937
g2586 not U3342 ; U4938
g2587 not U3226 ; U4939
g2588 nand U4517 U2486 ; U4940
g2589 nand U2498 U2358 ; U4941
g2590 nand U3307 U4941 ; U4942
g2591 nand U4938 U4942 ; U4943
g2592 nand U3340 STATE2_REG_3__SCAN_IN ; U4944
g2593 nand U3226 STATE2_REG_2__SCAN_IN ; U4945
g2594 nand U4943 U3638 ; U4946
g2595 nand U2498 U2388 ; U4947
g2596 nand U3307 U4947 ; U4948
g2597 nand U4948 U3342 ; U4949
g2598 nand U4939 STATE2_REG_2__SCAN_IN ; U4950
g2599 nand U4950 U4949 ; U4951
g2600 nand U4936 U2415 ; U4952
g2601 nand U2497 U2413 ; U4953
g2602 nand U4935 U2412 ; U4954
g2603 nand U2397 U4951 ; U4955
g2604 nand U4946 INSTQUEUE_REG_8__7__SCAN_IN ; U4956
g2605 nand U4936 U2416 ; U4957
g2606 nand U2497 U2411 ; U4958
g2607 nand U4935 U2410 ; U4959
g2608 nand U2396 U4951 ; U4960
g2609 nand U4946 INSTQUEUE_REG_8__6__SCAN_IN ; U4961
g2610 nand U4936 U2420 ; U4962
g2611 nand U2497 U2409 ; U4963
g2612 nand U4935 U2408 ; U4964
g2613 nand U2395 U4951 ; U4965
g2614 nand U4946 INSTQUEUE_REG_8__5__SCAN_IN ; U4966
g2615 nand U4936 U2419 ; U4967
g2616 nand U2497 U2407 ; U4968
g2617 nand U4935 U2406 ; U4969
g2618 nand U2394 U4951 ; U4970
g2619 nand U4946 INSTQUEUE_REG_8__4__SCAN_IN ; U4971
g2620 nand U4936 U2418 ; U4972
g2621 nand U2497 U2405 ; U4973
g2622 nand U4935 U2404 ; U4974
g2623 nand U2393 U4951 ; U4975
g2624 nand U4946 INSTQUEUE_REG_8__3__SCAN_IN ; U4976
g2625 nand U4936 U2421 ; U4977
g2626 nand U2497 U2403 ; U4978
g2627 nand U4935 U2402 ; U4979
g2628 nand U2392 U4951 ; U4980
g2629 nand U4946 INSTQUEUE_REG_8__2__SCAN_IN ; U4981
g2630 nand U4936 U2414 ; U4982
g2631 nand U2497 U2401 ; U4983
g2632 nand U4935 U2400 ; U4984
g2633 nand U2391 U4951 ; U4985
g2634 nand U4946 INSTQUEUE_REG_8__1__SCAN_IN ; U4986
g2635 nand U4936 U2417 ; U4987
g2636 nand U2497 U2399 ; U4988
g2637 nand U4935 U2398 ; U4989
g2638 nand U2390 U4951 ; U4990
g2639 nand U4946 INSTQUEUE_REG_8__0__SCAN_IN ; U4991
g2640 not U3346 ; U4992
g2641 nand U2439 U2442 ; U4993
g2642 not U3348 ; U4994
g2643 nand U2433 U2436 ; U4995
g2644 not U3349 ; U4996
g2645 nand U2500 U2358 ; U4997
g2646 nand U3307 U4997 ; U4998
g2647 nand U4994 U4998 ; U4999
g2648 nand U3343 STATE2_REG_3__SCAN_IN ; U5000
g2649 nand U4996 STATE2_REG_2__SCAN_IN ; U5001
g2650 nand U4999 U3647 ; U5002
g2651 nand U2500 U2388 ; U5003
g2652 nand U3307 U5003 ; U5004
g2653 nand U5004 U3348 ; U5005
g2654 nand U3349 STATE2_REG_2__SCAN_IN ; U5006
g2655 nand U5006 U5005 ; U5007
g2656 nand U4525 U2415 ; U5008
g2657 nand U4226 U2413 ; U5009
g2658 nand U4992 U2412 ; U5010
g2659 nand U2397 U5007 ; U5011
g2660 nand U5002 INSTQUEUE_REG_7__7__SCAN_IN ; U5012
g2661 nand U4525 U2416 ; U5013
g2662 nand U4226 U2411 ; U5014
g2663 nand U4992 U2410 ; U5015
g2664 nand U2396 U5007 ; U5016
g2665 nand U5002 INSTQUEUE_REG_7__6__SCAN_IN ; U5017
g2666 nand U4525 U2420 ; U5018
g2667 nand U4226 U2409 ; U5019
g2668 nand U4992 U2408 ; U5020
g2669 nand U2395 U5007 ; U5021
g2670 nand U5002 INSTQUEUE_REG_7__5__SCAN_IN ; U5022
g2671 nand U4525 U2419 ; U5023
g2672 nand U4226 U2407 ; U5024
g2673 nand U4992 U2406 ; U5025
g2674 nand U2394 U5007 ; U5026
g2675 nand U5002 INSTQUEUE_REG_7__4__SCAN_IN ; U5027
g2676 nand U4525 U2418 ; U5028
g2677 nand U4226 U2405 ; U5029
g2678 nand U4992 U2404 ; U5030
g2679 nand U2393 U5007 ; U5031
g2680 nand U5002 INSTQUEUE_REG_7__3__SCAN_IN ; U5032
g2681 nand U4525 U2421 ; U5033
g2682 nand U4226 U2403 ; U5034
g2683 nand U4992 U2402 ; U5035
g2684 nand U2392 U5007 ; U5036
g2685 nand U5002 INSTQUEUE_REG_7__2__SCAN_IN ; U5037
g2686 nand U4525 U2414 ; U5038
g2687 nand U4226 U2401 ; U5039
g2688 nand U4992 U2400 ; U5040
g2689 nand U2391 U5007 ; U5041
g2690 nand U5002 INSTQUEUE_REG_7__1__SCAN_IN ; U5042
g2691 nand U4525 U2417 ; U5043
g2692 nand U4226 U2399 ; U5044
g2693 nand U4992 U2398 ; U5045
g2694 nand U2390 U5007 ; U5046
g2695 nand U5002 INSTQUEUE_REG_7__0__SCAN_IN ; U5047
g2696 not U3351 ; U5048
g2697 not U3350 ; U5049
g2698 nand U2439 U2443 ; U5050
g2699 not U3352 ; U5051
g2700 not U3227 ; U5052
g2701 nand U4512 U2474 ; U5053
g2702 nand U2502 U2358 ; U5054
g2703 nand U3307 U5054 ; U5055
g2704 nand U5051 U5055 ; U5056
g2705 nand U3350 STATE2_REG_3__SCAN_IN ; U5057
g2706 nand U3227 STATE2_REG_2__SCAN_IN ; U5058
g2707 nand U5056 U3656 ; U5059
g2708 nand U2502 U2388 ; U5060
g2709 nand U3307 U5060 ; U5061
g2710 nand U5061 U3352 ; U5062
g2711 nand U5052 STATE2_REG_2__SCAN_IN ; U5063
g2712 nand U5063 U5062 ; U5064
g2713 nand U5049 U2415 ; U5065
g2714 nand U2501 U2413 ; U5066
g2715 nand U5048 U2412 ; U5067
g2716 nand U2397 U5064 ; U5068
g2717 nand U5059 INSTQUEUE_REG_6__7__SCAN_IN ; U5069
g2718 nand U5049 U2416 ; U5070
g2719 nand U2501 U2411 ; U5071
g2720 nand U5048 U2410 ; U5072
g2721 nand U2396 U5064 ; U5073
g2722 nand U5059 INSTQUEUE_REG_6__6__SCAN_IN ; U5074
g2723 nand U5049 U2420 ; U5075
g2724 nand U2501 U2409 ; U5076
g2725 nand U5048 U2408 ; U5077
g2726 nand U2395 U5064 ; U5078
g2727 nand U5059 INSTQUEUE_REG_6__5__SCAN_IN ; U5079
g2728 nand U5049 U2419 ; U5080
g2729 nand U2501 U2407 ; U5081
g2730 nand U5048 U2406 ; U5082
g2731 nand U2394 U5064 ; U5083
g2732 nand U5059 INSTQUEUE_REG_6__4__SCAN_IN ; U5084
g2733 nand U5049 U2418 ; U5085
g2734 nand U2501 U2405 ; U5086
g2735 nand U5048 U2404 ; U5087
g2736 nand U2393 U5064 ; U5088
g2737 nand U5059 INSTQUEUE_REG_6__3__SCAN_IN ; U5089
g2738 nand U5049 U2421 ; U5090
g2739 nand U2501 U2403 ; U5091
g2740 nand U5048 U2402 ; U5092
g2741 nand U2392 U5064 ; U5093
g2742 nand U5059 INSTQUEUE_REG_6__2__SCAN_IN ; U5094
g2743 nand U5049 U2414 ; U5095
g2744 nand U2501 U2401 ; U5096
g2745 nand U5048 U2400 ; U5097
g2746 nand U2391 U5064 ; U5098
g2747 nand U5059 INSTQUEUE_REG_6__1__SCAN_IN ; U5099
g2748 nand U5049 U2417 ; U5100
g2749 nand U2501 U2399 ; U5101
g2750 nand U5048 U2398 ; U5102
g2751 nand U2390 U5064 ; U5103
g2752 nand U5059 INSTQUEUE_REG_6__0__SCAN_IN ; U5104
g2753 not U3354 ; U5105
g2754 not U3353 ; U5106
g2755 nand U2439 U2444 ; U5107
g2756 not U3355 ; U5108
g2757 nand U2433 U2437 ; U5109
g2758 not U3356 ; U5110
g2759 nand U4513 U2474 ; U5111
g2760 nand U2504 U2358 ; U5112
g2761 nand U3307 U5112 ; U5113
g2762 nand U5108 U5113 ; U5114
g2763 nand U3353 STATE2_REG_3__SCAN_IN ; U5115
g2764 nand U5110 STATE2_REG_2__SCAN_IN ; U5116
g2765 nand U5114 U3665 ; U5117
g2766 nand U2504 U2388 ; U5118
g2767 nand U3307 U5118 ; U5119
g2768 nand U5119 U3355 ; U5120
g2769 nand U3356 STATE2_REG_2__SCAN_IN ; U5121
g2770 nand U5121 U5120 ; U5122
g2771 nand U5106 U2415 ; U5123
g2772 nand U2503 U2413 ; U5124
g2773 nand U5105 U2412 ; U5125
g2774 nand U2397 U5122 ; U5126
g2775 nand U5117 INSTQUEUE_REG_5__7__SCAN_IN ; U5127
g2776 nand U5106 U2416 ; U5128
g2777 nand U2503 U2411 ; U5129
g2778 nand U5105 U2410 ; U5130
g2779 nand U2396 U5122 ; U5131
g2780 nand U5117 INSTQUEUE_REG_5__6__SCAN_IN ; U5132
g2781 nand U5106 U2420 ; U5133
g2782 nand U2503 U2409 ; U5134
g2783 nand U5105 U2408 ; U5135
g2784 nand U2395 U5122 ; U5136
g2785 nand U5117 INSTQUEUE_REG_5__5__SCAN_IN ; U5137
g2786 nand U5106 U2419 ; U5138
g2787 nand U2503 U2407 ; U5139
g2788 nand U5105 U2406 ; U5140
g2789 nand U2394 U5122 ; U5141
g2790 nand U5117 INSTQUEUE_REG_5__4__SCAN_IN ; U5142
g2791 nand U5106 U2418 ; U5143
g2792 nand U2503 U2405 ; U5144
g2793 nand U5105 U2404 ; U5145
g2794 nand U2393 U5122 ; U5146
g2795 nand U5117 INSTQUEUE_REG_5__3__SCAN_IN ; U5147
g2796 nand U5106 U2421 ; U5148
g2797 nand U2503 U2403 ; U5149
g2798 nand U5105 U2402 ; U5150
g2799 nand U2392 U5122 ; U5151
g2800 nand U5117 INSTQUEUE_REG_5__2__SCAN_IN ; U5152
g2801 nand U5106 U2414 ; U5153
g2802 nand U2503 U2401 ; U5154
g2803 nand U5105 U2400 ; U5155
g2804 nand U2391 U5122 ; U5156
g2805 nand U5117 INSTQUEUE_REG_5__1__SCAN_IN ; U5157
g2806 nand U5106 U2417 ; U5158
g2807 nand U2503 U2399 ; U5159
g2808 nand U5105 U2398 ; U5160
g2809 nand U2390 U5122 ; U5161
g2810 nand U5117 INSTQUEUE_REG_5__0__SCAN_IN ; U5162
g2811 not U3358 ; U5163
g2812 not U3357 ; U5164
g2813 nand U2439 U2445 ; U5165
g2814 not U3359 ; U5166
g2815 not U3228 ; U5167
g2816 nand U2486 U2474 ; U5168
g2817 nand U2506 U2358 ; U5169
g2818 nand U3307 U5169 ; U5170
g2819 nand U5166 U5170 ; U5171
g2820 nand U3357 STATE2_REG_3__SCAN_IN ; U5172
g2821 nand U3228 STATE2_REG_2__SCAN_IN ; U5173
g2822 nand U5171 U3674 ; U5174
g2823 nand U2506 U2388 ; U5175
g2824 nand U3307 U5175 ; U5176
g2825 nand U5176 U3359 ; U5177
g2826 nand U5167 STATE2_REG_2__SCAN_IN ; U5178
g2827 nand U5178 U5177 ; U5179
g2828 nand U5164 U2415 ; U5180
g2829 nand U2505 U2413 ; U5181
g2830 nand U5163 U2412 ; U5182
g2831 nand U2397 U5179 ; U5183
g2832 nand U5174 INSTQUEUE_REG_4__7__SCAN_IN ; U5184
g2833 nand U5164 U2416 ; U5185
g2834 nand U2505 U2411 ; U5186
g2835 nand U5163 U2410 ; U5187
g2836 nand U2396 U5179 ; U5188
g2837 nand U5174 INSTQUEUE_REG_4__6__SCAN_IN ; U5189
g2838 nand U5164 U2420 ; U5190
g2839 nand U2505 U2409 ; U5191
g2840 nand U5163 U2408 ; U5192
g2841 nand U2395 U5179 ; U5193
g2842 nand U5174 INSTQUEUE_REG_4__5__SCAN_IN ; U5194
g2843 nand U5164 U2419 ; U5195
g2844 nand U2505 U2407 ; U5196
g2845 nand U5163 U2406 ; U5197
g2846 nand U2394 U5179 ; U5198
g2847 nand U5174 INSTQUEUE_REG_4__4__SCAN_IN ; U5199
g2848 nand U5164 U2418 ; U5200
g2849 nand U2505 U2405 ; U5201
g2850 nand U5163 U2404 ; U5202
g2851 nand U2393 U5179 ; U5203
g2852 nand U5174 INSTQUEUE_REG_4__3__SCAN_IN ; U5204
g2853 nand U5164 U2421 ; U5205
g2854 nand U2505 U2403 ; U5206
g2855 nand U5163 U2402 ; U5207
g2856 nand U2392 U5179 ; U5208
g2857 nand U5174 INSTQUEUE_REG_4__2__SCAN_IN ; U5209
g2858 nand U5164 U2414 ; U5210
g2859 nand U2505 U2401 ; U5211
g2860 nand U5163 U2400 ; U5212
g2861 nand U2391 U5179 ; U5213
g2862 nand U5174 INSTQUEUE_REG_4__1__SCAN_IN ; U5214
g2863 nand U5164 U2417 ; U5215
g2864 nand U2505 U2399 ; U5216
g2865 nand U5163 U2398 ; U5217
g2866 nand U2390 U5179 ; U5218
g2867 nand U5174 INSTQUEUE_REG_4__0__SCAN_IN ; U5219
g2868 not U3361 ; U5220
g2869 not U3360 ; U5221
g2870 nand U2441 U2442 ; U5222
g2871 not U3362 ; U5223
g2872 nand U2435 U2436 ; U5224
g2873 not U3363 ; U5225
g2874 nand U2508 U4516 ; U5226
g2875 nand U2511 U2358 ; U5227
g2876 nand U3307 U5227 ; U5228
g2877 nand U5223 U5228 ; U5229
g2878 nand U3360 STATE2_REG_3__SCAN_IN ; U5230
g2879 nand U5225 STATE2_REG_2__SCAN_IN ; U5231
g2880 nand U5229 U3683 ; U5232
g2881 nand U2511 U2388 ; U5233
g2882 nand U3307 U5233 ; U5234
g2883 nand U5234 U3362 ; U5235
g2884 nand U3363 STATE2_REG_2__SCAN_IN ; U5236
g2885 nand U5236 U5235 ; U5237
g2886 nand U5221 U2415 ; U5238
g2887 nand U2509 U2413 ; U5239
g2888 nand U5220 U2412 ; U5240
g2889 nand U2397 U5237 ; U5241
g2890 nand U5232 INSTQUEUE_REG_3__7__SCAN_IN ; U5242
g2891 nand U5221 U2416 ; U5243
g2892 nand U2509 U2411 ; U5244
g2893 nand U5220 U2410 ; U5245
g2894 nand U2396 U5237 ; U5246
g2895 nand U5232 INSTQUEUE_REG_3__6__SCAN_IN ; U5247
g2896 nand U5221 U2420 ; U5248
g2897 nand U2509 U2409 ; U5249
g2898 nand U5220 U2408 ; U5250
g2899 nand U2395 U5237 ; U5251
g2900 nand U5232 INSTQUEUE_REG_3__5__SCAN_IN ; U5252
g2901 nand U5221 U2419 ; U5253
g2902 nand U2509 U2407 ; U5254
g2903 nand U5220 U2406 ; U5255
g2904 nand U2394 U5237 ; U5256
g2905 nand U5232 INSTQUEUE_REG_3__4__SCAN_IN ; U5257
g2906 nand U5221 U2418 ; U5258
g2907 nand U2509 U2405 ; U5259
g2908 nand U5220 U2404 ; U5260
g2909 nand U2393 U5237 ; U5261
g2910 nand U5232 INSTQUEUE_REG_3__3__SCAN_IN ; U5262
g2911 nand U5221 U2421 ; U5263
g2912 nand U2509 U2403 ; U5264
g2913 nand U5220 U2402 ; U5265
g2914 nand U2392 U5237 ; U5266
g2915 nand U5232 INSTQUEUE_REG_3__2__SCAN_IN ; U5267
g2916 nand U5221 U2414 ; U5268
g2917 nand U2509 U2401 ; U5269
g2918 nand U5220 U2400 ; U5270
g2919 nand U2391 U5237 ; U5271
g2920 nand U5232 INSTQUEUE_REG_3__1__SCAN_IN ; U5272
g2921 nand U5221 U2417 ; U5273
g2922 nand U2509 U2399 ; U5274
g2923 nand U5220 U2398 ; U5275
g2924 nand U2390 U5237 ; U5276
g2925 nand U5232 INSTQUEUE_REG_3__0__SCAN_IN ; U5277
g2926 not U3365 ; U5278
g2927 not U3364 ; U5279
g2928 nand U2441 U2443 ; U5280
g2929 not U3366 ; U5281
g2930 not U3229 ; U5282
g2931 nand U2508 U4512 ; U5283
g2932 nand U2513 U2358 ; U5284
g2933 nand U3307 U5284 ; U5285
g2934 nand U5281 U5285 ; U5286
g2935 nand U3364 STATE2_REG_3__SCAN_IN ; U5287
g2936 nand U3229 STATE2_REG_2__SCAN_IN ; U5288
g2937 nand U5286 U3692 ; U5289
g2938 nand U2513 U2388 ; U5290
g2939 nand U3307 U5290 ; U5291
g2940 nand U5291 U3366 ; U5292
g2941 nand U5282 STATE2_REG_2__SCAN_IN ; U5293
g2942 nand U5293 U5292 ; U5294
g2943 nand U5279 U2415 ; U5295
g2944 nand U2512 U2413 ; U5296
g2945 nand U5278 U2412 ; U5297
g2946 nand U2397 U5294 ; U5298
g2947 nand U5289 INSTQUEUE_REG_2__7__SCAN_IN ; U5299
g2948 nand U5279 U2416 ; U5300
g2949 nand U2512 U2411 ; U5301
g2950 nand U5278 U2410 ; U5302
g2951 nand U2396 U5294 ; U5303
g2952 nand U5289 INSTQUEUE_REG_2__6__SCAN_IN ; U5304
g2953 nand U5279 U2420 ; U5305
g2954 nand U2512 U2409 ; U5306
g2955 nand U5278 U2408 ; U5307
g2956 nand U2395 U5294 ; U5308
g2957 nand U5289 INSTQUEUE_REG_2__5__SCAN_IN ; U5309
g2958 nand U5279 U2419 ; U5310
g2959 nand U2512 U2407 ; U5311
g2960 nand U5278 U2406 ; U5312
g2961 nand U2394 U5294 ; U5313
g2962 nand U5289 INSTQUEUE_REG_2__4__SCAN_IN ; U5314
g2963 nand U5279 U2418 ; U5315
g2964 nand U2512 U2405 ; U5316
g2965 nand U5278 U2404 ; U5317
g2966 nand U2393 U5294 ; U5318
g2967 nand U5289 INSTQUEUE_REG_2__3__SCAN_IN ; U5319
g2968 nand U5279 U2421 ; U5320
g2969 nand U2512 U2403 ; U5321
g2970 nand U5278 U2402 ; U5322
g2971 nand U2392 U5294 ; U5323
g2972 nand U5289 INSTQUEUE_REG_2__2__SCAN_IN ; U5324
g2973 nand U5279 U2414 ; U5325
g2974 nand U2512 U2401 ; U5326
g2975 nand U5278 U2400 ; U5327
g2976 nand U2391 U5294 ; U5328
g2977 nand U5289 INSTQUEUE_REG_2__1__SCAN_IN ; U5329
g2978 nand U5279 U2417 ; U5330
g2979 nand U2512 U2399 ; U5331
g2980 nand U5278 U2398 ; U5332
g2981 nand U2390 U5294 ; U5333
g2982 nand U5289 INSTQUEUE_REG_2__0__SCAN_IN ; U5334
g2983 not U3368 ; U5335
g2984 not U3367 ; U5336
g2985 nand U2441 U2444 ; U5337
g2986 not U3369 ; U5338
g2987 nand U2435 U2437 ; U5339
g2988 not U3370 ; U5340
g2989 nand U2508 U4513 ; U5341
g2990 nand U2515 U2358 ; U5342
g2991 nand U3307 U5342 ; U5343
g2992 nand U5338 U5343 ; U5344
g2993 nand U3367 STATE2_REG_3__SCAN_IN ; U5345
g2994 nand U5340 STATE2_REG_2__SCAN_IN ; U5346
g2995 nand U5344 U3701 ; U5347
g2996 nand U2515 U2388 ; U5348
g2997 nand U3307 U5348 ; U5349
g2998 nand U5349 U3369 ; U5350
g2999 nand U3370 STATE2_REG_2__SCAN_IN ; U5351
g3000 nand U5351 U5350 ; U5352
g3001 nand U5336 U2415 ; U5353
g3002 nand U2514 U2413 ; U5354
g3003 nand U5335 U2412 ; U5355
g3004 nand U2397 U5352 ; U5356
g3005 nand U5347 INSTQUEUE_REG_1__7__SCAN_IN ; U5357
g3006 nand U5336 U2416 ; U5358
g3007 nand U2514 U2411 ; U5359
g3008 nand U5335 U2410 ; U5360
g3009 nand U2396 U5352 ; U5361
g3010 nand U5347 INSTQUEUE_REG_1__6__SCAN_IN ; U5362
g3011 nand U5336 U2420 ; U5363
g3012 nand U2514 U2409 ; U5364
g3013 nand U5335 U2408 ; U5365
g3014 nand U2395 U5352 ; U5366
g3015 nand U5347 INSTQUEUE_REG_1__5__SCAN_IN ; U5367
g3016 nand U5336 U2419 ; U5368
g3017 nand U2514 U2407 ; U5369
g3018 nand U5335 U2406 ; U5370
g3019 nand U2394 U5352 ; U5371
g3020 nand U5347 INSTQUEUE_REG_1__4__SCAN_IN ; U5372
g3021 nand U5336 U2418 ; U5373
g3022 nand U2514 U2405 ; U5374
g3023 nand U5335 U2404 ; U5375
g3024 nand U2393 U5352 ; U5376
g3025 nand U5347 INSTQUEUE_REG_1__3__SCAN_IN ; U5377
g3026 nand U5336 U2421 ; U5378
g3027 nand U2514 U2403 ; U5379
g3028 nand U5335 U2402 ; U5380
g3029 nand U2392 U5352 ; U5381
g3030 nand U5347 INSTQUEUE_REG_1__2__SCAN_IN ; U5382
g3031 nand U5336 U2414 ; U5383
g3032 nand U2514 U2401 ; U5384
g3033 nand U5335 U2400 ; U5385
g3034 nand U2391 U5352 ; U5386
g3035 nand U5347 INSTQUEUE_REG_1__1__SCAN_IN ; U5387
g3036 nand U5336 U2417 ; U5388
g3037 nand U2514 U2399 ; U5389
g3038 nand U5335 U2398 ; U5390
g3039 nand U2390 U5352 ; U5391
g3040 nand U5347 INSTQUEUE_REG_1__0__SCAN_IN ; U5392
g3041 not U3372 ; U5393
g3042 not U3371 ; U5394
g3043 nand U2441 U2445 ; U5395
g3044 not U3373 ; U5396
g3045 not U3230 ; U5397
g3046 nand U2508 U2486 ; U5398
g3047 nand U2517 U2358 ; U5399
g3048 nand U3307 U5399 ; U5400
g3049 nand U5396 U5400 ; U5401
g3050 nand U3371 STATE2_REG_3__SCAN_IN ; U5402
g3051 nand U3230 STATE2_REG_2__SCAN_IN ; U5403
g3052 nand U5401 U3710 ; U5404
g3053 nand U2517 U2388 ; U5405
g3054 nand U3307 U5405 ; U5406
g3055 nand U5406 U3373 ; U5407
g3056 nand U5397 STATE2_REG_2__SCAN_IN ; U5408
g3057 nand U5408 U5407 ; U5409
g3058 nand U5394 U2415 ; U5410
g3059 nand U2516 U2413 ; U5411
g3060 nand U5393 U2412 ; U5412
g3061 nand U2397 U5409 ; U5413
g3062 nand U5404 INSTQUEUE_REG_0__7__SCAN_IN ; U5414
g3063 nand U5394 U2416 ; U5415
g3064 nand U2516 U2411 ; U5416
g3065 nand U5393 U2410 ; U5417
g3066 nand U2396 U5409 ; U5418
g3067 nand U5404 INSTQUEUE_REG_0__6__SCAN_IN ; U5419
g3068 nand U5394 U2420 ; U5420
g3069 nand U2516 U2409 ; U5421
g3070 nand U5393 U2408 ; U5422
g3071 nand U2395 U5409 ; U5423
g3072 nand U5404 INSTQUEUE_REG_0__5__SCAN_IN ; U5424
g3073 nand U5394 U2419 ; U5425
g3074 nand U2516 U2407 ; U5426
g3075 nand U5393 U2406 ; U5427
g3076 nand U2394 U5409 ; U5428
g3077 nand U5394 U2418 ; U5429
g3078 nand U2516 U2405 ; U5430
g3079 nand U5393 U2404 ; U5431
g3080 nand U2393 U5409 ; U5432
g3081 nand U5404 INSTQUEUE_REG_0__3__SCAN_IN ; U5433
g3082 nand U5394 U2421 ; U5434
g3083 nand U2516 U2403 ; U5435
g3084 nand U5393 U2402 ; U5436
g3085 nand U2392 U5409 ; U5437
g3086 nand U5404 INSTQUEUE_REG_0__2__SCAN_IN ; U5438
g3087 nand U5394 U2414 ; U5439
g3088 nand U2516 U2401 ; U5440
g3089 nand U5393 U2400 ; U5441
g3090 nand U2391 U5409 ; U5442
g3091 nand U5404 INSTQUEUE_REG_0__1__SCAN_IN ; U5443
g3092 nand U5394 U2417 ; U5444
g3093 nand U2516 U2399 ; U5445
g3094 nand U5393 U2398 ; U5446
g3095 nand U2390 U5409 ; U5447
g3096 nand U5404 INSTQUEUE_REG_0__0__SCAN_IN ; U5448
g3097 not U3410 ; U5449
g3098 nand U3378 U3381 U4491 ; U5450
g3099 nand U4388 U4161 U4448 ; U5451
g3100 not U3231 ; U5452
g3101 nand U4482 U3276 ; U5453
g3102 nand U5453 U3270 U5452 ; U5454
g3103 nand U3720 U2452 ; U5455
g3104 nand U4196 U5450 ; U5456
g3105 nand U3721 U7597 ; U5457
g3106 nand U4203 U3244 GTE_485_U6 ; U5458
g3107 nand U2449 U7482 ; U5459
g3108 nand U4245 U4491 ; U5460
g3109 not U4170 ; U5461
g3110 nand U2368 U4170 ; U5462
g3111 nand U3281 STATE2_REG_3__SCAN_IN ; U5463
g3112 not U4160 ; U5464
g3113 nand INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U5465
g3114 nand U5465 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U5466
g3115 nand U4369 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U5467
g3116 not U3429 ; U5468
g3117 nand U3486 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U5469
g3118 nand U5469 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U5470
g3119 not U3425 ; U5471
g3120 nand U3262 U3251 ; U5472
g3121 nand U5472 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U5473
g3122 nand U2469 U3262 ; U5474
g3123 nand U4482 U3277 ; U5475
g3124 nand U4388 U2605 ; U5476
g3125 nand U7692 U7691 U7482 ; U5477
g3126 nand U4437 U5476 ; U5478
g3127 nand U4388 U3381 U3396 ; U5479
g3128 nand U5479 U4159 ; U5480
g3129 nand U7617 U5480 ; U5481
g3130 nand U4448 U4159 ; U5482
g3131 nand U3382 U5482 ; U5483
g3132 nand U4196 U5450 ; U5484
g3133 nand U4245 U4491 ; U5485
g3134 nand U5483 U3258 ; U5486
g3135 nand U4482 U7695 ; U5487
g3136 nand U4178 U3231 ; U5488
g3137 nand U3279 U4205 ; U5489
g3138 nand U3728 U5489 ; U5490
g3139 nand R2182_U25 U7497 ; U5491
g3140 nand U4206 U3425 ; U5492
g3141 nand U4202 U3429 ; U5493
g3142 nand U5491 U3735 ; U5494
g3143 nand U4240 U3425 ; U5495
g3144 nand U2427 U5494 ; U5496
g3145 nand U5496 U5495 ; U5497
g3146 nand U3262 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U5498
g3147 not U3388 ; U5499
g3148 nand R2182_U42 U7497 ; U5500
g3149 nand U4202 U3443 ; U5501
g3150 nand U3737 U5500 ; U5502
g3151 nand U2446 U3457 ; U5503
g3152 nand U4240 U3388 ; U5504
g3153 nand U2427 U5502 ; U5505
g3154 nand U5505 U5503 U5504 ; U5506
g3155 not U3389 ; U5507
g3156 nand U2431 U4237 ; U5508
g3157 nand U3279 U5508 ; U5509
g3158 nand U5507 U5509 ; U5510
g3159 nand R2182_U33 U7497 ; U5511
g3160 nand U4202 U3252 ; U5512
g3161 nand U3738 U5511 ; U5513
g3162 nand U7700 U2446 ; U5514
g3163 nand U5507 U4240 ; U5515
g3164 nand U2427 U5513 ; U5516
g3165 nand U5516 U5514 U5515 ; U5517
g3166 nand R2182_U34 U7497 ; U5518
g3167 nand U4163 U5518 ; U5519
g3168 nand U4240 U3253 ; U5520
g3169 nand U2427 U5519 ; U5521
g3170 nand U7703 STATE2_REG_1__SCAN_IN ; U5522
g3171 nand U5521 U5522 U5520 ; U5523
g3172 nand U2428 LT_589_U6 STATE2_REG_0__SCAN_IN ; U5524
g3173 not U3391 ; U5525
g3174 nand U3283 STATE2_REG_1__SCAN_IN ; U5526
g3175 nand U4515 U3441 ; U5527
g3176 nand U3345 U5527 ; U5528
g3177 nand U3346 U5528 ; U5529
g3178 nand U2388 U5529 ; U5530
g3179 nand R2182_U25 U5526 ; U5531
g3180 nand U4214 R2144_U8 ; U5532
g3181 nand U3739 U5530 ; U5533
g3182 nand U2388 U7721 ; U5534
g3183 nand R2182_U42 U5526 ; U5535
g3184 nand U4214 R2144_U49 ; U5536
g3185 nand U3740 U5534 ; U5537
g3186 nand U3313 U3320 ; U5538
g3187 nand U2388 U5538 ; U5539
g3188 nand R2182_U33 U5526 ; U5540
g3189 nand U4214 R2144_U50 ; U5541
g3190 nand U3741 U5539 ; U5542
g3191 nand R2182_U34 U5526 ; U5543
g3192 nand R2144_U43 U4197 ; U5544
g3193 nand U5543 U5544 U4233 ; U5545
g3194 nand U4465 U3259 ; U5546
g3195 nand U4248 U2431 ; U5547
g3196 nand U2518 U5547 U7731 U7730 ; U5548
g3197 nand U4223 U4491 U4180 ; U5549
g3198 nand U2368 U5548 ; U5550
g3199 nand U4191 U3250 ; U5551
g3200 not U3401 ; U5552
g3201 nand U4250 U4196 ; U5553
g3202 nand U4244 U2389 ; U5554
g3203 nand U4254 U4238 ; U5555
g3204 nand U4252 U4482 ; U5556
g3205 nand U3746 U2519 ; U5557
g3206 nand R2099_U86 U2380 ; U5558
g3207 nand R2027_U5 U2378 ; U5559
g3208 nand R2278_U17 U2377 ; U5560
g3209 nand ADD_405_U4 U2375 ; U5561
g3210 nand U2374 INSTADDRPOINTER_REG_0__SCAN_IN ; U5562
g3211 nand U2370 REIP_REG_0__SCAN_IN ; U5563
g3212 nand U5552 INSTADDRPOINTER_REG_0__SCAN_IN ; U5564
g3213 nand R2099_U87 U2380 ; U5565
g3214 nand R2027_U71 U2378 ; U5566
g3215 nand R2278_U42 U2377 ; U5567
g3216 nand ADD_405_U81 U2375 ; U5568
g3217 nand ADD_515_U4 U2374 ; U5569
g3218 nand U2370 REIP_REG_1__SCAN_IN ; U5570
g3219 nand U5552 INSTADDRPOINTER_REG_1__SCAN_IN ; U5571
g3220 nand R2099_U138 U2380 ; U5572
g3221 nand R2027_U60 U2378 ; U5573
g3222 nand R2278_U101 U2377 ; U5574
g3223 nand ADD_405_U5 U2375 ; U5575
g3224 nand ADD_515_U71 U2374 ; U5576
g3225 nand U2370 REIP_REG_2__SCAN_IN ; U5577
g3226 nand U5552 INSTADDRPOINTER_REG_2__SCAN_IN ; U5578
g3227 nand R2099_U42 U2380 ; U5579
g3228 nand R2027_U57 U2378 ; U5580
g3229 nand R2278_U92 U2377 ; U5581
g3230 nand ADD_405_U93 U2375 ; U5582
g3231 nand ADD_515_U68 U2374 ; U5583
g3232 nand U2370 REIP_REG_3__SCAN_IN ; U5584
g3233 nand U5552 INSTADDRPOINTER_REG_3__SCAN_IN ; U5585
g3234 nand R2099_U41 U2380 ; U5586
g3235 nand R2027_U56 U2378 ; U5587
g3236 nand R2278_U89 U2377 ; U5588
g3237 nand ADD_405_U68 U2375 ; U5589
g3238 nand ADD_515_U67 U2374 ; U5590
g3239 nand U2370 REIP_REG_4__SCAN_IN ; U5591
g3240 nand U5552 INSTADDRPOINTER_REG_4__SCAN_IN ; U5592
g3241 nand R2099_U40 U2380 ; U5593
g3242 nand R2027_U55 U2378 ; U5594
g3243 nand R2278_U86 U2377 ; U5595
g3244 nand ADD_405_U67 U2375 ; U5596
g3245 nand ADD_515_U66 U2374 ; U5597
g3246 nand U2370 REIP_REG_5__SCAN_IN ; U5598
g3247 nand U5552 INSTADDRPOINTER_REG_5__SCAN_IN ; U5599
g3248 nand R2099_U39 U2380 ; U5600
g3249 nand R2027_U54 U2378 ; U5601
g3250 nand R2278_U83 U2377 ; U5602
g3251 nand ADD_405_U66 U2375 ; U5603
g3252 nand ADD_515_U65 U2374 ; U5604
g3253 nand U2370 REIP_REG_6__SCAN_IN ; U5605
g3254 nand U5552 INSTADDRPOINTER_REG_6__SCAN_IN ; U5606
g3255 nand R2099_U38 U2380 ; U5607
g3256 nand R2027_U53 U2378 ; U5608
g3257 nand R2278_U80 U2377 ; U5609
g3258 nand ADD_405_U65 U2375 ; U5610
g3259 nand ADD_515_U64 U2374 ; U5611
g3260 nand U2370 REIP_REG_7__SCAN_IN ; U5612
g3261 nand U5552 INSTADDRPOINTER_REG_7__SCAN_IN ; U5613
g3262 nand R2099_U37 U2380 ; U5614
g3263 nand R2027_U52 U2378 ; U5615
g3264 nand R2278_U77 U2377 ; U5616
g3265 nand ADD_405_U64 U2375 ; U5617
g3266 nand ADD_515_U63 U2374 ; U5618
g3267 nand U2370 REIP_REG_8__SCAN_IN ; U5619
g3268 nand U5552 INSTADDRPOINTER_REG_8__SCAN_IN ; U5620
g3269 nand R2099_U36 U2380 ; U5621
g3270 nand R2027_U51 U2378 ; U5622
g3271 nand R2278_U74 U2377 ; U5623
g3272 nand ADD_405_U63 U2375 ; U5624
g3273 nand ADD_515_U62 U2374 ; U5625
g3274 nand U2370 REIP_REG_9__SCAN_IN ; U5626
g3275 nand U5552 INSTADDRPOINTER_REG_9__SCAN_IN ; U5627
g3276 nand R2099_U85 U2380 ; U5628
g3277 nand R2027_U81 U2378 ; U5629
g3278 nand R2278_U160 U2377 ; U5630
g3279 nand ADD_405_U91 U2375 ; U5631
g3280 nand ADD_515_U91 U2374 ; U5632
g3281 nand U2370 REIP_REG_10__SCAN_IN ; U5633
g3282 nand U5552 INSTADDRPOINTER_REG_10__SCAN_IN ; U5634
g3283 nand R2099_U84 U2380 ; U5635
g3284 nand R2027_U80 U2378 ; U5636
g3285 nand R2278_U157 U2377 ; U5637
g3286 nand ADD_405_U90 U2375 ; U5638
g3287 nand ADD_515_U90 U2374 ; U5639
g3288 nand U2370 REIP_REG_11__SCAN_IN ; U5640
g3289 nand U5552 INSTADDRPOINTER_REG_11__SCAN_IN ; U5641
g3290 nand R2099_U83 U2380 ; U5642
g3291 nand R2027_U79 U2378 ; U5643
g3292 nand R2278_U154 U2377 ; U5644
g3293 nand ADD_405_U89 U2375 ; U5645
g3294 nand ADD_515_U89 U2374 ; U5646
g3295 nand U2370 REIP_REG_12__SCAN_IN ; U5647
g3296 nand U5552 INSTADDRPOINTER_REG_12__SCAN_IN ; U5648
g3297 nand R2099_U82 U2380 ; U5649
g3298 nand R2027_U78 U2378 ; U5650
g3299 nand R2278_U151 U2377 ; U5651
g3300 nand ADD_405_U88 U2375 ; U5652
g3301 nand ADD_515_U88 U2374 ; U5653
g3302 nand U2370 REIP_REG_13__SCAN_IN ; U5654
g3303 nand U5552 INSTADDRPOINTER_REG_13__SCAN_IN ; U5655
g3304 nand R2099_U81 U2380 ; U5656
g3305 nand R2027_U77 U2378 ; U5657
g3306 nand R2278_U148 U2377 ; U5658
g3307 nand ADD_405_U87 U2375 ; U5659
g3308 nand ADD_515_U87 U2374 ; U5660
g3309 nand U2370 REIP_REG_14__SCAN_IN ; U5661
g3310 nand U5552 INSTADDRPOINTER_REG_14__SCAN_IN ; U5662
g3311 nand R2099_U80 U2380 ; U5663
g3312 nand R2027_U76 U2378 ; U5664
g3313 nand R2278_U145 U2377 ; U5665
g3314 nand ADD_405_U86 U2375 ; U5666
g3315 nand ADD_515_U86 U2374 ; U5667
g3316 nand U2370 REIP_REG_15__SCAN_IN ; U5668
g3317 nand U5552 INSTADDRPOINTER_REG_15__SCAN_IN ; U5669
g3318 nand R2099_U79 U2380 ; U5670
g3319 nand R2027_U75 U2378 ; U5671
g3320 nand R2278_U142 U2377 ; U5672
g3321 nand ADD_405_U85 U2375 ; U5673
g3322 nand ADD_515_U85 U2374 ; U5674
g3323 nand U2370 REIP_REG_16__SCAN_IN ; U5675
g3324 nand U5552 INSTADDRPOINTER_REG_16__SCAN_IN ; U5676
g3325 nand R2099_U78 U2380 ; U5677
g3326 nand R2027_U74 U2378 ; U5678
g3327 nand R2278_U139 U2377 ; U5679
g3328 nand ADD_405_U84 U2375 ; U5680
g3329 nand ADD_515_U84 U2374 ; U5681
g3330 nand U2370 REIP_REG_17__SCAN_IN ; U5682
g3331 nand U5552 INSTADDRPOINTER_REG_17__SCAN_IN ; U5683
g3332 nand R2099_U77 U2380 ; U5684
g3333 nand R2027_U73 U2378 ; U5685
g3334 nand R2278_U136 U2377 ; U5686
g3335 nand ADD_405_U83 U2375 ; U5687
g3336 nand ADD_515_U83 U2374 ; U5688
g3337 nand U2370 REIP_REG_18__SCAN_IN ; U5689
g3338 nand U5552 INSTADDRPOINTER_REG_18__SCAN_IN ; U5690
g3339 nand R2099_U76 U2380 ; U5691
g3340 nand R2027_U72 U2378 ; U5692
g3341 nand R2278_U133 U2377 ; U5693
g3342 nand ADD_405_U82 U2375 ; U5694
g3343 nand ADD_515_U82 U2374 ; U5695
g3344 nand U2370 REIP_REG_19__SCAN_IN ; U5696
g3345 nand U5552 INSTADDRPOINTER_REG_19__SCAN_IN ; U5697
g3346 nand R2099_U75 U2380 ; U5698
g3347 nand R2027_U70 U2378 ; U5699
g3348 nand R2278_U129 U2377 ; U5700
g3349 nand ADD_405_U80 U2375 ; U5701
g3350 nand ADD_515_U81 U2374 ; U5702
g3351 nand U2370 REIP_REG_20__SCAN_IN ; U5703
g3352 nand U5552 INSTADDRPOINTER_REG_20__SCAN_IN ; U5704
g3353 nand R2099_U74 U2380 ; U5705
g3354 nand R2027_U69 U2378 ; U5706
g3355 nand R2278_U126 U2377 ; U5707
g3356 nand ADD_405_U79 U2375 ; U5708
g3357 nand ADD_515_U80 U2374 ; U5709
g3358 nand U2370 REIP_REG_21__SCAN_IN ; U5710
g3359 nand U5552 INSTADDRPOINTER_REG_21__SCAN_IN ; U5711
g3360 nand R2099_U73 U2380 ; U5712
g3361 nand R2027_U68 U2378 ; U5713
g3362 nand R2278_U123 U2377 ; U5714
g3363 nand ADD_405_U78 U2375 ; U5715
g3364 nand ADD_515_U79 U2374 ; U5716
g3365 nand U2370 REIP_REG_22__SCAN_IN ; U5717
g3366 nand U5552 INSTADDRPOINTER_REG_22__SCAN_IN ; U5718
g3367 nand R2099_U72 U2380 ; U5719
g3368 nand R2027_U67 U2378 ; U5720
g3369 nand R2278_U120 U2377 ; U5721
g3370 nand ADD_405_U77 U2375 ; U5722
g3371 nand ADD_515_U78 U2374 ; U5723
g3372 nand U2370 REIP_REG_23__SCAN_IN ; U5724
g3373 nand U5552 INSTADDRPOINTER_REG_23__SCAN_IN ; U5725
g3374 nand R2099_U71 U2380 ; U5726
g3375 nand R2027_U66 U2378 ; U5727
g3376 nand R2278_U117 U2377 ; U5728
g3377 nand ADD_405_U76 U2375 ; U5729
g3378 nand ADD_515_U77 U2374 ; U5730
g3379 nand U2370 REIP_REG_24__SCAN_IN ; U5731
g3380 nand U5552 INSTADDRPOINTER_REG_24__SCAN_IN ; U5732
g3381 nand R2099_U70 U2380 ; U5733
g3382 nand R2027_U65 U2378 ; U5734
g3383 nand R2278_U114 U2377 ; U5735
g3384 nand ADD_405_U75 U2375 ; U5736
g3385 nand ADD_515_U76 U2374 ; U5737
g3386 nand U2370 REIP_REG_25__SCAN_IN ; U5738
g3387 nand U5552 INSTADDRPOINTER_REG_25__SCAN_IN ; U5739
g3388 nand R2099_U69 U2380 ; U5740
g3389 nand R2027_U64 U2378 ; U5741
g3390 nand R2278_U111 U2377 ; U5742
g3391 nand ADD_405_U74 U2375 ; U5743
g3392 nand ADD_515_U75 U2374 ; U5744
g3393 nand U2370 REIP_REG_26__SCAN_IN ; U5745
g3394 nand U5552 INSTADDRPOINTER_REG_26__SCAN_IN ; U5746
g3395 nand R2099_U68 U2380 ; U5747
g3396 nand R2027_U63 U2378 ; U5748
g3397 nand R2278_U108 U2377 ; U5749
g3398 nand ADD_405_U73 U2375 ; U5750
g3399 nand ADD_515_U74 U2374 ; U5751
g3400 nand U2370 REIP_REG_27__SCAN_IN ; U5752
g3401 nand U5552 INSTADDRPOINTER_REG_27__SCAN_IN ; U5753
g3402 nand R2099_U67 U2380 ; U5754
g3403 nand R2027_U62 U2378 ; U5755
g3404 nand R2278_U105 U2377 ; U5756
g3405 nand ADD_405_U72 U2375 ; U5757
g3406 nand ADD_515_U73 U2374 ; U5758
g3407 nand U2370 REIP_REG_28__SCAN_IN ; U5759
g3408 nand U5552 INSTADDRPOINTER_REG_28__SCAN_IN ; U5760
g3409 nand R2099_U66 U2380 ; U5761
g3410 nand R2027_U61 U2378 ; U5762
g3411 nand R2278_U103 U2377 ; U5763
g3412 nand ADD_405_U71 U2375 ; U5764
g3413 nand ADD_515_U72 U2374 ; U5765
g3414 nand U2370 REIP_REG_29__SCAN_IN ; U5766
g3415 nand U5552 INSTADDRPOINTER_REG_29__SCAN_IN ; U5767
g3416 nand R2099_U65 U2380 ; U5768
g3417 nand R2027_U59 U2378 ; U5769
g3418 nand R2278_U98 U2377 ; U5770
g3419 nand ADD_405_U70 U2375 ; U5771
g3420 nand ADD_515_U70 U2374 ; U5772
g3421 nand U2370 REIP_REG_30__SCAN_IN ; U5773
g3422 nand U5552 INSTADDRPOINTER_REG_30__SCAN_IN ; U5774
g3423 nand R2099_U64 U2380 ; U5775
g3424 nand R2027_U58 U2378 ; U5776
g3425 nand R2278_U96 U2377 ; U5777
g3426 nand ADD_405_U69 U2375 ; U5778
g3427 nand ADD_515_U69 U2374 ; U5779
g3428 nand U2370 REIP_REG_31__SCAN_IN ; U5780
g3429 nand U5552 INSTADDRPOINTER_REG_31__SCAN_IN ; U5781
g3430 nand U4197 U3281 ; U5782
g3431 not U3403 ; U5783
g3432 nand U3281 STATE2_REG_2__SCAN_IN ; U5784
g3433 nand U3295 STATE2_REG_1__SCAN_IN ; U5785
g3434 nand U5785 U5784 ; U5786
g3435 nand U2376 PHYADDRPOINTER_REG_0__SCAN_IN ; U5787
g3436 nand U2372 R2278_U17 ; U5788
g3437 nand U2365 REIP_REG_0__SCAN_IN ; U5789
g3438 nand R2358_U82 U2364 ; U5790
g3439 nand U5783 PHYADDRPOINTER_REG_0__SCAN_IN ; U5791
g3440 nand R2337_U5 U2376 ; U5792
g3441 nand U2372 R2278_U42 ; U5793
g3442 nand U2365 REIP_REG_1__SCAN_IN ; U5794
g3443 nand R2358_U112 U2364 ; U5795
g3444 nand U5783 PHYADDRPOINTER_REG_1__SCAN_IN ; U5796
g3445 nand R2337_U60 U2376 ; U5797
g3446 nand U2372 R2278_U101 ; U5798
g3447 nand U2365 REIP_REG_2__SCAN_IN ; U5799
g3448 nand R2358_U19 U2364 ; U5800
g3449 nand U5783 PHYADDRPOINTER_REG_2__SCAN_IN ; U5801
g3450 nand R2337_U57 U2376 ; U5802
g3451 nand U2372 R2278_U92 ; U5803
g3452 nand U2365 REIP_REG_3__SCAN_IN ; U5804
g3453 nand R2358_U20 U2364 ; U5805
g3454 nand U5783 PHYADDRPOINTER_REG_3__SCAN_IN ; U5806
g3455 nand R2337_U56 U2376 ; U5807
g3456 nand U2372 R2278_U89 ; U5808
g3457 nand U2365 REIP_REG_4__SCAN_IN ; U5809
g3458 nand R2358_U90 U2364 ; U5810
g3459 nand U5783 PHYADDRPOINTER_REG_4__SCAN_IN ; U5811
g3460 nand R2337_U55 U2376 ; U5812
g3461 nand U2372 R2278_U86 ; U5813
g3462 nand U2365 REIP_REG_5__SCAN_IN ; U5814
g3463 nand R2358_U88 U2364 ; U5815
g3464 nand U5783 PHYADDRPOINTER_REG_5__SCAN_IN ; U5816
g3465 nand R2337_U54 U2376 ; U5817
g3466 nand U2372 R2278_U83 ; U5818
g3467 nand U2365 REIP_REG_6__SCAN_IN ; U5819
g3468 nand R2358_U86 U2364 ; U5820
g3469 nand U5783 PHYADDRPOINTER_REG_6__SCAN_IN ; U5821
g3470 nand R2337_U53 U2376 ; U5822
g3471 nand U2372 R2278_U80 ; U5823
g3472 nand U2365 REIP_REG_7__SCAN_IN ; U5824
g3473 nand R2358_U21 U2364 ; U5825
g3474 nand U5783 PHYADDRPOINTER_REG_7__SCAN_IN ; U5826
g3475 nand R2337_U52 U2376 ; U5827
g3476 nand U2372 R2278_U77 ; U5828
g3477 nand U2365 REIP_REG_8__SCAN_IN ; U5829
g3478 nand R2358_U85 U2364 ; U5830
g3479 nand U5783 PHYADDRPOINTER_REG_8__SCAN_IN ; U5831
g3480 nand R2337_U51 U2376 ; U5832
g3481 nand U2372 R2278_U74 ; U5833
g3482 nand U2365 REIP_REG_9__SCAN_IN ; U5834
g3483 nand R2358_U83 U2364 ; U5835
g3484 nand U5783 PHYADDRPOINTER_REG_9__SCAN_IN ; U5836
g3485 nand R2337_U80 U2376 ; U5837
g3486 nand U2372 R2278_U160 ; U5838
g3487 nand U2365 REIP_REG_10__SCAN_IN ; U5839
g3488 nand R2358_U14 U2364 ; U5840
g3489 nand U5783 PHYADDRPOINTER_REG_10__SCAN_IN ; U5841
g3490 nand R2337_U79 U2376 ; U5842
g3491 nand U2372 R2278_U157 ; U5843
g3492 nand U2365 REIP_REG_11__SCAN_IN ; U5844
g3493 nand R2358_U15 U2364 ; U5845
g3494 nand U5783 PHYADDRPOINTER_REG_11__SCAN_IN ; U5846
g3495 nand R2337_U78 U2376 ; U5847
g3496 nand U2372 R2278_U154 ; U5848
g3497 nand U2365 REIP_REG_12__SCAN_IN ; U5849
g3498 nand R2358_U122 U2364 ; U5850
g3499 nand U5783 PHYADDRPOINTER_REG_12__SCAN_IN ; U5851
g3500 nand R2337_U77 U2376 ; U5852
g3501 nand U2372 R2278_U151 ; U5853
g3502 nand U2365 REIP_REG_13__SCAN_IN ; U5854
g3503 nand R2358_U120 U2364 ; U5855
g3504 nand U5783 PHYADDRPOINTER_REG_13__SCAN_IN ; U5856
g3505 nand R2337_U76 U2376 ; U5857
g3506 nand U2372 R2278_U148 ; U5858
g3507 nand U2365 REIP_REG_14__SCAN_IN ; U5859
g3508 nand R2358_U119 U2364 ; U5860
g3509 nand U5783 PHYADDRPOINTER_REG_14__SCAN_IN ; U5861
g3510 nand R2337_U75 U2376 ; U5862
g3511 nand U2372 R2278_U145 ; U5863
g3512 nand U2365 REIP_REG_15__SCAN_IN ; U5864
g3513 nand R2358_U16 U2364 ; U5865
g3514 nand U5783 PHYADDRPOINTER_REG_15__SCAN_IN ; U5866
g3515 nand R2337_U74 U2376 ; U5867
g3516 nand U2372 R2278_U142 ; U5868
g3517 nand U2365 REIP_REG_16__SCAN_IN ; U5869
g3518 nand R2358_U17 U2364 ; U5870
g3519 nand U5783 PHYADDRPOINTER_REG_16__SCAN_IN ; U5871
g3520 nand R2337_U73 U2376 ; U5872
g3521 nand U2372 R2278_U139 ; U5873
g3522 nand U2365 REIP_REG_17__SCAN_IN ; U5874
g3523 nand R2358_U118 U2364 ; U5875
g3524 nand U5783 PHYADDRPOINTER_REG_17__SCAN_IN ; U5876
g3525 nand R2337_U72 U2376 ; U5877
g3526 nand U2372 R2278_U136 ; U5878
g3527 nand U2365 REIP_REG_18__SCAN_IN ; U5879
g3528 nand R2358_U116 U2364 ; U5880
g3529 nand U5783 PHYADDRPOINTER_REG_18__SCAN_IN ; U5881
g3530 nand R2337_U71 U2376 ; U5882
g3531 nand U2372 R2278_U133 ; U5883
g3532 nand U2365 REIP_REG_19__SCAN_IN ; U5884
g3533 nand R2358_U114 U2364 ; U5885
g3534 nand U5783 PHYADDRPOINTER_REG_19__SCAN_IN ; U5886
g3535 nand R2337_U70 U2376 ; U5887
g3536 nand U2372 R2278_U129 ; U5888
g3537 nand U2365 REIP_REG_20__SCAN_IN ; U5889
g3538 nand R2358_U110 U2364 ; U5890
g3539 nand U5783 PHYADDRPOINTER_REG_20__SCAN_IN ; U5891
g3540 nand R2337_U69 U2376 ; U5892
g3541 nand U2372 R2278_U126 ; U5893
g3542 nand U2365 REIP_REG_21__SCAN_IN ; U5894
g3543 nand R2358_U18 U2364 ; U5895
g3544 nand U5783 PHYADDRPOINTER_REG_21__SCAN_IN ; U5896
g3545 nand R2337_U68 U2376 ; U5897
g3546 nand U2372 R2278_U123 ; U5898
g3547 nand U2365 REIP_REG_22__SCAN_IN ; U5899
g3548 nand R2358_U109 U2364 ; U5900
g3549 nand U5783 PHYADDRPOINTER_REG_22__SCAN_IN ; U5901
g3550 nand R2337_U67 U2376 ; U5902
g3551 nand U2372 R2278_U120 ; U5903
g3552 nand U2365 REIP_REG_23__SCAN_IN ; U5904
g3553 nand R2358_U107 U2364 ; U5905
g3554 nand U5783 PHYADDRPOINTER_REG_23__SCAN_IN ; U5906
g3555 nand R2337_U66 U2376 ; U5907
g3556 nand U2372 R2278_U117 ; U5908
g3557 nand U2365 REIP_REG_24__SCAN_IN ; U5909
g3558 nand R2358_U105 U2364 ; U5910
g3559 nand U5783 PHYADDRPOINTER_REG_24__SCAN_IN ; U5911
g3560 nand R2337_U65 U2376 ; U5912
g3561 nand U2372 R2278_U114 ; U5913
g3562 nand U2365 REIP_REG_25__SCAN_IN ; U5914
g3563 nand R2358_U103 U2364 ; U5915
g3564 nand U5783 PHYADDRPOINTER_REG_25__SCAN_IN ; U5916
g3565 nand R2337_U64 U2376 ; U5917
g3566 nand U2372 R2278_U111 ; U5918
g3567 nand U2365 REIP_REG_26__SCAN_IN ; U5919
g3568 nand R2358_U101 U2364 ; U5920
g3569 nand U5783 PHYADDRPOINTER_REG_26__SCAN_IN ; U5921
g3570 nand R2337_U63 U2376 ; U5922
g3571 nand U2372 R2278_U108 ; U5923
g3572 nand U2365 REIP_REG_27__SCAN_IN ; U5924
g3573 nand R2358_U99 U2364 ; U5925
g3574 nand U5783 PHYADDRPOINTER_REG_27__SCAN_IN ; U5926
g3575 nand R2337_U62 U2376 ; U5927
g3576 nand U2372 R2278_U105 ; U5928
g3577 nand U2365 REIP_REG_28__SCAN_IN ; U5929
g3578 nand R2358_U97 U2364 ; U5930
g3579 nand U5783 PHYADDRPOINTER_REG_28__SCAN_IN ; U5931
g3580 nand R2337_U61 U2376 ; U5932
g3581 nand U2372 R2278_U103 ; U5933
g3582 nand U2365 REIP_REG_29__SCAN_IN ; U5934
g3583 nand R2358_U95 U2364 ; U5935
g3584 nand U5783 PHYADDRPOINTER_REG_29__SCAN_IN ; U5936
g3585 nand R2337_U59 U2376 ; U5937
g3586 nand U2372 R2278_U98 ; U5938
g3587 nand U2365 REIP_REG_30__SCAN_IN ; U5939
g3588 nand R2358_U93 U2364 ; U5940
g3589 nand U5783 PHYADDRPOINTER_REG_30__SCAN_IN ; U5941
g3590 nand R2337_U58 U2376 ; U5942
g3591 nand U2372 R2278_U96 ; U5943
g3592 nand U2365 REIP_REG_31__SCAN_IN ; U5944
g3593 nand R2358_U91 U2364 ; U5945
g3594 nand U5783 PHYADDRPOINTER_REG_31__SCAN_IN ; U5946
g3595 nand READY_N U3269 ; U5947
g3596 nand U2382 EAX_REG_15__SCAN_IN ; U5948
g3597 nand DATAI_15_ U2381 ; U5949
g3598 nand U5949 U5948 ; U5950
g3599 nand U2382 EAX_REG_14__SCAN_IN ; U5951
g3600 nand DATAI_14_ U2381 ; U5952
g3601 nand U5952 U5951 ; U5953
g3602 nand U2382 EAX_REG_13__SCAN_IN ; U5954
g3603 nand DATAI_13_ U2381 ; U5955
g3604 nand U5955 U5954 ; U5956
g3605 nand U2382 EAX_REG_12__SCAN_IN ; U5957
g3606 nand DATAI_12_ U2381 ; U5958
g3607 nand U5958 U5957 ; U5959
g3608 nand U2382 EAX_REG_11__SCAN_IN ; U5960
g3609 nand DATAI_11_ U2381 ; U5961
g3610 nand U5961 U5960 ; U5962
g3611 nand U2382 EAX_REG_10__SCAN_IN ; U5963
g3612 nand DATAI_10_ U2381 ; U5964
g3613 nand U5964 U5963 ; U5965
g3614 nand U2382 EAX_REG_9__SCAN_IN ; U5966
g3615 nand DATAI_9_ U2381 ; U5967
g3616 nand U5967 U5966 ; U5968
g3617 nand U2382 EAX_REG_8__SCAN_IN ; U5969
g3618 nand DATAI_8_ U2381 ; U5970
g3619 nand U5970 U5969 ; U5971
g3620 nand U2382 EAX_REG_7__SCAN_IN ; U5972
g3621 nand U2381 DATAI_7_ ; U5973
g3622 nand U5973 U5972 ; U5974
g3623 nand U2382 EAX_REG_6__SCAN_IN ; U5975
g3624 nand U2381 DATAI_6_ ; U5976
g3625 nand U5976 U5975 ; U5977
g3626 nand U2382 EAX_REG_5__SCAN_IN ; U5978
g3627 nand U2381 DATAI_5_ ; U5979
g3628 nand U5979 U5978 ; U5980
g3629 nand U2382 EAX_REG_4__SCAN_IN ; U5981
g3630 nand U2381 DATAI_4_ ; U5982
g3631 nand U5982 U5981 ; U5983
g3632 nand U2382 EAX_REG_3__SCAN_IN ; U5984
g3633 nand U2381 DATAI_3_ ; U5985
g3634 nand U5985 U5984 ; U5986
g3635 nand U2382 EAX_REG_2__SCAN_IN ; U5987
g3636 nand U2381 DATAI_2_ ; U5988
g3637 nand U5988 U5987 ; U5989
g3638 nand U2382 EAX_REG_1__SCAN_IN ; U5990
g3639 nand U2381 DATAI_1_ ; U5991
g3640 nand U5991 U5990 ; U5992
g3641 nand U2382 EAX_REG_0__SCAN_IN ; U5993
g3642 nand U2381 DATAI_0_ ; U5994
g3643 nand U5994 U5993 ; U5995
g3644 nand U2382 EAX_REG_30__SCAN_IN ; U5996
g3645 nand DATAI_14_ U2381 ; U5997
g3646 nand U5997 U5996 ; U5998
g3647 nand U2382 EAX_REG_29__SCAN_IN ; U5999
g3648 nand DATAI_13_ U2381 ; U6000
g3649 nand U6000 U5999 ; U6001
g3650 nand U2382 EAX_REG_28__SCAN_IN ; U6002
g3651 nand DATAI_12_ U2381 ; U6003
g3652 nand U6003 U6002 ; U6004
g3653 nand U2382 EAX_REG_27__SCAN_IN ; U6005
g3654 nand DATAI_11_ U2381 ; U6006
g3655 nand U6006 U6005 ; U6007
g3656 nand U2382 EAX_REG_26__SCAN_IN ; U6008
g3657 nand DATAI_10_ U2381 ; U6009
g3658 nand U6009 U6008 ; U6010
g3659 nand U2382 EAX_REG_25__SCAN_IN ; U6011
g3660 nand DATAI_9_ U2381 ; U6012
g3661 nand U6012 U6011 ; U6013
g3662 nand U2382 EAX_REG_24__SCAN_IN ; U6014
g3663 nand DATAI_8_ U2381 ; U6015
g3664 nand U6015 U6014 ; U6016
g3665 nand U2382 EAX_REG_23__SCAN_IN ; U6017
g3666 nand U2381 DATAI_7_ ; U6018
g3667 nand U6018 U6017 ; U6019
g3668 nand U2382 EAX_REG_22__SCAN_IN ; U6020
g3669 nand U2381 DATAI_6_ ; U6021
g3670 nand U6021 U6020 ; U6022
g3671 nand U2382 EAX_REG_21__SCAN_IN ; U6023
g3672 nand U2381 DATAI_5_ ; U6024
g3673 nand U6024 U6023 ; U6025
g3674 nand U2382 EAX_REG_20__SCAN_IN ; U6026
g3675 nand U2381 DATAI_4_ ; U6027
g3676 nand U6027 U6026 ; U6028
g3677 nand U2382 EAX_REG_19__SCAN_IN ; U6029
g3678 nand U2381 DATAI_3_ ; U6030
g3679 nand U6030 U6029 ; U6031
g3680 nand U2382 EAX_REG_18__SCAN_IN ; U6032
g3681 nand U2381 DATAI_2_ ; U6033
g3682 nand U6033 U6032 ; U6034
g3683 nand U2382 EAX_REG_17__SCAN_IN ; U6035
g3684 nand U2381 DATAI_1_ ; U6036
g3685 nand U6036 U6035 ; U6037
g3686 nand U2382 EAX_REG_16__SCAN_IN ; U6038
g3687 nand U2381 DATAI_0_ ; U6039
g3688 nand U6039 U6038 ; U6040
g3689 nand U4223 U7594 U4247 ; U6041
g3690 nand U2428 U3281 ; U6042
g3691 not U3404 ; U6043
g3692 nand U2385 LWORD_REG_0__SCAN_IN ; U6044
g3693 nand U2384 EAX_REG_0__SCAN_IN ; U6045
g3694 nand U6043 DATAO_REG_0__SCAN_IN ; U6046
g3695 nand U2385 LWORD_REG_1__SCAN_IN ; U6047
g3696 nand U2384 EAX_REG_1__SCAN_IN ; U6048
g3697 nand U6043 DATAO_REG_1__SCAN_IN ; U6049
g3698 nand U2385 LWORD_REG_2__SCAN_IN ; U6050
g3699 nand U2384 EAX_REG_2__SCAN_IN ; U6051
g3700 nand U6043 DATAO_REG_2__SCAN_IN ; U6052
g3701 nand U2385 LWORD_REG_3__SCAN_IN ; U6053
g3702 nand U2384 EAX_REG_3__SCAN_IN ; U6054
g3703 nand U6043 DATAO_REG_3__SCAN_IN ; U6055
g3704 nand U2385 LWORD_REG_4__SCAN_IN ; U6056
g3705 nand U2384 EAX_REG_4__SCAN_IN ; U6057
g3706 nand U6043 DATAO_REG_4__SCAN_IN ; U6058
g3707 nand U2385 LWORD_REG_5__SCAN_IN ; U6059
g3708 nand U2384 EAX_REG_5__SCAN_IN ; U6060
g3709 nand U6043 DATAO_REG_5__SCAN_IN ; U6061
g3710 nand U2385 LWORD_REG_6__SCAN_IN ; U6062
g3711 nand U2384 EAX_REG_6__SCAN_IN ; U6063
g3712 nand U6043 DATAO_REG_6__SCAN_IN ; U6064
g3713 nand U2385 LWORD_REG_7__SCAN_IN ; U6065
g3714 nand U2384 EAX_REG_7__SCAN_IN ; U6066
g3715 nand U6043 DATAO_REG_7__SCAN_IN ; U6067
g3716 nand U2385 LWORD_REG_8__SCAN_IN ; U6068
g3717 nand U2384 EAX_REG_8__SCAN_IN ; U6069
g3718 nand U6043 DATAO_REG_8__SCAN_IN ; U6070
g3719 nand U2385 LWORD_REG_9__SCAN_IN ; U6071
g3720 nand U2384 EAX_REG_9__SCAN_IN ; U6072
g3721 nand U6043 DATAO_REG_9__SCAN_IN ; U6073
g3722 nand U2385 LWORD_REG_10__SCAN_IN ; U6074
g3723 nand U2384 EAX_REG_10__SCAN_IN ; U6075
g3724 nand U6043 DATAO_REG_10__SCAN_IN ; U6076
g3725 nand U2385 LWORD_REG_11__SCAN_IN ; U6077
g3726 nand U2384 EAX_REG_11__SCAN_IN ; U6078
g3727 nand U6043 DATAO_REG_11__SCAN_IN ; U6079
g3728 nand U2385 LWORD_REG_12__SCAN_IN ; U6080
g3729 nand U2384 EAX_REG_12__SCAN_IN ; U6081
g3730 nand U6043 DATAO_REG_12__SCAN_IN ; U6082
g3731 nand U2385 LWORD_REG_13__SCAN_IN ; U6083
g3732 nand U2384 EAX_REG_13__SCAN_IN ; U6084
g3733 nand U6043 DATAO_REG_13__SCAN_IN ; U6085
g3734 nand U2385 LWORD_REG_14__SCAN_IN ; U6086
g3735 nand U2384 EAX_REG_14__SCAN_IN ; U6087
g3736 nand U6043 DATAO_REG_14__SCAN_IN ; U6088
g3737 nand U2385 LWORD_REG_15__SCAN_IN ; U6089
g3738 nand U2384 EAX_REG_15__SCAN_IN ; U6090
g3739 nand U6043 DATAO_REG_15__SCAN_IN ; U6091
g3740 nand U2424 EAX_REG_16__SCAN_IN ; U6092
g3741 nand U2385 UWORD_REG_0__SCAN_IN ; U6093
g3742 nand U6043 DATAO_REG_16__SCAN_IN ; U6094
g3743 nand U2424 EAX_REG_17__SCAN_IN ; U6095
g3744 nand U2385 UWORD_REG_1__SCAN_IN ; U6096
g3745 nand U6043 DATAO_REG_17__SCAN_IN ; U6097
g3746 nand U2424 EAX_REG_18__SCAN_IN ; U6098
g3747 nand U2385 UWORD_REG_2__SCAN_IN ; U6099
g3748 nand U6043 DATAO_REG_18__SCAN_IN ; U6100
g3749 nand U2424 EAX_REG_19__SCAN_IN ; U6101
g3750 nand U2385 UWORD_REG_3__SCAN_IN ; U6102
g3751 nand U6043 DATAO_REG_19__SCAN_IN ; U6103
g3752 nand U2424 EAX_REG_20__SCAN_IN ; U6104
g3753 nand U2385 UWORD_REG_4__SCAN_IN ; U6105
g3754 nand U6043 DATAO_REG_20__SCAN_IN ; U6106
g3755 nand U2424 EAX_REG_21__SCAN_IN ; U6107
g3756 nand U2385 UWORD_REG_5__SCAN_IN ; U6108
g3757 nand U6043 DATAO_REG_21__SCAN_IN ; U6109
g3758 nand U2424 EAX_REG_22__SCAN_IN ; U6110
g3759 nand U2385 UWORD_REG_6__SCAN_IN ; U6111
g3760 nand U6043 DATAO_REG_22__SCAN_IN ; U6112
g3761 nand U2424 EAX_REG_23__SCAN_IN ; U6113
g3762 nand U2385 UWORD_REG_7__SCAN_IN ; U6114
g3763 nand U6043 DATAO_REG_23__SCAN_IN ; U6115
g3764 nand U2424 EAX_REG_24__SCAN_IN ; U6116
g3765 nand U2385 UWORD_REG_8__SCAN_IN ; U6117
g3766 nand U6043 DATAO_REG_24__SCAN_IN ; U6118
g3767 nand U2424 EAX_REG_25__SCAN_IN ; U6119
g3768 nand U2385 UWORD_REG_9__SCAN_IN ; U6120
g3769 nand U6043 DATAO_REG_25__SCAN_IN ; U6121
g3770 nand U2424 EAX_REG_26__SCAN_IN ; U6122
g3771 nand U2385 UWORD_REG_10__SCAN_IN ; U6123
g3772 nand U6043 DATAO_REG_26__SCAN_IN ; U6124
g3773 nand U2424 EAX_REG_27__SCAN_IN ; U6125
g3774 nand U2385 UWORD_REG_11__SCAN_IN ; U6126
g3775 nand U6043 DATAO_REG_27__SCAN_IN ; U6127
g3776 nand U2424 EAX_REG_28__SCAN_IN ; U6128
g3777 nand U2385 UWORD_REG_12__SCAN_IN ; U6129
g3778 nand U6043 DATAO_REG_28__SCAN_IN ; U6130
g3779 nand U2424 EAX_REG_29__SCAN_IN ; U6131
g3780 nand U2385 UWORD_REG_13__SCAN_IN ; U6132
g3781 nand U6043 DATAO_REG_29__SCAN_IN ; U6133
g3782 nand U2424 EAX_REG_30__SCAN_IN ; U6134
g3783 nand U2385 UWORD_REG_14__SCAN_IN ; U6135
g3784 nand U6043 DATAO_REG_30__SCAN_IN ; U6136
g3785 nand U4182 U2447 GTE_485_U6 ; U6137
g3786 nand U4242 U4185 U4182 ; U6138
g3787 nand U4188 U3270 R2167_U17 ; U6139
g3788 nand U7491 U3244 ; U6140
g3789 nand U3871 U6140 ; U6141
g3790 nand U2422 DATAI_0_ ; U6142
g3791 nand U2386 R2358_U82 ; U6143
g3792 nand U3411 EAX_REG_0__SCAN_IN ; U6144
g3793 nand U2422 DATAI_1_ ; U6145
g3794 nand U2386 R2358_U112 ; U6146
g3795 nand U3411 EAX_REG_1__SCAN_IN ; U6147
g3796 nand U2422 DATAI_2_ ; U6148
g3797 nand U2386 R2358_U19 ; U6149
g3798 nand U3411 EAX_REG_2__SCAN_IN ; U6150
g3799 nand U2422 DATAI_3_ ; U6151
g3800 nand U2386 R2358_U20 ; U6152
g3801 nand U3411 EAX_REG_3__SCAN_IN ; U6153
g3802 nand U2422 DATAI_4_ ; U6154
g3803 nand U2386 R2358_U90 ; U6155
g3804 nand U3411 EAX_REG_4__SCAN_IN ; U6156
g3805 nand U2422 DATAI_5_ ; U6157
g3806 nand U2386 R2358_U88 ; U6158
g3807 nand U3411 EAX_REG_5__SCAN_IN ; U6159
g3808 nand U2422 DATAI_6_ ; U6160
g3809 nand U2386 R2358_U86 ; U6161
g3810 nand U3411 EAX_REG_6__SCAN_IN ; U6162
g3811 nand U2422 DATAI_7_ ; U6163
g3812 nand U2386 R2358_U21 ; U6164
g3813 nand U3411 EAX_REG_7__SCAN_IN ; U6165
g3814 nand U2422 DATAI_8_ ; U6166
g3815 nand U2386 R2358_U85 ; U6167
g3816 nand U3411 EAX_REG_8__SCAN_IN ; U6168
g3817 nand U2422 DATAI_9_ ; U6169
g3818 nand U2386 R2358_U83 ; U6170
g3819 nand U3411 EAX_REG_9__SCAN_IN ; U6171
g3820 nand U2422 DATAI_10_ ; U6172
g3821 nand U2386 R2358_U14 ; U6173
g3822 nand U3411 EAX_REG_10__SCAN_IN ; U6174
g3823 nand U2422 DATAI_11_ ; U6175
g3824 nand U2386 R2358_U15 ; U6176
g3825 nand U3411 EAX_REG_11__SCAN_IN ; U6177
g3826 nand U2422 DATAI_12_ ; U6178
g3827 nand U2386 R2358_U122 ; U6179
g3828 nand U3411 EAX_REG_12__SCAN_IN ; U6180
g3829 nand U2422 DATAI_13_ ; U6181
g3830 nand U2386 R2358_U120 ; U6182
g3831 nand U3411 EAX_REG_13__SCAN_IN ; U6183
g3832 nand U2422 DATAI_14_ ; U6184
g3833 nand U2386 R2358_U119 ; U6185
g3834 nand U3411 EAX_REG_14__SCAN_IN ; U6186
g3835 nand U2422 DATAI_15_ ; U6187
g3836 nand U2386 R2358_U16 ; U6188
g3837 nand U3411 EAX_REG_15__SCAN_IN ; U6189
g3838 nand U2423 DATAI_16_ ; U6190
g3839 nand U2387 DATAI_0_ ; U6191
g3840 nand U2386 R2358_U17 ; U6192
g3841 nand U3411 EAX_REG_16__SCAN_IN ; U6193
g3842 nand U2423 DATAI_17_ ; U6194
g3843 nand U2387 DATAI_1_ ; U6195
g3844 nand U2386 R2358_U118 ; U6196
g3845 nand U3411 EAX_REG_17__SCAN_IN ; U6197
g3846 nand U2423 DATAI_18_ ; U6198
g3847 nand U2387 DATAI_2_ ; U6199
g3848 nand U2386 R2358_U116 ; U6200
g3849 nand U3411 EAX_REG_18__SCAN_IN ; U6201
g3850 nand U2423 DATAI_19_ ; U6202
g3851 nand U2387 DATAI_3_ ; U6203
g3852 nand U2386 R2358_U114 ; U6204
g3853 nand U3411 EAX_REG_19__SCAN_IN ; U6205
g3854 nand U2423 DATAI_20_ ; U6206
g3855 nand U2387 DATAI_4_ ; U6207
g3856 nand U2386 R2358_U110 ; U6208
g3857 nand U3411 EAX_REG_20__SCAN_IN ; U6209
g3858 nand U2423 DATAI_21_ ; U6210
g3859 nand U2387 DATAI_5_ ; U6211
g3860 nand U2386 R2358_U18 ; U6212
g3861 nand U3411 EAX_REG_21__SCAN_IN ; U6213
g3862 nand U2423 DATAI_22_ ; U6214
g3863 nand U2387 DATAI_6_ ; U6215
g3864 nand U2386 R2358_U109 ; U6216
g3865 nand U3411 EAX_REG_22__SCAN_IN ; U6217
g3866 nand U2423 DATAI_23_ ; U6218
g3867 nand U2387 DATAI_7_ ; U6219
g3868 nand U2386 R2358_U107 ; U6220
g3869 nand U3411 EAX_REG_23__SCAN_IN ; U6221
g3870 nand U2423 DATAI_24_ ; U6222
g3871 nand U2387 DATAI_8_ ; U6223
g3872 nand U2386 R2358_U105 ; U6224
g3873 nand U3411 EAX_REG_24__SCAN_IN ; U6225
g3874 nand U2423 DATAI_25_ ; U6226
g3875 nand U2387 DATAI_9_ ; U6227
g3876 nand U2386 R2358_U103 ; U6228
g3877 nand U3411 EAX_REG_25__SCAN_IN ; U6229
g3878 nand U2423 DATAI_26_ ; U6230
g3879 nand U2387 DATAI_10_ ; U6231
g3880 nand U2386 R2358_U101 ; U6232
g3881 nand U3411 EAX_REG_26__SCAN_IN ; U6233
g3882 nand U2423 DATAI_27_ ; U6234
g3883 nand U2387 DATAI_11_ ; U6235
g3884 nand U2386 R2358_U99 ; U6236
g3885 nand U3411 EAX_REG_27__SCAN_IN ; U6237
g3886 nand U2423 DATAI_28_ ; U6238
g3887 nand U2387 DATAI_12_ ; U6239
g3888 nand U2386 R2358_U97 ; U6240
g3889 nand U3411 EAX_REG_28__SCAN_IN ; U6241
g3890 nand U2423 DATAI_29_ ; U6242
g3891 nand U2387 DATAI_13_ ; U6243
g3892 nand U2386 R2358_U95 ; U6244
g3893 nand U3411 EAX_REG_29__SCAN_IN ; U6245
g3894 nand U2423 DATAI_30_ ; U6246
g3895 nand U2387 DATAI_14_ ; U6247
g3896 nand U2386 R2358_U93 ; U6248
g3897 nand U3411 EAX_REG_30__SCAN_IN ; U6249
g3898 nand U2423 DATAI_31_ ; U6250
g3899 nand U4186 U3260 ; U6251
g3900 nand U4193 U6251 ; U6252
g3901 nand U2383 R2358_U82 ; U6253
g3902 nand U2371 R2099_U86 ; U6254
g3903 nand U3413 EBX_REG_0__SCAN_IN ; U6255
g3904 nand U2383 R2358_U112 ; U6256
g3905 nand U2371 R2099_U87 ; U6257
g3906 nand U3413 EBX_REG_1__SCAN_IN ; U6258
g3907 nand U2383 R2358_U19 ; U6259
g3908 nand U2371 R2099_U138 ; U6260
g3909 nand U3413 EBX_REG_2__SCAN_IN ; U6261
g3910 nand U2383 R2358_U20 ; U6262
g3911 nand U2371 R2099_U42 ; U6263
g3912 nand U3413 EBX_REG_3__SCAN_IN ; U6264
g3913 nand U2383 R2358_U90 ; U6265
g3914 nand U2371 R2099_U41 ; U6266
g3915 nand U3413 EBX_REG_4__SCAN_IN ; U6267
g3916 nand U2383 R2358_U88 ; U6268
g3917 nand U2371 R2099_U40 ; U6269
g3918 nand U3413 EBX_REG_5__SCAN_IN ; U6270
g3919 nand U2383 R2358_U86 ; U6271
g3920 nand U2371 R2099_U39 ; U6272
g3921 nand U3413 EBX_REG_6__SCAN_IN ; U6273
g3922 nand U2383 R2358_U21 ; U6274
g3923 nand U2371 R2099_U38 ; U6275
g3924 nand U3413 EBX_REG_7__SCAN_IN ; U6276
g3925 nand U2383 R2358_U85 ; U6277
g3926 nand U2371 R2099_U37 ; U6278
g3927 nand U3413 EBX_REG_8__SCAN_IN ; U6279
g3928 nand U2383 R2358_U83 ; U6280
g3929 nand U2371 R2099_U36 ; U6281
g3930 nand U3413 EBX_REG_9__SCAN_IN ; U6282
g3931 nand U2383 R2358_U14 ; U6283
g3932 nand U2371 R2099_U85 ; U6284
g3933 nand U3413 EBX_REG_10__SCAN_IN ; U6285
g3934 nand U2383 R2358_U15 ; U6286
g3935 nand U2371 R2099_U84 ; U6287
g3936 nand U3413 EBX_REG_11__SCAN_IN ; U6288
g3937 nand U2383 R2358_U122 ; U6289
g3938 nand U2371 R2099_U83 ; U6290
g3939 nand U3413 EBX_REG_12__SCAN_IN ; U6291
g3940 nand U2383 R2358_U120 ; U6292
g3941 nand U2371 R2099_U82 ; U6293
g3942 nand U3413 EBX_REG_13__SCAN_IN ; U6294
g3943 nand U2383 R2358_U119 ; U6295
g3944 nand U2371 R2099_U81 ; U6296
g3945 nand U3413 EBX_REG_14__SCAN_IN ; U6297
g3946 nand U2383 R2358_U16 ; U6298
g3947 nand U2371 R2099_U80 ; U6299
g3948 nand U3413 EBX_REG_15__SCAN_IN ; U6300
g3949 nand U2383 R2358_U17 ; U6301
g3950 nand U2371 R2099_U79 ; U6302
g3951 nand U3413 EBX_REG_16__SCAN_IN ; U6303
g3952 nand U2383 R2358_U118 ; U6304
g3953 nand U2371 R2099_U78 ; U6305
g3954 nand U3413 EBX_REG_17__SCAN_IN ; U6306
g3955 nand U2383 R2358_U116 ; U6307
g3956 nand U2371 R2099_U77 ; U6308
g3957 nand U3413 EBX_REG_18__SCAN_IN ; U6309
g3958 nand U2383 R2358_U114 ; U6310
g3959 nand U2371 R2099_U76 ; U6311
g3960 nand U3413 EBX_REG_19__SCAN_IN ; U6312
g3961 nand U2383 R2358_U110 ; U6313
g3962 nand U2371 R2099_U75 ; U6314
g3963 nand U3413 EBX_REG_20__SCAN_IN ; U6315
g3964 nand U2383 R2358_U18 ; U6316
g3965 nand U2371 R2099_U74 ; U6317
g3966 nand U3413 EBX_REG_21__SCAN_IN ; U6318
g3967 nand U2383 R2358_U109 ; U6319
g3968 nand U2371 R2099_U73 ; U6320
g3969 nand U3413 EBX_REG_22__SCAN_IN ; U6321
g3970 nand U2383 R2358_U107 ; U6322
g3971 nand U2371 R2099_U72 ; U6323
g3972 nand U3413 EBX_REG_23__SCAN_IN ; U6324
g3973 nand U2383 R2358_U105 ; U6325
g3974 nand U2371 R2099_U71 ; U6326
g3975 nand U3413 EBX_REG_24__SCAN_IN ; U6327
g3976 nand U2383 R2358_U103 ; U6328
g3977 nand U2371 R2099_U70 ; U6329
g3978 nand U3413 EBX_REG_25__SCAN_IN ; U6330
g3979 nand U2383 R2358_U101 ; U6331
g3980 nand U2371 R2099_U69 ; U6332
g3981 nand U3413 EBX_REG_26__SCAN_IN ; U6333
g3982 nand U2383 R2358_U99 ; U6334
g3983 nand U2371 R2099_U68 ; U6335
g3984 nand U3413 EBX_REG_27__SCAN_IN ; U6336
g3985 nand U2383 R2358_U97 ; U6337
g3986 nand U2371 R2099_U67 ; U6338
g3987 nand U3413 EBX_REG_28__SCAN_IN ; U6339
g3988 nand U2383 R2358_U95 ; U6340
g3989 nand U2371 R2099_U66 ; U6341
g3990 nand U3413 EBX_REG_29__SCAN_IN ; U6342
g3991 nand U2383 R2358_U93 ; U6343
g3992 nand U2371 R2099_U65 ; U6344
g3993 nand U3413 EBX_REG_30__SCAN_IN ; U6345
g3994 nand U2371 R2099_U64 ; U6346
g3995 nand U3413 EBX_REG_31__SCAN_IN ; U6347
g3996 nand U4192 GTE_485_U6 ; U6348
g3997 nand U4190 R2167_U17 ; U6349
g3998 nand U4191 U3250 ; U6350
g3999 not U3418 ; U6351
g4000 nand U4237 STATE2_REG_2__SCAN_IN ; U6352
g4001 nand R2337_U58 STATE2_REG_1__SCAN_IN ; U6353
g4002 nand U6353 U6352 ; U6354
g4003 or READY_N STATEBS16_REG_SCAN_IN ; U6355
g4004 nand U2604 R2099_U86 ; U6356
g4005 nand U7473 REIP_REG_0__SCAN_IN ; U6357
g4006 nand U7472 EBX_REG_0__SCAN_IN ; U6358
g4007 nand U2429 R2358_U82 ; U6359
g4008 nand U2426 R2182_U34 ; U6360
g4009 nand U2373 PHYADDRPOINTER_REG_0__SCAN_IN ; U6361
g4010 nand U2366 PHYADDRPOINTER_REG_0__SCAN_IN ; U6362
g4011 nand U6351 REIP_REG_0__SCAN_IN ; U6363
g4012 nand U2604 R2099_U87 ; U6364
g4013 nand R2096_U4 U7473 ; U6365
g4014 nand U7472 EBX_REG_1__SCAN_IN ; U6366
g4015 nand U2429 R2358_U112 ; U6367
g4016 nand U2426 R2182_U33 ; U6368
g4017 nand U2373 PHYADDRPOINTER_REG_1__SCAN_IN ; U6369
g4018 nand U2366 R2337_U5 ; U6370
g4019 nand U6351 REIP_REG_1__SCAN_IN ; U6371
g4020 nand U2604 R2099_U138 ; U6372
g4021 nand R2096_U71 U7473 ; U6373
g4022 nand U7472 EBX_REG_2__SCAN_IN ; U6374
g4023 nand U2429 R2358_U19 ; U6375
g4024 nand U2426 R2182_U42 ; U6376
g4025 nand U2373 PHYADDRPOINTER_REG_2__SCAN_IN ; U6377
g4026 nand U2366 R2337_U60 ; U6378
g4027 nand U6351 REIP_REG_2__SCAN_IN ; U6379
g4028 nand U2604 R2099_U42 ; U6380
g4029 nand R2096_U68 U7473 ; U6381
g4030 nand U7472 EBX_REG_3__SCAN_IN ; U6382
g4031 nand U2429 R2358_U20 ; U6383
g4032 nand U2426 R2182_U25 ; U6384
g4033 nand U2373 PHYADDRPOINTER_REG_3__SCAN_IN ; U6385
g4034 nand U2366 R2337_U57 ; U6386
g4035 nand U6351 REIP_REG_3__SCAN_IN ; U6387
g4036 nand U2604 R2099_U41 ; U6388
g4037 nand R2096_U67 U7473 ; U6389
g4038 nand U7472 EBX_REG_4__SCAN_IN ; U6390
g4039 nand U2429 R2358_U90 ; U6391
g4040 nand U2426 R2182_U24 ; U6392
g4041 nand U2373 PHYADDRPOINTER_REG_4__SCAN_IN ; U6393
g4042 nand U2366 R2337_U56 ; U6394
g4043 nand U6351 REIP_REG_4__SCAN_IN ; U6395
g4044 nand U2604 R2099_U40 ; U6396
g4045 nand R2096_U66 U7473 ; U6397
g4046 nand U7472 EBX_REG_5__SCAN_IN ; U6398
g4047 nand U2429 R2358_U88 ; U6399
g4048 nand R2182_U5 U2426 ; U6400
g4049 nand U2373 PHYADDRPOINTER_REG_5__SCAN_IN ; U6401
g4050 nand U2366 R2337_U55 ; U6402
g4051 nand U6351 REIP_REG_5__SCAN_IN ; U6403
g4052 nand U2604 R2099_U39 ; U6404
g4053 nand R2096_U65 U7473 ; U6405
g4054 nand U7472 EBX_REG_6__SCAN_IN ; U6406
g4055 nand U2373 PHYADDRPOINTER_REG_6__SCAN_IN ; U6407
g4056 nand U2367 R2358_U86 ; U6408
g4057 nand U2366 R2337_U54 ; U6409
g4058 nand U6351 REIP_REG_6__SCAN_IN ; U6410
g4059 nand U2604 R2099_U38 ; U6411
g4060 nand R2096_U64 U7473 ; U6412
g4061 nand U7472 EBX_REG_7__SCAN_IN ; U6413
g4062 nand U2373 PHYADDRPOINTER_REG_7__SCAN_IN ; U6414
g4063 nand U2367 R2358_U21 ; U6415
g4064 nand U2366 R2337_U53 ; U6416
g4065 nand U6351 REIP_REG_7__SCAN_IN ; U6417
g4066 nand U2604 R2099_U37 ; U6418
g4067 nand R2096_U63 U7473 ; U6419
g4068 nand U7472 EBX_REG_8__SCAN_IN ; U6420
g4069 nand U2373 PHYADDRPOINTER_REG_8__SCAN_IN ; U6421
g4070 nand U2367 R2358_U85 ; U6422
g4071 nand U2366 R2337_U52 ; U6423
g4072 nand U6351 REIP_REG_8__SCAN_IN ; U6424
g4073 nand U2604 R2099_U36 ; U6425
g4074 nand R2096_U62 U7473 ; U6426
g4075 nand U7472 EBX_REG_9__SCAN_IN ; U6427
g4076 nand U2373 PHYADDRPOINTER_REG_9__SCAN_IN ; U6428
g4077 nand U2367 R2358_U83 ; U6429
g4078 nand U2366 R2337_U51 ; U6430
g4079 nand U6351 REIP_REG_9__SCAN_IN ; U6431
g4080 nand U2604 R2099_U85 ; U6432
g4081 nand R2096_U91 U7473 ; U6433
g4082 nand U7472 EBX_REG_10__SCAN_IN ; U6434
g4083 nand U2373 PHYADDRPOINTER_REG_10__SCAN_IN ; U6435
g4084 nand U2367 R2358_U14 ; U6436
g4085 nand U2366 R2337_U80 ; U6437
g4086 nand U6351 REIP_REG_10__SCAN_IN ; U6438
g4087 nand U2604 R2099_U84 ; U6439
g4088 nand R2096_U90 U7473 ; U6440
g4089 nand U7472 EBX_REG_11__SCAN_IN ; U6441
g4090 nand U2373 PHYADDRPOINTER_REG_11__SCAN_IN ; U6442
g4091 nand U2367 R2358_U15 ; U6443
g4092 nand U2366 R2337_U79 ; U6444
g4093 nand U6351 REIP_REG_11__SCAN_IN ; U6445
g4094 nand U2604 R2099_U83 ; U6446
g4095 nand R2096_U89 U7473 ; U6447
g4096 nand U7472 EBX_REG_12__SCAN_IN ; U6448
g4097 nand U2373 PHYADDRPOINTER_REG_12__SCAN_IN ; U6449
g4098 nand U2367 R2358_U122 ; U6450
g4099 nand U2366 R2337_U78 ; U6451
g4100 nand U6351 REIP_REG_12__SCAN_IN ; U6452
g4101 nand U2604 R2099_U82 ; U6453
g4102 nand R2096_U88 U7473 ; U6454
g4103 nand U7472 EBX_REG_13__SCAN_IN ; U6455
g4104 nand U2373 PHYADDRPOINTER_REG_13__SCAN_IN ; U6456
g4105 nand U2367 R2358_U120 ; U6457
g4106 nand U2366 R2337_U77 ; U6458
g4107 nand U6351 REIP_REG_13__SCAN_IN ; U6459
g4108 nand U2604 R2099_U81 ; U6460
g4109 nand R2096_U87 U7473 ; U6461
g4110 nand U7472 EBX_REG_14__SCAN_IN ; U6462
g4111 nand U2373 PHYADDRPOINTER_REG_14__SCAN_IN ; U6463
g4112 nand U2367 R2358_U119 ; U6464
g4113 nand U2366 R2337_U76 ; U6465
g4114 nand U6351 REIP_REG_14__SCAN_IN ; U6466
g4115 nand U2604 R2099_U80 ; U6467
g4116 nand R2096_U86 U7473 ; U6468
g4117 nand U7472 EBX_REG_15__SCAN_IN ; U6469
g4118 nand U2373 PHYADDRPOINTER_REG_15__SCAN_IN ; U6470
g4119 nand U2367 R2358_U16 ; U6471
g4120 nand U2366 R2337_U75 ; U6472
g4121 nand U6351 REIP_REG_15__SCAN_IN ; U6473
g4122 nand U2604 R2099_U79 ; U6474
g4123 nand R2096_U85 U7473 ; U6475
g4124 nand U7472 EBX_REG_16__SCAN_IN ; U6476
g4125 nand U2373 PHYADDRPOINTER_REG_16__SCAN_IN ; U6477
g4126 nand U2367 R2358_U17 ; U6478
g4127 nand U2366 R2337_U74 ; U6479
g4128 nand U6351 REIP_REG_16__SCAN_IN ; U6480
g4129 nand U2604 R2099_U78 ; U6481
g4130 nand R2096_U84 U7473 ; U6482
g4131 nand U7472 EBX_REG_17__SCAN_IN ; U6483
g4132 nand U2373 PHYADDRPOINTER_REG_17__SCAN_IN ; U6484
g4133 nand U2367 R2358_U118 ; U6485
g4134 nand U2366 R2337_U73 ; U6486
g4135 nand U6351 REIP_REG_17__SCAN_IN ; U6487
g4136 nand U2604 R2099_U77 ; U6488
g4137 nand R2096_U83 U7473 ; U6489
g4138 nand U7472 EBX_REG_18__SCAN_IN ; U6490
g4139 nand U2373 PHYADDRPOINTER_REG_18__SCAN_IN ; U6491
g4140 nand U2367 R2358_U116 ; U6492
g4141 nand U2366 R2337_U72 ; U6493
g4142 nand U6351 REIP_REG_18__SCAN_IN ; U6494
g4143 nand U2604 R2099_U76 ; U6495
g4144 nand R2096_U82 U7473 ; U6496
g4145 nand U7472 EBX_REG_19__SCAN_IN ; U6497
g4146 nand U2373 PHYADDRPOINTER_REG_19__SCAN_IN ; U6498
g4147 nand U2367 R2358_U114 ; U6499
g4148 nand U2366 R2337_U71 ; U6500
g4149 nand U6351 REIP_REG_19__SCAN_IN ; U6501
g4150 nand U2604 R2099_U75 ; U6502
g4151 nand R2096_U81 U7473 ; U6503
g4152 nand U7472 EBX_REG_20__SCAN_IN ; U6504
g4153 nand U2373 PHYADDRPOINTER_REG_20__SCAN_IN ; U6505
g4154 nand U2367 R2358_U110 ; U6506
g4155 nand U2366 R2337_U70 ; U6507
g4156 nand U6351 REIP_REG_20__SCAN_IN ; U6508
g4157 nand U2604 R2099_U74 ; U6509
g4158 nand R2096_U80 U7473 ; U6510
g4159 nand U7472 EBX_REG_21__SCAN_IN ; U6511
g4160 nand U2373 PHYADDRPOINTER_REG_21__SCAN_IN ; U6512
g4161 nand U2367 R2358_U18 ; U6513
g4162 nand U2366 R2337_U69 ; U6514
g4163 nand U6351 REIP_REG_21__SCAN_IN ; U6515
g4164 nand U2604 R2099_U73 ; U6516
g4165 nand R2096_U79 U7473 ; U6517
g4166 nand U7472 EBX_REG_22__SCAN_IN ; U6518
g4167 nand U2373 PHYADDRPOINTER_REG_22__SCAN_IN ; U6519
g4168 nand U2367 R2358_U109 ; U6520
g4169 nand U2366 R2337_U68 ; U6521
g4170 nand U6351 REIP_REG_22__SCAN_IN ; U6522
g4171 nand U2604 R2099_U72 ; U6523
g4172 nand R2096_U78 U7473 ; U6524
g4173 nand U7472 EBX_REG_23__SCAN_IN ; U6525
g4174 nand U2373 PHYADDRPOINTER_REG_23__SCAN_IN ; U6526
g4175 nand U2367 R2358_U107 ; U6527
g4176 nand U2366 R2337_U67 ; U6528
g4177 nand U6351 REIP_REG_23__SCAN_IN ; U6529
g4178 nand U2604 R2099_U71 ; U6530
g4179 nand R2096_U77 U7473 ; U6531
g4180 nand U7472 EBX_REG_24__SCAN_IN ; U6532
g4181 nand U2373 PHYADDRPOINTER_REG_24__SCAN_IN ; U6533
g4182 nand U2367 R2358_U105 ; U6534
g4183 nand U2366 R2337_U66 ; U6535
g4184 nand U6351 REIP_REG_24__SCAN_IN ; U6536
g4185 nand U2604 R2099_U70 ; U6537
g4186 nand R2096_U76 U7473 ; U6538
g4187 nand U7472 EBX_REG_25__SCAN_IN ; U6539
g4188 nand U2373 PHYADDRPOINTER_REG_25__SCAN_IN ; U6540
g4189 nand U2367 R2358_U103 ; U6541
g4190 nand U2366 R2337_U65 ; U6542
g4191 nand U6351 REIP_REG_25__SCAN_IN ; U6543
g4192 nand U2604 R2099_U69 ; U6544
g4193 nand R2096_U75 U7473 ; U6545
g4194 nand U7472 EBX_REG_26__SCAN_IN ; U6546
g4195 nand U2373 PHYADDRPOINTER_REG_26__SCAN_IN ; U6547
g4196 nand U2367 R2358_U101 ; U6548
g4197 nand U2366 R2337_U64 ; U6549
g4198 nand U6351 REIP_REG_26__SCAN_IN ; U6550
g4199 nand U2604 R2099_U68 ; U6551
g4200 nand R2096_U74 U7473 ; U6552
g4201 nand U7472 EBX_REG_27__SCAN_IN ; U6553
g4202 nand U2373 PHYADDRPOINTER_REG_27__SCAN_IN ; U6554
g4203 nand U2367 R2358_U99 ; U6555
g4204 nand U2366 R2337_U63 ; U6556
g4205 nand U6351 REIP_REG_27__SCAN_IN ; U6557
g4206 nand U2604 R2099_U67 ; U6558
g4207 nand R2096_U73 U7473 ; U6559
g4208 nand U7472 EBX_REG_28__SCAN_IN ; U6560
g4209 nand U2373 PHYADDRPOINTER_REG_28__SCAN_IN ; U6561
g4210 nand U2367 R2358_U97 ; U6562
g4211 nand U2366 R2337_U62 ; U6563
g4212 nand U6351 REIP_REG_28__SCAN_IN ; U6564
g4213 nand U2604 R2099_U66 ; U6565
g4214 nand R2096_U72 U7473 ; U6566
g4215 nand U7472 EBX_REG_29__SCAN_IN ; U6567
g4216 nand U2373 PHYADDRPOINTER_REG_29__SCAN_IN ; U6568
g4217 nand U2367 R2358_U95 ; U6569
g4218 nand U2366 R2337_U61 ; U6570
g4219 nand U6351 REIP_REG_29__SCAN_IN ; U6571
g4220 nand U2604 R2099_U65 ; U6572
g4221 nand R2096_U70 U7473 ; U6573
g4222 nand U7472 EBX_REG_30__SCAN_IN ; U6574
g4223 nand U2373 PHYADDRPOINTER_REG_30__SCAN_IN ; U6575
g4224 nand U2367 R2358_U93 ; U6576
g4225 nand U2366 R2337_U59 ; U6577
g4226 nand U6351 REIP_REG_30__SCAN_IN ; U6578
g4227 nand U2604 R2099_U64 ; U6579
g4228 nand R2096_U69 U7473 ; U6580
g4229 nand U7472 EBX_REG_31__SCAN_IN ; U6581
g4230 nand U2373 PHYADDRPOINTER_REG_31__SCAN_IN ; U6582
g4231 nand U2367 R2358_U91 ; U6583
g4232 nand U2366 R2337_U58 ; U6584
g4233 nand U6351 REIP_REG_31__SCAN_IN ; U6585
g4234 nand DATAWIDTH_REG_0__SCAN_IN DATAWIDTH_REG_1__SCAN_IN ; U6586
g4235 or REIP_REG_0__SCAN_IN REIP_REG_1__SCAN_IN ; U6587
g4236 not U4165 ; U6588
g4237 nand U4165 FLUSH_REG_SCAN_IN ; U6589
g4238 nand U3954 U2428 ; U6590
g4239 not U4168 ; U6591
g4240 nand U4485 STATEBS16_REG_SCAN_IN ; U6592
g4241 nand U4196 U6592 ; U6593
g4242 nand U3952 U6593 ; U6594
g4243 nand U6594 STATE2_REG_0__SCAN_IN ; U6595
g4244 nand U4181 U3259 ; U6596
g4245 nand U3953 U6595 ; U6597
g4246 nand U2368 U2473 ; U6598
g4247 nand U6598 CODEFETCH_REG_SCAN_IN ; U6599
g4248 nand U4243 STATE2_REG_0__SCAN_IN ; U6600
g4249 nand STATE_REG_0__SCAN_IN ADS_N_REG_SCAN_IN ; U6601
g4250 not U4169 ; U6602
g4251 nand U3956 U3278 ; U6603
g4252 nand U4487 U3957 U3393 ; U6604
g4253 nand U6604 MEMORYFETCH_REG_SCAN_IN ; U6605
g4254 nand U2544 INSTQUEUE_REG_15__7__SCAN_IN ; U6606
g4255 nand U2543 INSTQUEUE_REG_14__7__SCAN_IN ; U6607
g4256 nand U2542 INSTQUEUE_REG_13__7__SCAN_IN ; U6608
g4257 nand U2541 INSTQUEUE_REG_12__7__SCAN_IN ; U6609
g4258 nand U2539 INSTQUEUE_REG_11__7__SCAN_IN ; U6610
g4259 nand U2538 INSTQUEUE_REG_10__7__SCAN_IN ; U6611
g4260 nand U2537 INSTQUEUE_REG_9__7__SCAN_IN ; U6612
g4261 nand U2536 INSTQUEUE_REG_8__7__SCAN_IN ; U6613
g4262 nand U2534 INSTQUEUE_REG_7__7__SCAN_IN ; U6614
g4263 nand U2533 INSTQUEUE_REG_6__7__SCAN_IN ; U6615
g4264 nand U2532 INSTQUEUE_REG_5__7__SCAN_IN ; U6616
g4265 nand U2531 INSTQUEUE_REG_4__7__SCAN_IN ; U6617
g4266 nand U2529 INSTQUEUE_REG_3__7__SCAN_IN ; U6618
g4267 nand U2527 INSTQUEUE_REG_2__7__SCAN_IN ; U6619
g4268 nand U2525 INSTQUEUE_REG_1__7__SCAN_IN ; U6620
g4269 nand U2523 INSTQUEUE_REG_0__7__SCAN_IN ; U6621
g4270 nand U2544 INSTQUEUE_REG_15__6__SCAN_IN ; U6622
g4271 nand U2543 INSTQUEUE_REG_14__6__SCAN_IN ; U6623
g4272 nand U2542 INSTQUEUE_REG_13__6__SCAN_IN ; U6624
g4273 nand U2541 INSTQUEUE_REG_12__6__SCAN_IN ; U6625
g4274 nand U2539 INSTQUEUE_REG_11__6__SCAN_IN ; U6626
g4275 nand U2538 INSTQUEUE_REG_10__6__SCAN_IN ; U6627
g4276 nand U2537 INSTQUEUE_REG_9__6__SCAN_IN ; U6628
g4277 nand U2536 INSTQUEUE_REG_8__6__SCAN_IN ; U6629
g4278 nand U2534 INSTQUEUE_REG_7__6__SCAN_IN ; U6630
g4279 nand U2533 INSTQUEUE_REG_6__6__SCAN_IN ; U6631
g4280 nand U2532 INSTQUEUE_REG_5__6__SCAN_IN ; U6632
g4281 nand U2531 INSTQUEUE_REG_4__6__SCAN_IN ; U6633
g4282 nand U2529 INSTQUEUE_REG_3__6__SCAN_IN ; U6634
g4283 nand U2527 INSTQUEUE_REG_2__6__SCAN_IN ; U6635
g4284 nand U2525 INSTQUEUE_REG_1__6__SCAN_IN ; U6636
g4285 nand U2523 INSTQUEUE_REG_0__6__SCAN_IN ; U6637
g4286 nand U2544 INSTQUEUE_REG_15__5__SCAN_IN ; U6638
g4287 nand U2543 INSTQUEUE_REG_14__5__SCAN_IN ; U6639
g4288 nand U2542 INSTQUEUE_REG_13__5__SCAN_IN ; U6640
g4289 nand U2541 INSTQUEUE_REG_12__5__SCAN_IN ; U6641
g4290 nand U2539 INSTQUEUE_REG_11__5__SCAN_IN ; U6642
g4291 nand U2538 INSTQUEUE_REG_10__5__SCAN_IN ; U6643
g4292 nand U2537 INSTQUEUE_REG_9__5__SCAN_IN ; U6644
g4293 nand U2536 INSTQUEUE_REG_8__5__SCAN_IN ; U6645
g4294 nand U2534 INSTQUEUE_REG_7__5__SCAN_IN ; U6646
g4295 nand U2533 INSTQUEUE_REG_6__5__SCAN_IN ; U6647
g4296 nand U2532 INSTQUEUE_REG_5__5__SCAN_IN ; U6648
g4297 nand U2531 INSTQUEUE_REG_4__5__SCAN_IN ; U6649
g4298 nand U2529 INSTQUEUE_REG_3__5__SCAN_IN ; U6650
g4299 nand U2527 INSTQUEUE_REG_2__5__SCAN_IN ; U6651
g4300 nand U2525 INSTQUEUE_REG_1__5__SCAN_IN ; U6652
g4301 nand U2523 INSTQUEUE_REG_0__5__SCAN_IN ; U6653
g4302 nand U2544 INSTQUEUE_REG_15__4__SCAN_IN ; U6654
g4303 nand U2543 INSTQUEUE_REG_14__4__SCAN_IN ; U6655
g4304 nand U2542 INSTQUEUE_REG_13__4__SCAN_IN ; U6656
g4305 nand U2541 INSTQUEUE_REG_12__4__SCAN_IN ; U6657
g4306 nand U2539 INSTQUEUE_REG_11__4__SCAN_IN ; U6658
g4307 nand U2538 INSTQUEUE_REG_10__4__SCAN_IN ; U6659
g4308 nand U2537 INSTQUEUE_REG_9__4__SCAN_IN ; U6660
g4309 nand U2536 INSTQUEUE_REG_8__4__SCAN_IN ; U6661
g4310 nand U2534 INSTQUEUE_REG_7__4__SCAN_IN ; U6662
g4311 nand U2533 INSTQUEUE_REG_6__4__SCAN_IN ; U6663
g4312 nand U2532 INSTQUEUE_REG_5__4__SCAN_IN ; U6664
g4313 nand U2531 INSTQUEUE_REG_4__4__SCAN_IN ; U6665
g4314 nand U2529 INSTQUEUE_REG_3__4__SCAN_IN ; U6666
g4315 nand U2527 INSTQUEUE_REG_2__4__SCAN_IN ; U6667
g4316 nand U2525 INSTQUEUE_REG_1__4__SCAN_IN ; U6668
g4317 nand U2544 INSTQUEUE_REG_15__3__SCAN_IN ; U6669
g4318 nand U2543 INSTQUEUE_REG_14__3__SCAN_IN ; U6670
g4319 nand U2542 INSTQUEUE_REG_13__3__SCAN_IN ; U6671
g4320 nand U2541 INSTQUEUE_REG_12__3__SCAN_IN ; U6672
g4321 nand U2539 INSTQUEUE_REG_11__3__SCAN_IN ; U6673
g4322 nand U2538 INSTQUEUE_REG_10__3__SCAN_IN ; U6674
g4323 nand U2537 INSTQUEUE_REG_9__3__SCAN_IN ; U6675
g4324 nand U2536 INSTQUEUE_REG_8__3__SCAN_IN ; U6676
g4325 nand U2534 INSTQUEUE_REG_7__3__SCAN_IN ; U6677
g4326 nand U2533 INSTQUEUE_REG_6__3__SCAN_IN ; U6678
g4327 nand U2532 INSTQUEUE_REG_5__3__SCAN_IN ; U6679
g4328 nand U2531 INSTQUEUE_REG_4__3__SCAN_IN ; U6680
g4329 nand U2529 INSTQUEUE_REG_3__3__SCAN_IN ; U6681
g4330 nand U2527 INSTQUEUE_REG_2__3__SCAN_IN ; U6682
g4331 nand U2525 INSTQUEUE_REG_1__3__SCAN_IN ; U6683
g4332 nand U2523 INSTQUEUE_REG_0__3__SCAN_IN ; U6684
g4333 nand U2544 INSTQUEUE_REG_15__2__SCAN_IN ; U6685
g4334 nand U2543 INSTQUEUE_REG_14__2__SCAN_IN ; U6686
g4335 nand U2542 INSTQUEUE_REG_13__2__SCAN_IN ; U6687
g4336 nand U2541 INSTQUEUE_REG_12__2__SCAN_IN ; U6688
g4337 nand U2539 INSTQUEUE_REG_11__2__SCAN_IN ; U6689
g4338 nand U2538 INSTQUEUE_REG_10__2__SCAN_IN ; U6690
g4339 nand U2537 INSTQUEUE_REG_9__2__SCAN_IN ; U6691
g4340 nand U2536 INSTQUEUE_REG_8__2__SCAN_IN ; U6692
g4341 nand U2534 INSTQUEUE_REG_7__2__SCAN_IN ; U6693
g4342 nand U2533 INSTQUEUE_REG_6__2__SCAN_IN ; U6694
g4343 nand U2532 INSTQUEUE_REG_5__2__SCAN_IN ; U6695
g4344 nand U2531 INSTQUEUE_REG_4__2__SCAN_IN ; U6696
g4345 nand U2529 INSTQUEUE_REG_3__2__SCAN_IN ; U6697
g4346 nand U2527 INSTQUEUE_REG_2__2__SCAN_IN ; U6698
g4347 nand U2525 INSTQUEUE_REG_1__2__SCAN_IN ; U6699
g4348 nand U2523 INSTQUEUE_REG_0__2__SCAN_IN ; U6700
g4349 nand U2544 INSTQUEUE_REG_15__1__SCAN_IN ; U6701
g4350 nand U2543 INSTQUEUE_REG_14__1__SCAN_IN ; U6702
g4351 nand U2542 INSTQUEUE_REG_13__1__SCAN_IN ; U6703
g4352 nand U2541 INSTQUEUE_REG_12__1__SCAN_IN ; U6704
g4353 nand U2539 INSTQUEUE_REG_11__1__SCAN_IN ; U6705
g4354 nand U2538 INSTQUEUE_REG_10__1__SCAN_IN ; U6706
g4355 nand U2537 INSTQUEUE_REG_9__1__SCAN_IN ; U6707
g4356 nand U2536 INSTQUEUE_REG_8__1__SCAN_IN ; U6708
g4357 nand U2534 INSTQUEUE_REG_7__1__SCAN_IN ; U6709
g4358 nand U2533 INSTQUEUE_REG_6__1__SCAN_IN ; U6710
g4359 nand U2532 INSTQUEUE_REG_5__1__SCAN_IN ; U6711
g4360 nand U2531 INSTQUEUE_REG_4__1__SCAN_IN ; U6712
g4361 nand U2529 INSTQUEUE_REG_3__1__SCAN_IN ; U6713
g4362 nand U2527 INSTQUEUE_REG_2__1__SCAN_IN ; U6714
g4363 nand U2525 INSTQUEUE_REG_1__1__SCAN_IN ; U6715
g4364 nand U2523 INSTQUEUE_REG_0__1__SCAN_IN ; U6716
g4365 nand U2544 INSTQUEUE_REG_15__0__SCAN_IN ; U6717
g4366 nand U2543 INSTQUEUE_REG_14__0__SCAN_IN ; U6718
g4367 nand U2542 INSTQUEUE_REG_13__0__SCAN_IN ; U6719
g4368 nand U2541 INSTQUEUE_REG_12__0__SCAN_IN ; U6720
g4369 nand U2539 INSTQUEUE_REG_11__0__SCAN_IN ; U6721
g4370 nand U2538 INSTQUEUE_REG_10__0__SCAN_IN ; U6722
g4371 nand U2537 INSTQUEUE_REG_9__0__SCAN_IN ; U6723
g4372 nand U2536 INSTQUEUE_REG_8__0__SCAN_IN ; U6724
g4373 nand U2534 INSTQUEUE_REG_7__0__SCAN_IN ; U6725
g4374 nand U2533 INSTQUEUE_REG_6__0__SCAN_IN ; U6726
g4375 nand U2532 INSTQUEUE_REG_5__0__SCAN_IN ; U6727
g4376 nand U2531 INSTQUEUE_REG_4__0__SCAN_IN ; U6728
g4377 nand U2529 INSTQUEUE_REG_3__0__SCAN_IN ; U6729
g4378 nand U2527 INSTQUEUE_REG_2__0__SCAN_IN ; U6730
g4379 nand U2525 INSTQUEUE_REG_1__0__SCAN_IN ; U6731
g4380 nand U2523 INSTQUEUE_REG_0__0__SCAN_IN ; U6732
g4381 nand U4448 STATE2_REG_2__SCAN_IN ; U6733
g4382 nand U3399 U6733 ; U6734
g4383 nand U4176 EAX_REG_9__SCAN_IN ; U6735
g4384 nand U4175 PHYADDRPOINTER_REG_9__SCAN_IN ; U6736
g4385 nand R2337_U51 U2352 ; U6737
g4386 nand U4176 EAX_REG_8__SCAN_IN ; U6738
g4387 nand U4175 PHYADDRPOINTER_REG_8__SCAN_IN ; U6739
g4388 nand R2337_U52 U2352 ; U6740
g4389 nand U4176 EAX_REG_7__SCAN_IN ; U6741
g4390 nand U4175 PHYADDRPOINTER_REG_7__SCAN_IN ; U6742
g4391 nand R2337_U53 U2352 ; U6743
g4392 nand U4176 EAX_REG_6__SCAN_IN ; U6744
g4393 nand U4175 PHYADDRPOINTER_REG_6__SCAN_IN ; U6745
g4394 nand R2337_U54 U2352 ; U6746
g4395 nand R2182_U5 U6734 ; U6747
g4396 nand U4176 EAX_REG_5__SCAN_IN ; U6748
g4397 nand U4175 PHYADDRPOINTER_REG_5__SCAN_IN ; U6749
g4398 nand R2337_U55 U2352 ; U6750
g4399 nand R2182_U24 U6734 ; U6751
g4400 nand U4176 EAX_REG_4__SCAN_IN ; U6752
g4401 nand U4175 PHYADDRPOINTER_REG_4__SCAN_IN ; U6753
g4402 nand R2337_U56 U2352 ; U6754
g4403 nand U2353 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; U6755
g4404 nand U4176 EAX_REG_31__SCAN_IN ; U6756
g4405 nand U4175 PHYADDRPOINTER_REG_31__SCAN_IN ; U6757
g4406 nand R2337_U58 U2352 ; U6758
g4407 nand R2182_U26 U6734 ; U6759
g4408 nand U4176 EAX_REG_30__SCAN_IN ; U6760
g4409 nand U4175 PHYADDRPOINTER_REG_30__SCAN_IN ; U6761
g4410 nand R2337_U59 U2352 ; U6762
g4411 nand R2182_U25 U6734 ; U6763
g4412 nand U4176 EAX_REG_3__SCAN_IN ; U6764
g4413 nand U4175 PHYADDRPOINTER_REG_3__SCAN_IN ; U6765
g4414 nand R2337_U57 U2352 ; U6766
g4415 nand U2353 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U6767
g4416 nand R2182_U27 U6734 ; U6768
g4417 nand U4176 EAX_REG_29__SCAN_IN ; U6769
g4418 nand U4175 PHYADDRPOINTER_REG_29__SCAN_IN ; U6770
g4419 nand R2337_U61 U2352 ; U6771
g4420 nand R2182_U28 U6734 ; U6772
g4421 nand U4176 EAX_REG_28__SCAN_IN ; U6773
g4422 nand U4175 PHYADDRPOINTER_REG_28__SCAN_IN ; U6774
g4423 nand R2337_U62 U2352 ; U6775
g4424 nand R2182_U29 U6734 ; U6776
g4425 nand U4176 EAX_REG_27__SCAN_IN ; U6777
g4426 nand U4175 PHYADDRPOINTER_REG_27__SCAN_IN ; U6778
g4427 nand R2337_U63 U2352 ; U6779
g4428 nand R2182_U30 U6734 ; U6780
g4429 nand U4176 EAX_REG_26__SCAN_IN ; U6781
g4430 nand U4175 PHYADDRPOINTER_REG_26__SCAN_IN ; U6782
g4431 nand R2337_U64 U2352 ; U6783
g4432 nand R2182_U31 U6734 ; U6784
g4433 nand U4176 EAX_REG_25__SCAN_IN ; U6785
g4434 nand U4175 PHYADDRPOINTER_REG_25__SCAN_IN ; U6786
g4435 nand R2337_U65 U2352 ; U6787
g4436 nand R2182_U32 U6734 ; U6788
g4437 nand U4176 EAX_REG_24__SCAN_IN ; U6789
g4438 nand U4175 PHYADDRPOINTER_REG_24__SCAN_IN ; U6790
g4439 nand R2337_U66 U2352 ; U6791
g4440 nand R2182_U6 U6734 ; U6792
g4441 nand U4176 EAX_REG_23__SCAN_IN ; U6793
g4442 nand U4175 PHYADDRPOINTER_REG_23__SCAN_IN ; U6794
g4443 nand R2337_U67 U2352 ; U6795
g4444 nand U2724 U6734 ; U6796
g4445 nand U4176 EAX_REG_22__SCAN_IN ; U6797
g4446 nand U4175 PHYADDRPOINTER_REG_22__SCAN_IN ; U6798
g4447 nand R2337_U68 U2352 ; U6799
g4448 nand U2725 U6734 ; U6800
g4449 nand U4176 EAX_REG_21__SCAN_IN ; U6801
g4450 nand U4175 PHYADDRPOINTER_REG_21__SCAN_IN ; U6802
g4451 nand R2337_U69 U2352 ; U6803
g4452 nand U2726 U6734 ; U6804
g4453 nand U4176 EAX_REG_20__SCAN_IN ; U6805
g4454 nand U4175 PHYADDRPOINTER_REG_20__SCAN_IN ; U6806
g4455 nand R2337_U70 U2352 ; U6807
g4456 nand R2182_U42 U6734 ; U6808
g4457 nand U4176 EAX_REG_2__SCAN_IN ; U6809
g4458 nand U4175 PHYADDRPOINTER_REG_2__SCAN_IN ; U6810
g4459 nand R2337_U60 U2352 ; U6811
g4460 nand U2353 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U6812
g4461 nand U2727 U6734 ; U6813
g4462 nand U4176 EAX_REG_19__SCAN_IN ; U6814
g4463 nand U4175 PHYADDRPOINTER_REG_19__SCAN_IN ; U6815
g4464 nand R2337_U71 U2352 ; U6816
g4465 nand U2728 U6734 ; U6817
g4466 nand U4176 EAX_REG_18__SCAN_IN ; U6818
g4467 nand U4175 PHYADDRPOINTER_REG_18__SCAN_IN ; U6819
g4468 nand R2337_U72 U2352 ; U6820
g4469 nand U2729 U6734 ; U6821
g4470 nand U4176 EAX_REG_17__SCAN_IN ; U6822
g4471 nand U4175 PHYADDRPOINTER_REG_17__SCAN_IN ; U6823
g4472 nand R2337_U73 U2352 ; U6824
g4473 nand U2730 U6734 ; U6825
g4474 nand U4176 EAX_REG_16__SCAN_IN ; U6826
g4475 nand U4175 PHYADDRPOINTER_REG_16__SCAN_IN ; U6827
g4476 nand R2337_U74 U2352 ; U6828
g4477 nand U4176 EAX_REG_15__SCAN_IN ; U6829
g4478 nand U4175 PHYADDRPOINTER_REG_15__SCAN_IN ; U6830
g4479 nand R2337_U75 U2352 ; U6831
g4480 nand U4176 EAX_REG_14__SCAN_IN ; U6832
g4481 nand U4175 PHYADDRPOINTER_REG_14__SCAN_IN ; U6833
g4482 nand R2337_U76 U2352 ; U6834
g4483 nand U4176 EAX_REG_13__SCAN_IN ; U6835
g4484 nand U4175 PHYADDRPOINTER_REG_13__SCAN_IN ; U6836
g4485 nand R2337_U77 U2352 ; U6837
g4486 nand U4176 EAX_REG_12__SCAN_IN ; U6838
g4487 nand U4175 PHYADDRPOINTER_REG_12__SCAN_IN ; U6839
g4488 nand R2337_U78 U2352 ; U6840
g4489 nand U4176 EAX_REG_11__SCAN_IN ; U6841
g4490 nand U4175 PHYADDRPOINTER_REG_11__SCAN_IN ; U6842
g4491 nand R2337_U79 U2352 ; U6843
g4492 nand U4176 EAX_REG_10__SCAN_IN ; U6844
g4493 nand U4175 PHYADDRPOINTER_REG_10__SCAN_IN ; U6845
g4494 nand R2337_U80 U2352 ; U6846
g4495 nand R2182_U33 U6734 ; U6847
g4496 nand U4176 EAX_REG_1__SCAN_IN ; U6848
g4497 nand U4175 PHYADDRPOINTER_REG_1__SCAN_IN ; U6849
g4498 nand R2337_U5 U2352 ; U6850
g4499 nand U2353 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U6851
g4500 nand R2182_U34 U6734 ; U6852
g4501 nand U4176 EAX_REG_0__SCAN_IN ; U6853
g4502 nand U4175 PHYADDRPOINTER_REG_0__SCAN_IN ; U6854
g4503 nand U2352 PHYADDRPOINTER_REG_0__SCAN_IN ; U6855
g4504 nand U2353 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U6856
g4505 nand R2144_U49 U6734 ; U6857
g4506 nand U3426 U4448 U3296 ; U6858
g4507 nand U4147 R2144_U80 ; U6859
g4508 nand ADD_371_U6 U4196 ; U6860
g4509 nand U4147 R2144_U10 ; U6861
g4510 nand ADD_371_U17 U4196 ; U6862
g4511 nand U4147 R2144_U9 ; U6863
g4512 nand ADD_371_U18 U4196 ; U6864
g4513 nand U4147 R2144_U45 ; U6865
g4514 nand ADD_371_U19 U4196 ; U6866
g4515 nand U4147 R2144_U47 ; U6867
g4516 nand ADD_371_U20 U4196 ; U6868
g4517 nand U4147 R2144_U8 ; U6869
g4518 nand ADD_371_U25 U4196 ; U6870
g4519 nand U4147 R2144_U49 ; U6871
g4520 nand ADD_371_U5 U4196 ; U6872
g4521 nand U4482 U3270 ; U6873
g4522 nand U4147 R2144_U50 ; U6874
g4523 nand ADD_371_U21 U4196 ; U6875
g4524 nand U2605 U3271 ; U6876
g4525 nand U4147 R2144_U43 ; U6877
g4526 nand ADD_371_U4 U4196 ; U6878
g4527 nand U4482 U3270 ; U6879
g4528 nand U2564 INSTQUEUE_REG_15__1__SCAN_IN ; U6880
g4529 nand U2563 INSTQUEUE_REG_14__1__SCAN_IN ; U6881
g4530 nand U2562 INSTQUEUE_REG_13__1__SCAN_IN ; U6882
g4531 nand U2561 INSTQUEUE_REG_12__1__SCAN_IN ; U6883
g4532 nand U2559 INSTQUEUE_REG_11__1__SCAN_IN ; U6884
g4533 nand U2558 INSTQUEUE_REG_10__1__SCAN_IN ; U6885
g4534 nand U2557 INSTQUEUE_REG_9__1__SCAN_IN ; U6886
g4535 nand U2556 INSTQUEUE_REG_8__1__SCAN_IN ; U6887
g4536 nand U2554 INSTQUEUE_REG_7__1__SCAN_IN ; U6888
g4537 nand U2553 INSTQUEUE_REG_6__1__SCAN_IN ; U6889
g4538 nand U2552 INSTQUEUE_REG_5__1__SCAN_IN ; U6890
g4539 nand U2551 INSTQUEUE_REG_4__1__SCAN_IN ; U6891
g4540 nand U2549 INSTQUEUE_REG_3__1__SCAN_IN ; U6892
g4541 nand U2548 INSTQUEUE_REG_2__1__SCAN_IN ; U6893
g4542 nand U2547 INSTQUEUE_REG_1__1__SCAN_IN ; U6894
g4543 nand U2546 INSTQUEUE_REG_0__1__SCAN_IN ; U6895
g4544 nand U4020 U4019 U4018 U4017 ; U6896
g4545 nand U3392 U3405 ; U6897
g4546 nand U2564 INSTQUEUE_REG_15__0__SCAN_IN ; U6898
g4547 nand U2563 INSTQUEUE_REG_14__0__SCAN_IN ; U6899
g4548 nand U2562 INSTQUEUE_REG_13__0__SCAN_IN ; U6900
g4549 nand U2561 INSTQUEUE_REG_12__0__SCAN_IN ; U6901
g4550 nand U2559 INSTQUEUE_REG_11__0__SCAN_IN ; U6902
g4551 nand U2558 INSTQUEUE_REG_10__0__SCAN_IN ; U6903
g4552 nand U2557 INSTQUEUE_REG_9__0__SCAN_IN ; U6904
g4553 nand U2556 INSTQUEUE_REG_8__0__SCAN_IN ; U6905
g4554 nand U2554 INSTQUEUE_REG_7__0__SCAN_IN ; U6906
g4555 nand U2553 INSTQUEUE_REG_6__0__SCAN_IN ; U6907
g4556 nand U2552 INSTQUEUE_REG_5__0__SCAN_IN ; U6908
g4557 nand U2551 INSTQUEUE_REG_4__0__SCAN_IN ; U6909
g4558 nand U2549 INSTQUEUE_REG_3__0__SCAN_IN ; U6910
g4559 nand U2548 INSTQUEUE_REG_2__0__SCAN_IN ; U6911
g4560 nand U2547 INSTQUEUE_REG_1__0__SCAN_IN ; U6912
g4561 nand U2546 INSTQUEUE_REG_0__0__SCAN_IN ; U6913
g4562 nand U4024 U4023 U4022 U4021 ; U6914
g4563 nand U4195 U3221 ; U6915
g4564 nand U2355 SUB_357_U8 ; U6916
g4565 nand U4195 U3220 ; U6917
g4566 nand SUB_357_U6 U2355 ; U6918
g4567 nand U4195 U3219 ; U6919
g4568 nand SUB_357_U9 U2355 ; U6920
g4569 nand U4195 U3218 ; U6921
g4570 nand SUB_357_U13 U2355 ; U6922
g4571 nand U4195 U3217 ; U6923
g4572 nand SUB_357_U11 U2355 ; U6924
g4573 nand R2182_U25 U3281 ; U6925
g4574 nand U4195 U3216 ; U6926
g4575 nand SUB_357_U12 U2355 ; U6927
g4576 nand R2182_U42 U3281 ; U6928
g4577 nand U2564 INSTQUEUE_REG_15__7__SCAN_IN ; U6929
g4578 nand U2563 INSTQUEUE_REG_14__7__SCAN_IN ; U6930
g4579 nand U2562 INSTQUEUE_REG_13__7__SCAN_IN ; U6931
g4580 nand U2561 INSTQUEUE_REG_12__7__SCAN_IN ; U6932
g4581 nand U2559 INSTQUEUE_REG_11__7__SCAN_IN ; U6933
g4582 nand U2558 INSTQUEUE_REG_10__7__SCAN_IN ; U6934
g4583 nand U2557 INSTQUEUE_REG_9__7__SCAN_IN ; U6935
g4584 nand U2556 INSTQUEUE_REG_8__7__SCAN_IN ; U6936
g4585 nand U2554 INSTQUEUE_REG_7__7__SCAN_IN ; U6937
g4586 nand U2553 INSTQUEUE_REG_6__7__SCAN_IN ; U6938
g4587 nand U2552 INSTQUEUE_REG_5__7__SCAN_IN ; U6939
g4588 nand U2551 INSTQUEUE_REG_4__7__SCAN_IN ; U6940
g4589 nand U2549 INSTQUEUE_REG_3__7__SCAN_IN ; U6941
g4590 nand U2548 INSTQUEUE_REG_2__7__SCAN_IN ; U6942
g4591 nand U2547 INSTQUEUE_REG_1__7__SCAN_IN ; U6943
g4592 nand U2546 INSTQUEUE_REG_0__7__SCAN_IN ; U6944
g4593 nand U4028 U4027 U4026 U4025 ; U6945
g4594 nand U2564 INSTQUEUE_REG_15__6__SCAN_IN ; U6946
g4595 nand U2563 INSTQUEUE_REG_14__6__SCAN_IN ; U6947
g4596 nand U2562 INSTQUEUE_REG_13__6__SCAN_IN ; U6948
g4597 nand U2561 INSTQUEUE_REG_12__6__SCAN_IN ; U6949
g4598 nand U2559 INSTQUEUE_REG_11__6__SCAN_IN ; U6950
g4599 nand U2558 INSTQUEUE_REG_10__6__SCAN_IN ; U6951
g4600 nand U2557 INSTQUEUE_REG_9__6__SCAN_IN ; U6952
g4601 nand U2556 INSTQUEUE_REG_8__6__SCAN_IN ; U6953
g4602 nand U2554 INSTQUEUE_REG_7__6__SCAN_IN ; U6954
g4603 nand U2553 INSTQUEUE_REG_6__6__SCAN_IN ; U6955
g4604 nand U2552 INSTQUEUE_REG_5__6__SCAN_IN ; U6956
g4605 nand U2551 INSTQUEUE_REG_4__6__SCAN_IN ; U6957
g4606 nand U2549 INSTQUEUE_REG_3__6__SCAN_IN ; U6958
g4607 nand U2548 INSTQUEUE_REG_2__6__SCAN_IN ; U6959
g4608 nand U2547 INSTQUEUE_REG_1__6__SCAN_IN ; U6960
g4609 nand U2546 INSTQUEUE_REG_0__6__SCAN_IN ; U6961
g4610 nand U4032 U4031 U4030 U4029 ; U6962
g4611 nand U2564 INSTQUEUE_REG_15__5__SCAN_IN ; U6963
g4612 nand U2563 INSTQUEUE_REG_14__5__SCAN_IN ; U6964
g4613 nand U2562 INSTQUEUE_REG_13__5__SCAN_IN ; U6965
g4614 nand U2561 INSTQUEUE_REG_12__5__SCAN_IN ; U6966
g4615 nand U2559 INSTQUEUE_REG_11__5__SCAN_IN ; U6967
g4616 nand U2558 INSTQUEUE_REG_10__5__SCAN_IN ; U6968
g4617 nand U2557 INSTQUEUE_REG_9__5__SCAN_IN ; U6969
g4618 nand U2556 INSTQUEUE_REG_8__5__SCAN_IN ; U6970
g4619 nand U2554 INSTQUEUE_REG_7__5__SCAN_IN ; U6971
g4620 nand U2553 INSTQUEUE_REG_6__5__SCAN_IN ; U6972
g4621 nand U2552 INSTQUEUE_REG_5__5__SCAN_IN ; U6973
g4622 nand U2551 INSTQUEUE_REG_4__5__SCAN_IN ; U6974
g4623 nand U2549 INSTQUEUE_REG_3__5__SCAN_IN ; U6975
g4624 nand U2548 INSTQUEUE_REG_2__5__SCAN_IN ; U6976
g4625 nand U2547 INSTQUEUE_REG_1__5__SCAN_IN ; U6977
g4626 nand U2546 INSTQUEUE_REG_0__5__SCAN_IN ; U6978
g4627 nand U4036 U4035 U4034 U4033 ; U6979
g4628 nand U2564 INSTQUEUE_REG_15__4__SCAN_IN ; U6980
g4629 nand U2563 INSTQUEUE_REG_14__4__SCAN_IN ; U6981
g4630 nand U2562 INSTQUEUE_REG_13__4__SCAN_IN ; U6982
g4631 nand U2561 INSTQUEUE_REG_12__4__SCAN_IN ; U6983
g4632 nand U2559 INSTQUEUE_REG_11__4__SCAN_IN ; U6984
g4633 nand U2558 INSTQUEUE_REG_10__4__SCAN_IN ; U6985
g4634 nand U2557 INSTQUEUE_REG_9__4__SCAN_IN ; U6986
g4635 nand U2556 INSTQUEUE_REG_8__4__SCAN_IN ; U6987
g4636 nand U2554 INSTQUEUE_REG_7__4__SCAN_IN ; U6988
g4637 nand U2553 INSTQUEUE_REG_6__4__SCAN_IN ; U6989
g4638 nand U2552 INSTQUEUE_REG_5__4__SCAN_IN ; U6990
g4639 nand U2551 INSTQUEUE_REG_4__4__SCAN_IN ; U6991
g4640 nand U2549 INSTQUEUE_REG_3__4__SCAN_IN ; U6992
g4641 nand U2548 INSTQUEUE_REG_2__4__SCAN_IN ; U6993
g4642 nand U2547 INSTQUEUE_REG_1__4__SCAN_IN ; U6994
g4643 nand U2564 INSTQUEUE_REG_15__3__SCAN_IN ; U6995
g4644 nand U2563 INSTQUEUE_REG_14__3__SCAN_IN ; U6996
g4645 nand U2562 INSTQUEUE_REG_13__3__SCAN_IN ; U6997
g4646 nand U2561 INSTQUEUE_REG_12__3__SCAN_IN ; U6998
g4647 nand U2559 INSTQUEUE_REG_11__3__SCAN_IN ; U6999
g4648 nand U2558 INSTQUEUE_REG_10__3__SCAN_IN ; U7000
g4649 nand U2557 INSTQUEUE_REG_9__3__SCAN_IN ; U7001
g4650 nand U2556 INSTQUEUE_REG_8__3__SCAN_IN ; U7002
g4651 nand U2554 INSTQUEUE_REG_7__3__SCAN_IN ; U7003
g4652 nand U2553 INSTQUEUE_REG_6__3__SCAN_IN ; U7004
g4653 nand U2552 INSTQUEUE_REG_5__3__SCAN_IN ; U7005
g4654 nand U2551 INSTQUEUE_REG_4__3__SCAN_IN ; U7006
g4655 nand U2549 INSTQUEUE_REG_3__3__SCAN_IN ; U7007
g4656 nand U2548 INSTQUEUE_REG_2__3__SCAN_IN ; U7008
g4657 nand U2547 INSTQUEUE_REG_1__3__SCAN_IN ; U7009
g4658 nand U2546 INSTQUEUE_REG_0__3__SCAN_IN ; U7010
g4659 nand U4044 U4043 U4042 U4041 ; U7011
g4660 nand U2564 INSTQUEUE_REG_15__2__SCAN_IN ; U7012
g4661 nand U2563 INSTQUEUE_REG_14__2__SCAN_IN ; U7013
g4662 nand U2562 INSTQUEUE_REG_13__2__SCAN_IN ; U7014
g4663 nand U2561 INSTQUEUE_REG_12__2__SCAN_IN ; U7015
g4664 nand U2559 INSTQUEUE_REG_11__2__SCAN_IN ; U7016
g4665 nand U2558 INSTQUEUE_REG_10__2__SCAN_IN ; U7017
g4666 nand U2557 INSTQUEUE_REG_9__2__SCAN_IN ; U7018
g4667 nand U2556 INSTQUEUE_REG_8__2__SCAN_IN ; U7019
g4668 nand U2554 INSTQUEUE_REG_7__2__SCAN_IN ; U7020
g4669 nand U2553 INSTQUEUE_REG_6__2__SCAN_IN ; U7021
g4670 nand U2552 INSTQUEUE_REG_5__2__SCAN_IN ; U7022
g4671 nand U2551 INSTQUEUE_REG_4__2__SCAN_IN ; U7023
g4672 nand U2549 INSTQUEUE_REG_3__2__SCAN_IN ; U7024
g4673 nand U2548 INSTQUEUE_REG_2__2__SCAN_IN ; U7025
g4674 nand U2547 INSTQUEUE_REG_1__2__SCAN_IN ; U7026
g4675 nand U2546 INSTQUEUE_REG_0__2__SCAN_IN ; U7027
g4676 nand U4048 U4047 U4046 U4045 ; U7028
g4677 nand U4195 U3215 ; U7029
g4678 nand SUB_357_U7 U2355 ; U7030
g4679 nand R2182_U33 U3281 ; U7031
g4680 nand U4195 U3214 ; U7032
g4681 nand SUB_357_U10 U2355 ; U7033
g4682 nand R2182_U34 U3281 ; U7034
g4683 nand U4194 U3221 ; U7035
g4684 nand U4180 INSTQUEUE_REG_0__7__SCAN_IN ; U7036
g4685 nand U4194 U3220 ; U7037
g4686 nand U4180 INSTQUEUE_REG_0__6__SCAN_IN ; U7038
g4687 nand U4194 U3219 ; U7039
g4688 nand U4180 INSTQUEUE_REG_0__5__SCAN_IN ; U7040
g4689 nand U4194 U3218 ; U7041
g4690 nand U4194 U3217 ; U7042
g4691 nand U4180 INSTQUEUE_REG_0__3__SCAN_IN ; U7043
g4692 nand U4194 U3216 ; U7044
g4693 nand U4180 INSTQUEUE_REG_0__2__SCAN_IN ; U7045
g4694 nand U4194 U3215 ; U7046
g4695 nand U4180 INSTQUEUE_REG_0__1__SCAN_IN ; U7047
g4696 nand U4194 U3214 ; U7048
g4697 nand U3221 U4388 ; U7049
g4698 nand U4180 INSTQUEUE_REG_0__0__SCAN_IN ; U7050
g4699 nand U3415 U3414 ; U7051
g4700 nand U3251 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7052
g4701 not U3432 ; U7053
g4702 nand U2582 INSTQUEUE_REG_8__7__SCAN_IN ; U7054
g4703 nand U2581 INSTQUEUE_REG_9__7__SCAN_IN ; U7055
g4704 nand U2580 INSTQUEUE_REG_10__7__SCAN_IN ; U7056
g4705 nand U2579 INSTQUEUE_REG_11__7__SCAN_IN ; U7057
g4706 nand U2577 INSTQUEUE_REG_12__7__SCAN_IN ; U7058
g4707 nand U2576 INSTQUEUE_REG_13__7__SCAN_IN ; U7059
g4708 nand U2575 INSTQUEUE_REG_14__7__SCAN_IN ; U7060
g4709 nand U2574 INSTQUEUE_REG_15__7__SCAN_IN ; U7061
g4710 nand U2573 INSTQUEUE_REG_0__7__SCAN_IN ; U7062
g4711 nand U2572 INSTQUEUE_REG_1__7__SCAN_IN ; U7063
g4712 nand U2571 INSTQUEUE_REG_2__7__SCAN_IN ; U7064
g4713 nand U2570 INSTQUEUE_REG_3__7__SCAN_IN ; U7065
g4714 nand U2568 INSTQUEUE_REG_4__7__SCAN_IN ; U7066
g4715 nand U2567 INSTQUEUE_REG_5__7__SCAN_IN ; U7067
g4716 nand U2566 INSTQUEUE_REG_6__7__SCAN_IN ; U7068
g4717 nand U2565 INSTQUEUE_REG_7__7__SCAN_IN ; U7069
g4718 nand U4054 U4053 U4052 U4051 ; U7070
g4719 nand U3412 U3408 ; U7071
g4720 nand U4061 U4179 ; U7072
g4721 nand U7072 U3409 ; U7073
g4722 nand U4491 U3265 ; U7074
g4723 not U3232 ; U7075
g4724 nand U4388 U4491 U4142 U3381 ; U7076
g4725 nand U4177 STATE2_REG_0__SCAN_IN ; U7077
g4726 nand U4055 U3232 ; U7078
g4727 not U3438 ; U7079
g4728 nand U3438 U5480 U7617 ; U7080
g4729 nand U4182 U7080 ; U7081
g4730 not U3437 ; U7082
g4731 nand U3284 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; U7083
g4732 nand U3437 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7084
g4733 nand U4191 U3347 ; U7085
g4734 nand U2582 INSTQUEUE_REG_8__6__SCAN_IN ; U7086
g4735 nand U2581 INSTQUEUE_REG_9__6__SCAN_IN ; U7087
g4736 nand U2580 INSTQUEUE_REG_10__6__SCAN_IN ; U7088
g4737 nand U2579 INSTQUEUE_REG_11__6__SCAN_IN ; U7089
g4738 nand U2577 INSTQUEUE_REG_12__6__SCAN_IN ; U7090
g4739 nand U2576 INSTQUEUE_REG_13__6__SCAN_IN ; U7091
g4740 nand U2575 INSTQUEUE_REG_14__6__SCAN_IN ; U7092
g4741 nand U2574 INSTQUEUE_REG_15__6__SCAN_IN ; U7093
g4742 nand U2573 INSTQUEUE_REG_0__6__SCAN_IN ; U7094
g4743 nand U2572 INSTQUEUE_REG_1__6__SCAN_IN ; U7095
g4744 nand U2571 INSTQUEUE_REG_2__6__SCAN_IN ; U7096
g4745 nand U2570 INSTQUEUE_REG_3__6__SCAN_IN ; U7097
g4746 nand U2568 INSTQUEUE_REG_4__6__SCAN_IN ; U7098
g4747 nand U2567 INSTQUEUE_REG_5__6__SCAN_IN ; U7099
g4748 nand U2566 INSTQUEUE_REG_6__6__SCAN_IN ; U7100
g4749 nand U2565 INSTQUEUE_REG_7__6__SCAN_IN ; U7101
g4750 nand U4070 U4069 U4068 U4067 ; U7102
g4751 nand U2582 INSTQUEUE_REG_8__5__SCAN_IN ; U7103
g4752 nand U2581 INSTQUEUE_REG_9__5__SCAN_IN ; U7104
g4753 nand U2580 INSTQUEUE_REG_10__5__SCAN_IN ; U7105
g4754 nand U2579 INSTQUEUE_REG_11__5__SCAN_IN ; U7106
g4755 nand U2577 INSTQUEUE_REG_12__5__SCAN_IN ; U7107
g4756 nand U2576 INSTQUEUE_REG_13__5__SCAN_IN ; U7108
g4757 nand U2575 INSTQUEUE_REG_14__5__SCAN_IN ; U7109
g4758 nand U2574 INSTQUEUE_REG_15__5__SCAN_IN ; U7110
g4759 nand U2573 INSTQUEUE_REG_0__5__SCAN_IN ; U7111
g4760 nand U2572 INSTQUEUE_REG_1__5__SCAN_IN ; U7112
g4761 nand U2571 INSTQUEUE_REG_2__5__SCAN_IN ; U7113
g4762 nand U2570 INSTQUEUE_REG_3__5__SCAN_IN ; U7114
g4763 nand U2568 INSTQUEUE_REG_4__5__SCAN_IN ; U7115
g4764 nand U2567 INSTQUEUE_REG_5__5__SCAN_IN ; U7116
g4765 nand U2566 INSTQUEUE_REG_6__5__SCAN_IN ; U7117
g4766 nand U2565 INSTQUEUE_REG_7__5__SCAN_IN ; U7118
g4767 nand U4074 U4073 U4072 U4071 ; U7119
g4768 nand U2582 INSTQUEUE_REG_8__4__SCAN_IN ; U7120
g4769 nand U2581 INSTQUEUE_REG_9__4__SCAN_IN ; U7121
g4770 nand U2580 INSTQUEUE_REG_10__4__SCAN_IN ; U7122
g4771 nand U2579 INSTQUEUE_REG_11__4__SCAN_IN ; U7123
g4772 nand U2577 INSTQUEUE_REG_12__4__SCAN_IN ; U7124
g4773 nand U2576 INSTQUEUE_REG_13__4__SCAN_IN ; U7125
g4774 nand U2575 INSTQUEUE_REG_14__4__SCAN_IN ; U7126
g4775 nand U2574 INSTQUEUE_REG_15__4__SCAN_IN ; U7127
g4776 nand U2572 INSTQUEUE_REG_1__4__SCAN_IN ; U7128
g4777 nand U2571 INSTQUEUE_REG_2__4__SCAN_IN ; U7129
g4778 nand U2570 INSTQUEUE_REG_3__4__SCAN_IN ; U7130
g4779 nand U2568 INSTQUEUE_REG_4__4__SCAN_IN ; U7131
g4780 nand U2567 INSTQUEUE_REG_5__4__SCAN_IN ; U7132
g4781 nand U2566 INSTQUEUE_REG_6__4__SCAN_IN ; U7133
g4782 nand U2565 INSTQUEUE_REG_7__4__SCAN_IN ; U7134
g4783 nand U2582 INSTQUEUE_REG_8__3__SCAN_IN ; U7135
g4784 nand U2581 INSTQUEUE_REG_9__3__SCAN_IN ; U7136
g4785 nand U2580 INSTQUEUE_REG_10__3__SCAN_IN ; U7137
g4786 nand U2579 INSTQUEUE_REG_11__3__SCAN_IN ; U7138
g4787 nand U2577 INSTQUEUE_REG_12__3__SCAN_IN ; U7139
g4788 nand U2576 INSTQUEUE_REG_13__3__SCAN_IN ; U7140
g4789 nand U2575 INSTQUEUE_REG_14__3__SCAN_IN ; U7141
g4790 nand U2574 INSTQUEUE_REG_15__3__SCAN_IN ; U7142
g4791 nand U2573 INSTQUEUE_REG_0__3__SCAN_IN ; U7143
g4792 nand U2572 INSTQUEUE_REG_1__3__SCAN_IN ; U7144
g4793 nand U2571 INSTQUEUE_REG_2__3__SCAN_IN ; U7145
g4794 nand U2570 INSTQUEUE_REG_3__3__SCAN_IN ; U7146
g4795 nand U2568 INSTQUEUE_REG_4__3__SCAN_IN ; U7147
g4796 nand U2567 INSTQUEUE_REG_5__3__SCAN_IN ; U7148
g4797 nand U2566 INSTQUEUE_REG_6__3__SCAN_IN ; U7149
g4798 nand U2565 INSTQUEUE_REG_7__3__SCAN_IN ; U7150
g4799 nand U4083 U4082 U4081 U4080 ; U7151
g4800 nand U2582 INSTQUEUE_REG_8__2__SCAN_IN ; U7152
g4801 nand U2581 INSTQUEUE_REG_9__2__SCAN_IN ; U7153
g4802 nand U2580 INSTQUEUE_REG_10__2__SCAN_IN ; U7154
g4803 nand U2579 INSTQUEUE_REG_11__2__SCAN_IN ; U7155
g4804 nand U2577 INSTQUEUE_REG_12__2__SCAN_IN ; U7156
g4805 nand U2576 INSTQUEUE_REG_13__2__SCAN_IN ; U7157
g4806 nand U2575 INSTQUEUE_REG_14__2__SCAN_IN ; U7158
g4807 nand U2574 INSTQUEUE_REG_15__2__SCAN_IN ; U7159
g4808 nand U2573 INSTQUEUE_REG_0__2__SCAN_IN ; U7160
g4809 nand U2572 INSTQUEUE_REG_1__2__SCAN_IN ; U7161
g4810 nand U2571 INSTQUEUE_REG_2__2__SCAN_IN ; U7162
g4811 nand U2570 INSTQUEUE_REG_3__2__SCAN_IN ; U7163
g4812 nand U2568 INSTQUEUE_REG_4__2__SCAN_IN ; U7164
g4813 nand U2567 INSTQUEUE_REG_5__2__SCAN_IN ; U7165
g4814 nand U2566 INSTQUEUE_REG_6__2__SCAN_IN ; U7166
g4815 nand U2565 INSTQUEUE_REG_7__2__SCAN_IN ; U7167
g4816 nand U4087 U4086 U4085 U4084 ; U7168
g4817 nand U2582 INSTQUEUE_REG_8__1__SCAN_IN ; U7169
g4818 nand U2581 INSTQUEUE_REG_9__1__SCAN_IN ; U7170
g4819 nand U2580 INSTQUEUE_REG_10__1__SCAN_IN ; U7171
g4820 nand U2579 INSTQUEUE_REG_11__1__SCAN_IN ; U7172
g4821 nand U2577 INSTQUEUE_REG_12__1__SCAN_IN ; U7173
g4822 nand U2576 INSTQUEUE_REG_13__1__SCAN_IN ; U7174
g4823 nand U2575 INSTQUEUE_REG_14__1__SCAN_IN ; U7175
g4824 nand U2574 INSTQUEUE_REG_15__1__SCAN_IN ; U7176
g4825 nand U2573 INSTQUEUE_REG_0__1__SCAN_IN ; U7177
g4826 nand U2572 INSTQUEUE_REG_1__1__SCAN_IN ; U7178
g4827 nand U2571 INSTQUEUE_REG_2__1__SCAN_IN ; U7179
g4828 nand U2570 INSTQUEUE_REG_3__1__SCAN_IN ; U7180
g4829 nand U2568 INSTQUEUE_REG_4__1__SCAN_IN ; U7181
g4830 nand U2567 INSTQUEUE_REG_5__1__SCAN_IN ; U7182
g4831 nand U2566 INSTQUEUE_REG_6__1__SCAN_IN ; U7183
g4832 nand U2565 INSTQUEUE_REG_7__1__SCAN_IN ; U7184
g4833 nand U4091 U4090 U4089 U4088 ; U7185
g4834 nand U2582 INSTQUEUE_REG_8__0__SCAN_IN ; U7186
g4835 nand U2581 INSTQUEUE_REG_9__0__SCAN_IN ; U7187
g4836 nand U2580 INSTQUEUE_REG_10__0__SCAN_IN ; U7188
g4837 nand U2579 INSTQUEUE_REG_11__0__SCAN_IN ; U7189
g4838 nand U2577 INSTQUEUE_REG_12__0__SCAN_IN ; U7190
g4839 nand U2576 INSTQUEUE_REG_13__0__SCAN_IN ; U7191
g4840 nand U2575 INSTQUEUE_REG_14__0__SCAN_IN ; U7192
g4841 nand U2574 INSTQUEUE_REG_15__0__SCAN_IN ; U7193
g4842 nand U2573 INSTQUEUE_REG_0__0__SCAN_IN ; U7194
g4843 nand U2572 INSTQUEUE_REG_1__0__SCAN_IN ; U7195
g4844 nand U2571 INSTQUEUE_REG_2__0__SCAN_IN ; U7196
g4845 nand U2570 INSTQUEUE_REG_3__0__SCAN_IN ; U7197
g4846 nand U2568 INSTQUEUE_REG_4__0__SCAN_IN ; U7198
g4847 nand U2567 INSTQUEUE_REG_5__0__SCAN_IN ; U7199
g4848 nand U2566 INSTQUEUE_REG_6__0__SCAN_IN ; U7200
g4849 nand U2565 INSTQUEUE_REG_7__0__SCAN_IN ; U7201
g4850 nand U4095 U4094 U4093 U4092 ; U7202
g4851 nand U3284 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U7203
g4852 nand U4191 U3442 ; U7204
g4853 nand U3284 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; U7205
g4854 nand U4191 U3222 ; U7206
g4855 not U4171 ; U7207
g4856 nand U2602 INSTQUEUE_REG_8__7__SCAN_IN ; U7208
g4857 nand U2601 INSTQUEUE_REG_9__7__SCAN_IN ; U7209
g4858 nand U2600 INSTQUEUE_REG_10__7__SCAN_IN ; U7210
g4859 nand U2599 INSTQUEUE_REG_11__7__SCAN_IN ; U7211
g4860 nand U2597 INSTQUEUE_REG_12__7__SCAN_IN ; U7212
g4861 nand U2596 INSTQUEUE_REG_13__7__SCAN_IN ; U7213
g4862 nand U2595 INSTQUEUE_REG_14__7__SCAN_IN ; U7214
g4863 nand U2594 INSTQUEUE_REG_15__7__SCAN_IN ; U7215
g4864 nand U2592 INSTQUEUE_REG_0__7__SCAN_IN ; U7216
g4865 nand U2591 INSTQUEUE_REG_1__7__SCAN_IN ; U7217
g4866 nand U2590 INSTQUEUE_REG_2__7__SCAN_IN ; U7218
g4867 nand U2589 INSTQUEUE_REG_3__7__SCAN_IN ; U7219
g4868 nand U2587 INSTQUEUE_REG_4__7__SCAN_IN ; U7220
g4869 nand U2586 INSTQUEUE_REG_5__7__SCAN_IN ; U7221
g4870 nand U2585 INSTQUEUE_REG_6__7__SCAN_IN ; U7222
g4871 nand U2584 INSTQUEUE_REG_7__7__SCAN_IN ; U7223
g4872 nand U4112 U4111 U4110 U4109 ; U7224
g4873 nand U2602 INSTQUEUE_REG_8__6__SCAN_IN ; U7225
g4874 nand U2601 INSTQUEUE_REG_9__6__SCAN_IN ; U7226
g4875 nand U2600 INSTQUEUE_REG_10__6__SCAN_IN ; U7227
g4876 nand U2599 INSTQUEUE_REG_11__6__SCAN_IN ; U7228
g4877 nand U2597 INSTQUEUE_REG_12__6__SCAN_IN ; U7229
g4878 nand U2596 INSTQUEUE_REG_13__6__SCAN_IN ; U7230
g4879 nand U2595 INSTQUEUE_REG_14__6__SCAN_IN ; U7231
g4880 nand U2594 INSTQUEUE_REG_15__6__SCAN_IN ; U7232
g4881 nand U2592 INSTQUEUE_REG_0__6__SCAN_IN ; U7233
g4882 nand U2591 INSTQUEUE_REG_1__6__SCAN_IN ; U7234
g4883 nand U2590 INSTQUEUE_REG_2__6__SCAN_IN ; U7235
g4884 nand U2589 INSTQUEUE_REG_3__6__SCAN_IN ; U7236
g4885 nand U2587 INSTQUEUE_REG_4__6__SCAN_IN ; U7237
g4886 nand U2586 INSTQUEUE_REG_5__6__SCAN_IN ; U7238
g4887 nand U2585 INSTQUEUE_REG_6__6__SCAN_IN ; U7239
g4888 nand U2584 INSTQUEUE_REG_7__6__SCAN_IN ; U7240
g4889 nand U4116 U4115 U4114 U4113 ; U7241
g4890 nand U2602 INSTQUEUE_REG_8__5__SCAN_IN ; U7242
g4891 nand U2601 INSTQUEUE_REG_9__5__SCAN_IN ; U7243
g4892 nand U2600 INSTQUEUE_REG_10__5__SCAN_IN ; U7244
g4893 nand U2599 INSTQUEUE_REG_11__5__SCAN_IN ; U7245
g4894 nand U2597 INSTQUEUE_REG_12__5__SCAN_IN ; U7246
g4895 nand U2596 INSTQUEUE_REG_13__5__SCAN_IN ; U7247
g4896 nand U2595 INSTQUEUE_REG_14__5__SCAN_IN ; U7248
g4897 nand U2594 INSTQUEUE_REG_15__5__SCAN_IN ; U7249
g4898 nand U2592 INSTQUEUE_REG_0__5__SCAN_IN ; U7250
g4899 nand U2591 INSTQUEUE_REG_1__5__SCAN_IN ; U7251
g4900 nand U2590 INSTQUEUE_REG_2__5__SCAN_IN ; U7252
g4901 nand U2589 INSTQUEUE_REG_3__5__SCAN_IN ; U7253
g4902 nand U2587 INSTQUEUE_REG_4__5__SCAN_IN ; U7254
g4903 nand U2586 INSTQUEUE_REG_5__5__SCAN_IN ; U7255
g4904 nand U2585 INSTQUEUE_REG_6__5__SCAN_IN ; U7256
g4905 nand U2584 INSTQUEUE_REG_7__5__SCAN_IN ; U7257
g4906 nand U4120 U4119 U4118 U4117 ; U7258
g4907 nand U2602 INSTQUEUE_REG_8__4__SCAN_IN ; U7259
g4908 nand U2601 INSTQUEUE_REG_9__4__SCAN_IN ; U7260
g4909 nand U2600 INSTQUEUE_REG_10__4__SCAN_IN ; U7261
g4910 nand U2599 INSTQUEUE_REG_11__4__SCAN_IN ; U7262
g4911 nand U2597 INSTQUEUE_REG_12__4__SCAN_IN ; U7263
g4912 nand U2596 INSTQUEUE_REG_13__4__SCAN_IN ; U7264
g4913 nand U2595 INSTQUEUE_REG_14__4__SCAN_IN ; U7265
g4914 nand U2594 INSTQUEUE_REG_15__4__SCAN_IN ; U7266
g4915 nand U2591 INSTQUEUE_REG_1__4__SCAN_IN ; U7267
g4916 nand U2590 INSTQUEUE_REG_2__4__SCAN_IN ; U7268
g4917 nand U2589 INSTQUEUE_REG_3__4__SCAN_IN ; U7269
g4918 nand U2587 INSTQUEUE_REG_4__4__SCAN_IN ; U7270
g4919 nand U2586 INSTQUEUE_REG_5__4__SCAN_IN ; U7271
g4920 nand U2585 INSTQUEUE_REG_6__4__SCAN_IN ; U7272
g4921 nand U2584 INSTQUEUE_REG_7__4__SCAN_IN ; U7273
g4922 nand U2602 INSTQUEUE_REG_8__3__SCAN_IN ; U7274
g4923 nand U2601 INSTQUEUE_REG_9__3__SCAN_IN ; U7275
g4924 nand U2600 INSTQUEUE_REG_10__3__SCAN_IN ; U7276
g4925 nand U2599 INSTQUEUE_REG_11__3__SCAN_IN ; U7277
g4926 nand U2597 INSTQUEUE_REG_12__3__SCAN_IN ; U7278
g4927 nand U2596 INSTQUEUE_REG_13__3__SCAN_IN ; U7279
g4928 nand U2595 INSTQUEUE_REG_14__3__SCAN_IN ; U7280
g4929 nand U2594 INSTQUEUE_REG_15__3__SCAN_IN ; U7281
g4930 nand U2592 INSTQUEUE_REG_0__3__SCAN_IN ; U7282
g4931 nand U2591 INSTQUEUE_REG_1__3__SCAN_IN ; U7283
g4932 nand U2590 INSTQUEUE_REG_2__3__SCAN_IN ; U7284
g4933 nand U2589 INSTQUEUE_REG_3__3__SCAN_IN ; U7285
g4934 nand U2587 INSTQUEUE_REG_4__3__SCAN_IN ; U7286
g4935 nand U2586 INSTQUEUE_REG_5__3__SCAN_IN ; U7287
g4936 nand U2585 INSTQUEUE_REG_6__3__SCAN_IN ; U7288
g4937 nand U2584 INSTQUEUE_REG_7__3__SCAN_IN ; U7289
g4938 nand U4128 U4127 U4126 U4125 ; U7290
g4939 nand U2602 INSTQUEUE_REG_8__2__SCAN_IN ; U7291
g4940 nand U2601 INSTQUEUE_REG_9__2__SCAN_IN ; U7292
g4941 nand U2600 INSTQUEUE_REG_10__2__SCAN_IN ; U7293
g4942 nand U2599 INSTQUEUE_REG_11__2__SCAN_IN ; U7294
g4943 nand U2597 INSTQUEUE_REG_12__2__SCAN_IN ; U7295
g4944 nand U2596 INSTQUEUE_REG_13__2__SCAN_IN ; U7296
g4945 nand U2595 INSTQUEUE_REG_14__2__SCAN_IN ; U7297
g4946 nand U2594 INSTQUEUE_REG_15__2__SCAN_IN ; U7298
g4947 nand U2592 INSTQUEUE_REG_0__2__SCAN_IN ; U7299
g4948 nand U2591 INSTQUEUE_REG_1__2__SCAN_IN ; U7300
g4949 nand U2590 INSTQUEUE_REG_2__2__SCAN_IN ; U7301
g4950 nand U2589 INSTQUEUE_REG_3__2__SCAN_IN ; U7302
g4951 nand U2587 INSTQUEUE_REG_4__2__SCAN_IN ; U7303
g4952 nand U2586 INSTQUEUE_REG_5__2__SCAN_IN ; U7304
g4953 nand U2585 INSTQUEUE_REG_6__2__SCAN_IN ; U7305
g4954 nand U2584 INSTQUEUE_REG_7__2__SCAN_IN ; U7306
g4955 nand U4132 U4131 U4130 U4129 ; U7307
g4956 nand U2602 INSTQUEUE_REG_8__1__SCAN_IN ; U7308
g4957 nand U2601 INSTQUEUE_REG_9__1__SCAN_IN ; U7309
g4958 nand U2600 INSTQUEUE_REG_10__1__SCAN_IN ; U7310
g4959 nand U2599 INSTQUEUE_REG_11__1__SCAN_IN ; U7311
g4960 nand U2597 INSTQUEUE_REG_12__1__SCAN_IN ; U7312
g4961 nand U2596 INSTQUEUE_REG_13__1__SCAN_IN ; U7313
g4962 nand U2595 INSTQUEUE_REG_14__1__SCAN_IN ; U7314
g4963 nand U2594 INSTQUEUE_REG_15__1__SCAN_IN ; U7315
g4964 nand U2592 INSTQUEUE_REG_0__1__SCAN_IN ; U7316
g4965 nand U2591 INSTQUEUE_REG_1__1__SCAN_IN ; U7317
g4966 nand U2590 INSTQUEUE_REG_2__1__SCAN_IN ; U7318
g4967 nand U2589 INSTQUEUE_REG_3__1__SCAN_IN ; U7319
g4968 nand U2587 INSTQUEUE_REG_4__1__SCAN_IN ; U7320
g4969 nand U2586 INSTQUEUE_REG_5__1__SCAN_IN ; U7321
g4970 nand U2585 INSTQUEUE_REG_6__1__SCAN_IN ; U7322
g4971 nand U2584 INSTQUEUE_REG_7__1__SCAN_IN ; U7323
g4972 nand U4136 U4135 U4134 U4133 ; U7324
g4973 nand U2602 INSTQUEUE_REG_8__0__SCAN_IN ; U7325
g4974 nand U2601 INSTQUEUE_REG_9__0__SCAN_IN ; U7326
g4975 nand U2600 INSTQUEUE_REG_10__0__SCAN_IN ; U7327
g4976 nand U2599 INSTQUEUE_REG_11__0__SCAN_IN ; U7328
g4977 nand U2597 INSTQUEUE_REG_12__0__SCAN_IN ; U7329
g4978 nand U2596 INSTQUEUE_REG_13__0__SCAN_IN ; U7330
g4979 nand U2595 INSTQUEUE_REG_14__0__SCAN_IN ; U7331
g4980 nand U2594 INSTQUEUE_REG_15__0__SCAN_IN ; U7332
g4981 nand U2592 INSTQUEUE_REG_0__0__SCAN_IN ; U7333
g4982 nand U2591 INSTQUEUE_REG_1__0__SCAN_IN ; U7334
g4983 nand U2590 INSTQUEUE_REG_2__0__SCAN_IN ; U7335
g4984 nand U2589 INSTQUEUE_REG_3__0__SCAN_IN ; U7336
g4985 nand U2587 INSTQUEUE_REG_4__0__SCAN_IN ; U7337
g4986 nand U2586 INSTQUEUE_REG_5__0__SCAN_IN ; U7338
g4987 nand U2585 INSTQUEUE_REG_6__0__SCAN_IN ; U7339
g4988 nand U2584 INSTQUEUE_REG_7__0__SCAN_IN ; U7340
g4989 nand U4140 U4139 U4138 U4137 ; U7341
g4990 nand U4219 U2354 U4222 ; U7342
g4991 nand U4141 U7075 ; U7343
g4992 nand U3383 U3397 ; U7344
g4993 nand U4222 U7344 ; U7345
g4994 nand U4178 U2452 ; U7346
g4995 nand U7343 U3258 ; U7347
g4996 nand U4196 U7076 ; U7348
g4997 nand U4148 U4196 ; U7349
g4998 nand U2451 U4198 ; U7350
g4999 nand U3407 U3421 U4183 U7350 U7349 ; U7351
g5000 nand R2238_U6 U7351 ; U7352
g5001 nand SUB_450_U6 U2354 ; U7353
g5002 nand R2238_U19 U7351 ; U7354
g5003 nand SUB_450_U19 U2354 ; U7355
g5004 nand R2238_U20 U7351 ; U7356
g5005 nand SUB_450_U20 U2354 ; U7357
g5006 nand R2238_U21 U7351 ; U7358
g5007 nand SUB_450_U21 U2354 ; U7359
g5008 nand R2238_U22 U7351 ; U7360
g5009 nand SUB_450_U22 U2354 ; U7361
g5010 nand R2238_U7 U7351 ; U7362
g5011 nand SUB_450_U7 U2354 ; U7363
g5012 nand R2238_U19 U4180 ; U7364
g5013 nand U3281 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; U7365
g5014 nand R2238_U20 U4180 ; U7366
g5015 nand U3281 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7367
g5016 nand U4161 STATE2_REG_0__SCAN_IN ; U7368
g5017 nand U3407 U7368 ; U7369
g5018 nand R2238_U21 U4180 ; U7370
g5019 nand U3281 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U7371
g5020 nand U2450 U3258 ; U7372
g5021 nand R2238_U22 U4180 ; U7373
g5022 nand U3281 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7374
g5023 nand U2451 U3271 ; U7375
g5024 nand R2238_U7 U4180 ; U7376
g5025 nand U3281 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7377
g5026 nand U3380 U3277 ; U7378
g5027 nand U3271 U3436 ; U7379
g5028 nand U7379 INSTADDRPOINTER_REG_9__SCAN_IN ; U7380
g5029 nand U7378 EBX_REG_9__SCAN_IN ; U7381
g5030 nand U7379 INSTADDRPOINTER_REG_8__SCAN_IN ; U7382
g5031 nand U7378 EBX_REG_8__SCAN_IN ; U7383
g5032 nand U7379 INSTADDRPOINTER_REG_7__SCAN_IN ; U7384
g5033 nand U7378 EBX_REG_7__SCAN_IN ; U7385
g5034 nand U7379 INSTADDRPOINTER_REG_6__SCAN_IN ; U7386
g5035 nand U7378 EBX_REG_6__SCAN_IN ; U7387
g5036 nand U7379 INSTADDRPOINTER_REG_5__SCAN_IN ; U7388
g5037 nand U7378 EBX_REG_5__SCAN_IN ; U7389
g5038 nand U7379 INSTADDRPOINTER_REG_4__SCAN_IN ; U7390
g5039 nand U7378 EBX_REG_4__SCAN_IN ; U7391
g5040 nand U7379 INSTADDRPOINTER_REG_31__SCAN_IN ; U7392
g5041 nand U7378 EBX_REG_31__SCAN_IN ; U7393
g5042 nand U7379 INSTADDRPOINTER_REG_30__SCAN_IN ; U7394
g5043 nand U7378 EBX_REG_30__SCAN_IN ; U7395
g5044 nand U7379 INSTADDRPOINTER_REG_3__SCAN_IN ; U7396
g5045 nand U7378 EBX_REG_3__SCAN_IN ; U7397
g5046 nand U7379 INSTADDRPOINTER_REG_29__SCAN_IN ; U7398
g5047 nand U7378 EBX_REG_29__SCAN_IN ; U7399
g5048 nand U7379 INSTADDRPOINTER_REG_28__SCAN_IN ; U7400
g5049 nand U7378 EBX_REG_28__SCAN_IN ; U7401
g5050 nand U7379 INSTADDRPOINTER_REG_27__SCAN_IN ; U7402
g5051 nand U7378 EBX_REG_27__SCAN_IN ; U7403
g5052 nand U7379 INSTADDRPOINTER_REG_26__SCAN_IN ; U7404
g5053 nand U7378 EBX_REG_26__SCAN_IN ; U7405
g5054 nand U7379 INSTADDRPOINTER_REG_25__SCAN_IN ; U7406
g5055 nand U7378 EBX_REG_25__SCAN_IN ; U7407
g5056 nand U7379 INSTADDRPOINTER_REG_24__SCAN_IN ; U7408
g5057 nand U7378 EBX_REG_24__SCAN_IN ; U7409
g5058 nand U7379 INSTADDRPOINTER_REG_23__SCAN_IN ; U7410
g5059 nand U7378 EBX_REG_23__SCAN_IN ; U7411
g5060 nand U7379 INSTADDRPOINTER_REG_22__SCAN_IN ; U7412
g5061 nand U7378 EBX_REG_22__SCAN_IN ; U7413
g5062 nand U7379 INSTADDRPOINTER_REG_21__SCAN_IN ; U7414
g5063 nand U7378 EBX_REG_21__SCAN_IN ; U7415
g5064 nand U7379 INSTADDRPOINTER_REG_20__SCAN_IN ; U7416
g5065 nand U7378 EBX_REG_20__SCAN_IN ; U7417
g5066 nand U7379 INSTADDRPOINTER_REG_2__SCAN_IN ; U7418
g5067 nand U7378 EBX_REG_2__SCAN_IN ; U7419
g5068 nand U7379 INSTADDRPOINTER_REG_19__SCAN_IN ; U7420
g5069 nand U7378 EBX_REG_19__SCAN_IN ; U7421
g5070 nand U7379 INSTADDRPOINTER_REG_18__SCAN_IN ; U7422
g5071 nand U7378 EBX_REG_18__SCAN_IN ; U7423
g5072 nand U7379 INSTADDRPOINTER_REG_17__SCAN_IN ; U7424
g5073 nand U7378 EBX_REG_17__SCAN_IN ; U7425
g5074 nand U7379 INSTADDRPOINTER_REG_16__SCAN_IN ; U7426
g5075 nand U7378 EBX_REG_16__SCAN_IN ; U7427
g5076 nand U7379 INSTADDRPOINTER_REG_15__SCAN_IN ; U7428
g5077 nand U7378 EBX_REG_15__SCAN_IN ; U7429
g5078 nand U7379 INSTADDRPOINTER_REG_14__SCAN_IN ; U7430
g5079 nand U7378 EBX_REG_14__SCAN_IN ; U7431
g5080 nand U7379 INSTADDRPOINTER_REG_13__SCAN_IN ; U7432
g5081 nand U7378 EBX_REG_13__SCAN_IN ; U7433
g5082 nand U7379 INSTADDRPOINTER_REG_12__SCAN_IN ; U7434
g5083 nand U7378 EBX_REG_12__SCAN_IN ; U7435
g5084 nand U7379 INSTADDRPOINTER_REG_11__SCAN_IN ; U7436
g5085 nand U7378 EBX_REG_11__SCAN_IN ; U7437
g5086 nand U7379 INSTADDRPOINTER_REG_10__SCAN_IN ; U7438
g5087 nand U7378 EBX_REG_10__SCAN_IN ; U7439
g5088 nand U7379 INSTADDRPOINTER_REG_1__SCAN_IN ; U7440
g5089 nand U7378 EBX_REG_1__SCAN_IN ; U7441
g5090 nand U7379 INSTADDRPOINTER_REG_0__SCAN_IN ; U7442
g5091 nand U7378 EBX_REG_0__SCAN_IN ; U7443
g5092 nand U4465 U4484 ; U7444
g5093 nand U2430 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; U7445
g5094 nand U3476 U3249 ; U7446
g5095 nand U2430 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7447
g5096 nand U3477 U3249 ; U7448
g5097 nand U2446 U3457 FLUSH_REG_SCAN_IN ; U7449
g5098 nand U2430 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U7450
g5099 nand U3478 U3249 ; U7451
g5100 nand U2446 U7700 FLUSH_REG_SCAN_IN ; U7452
g5101 nand U2430 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7453
g5102 nand U3479 U3249 ; U7454
g5103 nand U2430 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7455
g5104 nand U4173 STATE_REG_0__SCAN_IN ; U7456
g5105 or READY_N STATE2_REG_2__SCAN_IN ; U7457
g5106 nand U4098 U7206 ; U7458
g5107 nand U7072 U3409 ; U7459
g5108 nand U4199 STATE2_REG_0__SCAN_IN ; U7460
g5109 nand U4200 STATE2_REG_0__SCAN_IN ; U7461
g5110 nand U4201 STATE2_REG_0__SCAN_IN ; U7462
g5111 nand U4224 STATE2_REG_0__SCAN_IN ; U7463
g5112 nand U4252 STATE2_REG_0__SCAN_IN ; U7464
g5113 nand U7620 STATE2_REG_0__SCAN_IN ; U7465
g5114 nand U2608 U3253 ; U7466
g5115 nand U4105 U7081 U4106 U4108 ; U7467
g5116 nand U7620 STATE2_REG_0__SCAN_IN ; U7468
g5117 nand U2379 U3416 ; U7469
g5118 nand U2369 U6355 ; U7470
g5119 nand U3876 U2369 ; U7471
g5120 nand U7469 U4217 U7470 ; U7472
g5121 nand U7471 U4218 ; U7473
g5122 nand U5479 U4159 U4182 ; U7474
g5123 nand U7079 U4182 ; U7475
g5124 nand U4182 U3379 ; U7476
g5125 nand U4224 STATE2_REG_0__SCAN_IN ; U7477
g5126 nand U7773 U7772 U4060 ; U7478
g5127 nand U4096 U7204 ; U7479
g5128 nand U4097 U7082 ; U7480
g5129 not U3266 ; U7481
g5130 not U3263 ; U7482
g5131 nand U4059 U2607 U4058 U4057 U4056 ; U7483
g5132 nand U3722 U7481 ; U7484
g5133 nand U3723 U5457 ; U7485
g5134 nand U2425 U7481 ; U7486
g5135 nand U2425 U7481 ; U7487
g5136 nand U6349 U6348 U7487 ; U7488
g5137 nand U7481 R2167_U17 ; U7489
g5138 nand U7481 U4189 R2167_U17 ; U7490
g5139 nand U7490 U6137 ; U7491
g5140 nand U7481 U7073 ; U7492
g5141 nand U7481 U7459 ; U7493
g5142 nand U4104 U4103 U4102 ; U7494
g5143 nand U3747 U7481 ; U7495
g5144 nand U3749 U5553 U3748 ; U7496
g5145 nand U3734 U2519 ; U7497
g5146 nand U7481 U5950 ; U7498
g5147 nand U7481 U5953 ; U7499
g5148 nand U7481 U5956 ; U7500
g5149 nand U7481 U5959 ; U7501
g5150 nand U7481 U5962 ; U7502
g5151 nand U7481 U5965 ; U7503
g5152 nand U7481 U5968 ; U7504
g5153 nand U7481 U5971 ; U7505
g5154 nand U7481 U5974 ; U7506
g5155 nand U7481 U5977 ; U7507
g5156 nand U7481 U5980 ; U7508
g5157 nand U7481 U5983 ; U7509
g5158 nand U7481 U5986 ; U7510
g5159 nand U7481 U5989 ; U7511
g5160 nand U7481 U5992 ; U7512
g5161 nand U7481 U5995 ; U7513
g5162 nand U7481 U5998 ; U7514
g5163 nand U7481 U6001 ; U7515
g5164 nand U7481 U6004 ; U7516
g5165 nand U7481 U6007 ; U7517
g5166 nand U7481 U6010 ; U7518
g5167 nand U7481 U6013 ; U7519
g5168 nand U7481 U6016 ; U7520
g5169 nand U7481 U6019 ; U7521
g5170 nand U7481 U6022 ; U7522
g5171 nand U7481 U6025 ; U7523
g5172 nand U7481 U6028 ; U7524
g5173 nand U7481 U6031 ; U7525
g5174 nand U7481 U6034 ; U7526
g5175 nand U7481 U6037 ; U7527
g5176 nand U7481 U6040 ; U7528
g5177 nand U2357 U7481 ; U7529
g5178 nand U7529 UWORD_REG_0__SCAN_IN ; U7530
g5179 nand U2357 U7481 ; U7531
g5180 nand U7531 UWORD_REG_1__SCAN_IN ; U7532
g5181 nand U2357 U7481 ; U7533
g5182 nand U7533 UWORD_REG_2__SCAN_IN ; U7534
g5183 nand U2357 U7481 ; U7535
g5184 nand U7535 UWORD_REG_3__SCAN_IN ; U7536
g5185 nand U2357 U7481 ; U7537
g5186 nand U7537 UWORD_REG_4__SCAN_IN ; U7538
g5187 nand U2357 U7481 ; U7539
g5188 nand U7539 UWORD_REG_5__SCAN_IN ; U7540
g5189 nand U2357 U7481 ; U7541
g5190 nand U7541 UWORD_REG_6__SCAN_IN ; U7542
g5191 nand U2357 U7481 ; U7543
g5192 nand U7543 UWORD_REG_7__SCAN_IN ; U7544
g5193 nand U2357 U7481 ; U7545
g5194 nand U7545 UWORD_REG_8__SCAN_IN ; U7546
g5195 nand U2357 U7481 ; U7547
g5196 nand U7547 UWORD_REG_9__SCAN_IN ; U7548
g5197 nand U2357 U7481 ; U7549
g5198 nand U7549 UWORD_REG_10__SCAN_IN ; U7550
g5199 nand U2357 U7481 ; U7551
g5200 nand U7551 UWORD_REG_11__SCAN_IN ; U7552
g5201 nand U2357 U7481 ; U7553
g5202 nand U7553 UWORD_REG_12__SCAN_IN ; U7554
g5203 nand U2357 U7481 ; U7555
g5204 nand U7555 UWORD_REG_13__SCAN_IN ; U7556
g5205 nand U2357 U7481 ; U7557
g5206 nand U7557 UWORD_REG_14__SCAN_IN ; U7558
g5207 nand U2357 U7481 ; U7559
g5208 nand U7559 LWORD_REG_0__SCAN_IN ; U7560
g5209 nand U2357 U7481 ; U7561
g5210 nand U7561 LWORD_REG_1__SCAN_IN ; U7562
g5211 nand U2357 U7481 ; U7563
g5212 nand U7563 LWORD_REG_2__SCAN_IN ; U7564
g5213 nand U2357 U7481 ; U7565
g5214 nand U7565 LWORD_REG_3__SCAN_IN ; U7566
g5215 nand U2357 U7481 ; U7567
g5216 nand U7567 LWORD_REG_4__SCAN_IN ; U7568
g5217 nand U2357 U7481 ; U7569
g5218 nand U7569 LWORD_REG_5__SCAN_IN ; U7570
g5219 nand U2357 U7481 ; U7571
g5220 nand U7571 LWORD_REG_6__SCAN_IN ; U7572
g5221 nand U2357 U7481 ; U7573
g5222 nand U7573 LWORD_REG_7__SCAN_IN ; U7574
g5223 nand U2357 U7481 ; U7575
g5224 nand U7575 LWORD_REG_8__SCAN_IN ; U7576
g5225 nand U2357 U7481 ; U7577
g5226 nand U7577 LWORD_REG_9__SCAN_IN ; U7578
g5227 nand U2357 U7481 ; U7579
g5228 nand U7579 LWORD_REG_10__SCAN_IN ; U7580
g5229 nand U2357 U7481 ; U7581
g5230 nand U7581 LWORD_REG_11__SCAN_IN ; U7582
g5231 nand U2357 U7481 ; U7583
g5232 nand U7583 LWORD_REG_12__SCAN_IN ; U7584
g5233 nand U2357 U7481 ; U7585
g5234 nand U7585 LWORD_REG_13__SCAN_IN ; U7586
g5235 nand U2357 U7481 ; U7587
g5236 nand U7587 LWORD_REG_14__SCAN_IN ; U7588
g5237 nand U2357 U7481 ; U7589
g5238 nand U7589 LWORD_REG_15__SCAN_IN ; U7590
g5239 nand U7481 U3556 U4247 ; U7591
g5240 nand U7672 U7671 U3569 ; U7592
g5241 nand U3855 U7481 ; U7593
g5242 nand U7593 U3415 ; U7594
g5243 nand U4196 U7481 ; U7595
g5244 nand U7595 U3434 ; U7596
g5245 nand U3266 U3387 ; U7597
g5246 nand U3742 U7481 ; U7598
g5247 nand U3743 U7598 ; U7599
g5248 nand U5404 INSTQUEUE_REG_0__4__SCAN_IN ; U7600
g5249 nand U2523 INSTQUEUE_REG_0__4__SCAN_IN ; U7601
g5250 nand U2546 INSTQUEUE_REG_0__4__SCAN_IN ; U7602
g5251 nand U4040 U4039 U4038 U4037 ; U7603
g5252 nand U4180 INSTQUEUE_REG_0__4__SCAN_IN ; U7604
g5253 nand U2573 INSTQUEUE_REG_0__4__SCAN_IN ; U7605
g5254 nand U4079 U4077 U4076 U4075 ; U7606
g5255 nand U2592 INSTQUEUE_REG_0__4__SCAN_IN ; U7607
g5256 nand U4124 U4123 U4122 U4121 ; U7608
g5257 not U3246 ; U7609
g5258 nand U7609 U3248 ; U7610
g5259 nand U4349 U4346 STATE_REG_1__SCAN_IN ; U7611
g5260 nand U7456 STATE_REG_2__SCAN_IN ; U7612
g5261 nand U4346 STATE_REG_1__SCAN_IN ; U7613
g5262 nand U4490 U4498 ; U7614
g5263 nand U5475 U4159 ; U7615
g5264 nand U3270 U3276 ; U7616
g5265 not U3379 ; U7617
g5266 nand U4196 U7478 ; U7618
g5267 nand U5475 U4159 ; U7619
g5268 nand U7619 U7618 ; U7620
g5269 nand U3236 BE_N_REG_3__SCAN_IN ; U7621
g5270 nand U4209 BYTEENABLE_REG_3__SCAN_IN ; U7622
g5271 nand U3236 BE_N_REG_2__SCAN_IN ; U7623
g5272 nand U4209 BYTEENABLE_REG_2__SCAN_IN ; U7624
g5273 nand U3236 BE_N_REG_1__SCAN_IN ; U7625
g5274 nand U4209 BYTEENABLE_REG_1__SCAN_IN ; U7626
g5275 nand U3236 BE_N_REG_0__SCAN_IN ; U7627
g5276 nand U4209 BYTEENABLE_REG_0__SCAN_IN ; U7628
g5277 nand U3238 STATE_REG_0__SCAN_IN REQUESTPENDING_REG_SCAN_IN ; U7629
g5278 nand U3246 STATE_REG_2__SCAN_IN ; U7630
g5279 nand U7630 U7629 ; U7631
g5280 nand U7612 U4349 STATE_REG_1__SCAN_IN ; U7632
g5281 nand U7631 U3235 ; U7633
g5282 nand U3247 STATE_REG_2__SCAN_IN STATE_REG_0__SCAN_IN ; U7634
g5283 nand U4359 U3238 ; U7635
g5284 or STATE_REG_1__SCAN_IN STATE_REG_0__SCAN_IN ; U7636
g5285 nand U4246 STATE_REG_0__SCAN_IN ; U7637
g5286 not U3449 ; U7638
g5287 nand U7638 DATAWIDTH_REG_0__SCAN_IN ; U7639
g5288 nand U3450 U3449 ; U7640
g5289 nand U3449 U4364 ; U7641
g5290 nand U7638 DATAWIDTH_REG_1__SCAN_IN ; U7642
g5291 nand U3529 U3528 U3252 ; U7643
g5292 nand U3257 INSTQUEUE_REG_7__4__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7644
g5293 nand U3257 U3252 INSTQUEUE_REG_5__4__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7645
g5294 nand U3257 U3251 U3253 INSTQUEUE_REG_2__4__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7646
g5295 nand U3531 U3530 U3257 ; U7647
g5296 nand U3533 U3532 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7648
g5297 nand U3535 U3534 U3252 ; U7649
g5298 nand U3537 U3536 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7650
g5299 nand U3539 U3538 U3253 ; U7651
g5300 nand INSTQUEUE_REG_15__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_2__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7652
g5301 nand U3251 U3252 U3253 U3257 INSTQUEUE_REG_0__4__SCAN_IN ; U7653
g5302 nand U3251 U3252 U3253 INSTQUEUE_REG_8__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7654
g5303 nand U3251 U3253 INSTQUEUE_REG_10__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7655
g5304 nand U3541 U3540 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7656
g5305 nand U3251 U3257 INSTQUEUE_REG_3__4__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7657
g5306 nand U3251 INSTQUEUE_REG_11__4__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7658
g5307 nand U3251 U3257 INSTQUEUE_REG_3__5__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7659
g5308 nand U3517 U3516 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7660
g5309 nand U3251 U3252 INSTQUEUE_REG_9__6__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7661
g5310 nand U3523 U3522 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7662
g5311 nand U3251 U3253 INSTQUEUE_REG_10__6__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7663
g5312 nand U3251 INSTQUEUE_REG_11__6__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN INSTQUEUERD_ADDR_REG_1__SCAN_IN INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7664
g5313 nand U3251 U3252 U3253 U3257 INSTQUEUE_REG_0__6__SCAN_IN ; U7665
g5314 nand U3251 U3252 U3253 INSTQUEUE_REG_8__6__SCAN_IN INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7666
g5315 nand U4482 U3424 ; U7667
g5316 nand U7489 U3271 ; U7668
g5317 nand U4204 R2167_U17 ; U7669
g5318 nand U4494 U3260 ; U7670
g5319 nand U4500 STATE2_REG_0__SCAN_IN ; U7671
g5320 nand U4501 U3281 ; U7672
g5321 nand U3282 STATE2_REG_3__SCAN_IN ; U7673
g5322 nand U2428 U4502 ; U7674
g5323 or STATE2_REG_0__SCAN_IN STATEBS16_REG_SCAN_IN ; U7675
g5324 nand U7457 STATE2_REG_0__SCAN_IN ; U7676
g5325 nand U4510 STATE2_REG_0__SCAN_IN ; U7677
g5326 nand U7592 U4509 U3281 ; U7678
g5327 nand R2144_U49 U3300 ; U7679
g5328 nand U4516 U3298 ; U7680
g5329 not U3441 ; U7681
g5330 nand U3292 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U7682
g5331 nand U4521 U3291 ; U7683
g5332 not U3442 ; U7684
g5333 nand U4204 U3260 ; U7685
g5334 nand R2167_U17 U7485 ; U7686
g5335 nand U4420 U5454 ; U7687
g5336 nand U5455 U4159 ; U7688
g5337 nand U3454 U4160 ; U7689
g5338 nand U5464 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; U7690
g5339 nand U4448 U3265 ; U7691
g5340 nand U4403 U3264 ; U7692
g5341 nand U3258 U3402 ; U7693
g5342 nand U4465 U5481 ; U7694
g5343 nand U7694 U7693 ; U7695
g5344 nand U5464 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7696
g5345 nand U5497 U4160 ; U7697
g5346 nand U4162 INSTADDRPOINTER_REG_1__SCAN_IN ; U7698
g5347 nand SUB_580_U6 INSTADDRPOINTER_REG_31__SCAN_IN ; U7699
g5348 not U3457 ; U7700
g5349 nand U4162 INSTADDRPOINTER_REG_0__SCAN_IN ; U7701
g5350 nand INSTADDRPOINTER_REG_0__SCAN_IN INSTADDRPOINTER_REG_31__SCAN_IN ; U7702
g5351 not U3458 ; U7703
g5352 nand U5499 U5489 ; U7704
g5353 nand U4206 U3388 ; U7705
g5354 nand U3251 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7706
g5355 nand U3252 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U7707
g5356 not U3443 ; U7708
g5357 nand U5464 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U7709
g5358 nand U5506 U4160 ; U7710
g5359 nand U5464 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7711
g5360 nand U5517 U4160 ; U7712
g5361 nand U4202 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7713
g5362 nand U5509 U3253 ; U7714
g5363 nand U5464 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7715
g5364 nand U5523 U4160 ; U7716
g5365 nand U5525 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; U7717
g5366 nand U5533 U3391 ; U7718
g5367 nand U7681 U4515 ; U7719
g5368 nand U3441 U3301 ; U7720
g5369 nand U7720 U7719 ; U7721
g5370 nand U5525 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; U7722
g5371 nand U5537 U3391 ; U7723
g5372 nand U5525 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; U7724
g5373 nand U5542 U3391 ; U7725
g5374 nand U5525 INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; U7726
g5375 nand U5545 U3391 ; U7727
g5376 nand U4465 U3375 ; U7728
g5377 nand U3258 U3268 ; U7729
g5378 nand U7729 U7728 U3244 U4159 ; U7730
g5379 nand R2167_U17 U7599 U4420 ; U7731
g5380 nand U3411 EAX_REG_31__SCAN_IN ; U7732
g5381 nand U3466 U4211 ; U7733
g5382 nand U3420 BYTEENABLE_REG_3__SCAN_IN ; U7734
g5383 nand U3467 U4208 ; U7735
g5384 or DATAWIDTH_REG_0__SCAN_IN DATAWIDTH_REG_1__SCAN_IN ; U7736
g5385 nand U3400 DATAWIDTH_REG_0__SCAN_IN ; U7737
g5386 nand U7737 U7736 ; U7738
g5387 nand U7738 U3240 ; U7739
g5388 nand REIP_REG_0__SCAN_IN REIP_REG_1__SCAN_IN ; U7740
g5389 nand U7740 U7739 ; U7741
g5390 nand U3420 BYTEENABLE_REG_2__SCAN_IN ; U7742
g5391 nand U7741 U4208 ; U7743
g5392 nand U3420 BYTEENABLE_REG_1__SCAN_IN ; U7744
g5393 nand U4208 REIP_REG_1__SCAN_IN ; U7745
g5394 nand U3420 BYTEENABLE_REG_0__SCAN_IN ; U7746
g5395 nand U4208 U6587 ; U7747
g5396 nand U4209 U3423 ; U7748
g5397 nand U3236 W_R_N_REG_SCAN_IN ; U7749
g5398 nand U4165 MORE_REG_SCAN_IN ; U7750
g5399 nand U4225 U6588 ; U7751
g5400 nand U7638 STATEBS16_REG_SCAN_IN ; U7752
g5401 nand BS16_N U3449 ; U7753
g5402 nand U6591 REQUESTPENDING_REG_SCAN_IN ; U7754
g5403 nand U6597 U4168 ; U7755
g5404 nand U4209 U3422 ; U7756
g5405 nand U3236 D_C_N_REG_SCAN_IN ; U7757
g5406 nand U3236 M_IO_N_REG_SCAN_IN ; U7758
g5407 nand U4209 MEMORYFETCH_REG_SCAN_IN ; U7759
g5408 nand U6602 READREQUEST_REG_SCAN_IN ; U7760
g5409 nand U6603 U4169 ; U7761
g5410 nand U3475 U4170 ; U7762
g5411 nand U5461 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; U7763
g5412 nand U5461 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7764
g5413 nand U5494 U4170 ; U7765
g5414 nand U5461 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; U7766
g5415 nand U5502 U4170 ; U7767
g5416 nand U5461 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; U7768
g5417 nand U5513 U4170 ; U7769
g5418 nand U5461 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; U7770
g5419 nand U5519 U4170 ; U7771
g5420 nand U2605 U3264 ; U7772
g5421 nand U4448 U7483 ; U7773
g5422 nand U4191 U3288 ; U7774
g5423 nand U3284 INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; U7775
g5424 nand U4171 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; U7776
g5425 nand U7207 U3257 ; U7777
g5426 not U3444 ; U7778
g5427 nand U3263 U3271 ; U7779
g5428 nand U7695 U4482 ; U7780
g5429 nand U3480 U3249 ; U7781
g5430 nand U7703 STATE2_REG_1__SCAN_IN FLUSH_REG_SCAN_IN ; U7782
g5431 not INSTADDRPOINTER_REG_0__SCAN_IN ; R2027_U5
g5432 not INSTADDRPOINTER_REG_2__SCAN_IN ; R2027_U6
g5433 not INSTADDRPOINTER_REG_1__SCAN_IN ; R2027_U7
g5434 not INSTADDRPOINTER_REG_4__SCAN_IN ; R2027_U8
g5435 not INSTADDRPOINTER_REG_3__SCAN_IN ; R2027_U9
g5436 nand INSTADDRPOINTER_REG_0__SCAN_IN INSTADDRPOINTER_REG_1__SCAN_IN INSTADDRPOINTER_REG_2__SCAN_IN ; R2027_U10
g5437 not INSTADDRPOINTER_REG_6__SCAN_IN ; R2027_U11
g5438 not INSTADDRPOINTER_REG_5__SCAN_IN ; R2027_U12
g5439 nand R2027_U82 R2027_U111 ; R2027_U13
g5440 not INSTADDRPOINTER_REG_8__SCAN_IN ; R2027_U14
g5441 not INSTADDRPOINTER_REG_7__SCAN_IN ; R2027_U15
g5442 nand R2027_U83 R2027_U112 ; R2027_U16
g5443 nand R2027_U84 R2027_U118 ; R2027_U17
g5444 not INSTADDRPOINTER_REG_9__SCAN_IN ; R2027_U18
g5445 not INSTADDRPOINTER_REG_10__SCAN_IN ; R2027_U19
g5446 not INSTADDRPOINTER_REG_12__SCAN_IN ; R2027_U20
g5447 not INSTADDRPOINTER_REG_11__SCAN_IN ; R2027_U21
g5448 nand R2027_U85 R2027_U120 ; R2027_U22
g5449 not INSTADDRPOINTER_REG_14__SCAN_IN ; R2027_U23
g5450 not INSTADDRPOINTER_REG_13__SCAN_IN ; R2027_U24
g5451 nand R2027_U86 R2027_U113 ; R2027_U25
g5452 not INSTADDRPOINTER_REG_15__SCAN_IN ; R2027_U26
g5453 nand R2027_U87 R2027_U119 ; R2027_U27
g5454 not INSTADDRPOINTER_REG_16__SCAN_IN ; R2027_U28
g5455 not INSTADDRPOINTER_REG_18__SCAN_IN ; R2027_U29
g5456 not INSTADDRPOINTER_REG_17__SCAN_IN ; R2027_U30
g5457 nand R2027_U88 R2027_U124 ; R2027_U31
g5458 not INSTADDRPOINTER_REG_20__SCAN_IN ; R2027_U32
g5459 not INSTADDRPOINTER_REG_19__SCAN_IN ; R2027_U33
g5460 nand R2027_U89 R2027_U117 ; R2027_U34
g5461 not INSTADDRPOINTER_REG_21__SCAN_IN ; R2027_U35
g5462 nand R2027_U90 R2027_U114 ; R2027_U36
g5463 not INSTADDRPOINTER_REG_22__SCAN_IN ; R2027_U37
g5464 not INSTADDRPOINTER_REG_24__SCAN_IN ; R2027_U38
g5465 not INSTADDRPOINTER_REG_23__SCAN_IN ; R2027_U39
g5466 nand R2027_U91 R2027_U121 ; R2027_U40
g5467 not INSTADDRPOINTER_REG_26__SCAN_IN ; R2027_U41
g5468 not INSTADDRPOINTER_REG_25__SCAN_IN ; R2027_U42
g5469 nand R2027_U92 R2027_U115 ; R2027_U43
g5470 not INSTADDRPOINTER_REG_27__SCAN_IN ; R2027_U44
g5471 not INSTADDRPOINTER_REG_28__SCAN_IN ; R2027_U45
g5472 nand R2027_U93 R2027_U116 ; R2027_U46
g5473 not INSTADDRPOINTER_REG_29__SCAN_IN ; R2027_U47
g5474 nand R2027_U94 R2027_U122 ; R2027_U48
g5475 nand R2027_U123 INSTADDRPOINTER_REG_29__SCAN_IN ; R2027_U49
g5476 not INSTADDRPOINTER_REG_30__SCAN_IN ; R2027_U50
g5477 nand R2027_U142 R2027_U141 ; R2027_U51
g5478 nand R2027_U144 R2027_U143 ; R2027_U52
g5479 nand R2027_U146 R2027_U145 ; R2027_U53
g5480 nand R2027_U148 R2027_U147 ; R2027_U54
g5481 nand R2027_U150 R2027_U149 ; R2027_U55
g5482 nand R2027_U152 R2027_U151 ; R2027_U56
g5483 nand R2027_U154 R2027_U153 ; R2027_U57
g5484 nand R2027_U156 R2027_U155 ; R2027_U58
g5485 nand R2027_U158 R2027_U157 ; R2027_U59
g5486 nand R2027_U160 R2027_U159 ; R2027_U60
g5487 nand R2027_U162 R2027_U161 ; R2027_U61
g5488 nand R2027_U164 R2027_U163 ; R2027_U62
g5489 nand R2027_U166 R2027_U165 ; R2027_U63
g5490 nand R2027_U168 R2027_U167 ; R2027_U64
g5491 nand R2027_U170 R2027_U169 ; R2027_U65
g5492 nand R2027_U172 R2027_U171 ; R2027_U66
g5493 nand R2027_U174 R2027_U173 ; R2027_U67
g5494 nand R2027_U176 R2027_U175 ; R2027_U68
g5495 nand R2027_U178 R2027_U177 ; R2027_U69
g5496 nand R2027_U180 R2027_U179 ; R2027_U70
g5497 nand R2027_U182 R2027_U181 ; R2027_U71
g5498 nand R2027_U184 R2027_U183 ; R2027_U72
g5499 nand R2027_U186 R2027_U185 ; R2027_U73
g5500 nand R2027_U188 R2027_U187 ; R2027_U74
g5501 nand R2027_U190 R2027_U189 ; R2027_U75
g5502 nand R2027_U192 R2027_U191 ; R2027_U76
g5503 nand R2027_U194 R2027_U193 ; R2027_U77
g5504 nand R2027_U196 R2027_U195 ; R2027_U78
g5505 nand R2027_U198 R2027_U197 ; R2027_U79
g5506 nand R2027_U200 R2027_U199 ; R2027_U80
g5507 nand R2027_U202 R2027_U201 ; R2027_U81
g5508 and INSTADDRPOINTER_REG_3__SCAN_IN INSTADDRPOINTER_REG_4__SCAN_IN ; R2027_U82
g5509 and INSTADDRPOINTER_REG_5__SCAN_IN INSTADDRPOINTER_REG_6__SCAN_IN ; R2027_U83
g5510 and INSTADDRPOINTER_REG_7__SCAN_IN INSTADDRPOINTER_REG_8__SCAN_IN ; R2027_U84
g5511 and INSTADDRPOINTER_REG_9__SCAN_IN INSTADDRPOINTER_REG_10__SCAN_IN ; R2027_U85
g5512 and INSTADDRPOINTER_REG_11__SCAN_IN INSTADDRPOINTER_REG_12__SCAN_IN ; R2027_U86
g5513 and INSTADDRPOINTER_REG_13__SCAN_IN INSTADDRPOINTER_REG_14__SCAN_IN ; R2027_U87
g5514 and INSTADDRPOINTER_REG_15__SCAN_IN INSTADDRPOINTER_REG_16__SCAN_IN ; R2027_U88
g5515 and INSTADDRPOINTER_REG_17__SCAN_IN INSTADDRPOINTER_REG_18__SCAN_IN ; R2027_U89
g5516 and INSTADDRPOINTER_REG_19__SCAN_IN INSTADDRPOINTER_REG_20__SCAN_IN ; R2027_U90
g5517 and INSTADDRPOINTER_REG_21__SCAN_IN INSTADDRPOINTER_REG_22__SCAN_IN ; R2027_U91
g5518 and INSTADDRPOINTER_REG_23__SCAN_IN INSTADDRPOINTER_REG_24__SCAN_IN ; R2027_U92
g5519 and INSTADDRPOINTER_REG_25__SCAN_IN INSTADDRPOINTER_REG_26__SCAN_IN ; R2027_U93
g5520 and INSTADDRPOINTER_REG_27__SCAN_IN INSTADDRPOINTER_REG_28__SCAN_IN ; R2027_U94
g5521 nand R2027_U118 INSTADDRPOINTER_REG_7__SCAN_IN ; R2027_U95
g5522 nand R2027_U112 INSTADDRPOINTER_REG_5__SCAN_IN ; R2027_U96
g5523 nand R2027_U111 INSTADDRPOINTER_REG_3__SCAN_IN ; R2027_U97
g5524 not INSTADDRPOINTER_REG_31__SCAN_IN ; R2027_U98
g5525 nand R2027_U128 INSTADDRPOINTER_REG_30__SCAN_IN ; R2027_U99
g5526 nand INSTADDRPOINTER_REG_0__SCAN_IN INSTADDRPOINTER_REG_1__SCAN_IN ; R2027_U100
g5527 nand R2027_U122 INSTADDRPOINTER_REG_27__SCAN_IN ; R2027_U101
g5528 nand R2027_U116 INSTADDRPOINTER_REG_25__SCAN_IN ; R2027_U102
g5529 nand R2027_U115 INSTADDRPOINTER_REG_23__SCAN_IN ; R2027_U103
g5530 nand R2027_U121 INSTADDRPOINTER_REG_21__SCAN_IN ; R2027_U104
g5531 nand R2027_U114 INSTADDRPOINTER_REG_19__SCAN_IN ; R2027_U105
g5532 nand R2027_U117 INSTADDRPOINTER_REG_17__SCAN_IN ; R2027_U106
g5533 nand R2027_U124 INSTADDRPOINTER_REG_15__SCAN_IN ; R2027_U107
g5534 nand R2027_U119 INSTADDRPOINTER_REG_13__SCAN_IN ; R2027_U108
g5535 nand R2027_U113 INSTADDRPOINTER_REG_11__SCAN_IN ; R2027_U109
g5536 nand R2027_U120 INSTADDRPOINTER_REG_9__SCAN_IN ; R2027_U110
g5537 not R2027_U10 ; R2027_U111
g5538 not R2027_U13 ; R2027_U112
g5539 not R2027_U22 ; R2027_U113
g5540 not R2027_U34 ; R2027_U114
g5541 not R2027_U40 ; R2027_U115
g5542 not R2027_U43 ; R2027_U116
g5543 not R2027_U31 ; R2027_U117
g5544 not R2027_U16 ; R2027_U118
g5545 not R2027_U25 ; R2027_U119
g5546 not R2027_U17 ; R2027_U120
g5547 not R2027_U36 ; R2027_U121
g5548 not R2027_U46 ; R2027_U122
g5549 not R2027_U48 ; R2027_U123
g5550 not R2027_U27 ; R2027_U124
g5551 not R2027_U95 ; R2027_U125
g5552 not R2027_U96 ; R2027_U126
g5553 not R2027_U97 ; R2027_U127
g5554 not R2027_U49 ; R2027_U128
g5555 not R2027_U99 ; R2027_U129
g5556 not R2027_U100 ; R2027_U130
g5557 not R2027_U101 ; R2027_U131
g5558 not R2027_U102 ; R2027_U132
g5559 not R2027_U103 ; R2027_U133
g5560 not R2027_U104 ; R2027_U134
g5561 not R2027_U105 ; R2027_U135
g5562 not R2027_U106 ; R2027_U136
g5563 not R2027_U107 ; R2027_U137
g5564 not R2027_U108 ; R2027_U138
g5565 not R2027_U109 ; R2027_U139
g5566 not R2027_U110 ; R2027_U140
g5567 nand R2027_U120 R2027_U18 ; R2027_U141
g5568 nand R2027_U17 INSTADDRPOINTER_REG_9__SCAN_IN ; R2027_U142
g5569 nand R2027_U95 INSTADDRPOINTER_REG_8__SCAN_IN ; R2027_U143
g5570 nand R2027_U125 R2027_U14 ; R2027_U144
g5571 nand R2027_U118 R2027_U15 ; R2027_U145
g5572 nand R2027_U16 INSTADDRPOINTER_REG_7__SCAN_IN ; R2027_U146
g5573 nand R2027_U96 INSTADDRPOINTER_REG_6__SCAN_IN ; R2027_U147
g5574 nand R2027_U126 R2027_U11 ; R2027_U148
g5575 nand R2027_U112 R2027_U12 ; R2027_U149
g5576 nand R2027_U13 INSTADDRPOINTER_REG_5__SCAN_IN ; R2027_U150
g5577 nand R2027_U97 INSTADDRPOINTER_REG_4__SCAN_IN ; R2027_U151
g5578 nand R2027_U127 R2027_U8 ; R2027_U152
g5579 nand R2027_U111 R2027_U9 ; R2027_U153
g5580 nand R2027_U10 INSTADDRPOINTER_REG_3__SCAN_IN ; R2027_U154
g5581 nand R2027_U99 INSTADDRPOINTER_REG_31__SCAN_IN ; R2027_U155
g5582 nand R2027_U129 R2027_U98 ; R2027_U156
g5583 nand R2027_U49 INSTADDRPOINTER_REG_30__SCAN_IN ; R2027_U157
g5584 nand R2027_U128 R2027_U50 ; R2027_U158
g5585 nand R2027_U100 INSTADDRPOINTER_REG_2__SCAN_IN ; R2027_U159
g5586 nand R2027_U130 R2027_U6 ; R2027_U160
g5587 nand R2027_U123 R2027_U47 ; R2027_U161
g5588 nand R2027_U48 INSTADDRPOINTER_REG_29__SCAN_IN ; R2027_U162
g5589 nand R2027_U101 INSTADDRPOINTER_REG_28__SCAN_IN ; R2027_U163
g5590 nand R2027_U131 R2027_U45 ; R2027_U164
g5591 nand R2027_U122 R2027_U44 ; R2027_U165
g5592 nand R2027_U46 INSTADDRPOINTER_REG_27__SCAN_IN ; R2027_U166
g5593 nand R2027_U102 INSTADDRPOINTER_REG_26__SCAN_IN ; R2027_U167
g5594 nand R2027_U132 R2027_U41 ; R2027_U168
g5595 nand R2027_U116 R2027_U42 ; R2027_U169
g5596 nand R2027_U43 INSTADDRPOINTER_REG_25__SCAN_IN ; R2027_U170
g5597 nand R2027_U103 INSTADDRPOINTER_REG_24__SCAN_IN ; R2027_U171
g5598 nand R2027_U133 R2027_U38 ; R2027_U172
g5599 nand R2027_U115 R2027_U39 ; R2027_U173
g5600 nand R2027_U40 INSTADDRPOINTER_REG_23__SCAN_IN ; R2027_U174
g5601 nand R2027_U104 INSTADDRPOINTER_REG_22__SCAN_IN ; R2027_U175
g5602 nand R2027_U134 R2027_U37 ; R2027_U176
g5603 nand R2027_U121 R2027_U35 ; R2027_U177
g5604 nand R2027_U36 INSTADDRPOINTER_REG_21__SCAN_IN ; R2027_U178
g5605 nand R2027_U105 INSTADDRPOINTER_REG_20__SCAN_IN ; R2027_U179
g5606 nand R2027_U135 R2027_U32 ; R2027_U180
g5607 nand R2027_U7 INSTADDRPOINTER_REG_0__SCAN_IN ; R2027_U181
g5608 nand R2027_U5 INSTADDRPOINTER_REG_1__SCAN_IN ; R2027_U182
g5609 nand R2027_U114 R2027_U33 ; R2027_U183
g5610 nand R2027_U34 INSTADDRPOINTER_REG_19__SCAN_IN ; R2027_U184
g5611 nand R2027_U106 INSTADDRPOINTER_REG_18__SCAN_IN ; R2027_U185
g5612 nand R2027_U136 R2027_U29 ; R2027_U186
g5613 nand R2027_U117 R2027_U30 ; R2027_U187
g5614 nand R2027_U31 INSTADDRPOINTER_REG_17__SCAN_IN ; R2027_U188
g5615 nand R2027_U107 INSTADDRPOINTER_REG_16__SCAN_IN ; R2027_U189
g5616 nand R2027_U137 R2027_U28 ; R2027_U190
g5617 nand R2027_U124 R2027_U26 ; R2027_U191
g5618 nand R2027_U27 INSTADDRPOINTER_REG_15__SCAN_IN ; R2027_U192
g5619 nand R2027_U108 INSTADDRPOINTER_REG_14__SCAN_IN ; R2027_U193
g5620 nand R2027_U138 R2027_U23 ; R2027_U194
g5621 nand R2027_U119 R2027_U24 ; R2027_U195
g5622 nand R2027_U25 INSTADDRPOINTER_REG_13__SCAN_IN ; R2027_U196
g5623 nand R2027_U109 INSTADDRPOINTER_REG_12__SCAN_IN ; R2027_U197
g5624 nand R2027_U139 R2027_U20 ; R2027_U198
g5625 nand R2027_U113 R2027_U21 ; R2027_U199
g5626 nand R2027_U22 INSTADDRPOINTER_REG_11__SCAN_IN ; R2027_U200
g5627 nand R2027_U110 INSTADDRPOINTER_REG_10__SCAN_IN ; R2027_U201
g5628 nand R2027_U140 R2027_U19 ; R2027_U202
g5629 and R2278_U217 R2278_U215 ; R2278_U5
g5630 and R2278_U227 R2278_U225 ; R2278_U6
g5631 and R2278_U6 R2278_U208 ; R2278_U7
g5632 and R2278_U7 R2278_U207 ; R2278_U8
g5633 and R2278_U235 R2278_U231 ; R2278_U9
g5634 and R2278_U9 R2278_U206 ; R2278_U10
g5635 and R2278_U10 R2278_U205 ; R2278_U11
g5636 and R2278_U11 R2278_U242 ; R2278_U12
g5637 and R2278_U12 R2278_U204 ; R2278_U13
g5638 and R2278_U250 R2278_U246 ; R2278_U14
g5639 and R2278_U14 R2278_U253 ; R2278_U15
g5640 and R2278_U15 R2278_U256 ; R2278_U16
g5641 and R2278_U292 R2278_U19 ; R2278_U17
g5642 nand U2783 INSTADDRPOINTER_REG_4__SCAN_IN ; R2278_U18
g5643 nand U2787 INSTADDRPOINTER_REG_0__SCAN_IN ; R2278_U19
g5644 nand U2782 INSTADDRPOINTER_REG_5__SCAN_IN ; R2278_U20
g5645 not INSTADDRPOINTER_REG_30__SCAN_IN ; R2278_U21
g5646 not U2770 ; R2278_U22
g5647 nand U2770 INSTADDRPOINTER_REG_19__SCAN_IN ; R2278_U23
g5648 nand U2771 INSTADDRPOINTER_REG_16__SCAN_IN ; R2278_U24
g5649 nand R2278_U40 R2278_U207 ; R2278_U25
g5650 nand U2779 INSTADDRPOINTER_REG_8__SCAN_IN ; R2278_U26
g5651 nand U2778 INSTADDRPOINTER_REG_9__SCAN_IN ; R2278_U27
g5652 nand U2777 INSTADDRPOINTER_REG_10__SCAN_IN ; R2278_U28
g5653 nand U2775 INSTADDRPOINTER_REG_12__SCAN_IN ; R2278_U29
g5654 nand U2773 INSTADDRPOINTER_REG_14__SCAN_IN ; R2278_U30
g5655 nand U2774 INSTADDRPOINTER_REG_13__SCAN_IN ; R2278_U31
g5656 not INSTADDRPOINTER_REG_29__SCAN_IN ; R2278_U32
g5657 not U2770 ; R2278_U33
g5658 not INSTADDRPOINTER_REG_28__SCAN_IN ; R2278_U34
g5659 not U2770 ; R2278_U35
g5660 nand U2770 INSTADDRPOINTER_REG_26__SCAN_IN ; R2278_U36
g5661 nand R2278_U328 R2278_U257 ; R2278_U37
g5662 nand R2278_U325 R2278_U254 ; R2278_U38
g5663 nand R2278_U322 R2278_U251 ; R2278_U39
g5664 nand R2278_U306 R2278_U229 ; R2278_U40
g5665 nand R2278_U304 R2278_U228 ; R2278_U41
g5666 nand R2278_U402 R2278_U401 ; R2278_U42
g5667 and R2278_U178 R2278_U162 ; R2278_U43
g5668 and R2278_U303 R2278_U179 ; R2278_U44
g5669 and R2278_U182 R2278_U163 ; R2278_U45
g5670 and R2278_U302 R2278_U301 ; R2278_U46
g5671 and U2770 INSTADDRPOINTER_REG_20__SCAN_IN ; R2278_U47
g5672 and R2278_U178 R2278_U162 ; R2278_U48
g5673 and R2278_U337 R2278_U179 ; R2278_U49
g5674 and R2278_U301 R2278_U163 R2278_U182 ; R2278_U50
g5675 and R2278_U189 R2278_U185 ; R2278_U51
g5676 and R2278_U5 R2278_U51 ; R2278_U52
g5677 and R2278_U186 R2278_U189 ; R2278_U53
g5678 and R2278_U293 R2278_U216 R2278_U296 R2278_U295 ; R2278_U54
g5679 and R2278_U211 R2278_U213 R2278_U221 R2278_U209 ; R2278_U55
g5680 and R2278_U294 R2278_U210 R2278_U298 R2278_U297 ; R2278_U56
g5681 and R2278_U13 R2278_U8 ; R2278_U57
g5682 and R2278_U332 R2278_U245 ; R2278_U58
g5683 and R2278_U333 R2278_U320 R2278_U58 ; R2278_U59
g5684 and R2278_U16 R2278_U259 ; R2278_U60
g5685 and R2278_U331 R2278_U260 ; R2278_U61
g5686 nand R2278_U364 R2278_U363 ; R2278_U62
g5687 nand R2278_U369 R2278_U368 ; R2278_U63
g5688 nand R2278_U376 R2278_U375 ; R2278_U64
g5689 nand R2278_U381 R2278_U380 ; R2278_U65
g5690 and R2278_U25 R2278_U23 ; R2278_U66
g5691 and R2278_U318 R2278_U243 ; R2278_U67
g5692 and R2278_U315 R2278_U240 ; R2278_U68
g5693 and R2278_U312 R2278_U238 ; R2278_U69
g5694 and R2278_U310 R2278_U236 ; R2278_U70
g5695 and R2278_U293 R2278_U216 R2278_U296 R2278_U295 ; R2278_U71
g5696 nand R2278_U26 R2278_U187 ; R2278_U72
g5697 nand R2278_U189 R2278_U27 ; R2278_U73
g5698 and R2278_U350 R2278_U349 ; R2278_U74
g5699 nand R2278_U46 R2278_U183 R2278_U45 ; R2278_U75
g5700 nand R2278_U185 R2278_U26 ; R2278_U76
g5701 and R2278_U352 R2278_U351 ; R2278_U77
g5702 nand R2278_U197 R2278_U165 ; R2278_U78
g5703 nand R2278_U162 R2278_U163 ; R2278_U79
g5704 and R2278_U354 R2278_U353 ; R2278_U80
g5705 nand R2278_U20 R2278_U195 ; R2278_U81
g5706 nand R2278_U165 R2278_U164 ; R2278_U82
g5707 and R2278_U356 R2278_U355 ; R2278_U83
g5708 nand R2278_U18 R2278_U193 ; R2278_U84
g5709 nand R2278_U179 R2278_U20 ; R2278_U85
g5710 and R2278_U358 R2278_U357 ; R2278_U86
g5711 nand R2278_U175 R2278_U176 ; R2278_U87
g5712 nand R2278_U178 R2278_U18 ; R2278_U88
g5713 and R2278_U360 R2278_U359 ; R2278_U89
g5714 nand R2278_U172 R2278_U173 ; R2278_U90
g5715 nand R2278_U166 R2278_U175 ; R2278_U91
g5716 and R2278_U362 R2278_U361 ; R2278_U92
g5717 not U2769 ; R2278_U93
g5718 not INSTADDRPOINTER_REG_31__SCAN_IN ; R2278_U94
g5719 nand R2278_U61 R2278_U330 ; R2278_U95
g5720 and R2278_U367 R2278_U366 ; R2278_U96
g5721 nand R2278_U329 R2278_U327 ; R2278_U97
g5722 and R2278_U372 R2278_U371 ; R2278_U98
g5723 nand R2278_U169 R2278_U170 ; R2278_U99
g5724 nand R2278_U167 R2278_U172 ; R2278_U100
g5725 and R2278_U374 R2278_U373 ; R2278_U101
g5726 nand R2278_U326 R2278_U324 ; R2278_U102
g5727 and R2278_U379 R2278_U378 ; R2278_U103
g5728 nand R2278_U323 R2278_U321 ; R2278_U104
g5729 and R2278_U384 R2278_U383 ; R2278_U105
g5730 nand R2278_U36 R2278_U248 ; R2278_U106
g5731 nand R2278_U250 R2278_U251 ; R2278_U107
g5732 and R2278_U386 R2278_U385 ; R2278_U108
g5733 nand R2278_U246 R2278_U36 ; R2278_U109
g5734 nand R2278_U59 R2278_U347 ; R2278_U110
g5735 and R2278_U388 R2278_U387 ; R2278_U111
g5736 nand R2278_U67 R2278_U316 ; R2278_U112
g5737 nand R2278_U204 R2278_U245 ; R2278_U113
g5738 and R2278_U390 R2278_U389 ; R2278_U114
g5739 nand R2278_U68 R2278_U313 ; R2278_U115
g5740 nand R2278_U243 R2278_U242 ; R2278_U116
g5741 and R2278_U392 R2278_U391 ; R2278_U117
g5742 nand R2278_U69 R2278_U311 ; R2278_U118
g5743 nand R2278_U240 R2278_U205 ; R2278_U119
g5744 and R2278_U394 R2278_U393 ; R2278_U120
g5745 nand R2278_U70 R2278_U309 ; R2278_U121
g5746 nand R2278_U238 R2278_U206 ; R2278_U122
g5747 and R2278_U396 R2278_U395 ; R2278_U123
g5748 nand R2278_U232 R2278_U233 ; R2278_U124
g5749 nand R2278_U236 R2278_U235 ; R2278_U125
g5750 and R2278_U398 R2278_U397 ; R2278_U126
g5751 nand R2278_U231 R2278_U232 ; R2278_U127
g5752 nand R2278_U66 R2278_U345 ; R2278_U128
g5753 and R2278_U400 R2278_U399 ; R2278_U129
g5754 nand R2278_U168 R2278_U169 ; R2278_U130
g5755 nand R2278_U207 R2278_U23 ; R2278_U131
g5756 nand R2278_U307 R2278_U343 ; R2278_U132
g5757 and R2278_U404 R2278_U403 ; R2278_U133
g5758 nand R2278_U208 R2278_U229 ; R2278_U134
g5759 nand R2278_U305 R2278_U341 ; R2278_U135
g5760 and R2278_U406 R2278_U405 ; R2278_U136
g5761 nand R2278_U227 R2278_U228 ; R2278_U137
g5762 nand R2278_U339 R2278_U24 ; R2278_U138
g5763 and R2278_U408 R2278_U407 ; R2278_U139
g5764 nand R2278_U223 R2278_U56 ; R2278_U140
g5765 nand R2278_U225 R2278_U24 ; R2278_U141
g5766 and R2278_U410 R2278_U409 ; R2278_U142
g5767 nand R2278_U280 R2278_U30 ; R2278_U143
g5768 nand R2278_U209 R2278_U210 ; R2278_U144
g5769 and R2278_U412 R2278_U411 ; R2278_U145
g5770 nand R2278_U31 R2278_U278 ; R2278_U146
g5771 nand R2278_U30 R2278_U211 ; R2278_U147
g5772 and R2278_U414 R2278_U413 ; R2278_U148
g5773 nand R2278_U29 R2278_U276 ; R2278_U149
g5774 nand R2278_U213 R2278_U31 ; R2278_U150
g5775 and R2278_U416 R2278_U415 ; R2278_U151
g5776 nand R2278_U219 R2278_U71 ; R2278_U152
g5777 nand R2278_U221 R2278_U29 ; R2278_U153
g5778 and R2278_U418 R2278_U417 ; R2278_U154
g5779 nand R2278_U288 R2278_U28 ; R2278_U155
g5780 nand R2278_U215 R2278_U216 ; R2278_U156
g5781 and R2278_U420 R2278_U419 ; R2278_U157
g5782 nand R2278_U27 R2278_U286 ; R2278_U158
g5783 nand R2278_U28 R2278_U217 ; R2278_U159
g5784 and R2278_U422 R2278_U421 ; R2278_U160
g5785 not R2278_U19 ; R2278_U161
g5786 or U2780 INSTADDRPOINTER_REG_7__SCAN_IN ; R2278_U162
g5787 nand U2780 INSTADDRPOINTER_REG_7__SCAN_IN ; R2278_U163
g5788 or U2781 INSTADDRPOINTER_REG_6__SCAN_IN ; R2278_U164
g5789 nand U2781 INSTADDRPOINTER_REG_6__SCAN_IN ; R2278_U165
g5790 or U2784 INSTADDRPOINTER_REG_3__SCAN_IN ; R2278_U166
g5791 or U2785 INSTADDRPOINTER_REG_2__SCAN_IN ; R2278_U167
g5792 or U2786 INSTADDRPOINTER_REG_1__SCAN_IN ; R2278_U168
g5793 nand U2786 INSTADDRPOINTER_REG_1__SCAN_IN ; R2278_U169
g5794 nand R2278_U161 R2278_U168 ; R2278_U170
g5795 not R2278_U99 ; R2278_U171
g5796 nand U2785 INSTADDRPOINTER_REG_2__SCAN_IN ; R2278_U172
g5797 nand R2278_U99 R2278_U299 ; R2278_U173
g5798 not R2278_U90 ; R2278_U174
g5799 nand U2784 INSTADDRPOINTER_REG_3__SCAN_IN ; R2278_U175
g5800 nand R2278_U300 R2278_U166 ; R2278_U176
g5801 not R2278_U87 ; R2278_U177
g5802 or U2783 INSTADDRPOINTER_REG_4__SCAN_IN ; R2278_U178
g5803 or U2782 INSTADDRPOINTER_REG_5__SCAN_IN ; R2278_U179
g5804 not R2278_U20 ; R2278_U180
g5805 not R2278_U18 ; R2278_U181
g5806 nand R2278_U181 R2278_U179 R2278_U164 R2278_U162 ; R2278_U182
g5807 nand R2278_U43 R2278_U87 R2278_U44 ; R2278_U183
g5808 not R2278_U75 ; R2278_U184
g5809 or U2779 INSTADDRPOINTER_REG_8__SCAN_IN ; R2278_U185
g5810 not R2278_U26 ; R2278_U186
g5811 nand R2278_U185 R2278_U75 ; R2278_U187
g5812 not R2278_U72 ; R2278_U188
g5813 or U2778 INSTADDRPOINTER_REG_9__SCAN_IN ; R2278_U189
g5814 not R2278_U27 ; R2278_U190
g5815 not R2278_U73 ; R2278_U191
g5816 not R2278_U76 ; R2278_U192
g5817 nand R2278_U178 R2278_U87 ; R2278_U193
g5818 not R2278_U84 ; R2278_U194
g5819 nand R2278_U84 R2278_U179 ; R2278_U195
g5820 not R2278_U81 ; R2278_U196
g5821 nand R2278_U81 R2278_U164 ; R2278_U197
g5822 not R2278_U78 ; R2278_U198
g5823 not R2278_U79 ; R2278_U199
g5824 not R2278_U82 ; R2278_U200
g5825 not R2278_U85 ; R2278_U201
g5826 not R2278_U88 ; R2278_U202
g5827 not R2278_U91 ; R2278_U203
g5828 or U2770 INSTADDRPOINTER_REG_25__SCAN_IN ; R2278_U204
g5829 or U2770 INSTADDRPOINTER_REG_23__SCAN_IN ; R2278_U205
g5830 or U2770 INSTADDRPOINTER_REG_22__SCAN_IN ; R2278_U206
g5831 or U2770 INSTADDRPOINTER_REG_19__SCAN_IN ; R2278_U207
g5832 or U2770 INSTADDRPOINTER_REG_18__SCAN_IN ; R2278_U208
g5833 or U2772 INSTADDRPOINTER_REG_15__SCAN_IN ; R2278_U209
g5834 nand U2772 INSTADDRPOINTER_REG_15__SCAN_IN ; R2278_U210
g5835 or U2773 INSTADDRPOINTER_REG_14__SCAN_IN ; R2278_U211
g5836 not R2278_U30 ; R2278_U212
g5837 or U2774 INSTADDRPOINTER_REG_13__SCAN_IN ; R2278_U213
g5838 not R2278_U31 ; R2278_U214
g5839 or U2776 INSTADDRPOINTER_REG_11__SCAN_IN ; R2278_U215
g5840 nand U2776 INSTADDRPOINTER_REG_11__SCAN_IN ; R2278_U216
g5841 or U2777 INSTADDRPOINTER_REG_10__SCAN_IN ; R2278_U217
g5842 not R2278_U28 ; R2278_U218
g5843 nand R2278_U52 R2278_U335 ; R2278_U219
g5844 not R2278_U152 ; R2278_U220
g5845 or U2775 INSTADDRPOINTER_REG_12__SCAN_IN ; R2278_U221
g5846 not R2278_U29 ; R2278_U222
g5847 nand R2278_U55 R2278_U338 ; R2278_U223
g5848 not R2278_U140 ; R2278_U224
g5849 or U2771 INSTADDRPOINTER_REG_16__SCAN_IN ; R2278_U225
g5850 not R2278_U24 ; R2278_U226
g5851 or U2770 INSTADDRPOINTER_REG_17__SCAN_IN ; R2278_U227
g5852 nand U2770 INSTADDRPOINTER_REG_17__SCAN_IN ; R2278_U228
g5853 nand U2770 INSTADDRPOINTER_REG_18__SCAN_IN ; R2278_U229
g5854 not R2278_U23 ; R2278_U230
g5855 or U2770 INSTADDRPOINTER_REG_20__SCAN_IN ; R2278_U231
g5856 nand U2770 INSTADDRPOINTER_REG_20__SCAN_IN ; R2278_U232
g5857 nand R2278_U231 R2278_U128 ; R2278_U233
g5858 not R2278_U124 ; R2278_U234
g5859 or U2770 INSTADDRPOINTER_REG_21__SCAN_IN ; R2278_U235
g5860 nand U2770 INSTADDRPOINTER_REG_21__SCAN_IN ; R2278_U236
g5861 not R2278_U121 ; R2278_U237
g5862 nand U2770 INSTADDRPOINTER_REG_22__SCAN_IN ; R2278_U238
g5863 not R2278_U118 ; R2278_U239
g5864 nand U2770 INSTADDRPOINTER_REG_23__SCAN_IN ; R2278_U240
g5865 not R2278_U115 ; R2278_U241
g5866 or U2770 INSTADDRPOINTER_REG_24__SCAN_IN ; R2278_U242
g5867 nand U2770 INSTADDRPOINTER_REG_24__SCAN_IN ; R2278_U243
g5868 not R2278_U112 ; R2278_U244
g5869 nand U2770 INSTADDRPOINTER_REG_25__SCAN_IN ; R2278_U245
g5870 or U2770 INSTADDRPOINTER_REG_26__SCAN_IN ; R2278_U246
g5871 not R2278_U36 ; R2278_U247
g5872 nand R2278_U246 R2278_U110 ; R2278_U248
g5873 not R2278_U106 ; R2278_U249
g5874 or U2770 INSTADDRPOINTER_REG_27__SCAN_IN ; R2278_U250
g5875 nand U2770 INSTADDRPOINTER_REG_27__SCAN_IN ; R2278_U251
g5876 not R2278_U104 ; R2278_U252
g5877 or U2770 INSTADDRPOINTER_REG_28__SCAN_IN ; R2278_U253
g5878 nand U2770 INSTADDRPOINTER_REG_28__SCAN_IN ; R2278_U254
g5879 not R2278_U102 ; R2278_U255
g5880 or U2770 INSTADDRPOINTER_REG_29__SCAN_IN ; R2278_U256
g5881 nand U2770 INSTADDRPOINTER_REG_29__SCAN_IN ; R2278_U257
g5882 not R2278_U97 ; R2278_U258
g5883 or U2770 INSTADDRPOINTER_REG_30__SCAN_IN ; R2278_U259
g5884 nand U2770 INSTADDRPOINTER_REG_30__SCAN_IN ; R2278_U260
g5885 not R2278_U95 ; R2278_U261
g5886 not R2278_U100 ; R2278_U262
g5887 not R2278_U107 ; R2278_U263
g5888 not R2278_U109 ; R2278_U264
g5889 not R2278_U113 ; R2278_U265
g5890 not R2278_U116 ; R2278_U266
g5891 not R2278_U119 ; R2278_U267
g5892 not R2278_U122 ; R2278_U268
g5893 not R2278_U125 ; R2278_U269
g5894 not R2278_U127 ; R2278_U270
g5895 not R2278_U130 ; R2278_U271
g5896 not R2278_U131 ; R2278_U272
g5897 not R2278_U134 ; R2278_U273
g5898 not R2278_U137 ; R2278_U274
g5899 not R2278_U141 ; R2278_U275
g5900 nand R2278_U221 R2278_U152 ; R2278_U276
g5901 not R2278_U149 ; R2278_U277
g5902 nand R2278_U149 R2278_U213 ; R2278_U278
g5903 not R2278_U146 ; R2278_U279
g5904 nand R2278_U146 R2278_U211 ; R2278_U280
g5905 not R2278_U143 ; R2278_U281
g5906 not R2278_U144 ; R2278_U282
g5907 not R2278_U147 ; R2278_U283
g5908 not R2278_U150 ; R2278_U284
g5909 not R2278_U153 ; R2278_U285
g5910 nand R2278_U189 R2278_U72 ; R2278_U286
g5911 not R2278_U158 ; R2278_U287
g5912 nand R2278_U158 R2278_U217 ; R2278_U288
g5913 not R2278_U155 ; R2278_U289
g5914 not R2278_U156 ; R2278_U290
g5915 not R2278_U159 ; R2278_U291
g5916 or U2787 INSTADDRPOINTER_REG_0__SCAN_IN ; R2278_U292
g5917 nand R2278_U53 R2278_U5 ; R2278_U293
g5918 nand R2278_U222 R2278_U213 R2278_U211 R2278_U209 ; R2278_U294
g5919 nand R2278_U190 R2278_U5 ; R2278_U295
g5920 nand R2278_U218 R2278_U5 ; R2278_U296
g5921 nand R2278_U212 R2278_U209 ; R2278_U297
g5922 nand R2278_U211 R2278_U214 R2278_U209 ; R2278_U298
g5923 or U2785 INSTADDRPOINTER_REG_2__SCAN_IN ; R2278_U299
g5924 nand R2278_U172 R2278_U173 ; R2278_U300
g5925 nand R2278_U162 U2781 INSTADDRPOINTER_REG_6__SCAN_IN ; R2278_U301
g5926 nand R2278_U180 R2278_U162 R2278_U164 ; R2278_U302
g5927 or U2781 INSTADDRPOINTER_REG_6__SCAN_IN ; R2278_U303
g5928 nand R2278_U226 R2278_U227 ; R2278_U304
g5929 not R2278_U41 ; R2278_U305
g5930 nand R2278_U41 R2278_U208 ; R2278_U306
g5931 not R2278_U40 ; R2278_U307
g5932 not R2278_U25 ; R2278_U308
g5933 nand R2278_U9 R2278_U128 ; R2278_U309
g5934 nand R2278_U47 R2278_U235 ; R2278_U310
g5935 nand R2278_U10 R2278_U128 ; R2278_U311
g5936 nand R2278_U334 R2278_U206 ; R2278_U312
g5937 nand R2278_U11 R2278_U128 ; R2278_U313
g5938 nand R2278_U312 R2278_U238 ; R2278_U314
g5939 nand R2278_U314 R2278_U205 ; R2278_U315
g5940 nand R2278_U12 R2278_U128 ; R2278_U316
g5941 nand R2278_U315 R2278_U240 ; R2278_U317
g5942 nand R2278_U317 R2278_U242 ; R2278_U318
g5943 nand R2278_U318 R2278_U243 ; R2278_U319
g5944 nand R2278_U319 R2278_U204 ; R2278_U320
g5945 nand R2278_U14 R2278_U110 ; R2278_U321
g5946 nand R2278_U247 R2278_U250 ; R2278_U322
g5947 not R2278_U39 ; R2278_U323
g5948 nand R2278_U15 R2278_U110 ; R2278_U324
g5949 nand R2278_U39 R2278_U253 ; R2278_U325
g5950 not R2278_U38 ; R2278_U326
g5951 nand R2278_U16 R2278_U110 ; R2278_U327
g5952 nand R2278_U38 R2278_U256 ; R2278_U328
g5953 not R2278_U37 ; R2278_U329
g5954 nand R2278_U60 R2278_U110 ; R2278_U330
g5955 nand R2278_U37 R2278_U259 ; R2278_U331
g5956 nand R2278_U230 R2278_U13 ; R2278_U332
g5957 nand R2278_U308 R2278_U13 ; R2278_U333
g5958 nand R2278_U310 R2278_U236 ; R2278_U334
g5959 nand R2278_U336 R2278_U302 R2278_U50 ; R2278_U335
g5960 nand R2278_U48 R2278_U87 R2278_U49 ; R2278_U336
g5961 or U2781 INSTADDRPOINTER_REG_6__SCAN_IN ; R2278_U337
g5962 nand R2278_U219 R2278_U54 ; R2278_U338
g5963 nand R2278_U225 R2278_U140 ; R2278_U339
g5964 not R2278_U138 ; R2278_U340
g5965 nand R2278_U6 R2278_U140 ; R2278_U341
g5966 not R2278_U135 ; R2278_U342
g5967 nand R2278_U7 R2278_U140 ; R2278_U343
g5968 not R2278_U132 ; R2278_U344
g5969 nand R2278_U8 R2278_U140 ; R2278_U345
g5970 not R2278_U128 ; R2278_U346
g5971 nand R2278_U57 R2278_U140 ; R2278_U347
g5972 not R2278_U110 ; R2278_U348
g5973 nand R2278_U188 R2278_U73 ; R2278_U349
g5974 nand R2278_U191 R2278_U72 ; R2278_U350
g5975 nand R2278_U184 R2278_U76 ; R2278_U351
g5976 nand R2278_U192 R2278_U75 ; R2278_U352
g5977 nand R2278_U198 R2278_U79 ; R2278_U353
g5978 nand R2278_U199 R2278_U78 ; R2278_U354
g5979 nand R2278_U196 R2278_U82 ; R2278_U355
g5980 nand R2278_U200 R2278_U81 ; R2278_U356
g5981 nand R2278_U194 R2278_U85 ; R2278_U357
g5982 nand R2278_U201 R2278_U84 ; R2278_U358
g5983 nand R2278_U177 R2278_U88 ; R2278_U359
g5984 nand R2278_U202 R2278_U87 ; R2278_U360
g5985 nand R2278_U174 R2278_U91 ; R2278_U361
g5986 nand R2278_U203 R2278_U90 ; R2278_U362
g5987 nand U2769 R2278_U94 ; R2278_U363
g5988 nand R2278_U93 INSTADDRPOINTER_REG_31__SCAN_IN ; R2278_U364
g5989 not R2278_U62 ; R2278_U365
g5990 nand R2278_U261 R2278_U365 ; R2278_U366
g5991 nand R2278_U62 R2278_U95 ; R2278_U367
g5992 nand U2770 R2278_U21 ; R2278_U368
g5993 nand R2278_U22 INSTADDRPOINTER_REG_30__SCAN_IN ; R2278_U369
g5994 not R2278_U63 ; R2278_U370
g5995 nand R2278_U258 R2278_U370 ; R2278_U371
g5996 nand R2278_U63 R2278_U97 ; R2278_U372
g5997 nand R2278_U171 R2278_U100 ; R2278_U373
g5998 nand R2278_U262 R2278_U99 ; R2278_U374
g5999 nand U2770 R2278_U32 ; R2278_U375
g6000 nand R2278_U33 INSTADDRPOINTER_REG_29__SCAN_IN ; R2278_U376
g6001 not R2278_U64 ; R2278_U377
g6002 nand R2278_U255 R2278_U377 ; R2278_U378
g6003 nand R2278_U64 R2278_U102 ; R2278_U379
g6004 nand U2770 R2278_U34 ; R2278_U380
g6005 nand R2278_U35 INSTADDRPOINTER_REG_28__SCAN_IN ; R2278_U381
g6006 not R2278_U65 ; R2278_U382
g6007 nand R2278_U252 R2278_U382 ; R2278_U383
g6008 nand R2278_U65 R2278_U104 ; R2278_U384
g6009 nand R2278_U249 R2278_U107 ; R2278_U385
g6010 nand R2278_U263 R2278_U106 ; R2278_U386
g6011 nand R2278_U264 R2278_U110 ; R2278_U387
g6012 nand R2278_U348 R2278_U109 ; R2278_U388
g6013 nand R2278_U244 R2278_U113 ; R2278_U389
g6014 nand R2278_U265 R2278_U112 ; R2278_U390
g6015 nand R2278_U241 R2278_U116 ; R2278_U391
g6016 nand R2278_U266 R2278_U115 ; R2278_U392
g6017 nand R2278_U239 R2278_U119 ; R2278_U393
g6018 nand R2278_U267 R2278_U118 ; R2278_U394
g6019 nand R2278_U237 R2278_U122 ; R2278_U395
g6020 nand R2278_U268 R2278_U121 ; R2278_U396
g6021 nand R2278_U234 R2278_U125 ; R2278_U397
g6022 nand R2278_U269 R2278_U124 ; R2278_U398
g6023 nand R2278_U270 R2278_U128 ; R2278_U399
g6024 nand R2278_U346 R2278_U127 ; R2278_U400
g6025 nand R2278_U161 R2278_U130 ; R2278_U401
g6026 nand R2278_U271 R2278_U19 ; R2278_U402
g6027 nand R2278_U272 R2278_U132 ; R2278_U403
g6028 nand R2278_U344 R2278_U131 ; R2278_U404
g6029 nand R2278_U273 R2278_U135 ; R2278_U405
g6030 nand R2278_U342 R2278_U134 ; R2278_U406
g6031 nand R2278_U274 R2278_U138 ; R2278_U407
g6032 nand R2278_U340 R2278_U137 ; R2278_U408
g6033 nand R2278_U224 R2278_U141 ; R2278_U409
g6034 nand R2278_U275 R2278_U140 ; R2278_U410
g6035 nand R2278_U281 R2278_U144 ; R2278_U411
g6036 nand R2278_U282 R2278_U143 ; R2278_U412
g6037 nand R2278_U279 R2278_U147 ; R2278_U413
g6038 nand R2278_U283 R2278_U146 ; R2278_U414
g6039 nand R2278_U277 R2278_U150 ; R2278_U415
g6040 nand R2278_U284 R2278_U149 ; R2278_U416
g6041 nand R2278_U220 R2278_U153 ; R2278_U417
g6042 nand R2278_U285 R2278_U152 ; R2278_U418
g6043 nand R2278_U289 R2278_U156 ; R2278_U419
g6044 nand R2278_U290 R2278_U155 ; R2278_U420
g6045 nand R2278_U287 R2278_U159 ; R2278_U421
g6046 nand R2278_U291 R2278_U158 ; R2278_U422
g6047 and R2358_U293 R2358_U285 R2358_U282 R2358_U281 ; R2358_U5
g6048 and R2358_U329 R2358_U325 ; R2358_U6
g6049 and R2358_U6 R2358_U324 R2358_U141 ; R2358_U7
g6050 and R2358_U135 R2358_U5 ; R2358_U8
g6051 and R2358_U296 R2358_U294 ; R2358_U9
g6052 and R2358_U304 R2358_U253 ; R2358_U10
g6053 and R2358_U303 R2358_U301 ; R2358_U11
g6054 and R2358_U8 R2358_U7 ; R2358_U12
g6055 and R2358_U528 R2358_U527 ; R2358_U13
g6056 and R2358_U379 R2358_U378 ; R2358_U14
g6057 and R2358_U376 R2358_U374 ; R2358_U15
g6058 and R2358_U370 R2358_U367 ; R2358_U16
g6059 and R2358_U360 R2358_U359 ; R2358_U17
g6060 and R2358_U354 R2358_U352 ; R2358_U18
g6061 and R2358_U336 R2358_U335 ; R2358_U19
g6062 and R2358_U276 R2358_U274 ; R2358_U20
g6063 and R2358_U266 R2358_U262 ; R2358_U21
g6064 not U2352 ; R2358_U22
g6065 not U2643 ; R2358_U23
g6066 not U2644 ; R2358_U24
g6067 not U2645 ; R2358_U25
g6068 not U2646 ; R2358_U26
g6069 not U2649 ; R2358_U27
g6070 not U2648 ; R2358_U28
g6071 not U2650 ; R2358_U29
g6072 not U2647 ; R2358_U30
g6073 nand U2644 R2358_U77 ; R2358_U31
g6074 not U2642 ; R2358_U32
g6075 not U2641 ; R2358_U33
g6076 nand R2358_U246 R2358_U259 ; R2358_U34
g6077 not U2620 ; R2358_U35
g6078 not U2625 ; R2358_U36
g6079 not U2624 ; R2358_U37
g6080 not U2622 ; R2358_U38
g6081 not U2623 ; R2358_U39
g6082 not U2621 ; R2358_U40
g6083 not U2626 ; R2358_U41
g6084 not U2627 ; R2358_U42
g6085 not U2628 ; R2358_U43
g6086 not U2629 ; R2358_U44
g6087 not U2630 ; R2358_U45
g6088 nand U2630 R2358_U78 ; R2358_U46
g6089 not U2639 ; R2358_U47
g6090 not U2640 ; R2358_U48
g6091 nand U2642 R2358_U490 ; R2358_U49
g6092 not U2637 ; R2358_U50
g6093 nand U2637 R2358_U80 ; R2358_U51
g6094 not U2638 ; R2358_U52
g6095 nand U2638 R2358_U531 ; R2358_U53
g6096 not U2636 ; R2358_U54
g6097 nand R2358_U142 R2358_U9 ; R2358_U55
g6098 not U2631 ; R2358_U56
g6099 not U2632 ; R2358_U57
g6100 not U2633 ; R2358_U58
g6101 nand U2633 R2358_U607 ; R2358_U59
g6102 not U2634 ; R2358_U60
g6103 nand U2634 R2358_U601 ; R2358_U61
g6104 nand R2358_U438 R2358_U320 ; R2358_U62
g6105 nand R2358_U280 R2358_U291 ; R2358_U63
g6106 nand R2358_U233 R2358_U270 ; R2358_U64
g6107 nand R2358_U64 R2358_U229 ; R2358_U65
g6108 nand R2358_U417 R2358_U316 ; R2358_U66
g6109 nand R2358_U410 R2358_U219 R2358_U146 ; R2358_U67
g6110 nand R2358_U418 R2358_U416 ; R2358_U68
g6111 nand R2358_U407 R2358_U295 R2358_U408 ; R2358_U69
g6112 nand R2358_U313 R2358_U67 ; R2358_U70
g6113 not U2635 ; R2358_U71
g6114 nand R2358_U51 R2358_U364 ; R2358_U72
g6115 nand R2358_U414 R2358_U305 ; R2358_U73
g6116 nand R2358_U423 R2358_U413 ; R2358_U74
g6117 nand R2358_U74 R2358_U301 ; R2358_U75
g6118 nand R2358_U441 R2358_U440 ; R2358_U76
g6119 nand R2358_U454 R2358_U453 ; R2358_U77
g6120 nand R2358_U552 R2358_U551 ; R2358_U78
g6121 nand R2358_U520 R2358_U519 ; R2358_U79
g6122 nand R2358_U525 R2358_U524 ; R2358_U80
g6123 nand R2358_U533 R2358_U532 ; R2358_U81
g6124 nand R2358_U654 R2358_U653 ; R2358_U82
g6125 nand R2358_U492 R2358_U491 ; R2358_U83
g6126 and R2358_U49 R2358_U253 ; R2358_U84
g6127 nand R2358_U494 R2358_U493 ; R2358_U85
g6128 nand R2358_U499 R2358_U498 ; R2358_U86
g6129 and R2358_U246 R2358_U243 ; R2358_U87
g6130 nand R2358_U501 R2358_U500 ; R2358_U88
g6131 and R2358_U247 R2358_U244 ; R2358_U89
g6132 nand R2358_U503 R2358_U502 ; R2358_U90
g6133 nand R2358_U609 R2358_U608 ; R2358_U91
g6134 and R2358_U278 R2358_U277 ; R2358_U92
g6135 nand R2358_U611 R2358_U610 ; R2358_U93
g6136 and R2358_U280 R2358_U279 ; R2358_U94
g6137 nand R2358_U613 R2358_U612 ; R2358_U95
g6138 and R2358_U288 R2358_U281 ; R2358_U96
g6139 nand R2358_U615 R2358_U614 ; R2358_U97
g6140 and R2358_U289 R2358_U282 ; R2358_U98
g6141 nand R2358_U617 R2358_U616 ; R2358_U99
g6142 and R2358_U285 R2358_U284 ; R2358_U100
g6143 nand R2358_U619 R2358_U618 ; R2358_U101
g6144 and R2358_U293 R2358_U283 ; R2358_U102
g6145 nand R2358_U621 R2358_U620 ; R2358_U103
g6146 and R2358_U320 R2358_U319 ; R2358_U104
g6147 nand R2358_U623 R2358_U622 ; R2358_U105
g6148 and R2358_U322 R2358_U321 ; R2358_U106
g6149 nand R2358_U625 R2358_U624 ; R2358_U107
g6150 and R2358_U324 R2358_U323 ; R2358_U108
g6151 nand R2358_U627 R2358_U626 ; R2358_U109
g6152 nand R2358_U632 R2358_U631 ; R2358_U110
g6153 and R2358_U233 R2358_U232 ; R2358_U111
g6154 nand R2358_U634 R2358_U633 ; R2358_U112
g6155 and R2358_U317 R2358_U316 ; R2358_U113
g6156 nand R2358_U636 R2358_U635 ; R2358_U114
g6157 and R2358_U295 R2358_U294 ; R2358_U115
g6158 nand R2358_U638 R2358_U637 ; R2358_U116
g6159 and R2358_U59 R2358_U296 ; R2358_U117
g6160 nand R2358_U640 R2358_U639 ; R2358_U118
g6161 nand R2358_U645 R2358_U644 ; R2358_U119
g6162 nand R2358_U650 R2358_U649 ; R2358_U120
g6163 and R2358_U310 R2358_U53 ; R2358_U121
g6164 nand R2358_U652 R2358_U651 ; R2358_U122
g6165 and R2358_U235 R2358_U232 ; R2358_U123
g6166 and R2358_U231 R2358_U229 ; R2358_U124
g6167 and R2358_U244 R2358_U243 ; R2358_U125
g6168 and R2358_U249 R2358_U245 ; R2358_U126
g6169 and R2358_U245 R2358_U222 ; R2358_U127
g6170 and R2358_U265 R2358_U31 ; R2358_U128
g6171 and R2358_U231 R2358_U230 ; R2358_U129
g6172 and R2358_U285 R2358_U282 ; R2358_U130
g6173 and R2358_U288 R2358_U289 ; R2358_U131
g6174 and R2358_U281 R2358_U279 ; R2358_U132
g6175 and R2358_U326 R2358_U323 ; R2358_U133
g6176 and R2358_U322 R2358_U319 ; R2358_U134
g6177 and R2358_U279 R2358_U277 ; R2358_U135
g6178 and R2358_U11 R2358_U10 ; R2358_U136
g6179 and R2358_U432 R2358_U425 ; R2358_U137
g6180 and R2358_U310 R2358_U224 ; R2358_U138
g6181 and R2358_U415 R2358_U311 ; R2358_U139
g6182 and R2358_U420 R2358_U411 ; R2358_U140
g6183 and R2358_U322 R2358_U319 ; R2358_U141
g6184 and R2358_U317 R2358_U313 ; R2358_U142
g6185 and R2358_U12 R2358_U426 ; R2358_U143
g6186 and R2358_U402 R2358_U278 ; R2358_U144
g6187 and R2358_U144 R2358_U406 R2358_U430 ; R2358_U145
g6188 and R2358_U420 R2358_U411 ; R2358_U146
g6189 and R2358_U313 R2358_U317 ; R2358_U147
g6190 and R2358_U7 R2358_U149 ; R2358_U148
g6191 and R2358_U9 R2358_U147 ; R2358_U149
g6192 and R2358_U422 R2358_U439 ; R2358_U150
g6193 and R2358_U5 R2358_U279 ; R2358_U151
g6194 and R2358_U285 R2358_U282 R2358_U293 ; R2358_U152
g6195 and R2358_U289 R2358_U287 ; R2358_U153
g6196 and R2358_U284 R2358_U283 ; R2358_U154
g6197 and R2358_U156 R2358_U434 ; R2358_U155
g6198 and R2358_U6 R2358_U324 ; R2358_U156
g6199 and R2358_U418 R2358_U46 ; R2358_U157
g6200 and R2358_U6 R2358_U326 ; R2358_U158
g6201 and R2358_U313 R2358_U9 ; R2358_U159
g6202 and R2358_U299 R2358_U224 R2358_U300 ; R2358_U160
g6203 and R2358_U369 R2358_U227 ; R2358_U161
g6204 and R2358_U303 R2358_U302 ; R2358_U162
g6205 and R2358_U375 R2358_U307 ; R2358_U163
g6206 not U2612 ; R2358_U164
g6207 and R2358_U444 R2358_U443 ; R2358_U165
g6208 not U2610 ; R2358_U166
g6209 not U2609 ; R2358_U167
g6210 not U2667 ; R2358_U168
g6211 not U2668 ; R2358_U169
g6212 not U2670 ; R2358_U170
g6213 not U2671 ; R2358_U171
g6214 not U2672 ; R2358_U172
g6215 not U2669 ; R2358_U173
g6216 not U2611 ; R2358_U174
g6217 nand R2358_U49 R2358_U255 ; R2358_U175
g6218 nand R2358_U251 R2358_U250 R2358_U126 ; R2358_U176
g6219 nand R2358_U247 R2358_U257 ; R2358_U177
g6220 nand R2358_U230 R2358_U240 ; R2358_U178
g6221 not U2651 ; R2358_U179
g6222 and R2358_U505 R2358_U504 ; R2358_U180
g6223 not U2613 ; R2358_U181
g6224 not U2614 ; R2358_U182
g6225 not U2617 ; R2358_U183
g6226 not U2615 ; R2358_U184
g6227 not U2616 ; R2358_U185
g6228 not U2618 ; R2358_U186
g6229 not U2664 ; R2358_U187
g6230 not U2665 ; R2358_U188
g6231 not U2666 ; R2358_U189
g6232 not U2663 ; R2358_U190
g6233 not U2658 ; R2358_U191
g6234 not U2659 ; R2358_U192
g6235 not U2660 ; R2358_U193
g6236 not U2661 ; R2358_U194
g6237 not U2662 ; R2358_U195
g6238 not U2654 ; R2358_U196
g6239 not U2655 ; R2358_U197
g6240 not U2656 ; R2358_U198
g6241 not U2657 ; R2358_U199
g6242 not U2652 ; R2358_U200
g6243 not U2653 ; R2358_U201
g6244 nand R2358_U145 R2358_U429 ; R2358_U202
g6245 nand R2358_U292 R2358_U332 ; R2358_U203
g6246 nand R2358_U338 R2358_U337 ; R2358_U204
g6247 nand R2358_U153 R2358_U340 ; R2358_U205
g6248 nand R2358_U344 R2358_U285 ; R2358_U206
g6249 nand R2358_U283 R2358_U342 ; R2358_U207
g6250 nand R2358_U150 R2358_U421 ; R2358_U208
g6251 nand R2358_U321 R2358_U347 ; R2358_U209
g6252 nand R2358_U345 R2358_U437 ; R2358_U210
g6253 nand R2358_U350 R2358_U325 ; R2358_U211
g6254 nand R2358_U236 R2358_U268 ; R2358_U212
g6255 nand R2358_U412 R2358_U409 ; R2358_U213
g6256 nand R2358_U356 R2358_U59 ; R2358_U214
g6257 nand R2358_U61 R2358_U70 ; R2358_U215
g6258 nand R2358_U53 R2358_U361 ; R2358_U216
g6259 nand R2358_U137 R2358_U431 ; R2358_U217
g6260 nand R2358_U236 R2358_U235 ; R2358_U218
g6261 nand R2358_U138 R2358_U217 R2358_U139 ; R2358_U219
g6262 not R2358_U211 ; R2358_U220
g6263 not R2358_U206 ; R2358_U221
g6264 nand R2358_U404 R2358_U403 ; R2358_U222
g6265 not R2358_U51 ; R2358_U223
g6266 nand R2358_U521 R2358_U54 ; R2358_U224
g6267 not R2358_U46 ; R2358_U225
g6268 nand R2358_U349 R2358_U329 ; R2358_U226
g6269 nand U2636 R2358_U79 ; R2358_U227
g6270 not R2358_U31 ; R2358_U228
g6271 nand R2358_U480 R2358_U479 R2358_U28 ; R2358_U229
g6272 nand U2647 R2358_U485 ; R2358_U230
g6273 nand R2358_U482 R2358_U481 R2358_U30 ; R2358_U231
g6274 nand R2358_U476 R2358_U475 R2358_U27 ; R2358_U232
g6275 nand U2649 R2358_U471 ; R2358_U233
g6276 nand U2648 R2358_U468 ; R2358_U234
g6277 nand R2358_U478 R2358_U477 R2358_U29 ; R2358_U235
g6278 nand U2650 R2358_U474 ; R2358_U236
g6279 nand R2358_U236 R2358_U22 ; R2358_U237
g6280 nand R2358_U123 R2358_U237 ; R2358_U238
g6281 nand R2358_U238 R2358_U233 R2358_U234 ; R2358_U239
g6282 nand R2358_U124 R2358_U239 ; R2358_U240
g6283 not R2358_U178 ; R2358_U241
g6284 nand R2358_U452 R2358_U451 R2358_U23 ; R2358_U242
g6285 nand R2358_U463 R2358_U462 R2358_U25 ; R2358_U243
g6286 nand R2358_U465 R2358_U464 R2358_U26 ; R2358_U244
g6287 nand U2643 R2358_U450 ; R2358_U245
g6288 nand U2645 R2358_U458 ; R2358_U246
g6289 nand U2646 R2358_U461 ; R2358_U247
g6290 nand R2358_U247 R2358_U246 ; R2358_U248
g6291 nand R2358_U243 R2358_U248 R2358_U222 ; R2358_U249
g6292 nand R2358_U178 R2358_U125 R2358_U222 ; R2358_U250
g6293 nand R2358_U228 R2358_U242 ; R2358_U251
g6294 not R2358_U176 ; R2358_U252
g6295 nand R2358_U487 R2358_U486 R2358_U32 ; R2358_U253
g6296 not R2358_U49 ; R2358_U254
g6297 nand R2358_U253 R2358_U176 ; R2358_U255
g6298 not R2358_U175 ; R2358_U256
g6299 nand R2358_U244 R2358_U178 ; R2358_U257
g6300 not R2358_U177 ; R2358_U258
g6301 nand R2358_U177 R2358_U243 ; R2358_U259
g6302 not R2358_U34 ; R2358_U260
g6303 nand R2358_U260 R2358_U31 ; R2358_U261
g6304 nand R2358_U127 R2358_U261 ; R2358_U262
g6305 nand R2358_U455 R2358_U24 ; R2358_U263
g6306 nand R2358_U263 R2358_U34 ; R2358_U264
g6307 nand R2358_U245 R2358_U242 ; R2358_U265
g6308 nand R2358_U128 R2358_U264 ; R2358_U266
g6309 nand R2358_U455 R2358_U24 ; R2358_U267
g6310 nand U2352 R2358_U235 ; R2358_U268
g6311 not R2358_U212 ; R2358_U269
g6312 nand R2358_U212 R2358_U232 ; R2358_U270
g6313 not R2358_U64 ; R2358_U271
g6314 not R2358_U65 ; R2358_U272
g6315 nand R2358_U65 R2358_U234 ; R2358_U273
g6316 nand R2358_U129 R2358_U273 ; R2358_U274
g6317 nand R2358_U231 R2358_U230 ; R2358_U275
g6318 nand R2358_U65 R2358_U234 R2358_U275 ; R2358_U276
g6319 nand R2358_U563 R2358_U562 R2358_U35 ; R2358_U277
g6320 nand U2620 R2358_U580 ; R2358_U278
g6321 nand R2358_U565 R2358_U564 R2358_U40 ; R2358_U279
g6322 nand U2621 R2358_U595 ; R2358_U280
g6323 nand R2358_U555 R2358_U554 R2358_U38 ; R2358_U281
g6324 nand R2358_U557 R2358_U556 R2358_U39 ; R2358_U282
g6325 nand U2625 R2358_U583 ; R2358_U283
g6326 nand U2624 R2358_U586 ; R2358_U284
g6327 nand R2358_U559 R2358_U558 R2358_U37 ; R2358_U285
g6328 nand R2358_U284 R2358_U283 ; R2358_U286
g6329 nand R2358_U130 R2358_U286 ; R2358_U287
g6330 nand U2622 R2358_U592 ; R2358_U288
g6331 nand U2623 R2358_U589 ; R2358_U289
g6332 nand R2358_U131 R2358_U287 ; R2358_U290
g6333 nand R2358_U132 R2358_U290 ; R2358_U291
g6334 not R2358_U63 ; R2358_U292
g6335 nand R2358_U561 R2358_U560 R2358_U36 ; R2358_U293
g6336 nand R2358_U536 R2358_U535 R2358_U57 ; R2358_U294
g6337 nand U2632 R2358_U604 ; R2358_U295
g6338 nand R2358_U538 R2358_U537 R2358_U58 ; R2358_U296
g6339 not R2358_U59 ; R2358_U297
g6340 not R2358_U61 ; R2358_U298
g6341 nand R2358_U13 R2358_U71 ; R2358_U299
g6342 nand U2635 R2358_U81 ; R2358_U300
g6343 nand R2358_U510 R2358_U509 R2358_U48 ; R2358_U301
g6344 nand U2639 R2358_U515 ; R2358_U302
g6345 nand R2358_U512 R2358_U511 R2358_U47 ; R2358_U303
g6346 nand R2358_U442 R2358_U33 ; R2358_U304
g6347 nand U2641 R2358_U76 ; R2358_U305
g6348 not R2358_U74 ; R2358_U306
g6349 nand U2640 R2358_U518 ; R2358_U307
g6350 not R2358_U217 ; R2358_U308
g6351 not R2358_U53 ; R2358_U309
g6352 nand R2358_U523 R2358_U522 R2358_U52 ; R2358_U310
g6353 nand R2358_U526 R2358_U50 ; R2358_U311
g6354 not R2358_U67 ; R2358_U312
g6355 nand R2358_U540 R2358_U539 R2358_U60 ; R2358_U313
g6356 not R2358_U70 ; R2358_U314
g6357 not R2358_U213 ; R2358_U315
g6358 nand U2631 R2358_U598 ; R2358_U316
g6359 nand R2358_U542 R2358_U541 R2358_U56 ; R2358_U317
g6360 not R2358_U68 ; R2358_U318
g6361 nand R2358_U544 R2358_U543 R2358_U41 ; R2358_U319
g6362 nand U2626 R2358_U568 ; R2358_U320
g6363 nand U2627 R2358_U571 ; R2358_U321
g6364 nand R2358_U546 R2358_U545 R2358_U42 ; R2358_U322
g6365 nand U2628 R2358_U574 ; R2358_U323
g6366 nand R2358_U548 R2358_U547 R2358_U43 ; R2358_U324
g6367 nand R2358_U550 R2358_U549 R2358_U44 ; R2358_U325
g6368 nand U2629 R2358_U577 ; R2358_U326
g6369 nand R2358_U225 R2358_U325 ; R2358_U327
g6370 nand R2358_U437 R2358_U321 ; R2358_U328
g6371 nand R2358_U553 R2358_U45 ; R2358_U329
g6372 not R2358_U202 ; R2358_U330
g6373 not R2358_U208 ; R2358_U331
g6374 nand R2358_U151 R2358_U208 ; R2358_U332
g6375 not R2358_U203 ; R2358_U333
g6376 nand R2358_U234 R2358_U229 ; R2358_U334
g6377 nand R2358_U271 R2358_U334 ; R2358_U335
g6378 nand R2358_U272 R2358_U234 ; R2358_U336
g6379 nand R2358_U290 R2358_U281 ; R2358_U337
g6380 nand R2358_U5 R2358_U208 ; R2358_U338
g6381 not R2358_U204 ; R2358_U339
g6382 nand R2358_U152 R2358_U208 ; R2358_U340
g6383 not R2358_U205 ; R2358_U341
g6384 nand R2358_U208 R2358_U293 ; R2358_U342
g6385 not R2358_U207 ; R2358_U343
g6386 nand R2358_U154 R2358_U342 ; R2358_U344
g6387 nand R2358_U433 R2358_U155 ; R2358_U345
g6388 not R2358_U210 ; R2358_U346
g6389 nand R2358_U210 R2358_U322 ; R2358_U347
g6390 not R2358_U209 ; R2358_U348
g6391 nand R2358_U157 R2358_U416 ; R2358_U349
g6392 nand R2358_U326 R2358_U226 ; R2358_U350
g6393 nand R2358_U318 R2358_U46 ; R2358_U351
g6394 nand R2358_U158 R2358_U351 ; R2358_U352
g6395 nand R2358_U326 R2358_U325 ; R2358_U353
g6396 nand R2358_U226 R2358_U353 ; R2358_U354
g6397 not R2358_U215 ; R2358_U355
g6398 nand R2358_U215 R2358_U296 ; R2358_U356
g6399 not R2358_U214 ; R2358_U357
g6400 nand R2358_U313 R2358_U61 ; R2358_U358
g6401 nand R2358_U312 R2358_U358 ; R2358_U359
g6402 nand R2358_U314 R2358_U61 ; R2358_U360
g6403 nand R2358_U310 R2358_U217 ; R2358_U361
g6404 not R2358_U216 ; R2358_U362
g6405 nand R2358_U526 R2358_U50 ; R2358_U363
g6406 nand R2358_U363 R2358_U216 ; R2358_U364
g6407 not R2358_U72 ; R2358_U365
g6408 nand R2358_U365 R2358_U227 ; R2358_U366
g6409 nand R2358_U160 R2358_U366 ; R2358_U367
g6410 nand R2358_U72 R2358_U224 ; R2358_U368
g6411 nand R2358_U300 R2358_U299 ; R2358_U369
g6412 nand R2358_U161 R2358_U368 ; R2358_U370
g6413 nand R2358_U526 R2358_U50 ; R2358_U371
g6414 not R2358_U75 ; R2358_U372
g6415 nand R2358_U75 R2358_U307 ; R2358_U373
g6416 nand R2358_U162 R2358_U373 ; R2358_U374
g6417 nand R2358_U303 R2358_U302 ; R2358_U375
g6418 nand R2358_U163 R2358_U75 ; R2358_U376
g6419 nand R2358_U307 R2358_U301 ; R2358_U377
g6420 nand R2358_U306 R2358_U377 ; R2358_U378
g6421 nand R2358_U372 R2358_U307 ; R2358_U379
g6422 not R2358_U218 ; R2358_U380
g6423 nand R2358_U49 R2358_U253 ; R2358_U381
g6424 nand R2358_U267 R2358_U31 ; R2358_U382
g6425 nand R2358_U246 R2358_U243 ; R2358_U383
g6426 nand R2358_U247 R2358_U244 ; R2358_U384
g6427 nand R2358_U278 R2358_U277 ; R2358_U385
g6428 nand R2358_U280 R2358_U279 ; R2358_U386
g6429 nand R2358_U288 R2358_U281 ; R2358_U387
g6430 nand R2358_U289 R2358_U282 ; R2358_U388
g6431 nand R2358_U285 R2358_U284 ; R2358_U389
g6432 nand R2358_U293 R2358_U283 ; R2358_U390
g6433 nand R2358_U320 R2358_U319 ; R2358_U391
g6434 nand R2358_U322 R2358_U321 ; R2358_U392
g6435 nand R2358_U324 R2358_U323 ; R2358_U393
g6436 nand R2358_U329 R2358_U46 ; R2358_U394
g6437 nand R2358_U233 R2358_U232 ; R2358_U395
g6438 nand R2358_U317 R2358_U316 ; R2358_U396
g6439 nand R2358_U295 R2358_U294 ; R2358_U397
g6440 nand R2358_U59 R2358_U296 ; R2358_U398
g6441 nand R2358_U227 R2358_U224 ; R2358_U399
g6442 nand R2358_U371 R2358_U51 ; R2358_U400
g6443 nand R2358_U310 R2358_U53 ; R2358_U401
g6444 nand R2358_U63 R2358_U277 ; R2358_U402
g6445 nand R2358_U77 R2358_U242 ; R2358_U403
g6446 nand U2644 R2358_U242 ; R2358_U404
g6447 nand U2640 R2358_U518 ; R2358_U405
g6448 nand R2358_U8 R2358_U62 ; R2358_U406
g6449 nand R2358_U297 R2358_U9 ; R2358_U407
g6450 nand R2358_U298 R2358_U9 ; R2358_U408
g6451 nand R2358_U159 R2358_U67 ; R2358_U409
g6452 nand R2358_U223 R2358_U224 R2358_U299 ; R2358_U410
g6453 nand R2358_U309 R2358_U311 R2358_U224 R2358_U299 ; R2358_U411
g6454 not R2358_U69 ; R2358_U412
g6455 nand R2358_U10 R2358_U176 ; R2358_U413
g6456 nand R2358_U254 R2358_U304 ; R2358_U414
g6457 nand R2358_U13 R2358_U71 ; R2358_U415
g6458 nand R2358_U426 R2358_U67 ; R2358_U416
g6459 nand R2358_U69 R2358_U317 ; R2358_U417
g6460 not R2358_U66 ; R2358_U418
g6461 nand R2358_U13 R2358_U71 ; R2358_U419
g6462 nand R2358_U427 R2358_U419 R2358_U428 ; R2358_U420
g6463 nand R2358_U67 R2358_U148 ; R2358_U421
g6464 nand R2358_U66 R2358_U7 ; R2358_U422
g6465 not R2358_U73 ; R2358_U423
g6466 nand R2358_U405 R2358_U302 ; R2358_U424
g6467 nand R2358_U424 R2358_U303 ; R2358_U425
g6468 not R2358_U55 ; R2358_U426
g6469 nand R2358_U227 R2358_U71 ; R2358_U427
g6470 nand R2358_U534 R2358_U227 ; R2358_U428
g6471 nand R2358_U143 R2358_U435 ; R2358_U429
g6472 nand R2358_U12 R2358_U66 ; R2358_U430
g6473 nand R2358_U136 R2358_U176 ; R2358_U431
g6474 nand R2358_U11 R2358_U73 ; R2358_U432
g6475 nand R2358_U312 R2358_U418 ; R2358_U433
g6476 nand R2358_U418 R2358_U55 ; R2358_U434
g6477 nand R2358_U410 R2358_U219 R2358_U140 ; R2358_U435
g6478 nand R2358_U133 R2358_U327 ; R2358_U436
g6479 nand R2358_U436 R2358_U324 ; R2358_U437
g6480 nand R2358_U134 R2358_U328 ; R2358_U438
g6481 not R2358_U62 ; R2358_U439
g6482 nand U2352 R2358_U164 ; R2358_U440
g6483 nand U2612 R2358_U22 ; R2358_U441
g6484 not R2358_U76 ; R2358_U442
g6485 nand R2358_U442 U2641 ; R2358_U443
g6486 nand R2358_U76 R2358_U33 ; R2358_U444
g6487 nand R2358_U442 U2641 ; R2358_U445
g6488 nand R2358_U76 R2358_U33 ; R2358_U446
g6489 nand R2358_U446 R2358_U445 ; R2358_U447
g6490 nand U2352 R2358_U166 ; R2358_U448
g6491 nand U2610 R2358_U22 ; R2358_U449
g6492 nand R2358_U449 R2358_U448 ; R2358_U450
g6493 nand U2352 R2358_U166 ; R2358_U451
g6494 nand U2610 R2358_U22 ; R2358_U452
g6495 nand U2352 R2358_U167 ; R2358_U453
g6496 nand U2609 R2358_U22 ; R2358_U454
g6497 not R2358_U77 ; R2358_U455
g6498 nand U2352 R2358_U168 ; R2358_U456
g6499 nand U2667 R2358_U22 ; R2358_U457
g6500 nand R2358_U457 R2358_U456 ; R2358_U458
g6501 nand U2352 R2358_U169 ; R2358_U459
g6502 nand U2668 R2358_U22 ; R2358_U460
g6503 nand R2358_U460 R2358_U459 ; R2358_U461
g6504 nand U2352 R2358_U168 ; R2358_U462
g6505 nand U2667 R2358_U22 ; R2358_U463
g6506 nand U2352 R2358_U169 ; R2358_U464
g6507 nand U2668 R2358_U22 ; R2358_U465
g6508 nand U2352 R2358_U170 ; R2358_U466
g6509 nand U2670 R2358_U22 ; R2358_U467
g6510 nand R2358_U467 R2358_U466 ; R2358_U468
g6511 nand U2352 R2358_U171 ; R2358_U469
g6512 nand U2671 R2358_U22 ; R2358_U470
g6513 nand R2358_U470 R2358_U469 ; R2358_U471
g6514 nand U2352 R2358_U172 ; R2358_U472
g6515 nand U2672 R2358_U22 ; R2358_U473
g6516 nand R2358_U473 R2358_U472 ; R2358_U474
g6517 nand U2352 R2358_U171 ; R2358_U475
g6518 nand U2671 R2358_U22 ; R2358_U476
g6519 nand U2352 R2358_U172 ; R2358_U477
g6520 nand U2672 R2358_U22 ; R2358_U478
g6521 nand U2352 R2358_U170 ; R2358_U479
g6522 nand U2670 R2358_U22 ; R2358_U480
g6523 nand U2352 R2358_U173 ; R2358_U481
g6524 nand U2669 R2358_U22 ; R2358_U482
g6525 nand U2352 R2358_U173 ; R2358_U483
g6526 nand U2669 R2358_U22 ; R2358_U484
g6527 nand R2358_U484 R2358_U483 ; R2358_U485
g6528 nand U2352 R2358_U174 ; R2358_U486
g6529 nand U2611 R2358_U22 ; R2358_U487
g6530 nand U2352 R2358_U174 ; R2358_U488
g6531 nand U2611 R2358_U22 ; R2358_U489
g6532 nand R2358_U489 R2358_U488 ; R2358_U490
g6533 nand R2358_U165 R2358_U175 ; R2358_U491
g6534 nand R2358_U256 R2358_U447 ; R2358_U492
g6535 nand R2358_U381 R2358_U176 ; R2358_U493
g6536 nand R2358_U84 R2358_U252 ; R2358_U494
g6537 nand R2358_U455 U2644 ; R2358_U495
g6538 nand R2358_U77 R2358_U24 ; R2358_U496
g6539 nand R2358_U496 R2358_U495 ; R2358_U497
g6540 nand R2358_U382 R2358_U34 ; R2358_U498
g6541 nand R2358_U497 R2358_U260 ; R2358_U499
g6542 nand R2358_U383 R2358_U177 ; R2358_U500
g6543 nand R2358_U87 R2358_U258 ; R2358_U501
g6544 nand R2358_U384 R2358_U178 ; R2358_U502
g6545 nand R2358_U89 R2358_U241 ; R2358_U503
g6546 nand U2352 R2358_U179 ; R2358_U504
g6547 nand U2651 R2358_U22 ; R2358_U505
g6548 nand U2352 R2358_U179 ; R2358_U506
g6549 nand U2651 R2358_U22 ; R2358_U507
g6550 nand R2358_U507 R2358_U506 ; R2358_U508
g6551 nand U2352 R2358_U181 ; R2358_U509
g6552 nand U2613 R2358_U22 ; R2358_U510
g6553 nand U2352 R2358_U182 ; R2358_U511
g6554 nand U2614 R2358_U22 ; R2358_U512
g6555 nand U2352 R2358_U182 ; R2358_U513
g6556 nand U2614 R2358_U22 ; R2358_U514
g6557 nand R2358_U514 R2358_U513 ; R2358_U515
g6558 nand U2352 R2358_U181 ; R2358_U516
g6559 nand U2613 R2358_U22 ; R2358_U517
g6560 nand R2358_U517 R2358_U516 ; R2358_U518
g6561 nand U2352 R2358_U183 ; R2358_U519
g6562 nand U2617 R2358_U22 ; R2358_U520
g6563 not R2358_U79 ; R2358_U521
g6564 nand U2352 R2358_U184 ; R2358_U522
g6565 nand U2615 R2358_U22 ; R2358_U523
g6566 nand U2352 R2358_U185 ; R2358_U524
g6567 nand U2616 R2358_U22 ; R2358_U525
g6568 not R2358_U80 ; R2358_U526
g6569 nand U2352 R2358_U186 ; R2358_U527
g6570 nand U2618 R2358_U22 ; R2358_U528
g6571 nand U2352 R2358_U184 ; R2358_U529
g6572 nand U2615 R2358_U22 ; R2358_U530
g6573 nand R2358_U530 R2358_U529 ; R2358_U531
g6574 nand U2352 R2358_U186 ; R2358_U532
g6575 nand U2618 R2358_U22 ; R2358_U533
g6576 not R2358_U81 ; R2358_U534
g6577 nand U2352 R2358_U187 ; R2358_U535
g6578 nand U2664 R2358_U22 ; R2358_U536
g6579 nand U2352 R2358_U188 ; R2358_U537
g6580 nand U2665 R2358_U22 ; R2358_U538
g6581 nand U2352 R2358_U189 ; R2358_U539
g6582 nand U2666 R2358_U22 ; R2358_U540
g6583 nand U2352 R2358_U190 ; R2358_U541
g6584 nand U2663 R2358_U22 ; R2358_U542
g6585 nand U2352 R2358_U191 ; R2358_U543
g6586 nand U2658 R2358_U22 ; R2358_U544
g6587 nand U2352 R2358_U192 ; R2358_U545
g6588 nand U2659 R2358_U22 ; R2358_U546
g6589 nand U2352 R2358_U193 ; R2358_U547
g6590 nand U2660 R2358_U22 ; R2358_U548
g6591 nand U2352 R2358_U194 ; R2358_U549
g6592 nand U2661 R2358_U22 ; R2358_U550
g6593 nand U2352 R2358_U195 ; R2358_U551
g6594 nand U2662 R2358_U22 ; R2358_U552
g6595 not R2358_U78 ; R2358_U553
g6596 nand U2352 R2358_U196 ; R2358_U554
g6597 nand U2654 R2358_U22 ; R2358_U555
g6598 nand U2352 R2358_U197 ; R2358_U556
g6599 nand U2655 R2358_U22 ; R2358_U557
g6600 nand U2352 R2358_U198 ; R2358_U558
g6601 nand U2656 R2358_U22 ; R2358_U559
g6602 nand U2352 R2358_U199 ; R2358_U560
g6603 nand U2657 R2358_U22 ; R2358_U561
g6604 nand U2352 R2358_U200 ; R2358_U562
g6605 nand U2652 R2358_U22 ; R2358_U563
g6606 nand U2352 R2358_U201 ; R2358_U564
g6607 nand U2653 R2358_U22 ; R2358_U565
g6608 nand U2352 R2358_U191 ; R2358_U566
g6609 nand U2658 R2358_U22 ; R2358_U567
g6610 nand R2358_U567 R2358_U566 ; R2358_U568
g6611 nand U2352 R2358_U192 ; R2358_U569
g6612 nand U2659 R2358_U22 ; R2358_U570
g6613 nand R2358_U570 R2358_U569 ; R2358_U571
g6614 nand U2352 R2358_U193 ; R2358_U572
g6615 nand U2660 R2358_U22 ; R2358_U573
g6616 nand R2358_U573 R2358_U572 ; R2358_U574
g6617 nand U2352 R2358_U194 ; R2358_U575
g6618 nand U2661 R2358_U22 ; R2358_U576
g6619 nand R2358_U576 R2358_U575 ; R2358_U577
g6620 nand U2352 R2358_U200 ; R2358_U578
g6621 nand U2652 R2358_U22 ; R2358_U579
g6622 nand R2358_U579 R2358_U578 ; R2358_U580
g6623 nand U2352 R2358_U199 ; R2358_U581
g6624 nand U2657 R2358_U22 ; R2358_U582
g6625 nand R2358_U582 R2358_U581 ; R2358_U583
g6626 nand U2352 R2358_U198 ; R2358_U584
g6627 nand U2656 R2358_U22 ; R2358_U585
g6628 nand R2358_U585 R2358_U584 ; R2358_U586
g6629 nand U2352 R2358_U197 ; R2358_U587
g6630 nand U2655 R2358_U22 ; R2358_U588
g6631 nand R2358_U588 R2358_U587 ; R2358_U589
g6632 nand U2352 R2358_U196 ; R2358_U590
g6633 nand U2654 R2358_U22 ; R2358_U591
g6634 nand R2358_U591 R2358_U590 ; R2358_U592
g6635 nand U2352 R2358_U201 ; R2358_U593
g6636 nand U2653 R2358_U22 ; R2358_U594
g6637 nand R2358_U594 R2358_U593 ; R2358_U595
g6638 nand U2352 R2358_U190 ; R2358_U596
g6639 nand U2663 R2358_U22 ; R2358_U597
g6640 nand R2358_U597 R2358_U596 ; R2358_U598
g6641 nand U2352 R2358_U189 ; R2358_U599
g6642 nand U2666 R2358_U22 ; R2358_U600
g6643 nand R2358_U600 R2358_U599 ; R2358_U601
g6644 nand U2352 R2358_U187 ; R2358_U602
g6645 nand U2664 R2358_U22 ; R2358_U603
g6646 nand R2358_U603 R2358_U602 ; R2358_U604
g6647 nand U2352 R2358_U188 ; R2358_U605
g6648 nand U2665 R2358_U22 ; R2358_U606
g6649 nand R2358_U606 R2358_U605 ; R2358_U607
g6650 nand R2358_U180 R2358_U202 ; R2358_U608
g6651 nand R2358_U330 R2358_U508 ; R2358_U609
g6652 nand R2358_U385 R2358_U203 ; R2358_U610
g6653 nand R2358_U92 R2358_U333 ; R2358_U611
g6654 nand R2358_U386 R2358_U204 ; R2358_U612
g6655 nand R2358_U94 R2358_U339 ; R2358_U613
g6656 nand R2358_U387 R2358_U205 ; R2358_U614
g6657 nand R2358_U96 R2358_U341 ; R2358_U615
g6658 nand R2358_U221 R2358_U388 ; R2358_U616
g6659 nand R2358_U98 R2358_U206 ; R2358_U617
g6660 nand R2358_U389 R2358_U207 ; R2358_U618
g6661 nand R2358_U100 R2358_U343 ; R2358_U619
g6662 nand R2358_U390 R2358_U208 ; R2358_U620
g6663 nand R2358_U102 R2358_U331 ; R2358_U621
g6664 nand R2358_U391 R2358_U209 ; R2358_U622
g6665 nand R2358_U104 R2358_U348 ; R2358_U623
g6666 nand R2358_U392 R2358_U210 ; R2358_U624
g6667 nand R2358_U106 R2358_U346 ; R2358_U625
g6668 nand R2358_U220 R2358_U393 ; R2358_U626
g6669 nand R2358_U108 R2358_U211 ; R2358_U627
g6670 nand R2358_U553 U2630 ; R2358_U628
g6671 nand R2358_U78 R2358_U45 ; R2358_U629
g6672 nand R2358_U629 R2358_U628 ; R2358_U630
g6673 nand R2358_U394 R2358_U68 ; R2358_U631
g6674 nand R2358_U630 R2358_U318 ; R2358_U632
g6675 nand R2358_U395 R2358_U212 ; R2358_U633
g6676 nand R2358_U111 R2358_U269 ; R2358_U634
g6677 nand R2358_U396 R2358_U213 ; R2358_U635
g6678 nand R2358_U113 R2358_U315 ; R2358_U636
g6679 nand R2358_U397 R2358_U214 ; R2358_U637
g6680 nand R2358_U115 R2358_U357 ; R2358_U638
g6681 nand R2358_U398 R2358_U215 ; R2358_U639
g6682 nand R2358_U117 R2358_U355 ; R2358_U640
g6683 nand R2358_U521 U2636 ; R2358_U641
g6684 nand R2358_U79 R2358_U54 ; R2358_U642
g6685 nand R2358_U642 R2358_U641 ; R2358_U643
g6686 nand R2358_U399 R2358_U72 ; R2358_U644
g6687 nand R2358_U643 R2358_U365 ; R2358_U645
g6688 nand R2358_U526 U2637 ; R2358_U646
g6689 nand R2358_U80 R2358_U50 ; R2358_U647
g6690 nand R2358_U647 R2358_U646 ; R2358_U648
g6691 nand R2358_U400 R2358_U216 ; R2358_U649
g6692 nand R2358_U362 R2358_U648 ; R2358_U650
g6693 nand R2358_U401 R2358_U217 ; R2358_U651
g6694 nand R2358_U121 R2358_U308 ; R2358_U652
g6695 nand U2352 R2358_U218 ; R2358_U653
g6696 nand R2358_U380 R2358_U22 ; R2358_U654
g6697 not PHYADDRPOINTER_REG_1__SCAN_IN ; R2337_U5
g6698 not PHYADDRPOINTER_REG_5__SCAN_IN ; R2337_U6
g6699 not PHYADDRPOINTER_REG_4__SCAN_IN ; R2337_U7
g6700 not PHYADDRPOINTER_REG_3__SCAN_IN ; R2337_U8
g6701 not PHYADDRPOINTER_REG_2__SCAN_IN ; R2337_U9
g6702 nand PHYADDRPOINTER_REG_1__SCAN_IN PHYADDRPOINTER_REG_2__SCAN_IN PHYADDRPOINTER_REG_3__SCAN_IN PHYADDRPOINTER_REG_4__SCAN_IN PHYADDRPOINTER_REG_5__SCAN_IN ; R2337_U10
g6703 not PHYADDRPOINTER_REG_7__SCAN_IN ; R2337_U11
g6704 not PHYADDRPOINTER_REG_6__SCAN_IN ; R2337_U12
g6705 nand R2337_U81 R2337_U108 ; R2337_U13
g6706 not PHYADDRPOINTER_REG_8__SCAN_IN ; R2337_U14
g6707 not PHYADDRPOINTER_REG_9__SCAN_IN ; R2337_U15
g6708 nand PHYADDRPOINTER_REG_1__SCAN_IN PHYADDRPOINTER_REG_2__SCAN_IN PHYADDRPOINTER_REG_3__SCAN_IN ; R2337_U16
g6709 nand R2337_U82 R2337_U110 ; R2337_U17
g6710 not PHYADDRPOINTER_REG_11__SCAN_IN ; R2337_U18
g6711 not PHYADDRPOINTER_REG_10__SCAN_IN ; R2337_U19
g6712 nand R2337_U83 R2337_U112 ; R2337_U20
g6713 not PHYADDRPOINTER_REG_13__SCAN_IN ; R2337_U21
g6714 not PHYADDRPOINTER_REG_12__SCAN_IN ; R2337_U22
g6715 nand R2337_U84 R2337_U114 ; R2337_U23
g6716 not PHYADDRPOINTER_REG_15__SCAN_IN ; R2337_U24
g6717 not PHYADDRPOINTER_REG_14__SCAN_IN ; R2337_U25
g6718 nand R2337_U85 R2337_U116 ; R2337_U26
g6719 not PHYADDRPOINTER_REG_17__SCAN_IN ; R2337_U27
g6720 not PHYADDRPOINTER_REG_16__SCAN_IN ; R2337_U28
g6721 nand R2337_U86 R2337_U118 ; R2337_U29
g6722 not PHYADDRPOINTER_REG_19__SCAN_IN ; R2337_U30
g6723 not PHYADDRPOINTER_REG_18__SCAN_IN ; R2337_U31
g6724 nand R2337_U87 R2337_U120 ; R2337_U32
g6725 not PHYADDRPOINTER_REG_21__SCAN_IN ; R2337_U33
g6726 not PHYADDRPOINTER_REG_20__SCAN_IN ; R2337_U34
g6727 nand R2337_U88 R2337_U122 ; R2337_U35
g6728 not PHYADDRPOINTER_REG_23__SCAN_IN ; R2337_U36
g6729 not PHYADDRPOINTER_REG_22__SCAN_IN ; R2337_U37
g6730 nand R2337_U89 R2337_U124 ; R2337_U38
g6731 not PHYADDRPOINTER_REG_25__SCAN_IN ; R2337_U39
g6732 not PHYADDRPOINTER_REG_24__SCAN_IN ; R2337_U40
g6733 nand R2337_U90 R2337_U126 ; R2337_U41
g6734 not PHYADDRPOINTER_REG_26__SCAN_IN ; R2337_U42
g6735 nand R2337_U128 PHYADDRPOINTER_REG_26__SCAN_IN ; R2337_U43
g6736 not PHYADDRPOINTER_REG_27__SCAN_IN ; R2337_U44
g6737 nand R2337_U129 PHYADDRPOINTER_REG_27__SCAN_IN ; R2337_U45
g6738 not PHYADDRPOINTER_REG_28__SCAN_IN ; R2337_U46
g6739 nand R2337_U130 PHYADDRPOINTER_REG_28__SCAN_IN ; R2337_U47
g6740 not PHYADDRPOINTER_REG_29__SCAN_IN ; R2337_U48
g6741 nand R2337_U131 PHYADDRPOINTER_REG_29__SCAN_IN ; R2337_U49
g6742 not PHYADDRPOINTER_REG_30__SCAN_IN ; R2337_U50
g6743 nand R2337_U135 R2337_U134 ; R2337_U51
g6744 nand R2337_U137 R2337_U136 ; R2337_U52
g6745 nand R2337_U139 R2337_U138 ; R2337_U53
g6746 nand R2337_U141 R2337_U140 ; R2337_U54
g6747 nand R2337_U143 R2337_U142 ; R2337_U55
g6748 nand R2337_U145 R2337_U144 ; R2337_U56
g6749 nand R2337_U147 R2337_U146 ; R2337_U57
g6750 nand R2337_U149 R2337_U148 ; R2337_U58
g6751 nand R2337_U151 R2337_U150 ; R2337_U59
g6752 nand R2337_U153 R2337_U152 ; R2337_U60
g6753 nand R2337_U155 R2337_U154 ; R2337_U61
g6754 nand R2337_U157 R2337_U156 ; R2337_U62
g6755 nand R2337_U159 R2337_U158 ; R2337_U63
g6756 nand R2337_U161 R2337_U160 ; R2337_U64
g6757 nand R2337_U163 R2337_U162 ; R2337_U65
g6758 nand R2337_U165 R2337_U164 ; R2337_U66
g6759 nand R2337_U167 R2337_U166 ; R2337_U67
g6760 nand R2337_U169 R2337_U168 ; R2337_U68
g6761 nand R2337_U171 R2337_U170 ; R2337_U69
g6762 nand R2337_U173 R2337_U172 ; R2337_U70
g6763 nand R2337_U175 R2337_U174 ; R2337_U71
g6764 nand R2337_U177 R2337_U176 ; R2337_U72
g6765 nand R2337_U179 R2337_U178 ; R2337_U73
g6766 nand R2337_U181 R2337_U180 ; R2337_U74
g6767 nand R2337_U183 R2337_U182 ; R2337_U75
g6768 nand R2337_U185 R2337_U184 ; R2337_U76
g6769 nand R2337_U187 R2337_U186 ; R2337_U77
g6770 nand R2337_U189 R2337_U188 ; R2337_U78
g6771 nand R2337_U191 R2337_U190 ; R2337_U79
g6772 nand R2337_U193 R2337_U192 ; R2337_U80
g6773 and PHYADDRPOINTER_REG_6__SCAN_IN PHYADDRPOINTER_REG_7__SCAN_IN ; R2337_U81
g6774 and PHYADDRPOINTER_REG_8__SCAN_IN PHYADDRPOINTER_REG_9__SCAN_IN ; R2337_U82
g6775 and PHYADDRPOINTER_REG_10__SCAN_IN PHYADDRPOINTER_REG_11__SCAN_IN ; R2337_U83
g6776 and PHYADDRPOINTER_REG_12__SCAN_IN PHYADDRPOINTER_REG_13__SCAN_IN ; R2337_U84
g6777 and PHYADDRPOINTER_REG_14__SCAN_IN PHYADDRPOINTER_REG_15__SCAN_IN ; R2337_U85
g6778 and PHYADDRPOINTER_REG_16__SCAN_IN PHYADDRPOINTER_REG_17__SCAN_IN ; R2337_U86
g6779 and PHYADDRPOINTER_REG_18__SCAN_IN PHYADDRPOINTER_REG_19__SCAN_IN ; R2337_U87
g6780 and PHYADDRPOINTER_REG_20__SCAN_IN PHYADDRPOINTER_REG_21__SCAN_IN ; R2337_U88
g6781 and PHYADDRPOINTER_REG_22__SCAN_IN PHYADDRPOINTER_REG_23__SCAN_IN ; R2337_U89
g6782 and PHYADDRPOINTER_REG_24__SCAN_IN PHYADDRPOINTER_REG_25__SCAN_IN ; R2337_U90
g6783 nand R2337_U110 PHYADDRPOINTER_REG_8__SCAN_IN ; R2337_U91
g6784 nand R2337_U108 PHYADDRPOINTER_REG_6__SCAN_IN ; R2337_U92
g6785 nand R2337_U106 PHYADDRPOINTER_REG_4__SCAN_IN ; R2337_U93
g6786 nand PHYADDRPOINTER_REG_1__SCAN_IN PHYADDRPOINTER_REG_2__SCAN_IN ; R2337_U94
g6787 not PHYADDRPOINTER_REG_31__SCAN_IN ; R2337_U95
g6788 nand R2337_U132 PHYADDRPOINTER_REG_30__SCAN_IN ; R2337_U96
g6789 nand R2337_U126 PHYADDRPOINTER_REG_24__SCAN_IN ; R2337_U97
g6790 nand R2337_U124 PHYADDRPOINTER_REG_22__SCAN_IN ; R2337_U98
g6791 nand R2337_U122 PHYADDRPOINTER_REG_20__SCAN_IN ; R2337_U99
g6792 nand R2337_U120 PHYADDRPOINTER_REG_18__SCAN_IN ; R2337_U100
g6793 nand R2337_U118 PHYADDRPOINTER_REG_16__SCAN_IN ; R2337_U101
g6794 nand R2337_U116 PHYADDRPOINTER_REG_14__SCAN_IN ; R2337_U102
g6795 nand R2337_U114 PHYADDRPOINTER_REG_12__SCAN_IN ; R2337_U103
g6796 nand R2337_U112 PHYADDRPOINTER_REG_10__SCAN_IN ; R2337_U104
g6797 not R2337_U94 ; R2337_U105
g6798 not R2337_U16 ; R2337_U106
g6799 not R2337_U93 ; R2337_U107
g6800 not R2337_U10 ; R2337_U108
g6801 not R2337_U92 ; R2337_U109
g6802 not R2337_U13 ; R2337_U110
g6803 not R2337_U91 ; R2337_U111
g6804 not R2337_U17 ; R2337_U112
g6805 not R2337_U104 ; R2337_U113
g6806 not R2337_U20 ; R2337_U114
g6807 not R2337_U103 ; R2337_U115
g6808 not R2337_U23 ; R2337_U116
g6809 not R2337_U102 ; R2337_U117
g6810 not R2337_U26 ; R2337_U118
g6811 not R2337_U101 ; R2337_U119
g6812 not R2337_U29 ; R2337_U120
g6813 not R2337_U100 ; R2337_U121
g6814 not R2337_U32 ; R2337_U122
g6815 not R2337_U99 ; R2337_U123
g6816 not R2337_U35 ; R2337_U124
g6817 not R2337_U98 ; R2337_U125
g6818 not R2337_U38 ; R2337_U126
g6819 not R2337_U97 ; R2337_U127
g6820 not R2337_U41 ; R2337_U128
g6821 not R2337_U43 ; R2337_U129
g6822 not R2337_U45 ; R2337_U130
g6823 not R2337_U47 ; R2337_U131
g6824 not R2337_U49 ; R2337_U132
g6825 not R2337_U96 ; R2337_U133
g6826 nand R2337_U91 PHYADDRPOINTER_REG_9__SCAN_IN ; R2337_U134
g6827 nand R2337_U111 R2337_U15 ; R2337_U135
g6828 nand R2337_U13 PHYADDRPOINTER_REG_8__SCAN_IN ; R2337_U136
g6829 nand R2337_U110 R2337_U14 ; R2337_U137
g6830 nand R2337_U92 PHYADDRPOINTER_REG_7__SCAN_IN ; R2337_U138
g6831 nand R2337_U109 R2337_U11 ; R2337_U139
g6832 nand R2337_U10 PHYADDRPOINTER_REG_6__SCAN_IN ; R2337_U140
g6833 nand R2337_U108 R2337_U12 ; R2337_U141
g6834 nand R2337_U93 PHYADDRPOINTER_REG_5__SCAN_IN ; R2337_U142
g6835 nand R2337_U107 R2337_U6 ; R2337_U143
g6836 nand R2337_U16 PHYADDRPOINTER_REG_4__SCAN_IN ; R2337_U144
g6837 nand R2337_U106 R2337_U7 ; R2337_U145
g6838 nand R2337_U94 PHYADDRPOINTER_REG_3__SCAN_IN ; R2337_U146
g6839 nand R2337_U105 R2337_U8 ; R2337_U147
g6840 nand R2337_U96 PHYADDRPOINTER_REG_31__SCAN_IN ; R2337_U148
g6841 nand R2337_U133 R2337_U95 ; R2337_U149
g6842 nand R2337_U49 PHYADDRPOINTER_REG_30__SCAN_IN ; R2337_U150
g6843 nand R2337_U132 R2337_U50 ; R2337_U151
g6844 nand R2337_U9 PHYADDRPOINTER_REG_1__SCAN_IN ; R2337_U152
g6845 nand R2337_U5 PHYADDRPOINTER_REG_2__SCAN_IN ; R2337_U153
g6846 nand R2337_U47 PHYADDRPOINTER_REG_29__SCAN_IN ; R2337_U154
g6847 nand R2337_U131 R2337_U48 ; R2337_U155
g6848 nand R2337_U45 PHYADDRPOINTER_REG_28__SCAN_IN ; R2337_U156
g6849 nand R2337_U130 R2337_U46 ; R2337_U157
g6850 nand R2337_U43 PHYADDRPOINTER_REG_27__SCAN_IN ; R2337_U158
g6851 nand R2337_U129 R2337_U44 ; R2337_U159
g6852 nand R2337_U41 PHYADDRPOINTER_REG_26__SCAN_IN ; R2337_U160
g6853 nand R2337_U128 R2337_U42 ; R2337_U161
g6854 nand R2337_U97 PHYADDRPOINTER_REG_25__SCAN_IN ; R2337_U162
g6855 nand R2337_U127 R2337_U39 ; R2337_U163
g6856 nand R2337_U38 PHYADDRPOINTER_REG_24__SCAN_IN ; R2337_U164
g6857 nand R2337_U126 R2337_U40 ; R2337_U165
g6858 nand R2337_U98 PHYADDRPOINTER_REG_23__SCAN_IN ; R2337_U166
g6859 nand R2337_U125 R2337_U36 ; R2337_U167
g6860 nand R2337_U35 PHYADDRPOINTER_REG_22__SCAN_IN ; R2337_U168
g6861 nand R2337_U124 R2337_U37 ; R2337_U169
g6862 nand R2337_U99 PHYADDRPOINTER_REG_21__SCAN_IN ; R2337_U170
g6863 nand R2337_U123 R2337_U33 ; R2337_U171
g6864 nand R2337_U32 PHYADDRPOINTER_REG_20__SCAN_IN ; R2337_U172
g6865 nand R2337_U122 R2337_U34 ; R2337_U173
g6866 nand R2337_U100 PHYADDRPOINTER_REG_19__SCAN_IN ; R2337_U174
g6867 nand R2337_U121 R2337_U30 ; R2337_U175
g6868 nand R2337_U29 PHYADDRPOINTER_REG_18__SCAN_IN ; R2337_U176
g6869 nand R2337_U120 R2337_U31 ; R2337_U177
g6870 nand R2337_U101 PHYADDRPOINTER_REG_17__SCAN_IN ; R2337_U178
g6871 nand R2337_U119 R2337_U27 ; R2337_U179
g6872 nand R2337_U26 PHYADDRPOINTER_REG_16__SCAN_IN ; R2337_U180
g6873 nand R2337_U118 R2337_U28 ; R2337_U181
g6874 nand R2337_U102 PHYADDRPOINTER_REG_15__SCAN_IN ; R2337_U182
g6875 nand R2337_U117 R2337_U24 ; R2337_U183
g6876 nand R2337_U23 PHYADDRPOINTER_REG_14__SCAN_IN ; R2337_U184
g6877 nand R2337_U116 R2337_U25 ; R2337_U185
g6878 nand R2337_U103 PHYADDRPOINTER_REG_13__SCAN_IN ; R2337_U186
g6879 nand R2337_U115 R2337_U21 ; R2337_U187
g6880 nand R2337_U20 PHYADDRPOINTER_REG_12__SCAN_IN ; R2337_U188
g6881 nand R2337_U114 R2337_U22 ; R2337_U189
g6882 nand R2337_U104 PHYADDRPOINTER_REG_11__SCAN_IN ; R2337_U190
g6883 nand R2337_U113 R2337_U18 ; R2337_U191
g6884 nand R2337_U17 PHYADDRPOINTER_REG_10__SCAN_IN ; R2337_U192
g6885 nand R2337_U112 R2337_U19 ; R2337_U193
g6886 and R2182_U47 U2740 ; R2182_U5
g6887 and R2182_U60 R2182_U16 ; R2182_U6
g6888 not U2744 ; R2182_U7
g6889 not U3233 ; R2182_U8
g6890 nand U3233 U2744 ; R2182_U9
g6891 not U2742 ; R2182_U10
g6892 not U2741 ; R2182_U11
g6893 not U2740 ; R2182_U12
g6894 nand R2182_U35 R2182_U41 ; R2182_U13
g6895 not U2737 ; R2182_U14
g6896 not U2738 ; R2182_U15
g6897 nand U2723 U2739 ; R2182_U16
g6898 not U2736 ; R2182_U17
g6899 not U2735 ; R2182_U18
g6900 nand R2182_U36 R2182_U49 ; R2182_U19
g6901 not U2734 ; R2182_U20
g6902 nand R2182_U37 R2182_U46 ; R2182_U21
g6903 nand R2182_U48 U2734 ; R2182_U22
g6904 not U2733 ; R2182_U23
g6905 nand R2182_U64 R2182_U63 ; R2182_U24
g6906 nand R2182_U66 R2182_U65 ; R2182_U25
g6907 nand R2182_U68 R2182_U67 ; R2182_U26
g6908 nand R2182_U72 R2182_U71 ; R2182_U27
g6909 nand R2182_U74 R2182_U73 ; R2182_U28
g6910 nand R2182_U76 R2182_U75 ; R2182_U29
g6911 nand R2182_U78 R2182_U77 ; R2182_U30
g6912 nand R2182_U80 R2182_U79 ; R2182_U31
g6913 nand R2182_U82 R2182_U81 ; R2182_U32
g6914 nand R2182_U84 R2182_U83 ; R2182_U33
g6915 nand R2182_U86 R2182_U85 ; R2182_U34
g6916 and U2742 U2741 ; R2182_U35
g6917 and U2738 U2737 ; R2182_U36
g6918 and U2735 U2736 ; R2182_U37
g6919 nand U2742 R2182_U41 ; R2182_U38
g6920 not U2732 ; R2182_U39
g6921 nand U2733 R2182_U56 ; R2182_U40
g6922 nand R2182_U52 R2182_U53 ; R2182_U41
g6923 and R2182_U70 R2182_U69 ; R2182_U42
g6924 nand R2182_U46 U2736 ; R2182_U43
g6925 nand R2182_U49 U2738 ; R2182_U44
g6926 nand R2182_U51 R2182_U62 ; R2182_U45
g6927 not R2182_U19 ; R2182_U46
g6928 not R2182_U13 ; R2182_U47
g6929 not R2182_U21 ; R2182_U48
g6930 not R2182_U16 ; R2182_U49
g6931 not R2182_U9 ; R2182_U50
g6932 or U2743 U2731 ; R2182_U51
g6933 nand U2731 U2743 ; R2182_U52
g6934 nand R2182_U50 R2182_U51 ; R2182_U53
g6935 not R2182_U41 ; R2182_U54
g6936 not R2182_U38 ; R2182_U55
g6937 not R2182_U22 ; R2182_U56
g6938 not R2182_U40 ; R2182_U57
g6939 not R2182_U43 ; R2182_U58
g6940 not R2182_U44 ; R2182_U59
g6941 or U2739 U2723 ; R2182_U60
g6942 not R2182_U45 ; R2182_U61
g6943 nand U2731 U2743 ; R2182_U62
g6944 nand R2182_U47 R2182_U12 ; R2182_U63
g6945 nand U2740 R2182_U13 ; R2182_U64
g6946 nand U2741 R2182_U38 ; R2182_U65
g6947 nand R2182_U55 R2182_U11 ; R2182_U66
g6948 nand U2732 R2182_U40 ; R2182_U67
g6949 nand R2182_U57 R2182_U39 ; R2182_U68
g6950 nand U2742 R2182_U41 ; R2182_U69
g6951 nand R2182_U54 R2182_U10 ; R2182_U70
g6952 nand U2733 R2182_U22 ; R2182_U71
g6953 nand R2182_U56 R2182_U23 ; R2182_U72
g6954 nand R2182_U48 R2182_U20 ; R2182_U73
g6955 nand U2734 R2182_U21 ; R2182_U74
g6956 nand U2735 R2182_U43 ; R2182_U75
g6957 nand R2182_U58 R2182_U18 ; R2182_U76
g6958 nand R2182_U46 R2182_U17 ; R2182_U77
g6959 nand U2736 R2182_U19 ; R2182_U78
g6960 nand U2737 R2182_U44 ; R2182_U79
g6961 nand R2182_U59 R2182_U14 ; R2182_U80
g6962 nand R2182_U49 R2182_U15 ; R2182_U81
g6963 nand U2738 R2182_U16 ; R2182_U82
g6964 nand R2182_U50 R2182_U45 ; R2182_U83
g6965 nand R2182_U61 R2182_U9 ; R2182_U84
g6966 nand U3233 R2182_U7 ; R2182_U85
g6967 nand U2744 R2182_U8 ; R2182_U86
g6968 and R2144_U104 R2144_U103 ; R2144_U5
g6969 and R2144_U36 R2144_U35 R2144_U27 R2144_U29 ; R2144_U6
g6970 and R2144_U104 R2144_U81 ; R2144_U7
g6971 and R2144_U138 R2144_U136 ; R2144_U8
g6972 and R2144_U128 R2144_U127 ; R2144_U9
g6973 and R2144_U213 R2144_U212 R2144_U82 ; R2144_U10
g6974 nand R2144_U144 R2144_U146 ; R2144_U11
g6975 not U2355 ; R2144_U12
g6976 not U2750 ; R2144_U13
g6977 not U2751 ; R2144_U14
g6978 not U2752 ; R2144_U15
g6979 not U2749 ; R2144_U16
g6980 not U2745 ; R2144_U17
g6981 not U2748 ; R2144_U18
g6982 nand U2748 R2144_U178 ; R2144_U19
g6983 not U2747 ; R2144_U20
g6984 nand U2747 R2144_U170 ; R2144_U21
g6985 not U2746 ; R2144_U22
g6986 nand U2746 R2144_U173 ; R2144_U23
g6987 nand R2144_U79 R2144_U63 ; R2144_U24
g6988 nand R2144_U6 R2144_U79 ; R2144_U25
g6989 nand R2144_U65 R2144_U141 ; R2144_U26
g6990 nand R2144_U206 R2144_U205 ; R2144_U27
g6991 nand R2144_U186 R2144_U185 ; R2144_U28
g6992 nand R2144_U203 R2144_U202 ; R2144_U29
g6993 nand R2144_U209 R2144_U208 ; R2144_U30
g6994 nand R2144_U224 R2144_U223 ; R2144_U31
g6995 nand R2144_U221 R2144_U220 ; R2144_U32
g6996 nand R2144_U227 R2144_U226 ; R2144_U33
g6997 nand R2144_U230 R2144_U229 ; R2144_U34
g6998 nand R2144_U233 R2144_U232 ; R2144_U35
g6999 nand R2144_U236 R2144_U235 ; R2144_U36
g7000 nand R2144_U248 R2144_U247 ; R2144_U37
g7001 nand R2144_U250 R2144_U249 ; R2144_U38
g7002 nand R2144_U252 R2144_U251 ; R2144_U39
g7003 nand R2144_U254 R2144_U253 ; R2144_U40
g7004 nand R2144_U256 R2144_U255 ; R2144_U41
g7005 nand R2144_U258 R2144_U257 ; R2144_U42
g7006 nand R2144_U260 R2144_U259 ; R2144_U43
g7007 and R2144_U21 R2144_U105 ; R2144_U44
g7008 nand R2144_U217 R2144_U216 ; R2144_U45
g7009 and R2144_U19 R2144_U106 ; R2144_U46
g7010 nand R2144_U219 R2144_U218 ; R2144_U47
g7011 and R2144_U162 R2144_U109 ; R2144_U48
g7012 nand R2144_U239 R2144_U238 ; R2144_U49
g7013 nand R2144_U246 R2144_U245 ; R2144_U50
g7014 and R2144_U110 R2144_U109 ; R2144_U51
g7015 and R2144_U106 R2144_U105 ; R2144_U52
g7016 and R2144_U7 R2144_U52 ; R2144_U53
g7017 and R2144_U103 R2144_U151 R2144_U153 R2144_U152 ; R2144_U54
g7018 and R2144_U109 R2144_U106 ; R2144_U55
g7019 and R2144_U159 R2144_U19 ; R2144_U56
g7020 and R2144_U156 R2144_U21 ; R2144_U57
g7021 and R2144_U19 R2144_U21 R2144_U159 ; R2144_U58
g7022 and R2144_U5 R2144_U105 ; R2144_U59
g7023 and R2144_U126 R2144_U21 ; R2144_U60
g7024 and R2144_U23 R2144_U81 ; R2144_U61
g7025 and R2144_U111 R2144_U110 ; R2144_U62
g7026 and R2144_U6 R2144_U64 ; R2144_U63
g7027 and R2144_U34 R2144_U33 R2144_U31 R2144_U32 ; R2144_U64
g7028 and R2144_U34 R2144_U33 ; R2144_U65
g7029 and R2144_U36 R2144_U27 R2144_U29 ; R2144_U66
g7030 and R2144_U29 R2144_U27 ; R2144_U67
g7031 not U2762 ; R2144_U68
g7032 not U2761 ; R2144_U69
g7033 not U2763 ; R2144_U70
g7034 not U2764 ; R2144_U71
g7035 not U2766 ; R2144_U72
g7036 not U2767 ; R2144_U73
g7037 not U2768 ; R2144_U74
g7038 not U2765 ; R2144_U75
g7039 not U2760 ; R2144_U76
g7040 not U2759 ; R2144_U77
g7041 nand R2144_U29 R2144_U79 ; R2144_U78
g7042 nand R2144_U99 R2144_U54 ; R2144_U79
g7043 and R2144_U211 R2144_U210 ; R2144_U80
g7044 nand R2144_U165 R2144_U164 R2144_U22 ; R2144_U81
g7045 and R2144_U215 R2144_U214 ; R2144_U82
g7046 nand R2144_U56 R2144_U158 ; R2144_U83
g7047 nand R2144_U111 R2144_U118 ; R2144_U84
g7048 not U2754 ; R2144_U85
g7049 not U2753 ; R2144_U86
g7050 not U2755 ; R2144_U87
g7051 not U2756 ; R2144_U88
g7052 not U2757 ; R2144_U89
g7053 not U2758 ; R2144_U90
g7054 nand R2144_U100 R2144_U132 ; R2144_U91
g7055 and R2144_U241 R2144_U240 ; R2144_U92
g7056 nand R2144_U129 R2144_U113 ; R2144_U93
g7057 nand R2144_U143 R2144_U32 ; R2144_U94
g7058 nand R2144_U141 R2144_U34 ; R2144_U95
g7059 nand R2144_U79 R2144_U66 ; R2144_U96
g7060 nand R2144_U67 R2144_U79 ; R2144_U97
g7061 nand R2144_U113 R2144_U112 ; R2144_U98
g7062 nand R2144_U53 R2144_U84 ; R2144_U99
g7063 nand U2751 R2144_U28 ; R2144_U100
g7064 not R2144_U24 ; R2144_U101
g7065 not R2144_U81 ; R2144_U102
g7066 nand U2745 R2144_U181 ; R2144_U103
g7067 nand R2144_U167 R2144_U166 R2144_U17 ; R2144_U104
g7068 nand R2144_U175 R2144_U174 R2144_U20 ; R2144_U105
g7069 nand R2144_U201 R2144_U200 R2144_U18 ; R2144_U106
g7070 not R2144_U21 ; R2144_U107
g7071 not R2144_U23 ; R2144_U108
g7072 nand R2144_U194 R2144_U193 R2144_U13 ; R2144_U109
g7073 nand R2144_U196 R2144_U195 R2144_U16 ; R2144_U110
g7074 nand U2749 R2144_U199 ; R2144_U111
g7075 nand R2144_U189 R2144_U188 R2144_U15 ; R2144_U112
g7076 nand U2752 R2144_U192 ; R2144_U113
g7077 nand R2144_U187 R2144_U14 ; R2144_U114
g7078 nand U2355 R2144_U112 ; R2144_U115
g7079 nand U2750 R2144_U184 ; R2144_U116
g7080 nand R2144_U155 R2144_U157 ; R2144_U117
g7081 nand R2144_U51 R2144_U117 ; R2144_U118
g7082 not R2144_U84 ; R2144_U119
g7083 not R2144_U19 ; R2144_U120
g7084 not R2144_U79 ; R2144_U121
g7085 not R2144_U78 ; R2144_U122
g7086 not R2144_U83 ; R2144_U123
g7087 nand R2144_U83 R2144_U105 ; R2144_U124
g7088 nand R2144_U21 R2144_U124 ; R2144_U125
g7089 nand R2144_U23 R2144_U81 ; R2144_U126
g7090 nand R2144_U60 R2144_U124 ; R2144_U127
g7091 nand R2144_U61 R2144_U125 ; R2144_U128
g7092 nand U2355 R2144_U112 ; R2144_U129
g7093 not R2144_U93 ; R2144_U130
g7094 nand R2144_U187 R2144_U14 ; R2144_U131
g7095 nand R2144_U131 R2144_U93 ; R2144_U132
g7096 not R2144_U91 ; R2144_U133
g7097 nand R2144_U91 R2144_U109 ; R2144_U134
g7098 nand R2144_U134 R2144_U116 ; R2144_U135
g7099 nand R2144_U62 R2144_U135 ; R2144_U136
g7100 nand R2144_U161 R2144_U110 ; R2144_U137
g7101 nand R2144_U134 R2144_U116 R2144_U137 ; R2144_U138
g7102 not R2144_U97 ; R2144_U139
g7103 not R2144_U96 ; R2144_U140
g7104 not R2144_U25 ; R2144_U141
g7105 not R2144_U95 ; R2144_U142
g7106 not R2144_U26 ; R2144_U143
g7107 nand U2355 R2144_U24 ; R2144_U144
g7108 not R2144_U144 ; R2144_U145
g7109 nand R2144_U101 R2144_U12 ; R2144_U146
g7110 not R2144_U94 ; R2144_U147
g7111 not R2144_U98 ; R2144_U148
g7112 nand R2144_U21 R2144_U105 ; R2144_U149
g7113 nand R2144_U19 R2144_U106 ; R2144_U150
g7114 nand R2144_U120 R2144_U105 R2144_U7 ; R2144_U151
g7115 nand R2144_U107 R2144_U7 ; R2144_U152
g7116 nand R2144_U108 R2144_U7 ; R2144_U153
g7117 nand R2144_U113 R2144_U115 R2144_U100 ; R2144_U154
g7118 nand R2144_U154 R2144_U114 ; R2144_U155
g7119 nand R2144_U104 R2144_U103 ; R2144_U156
g7120 nand U2750 R2144_U184 ; R2144_U157
g7121 nand R2144_U117 R2144_U110 R2144_U55 ; R2144_U158
g7122 nand U2749 R2144_U106 R2144_U199 ; R2144_U159
g7123 nand R2144_U58 R2144_U158 ; R2144_U160
g7124 nand U2749 R2144_U199 ; R2144_U161
g7125 nand U2750 R2144_U184 ; R2144_U162
g7126 nand R2144_U116 R2144_U109 ; R2144_U163
g7127 nand U2355 R2144_U68 ; R2144_U164
g7128 nand U2762 R2144_U12 ; R2144_U165
g7129 nand U2355 R2144_U69 ; R2144_U166
g7130 nand U2761 R2144_U12 ; R2144_U167
g7131 nand U2355 R2144_U70 ; R2144_U168
g7132 nand U2763 R2144_U12 ; R2144_U169
g7133 nand R2144_U169 R2144_U168 ; R2144_U170
g7134 nand U2355 R2144_U68 ; R2144_U171
g7135 nand U2762 R2144_U12 ; R2144_U172
g7136 nand R2144_U172 R2144_U171 ; R2144_U173
g7137 nand U2355 R2144_U70 ; R2144_U174
g7138 nand U2763 R2144_U12 ; R2144_U175
g7139 nand U2355 R2144_U71 ; R2144_U176
g7140 nand U2764 R2144_U12 ; R2144_U177
g7141 nand R2144_U177 R2144_U176 ; R2144_U178
g7142 nand U2355 R2144_U69 ; R2144_U179
g7143 nand U2761 R2144_U12 ; R2144_U180
g7144 nand R2144_U180 R2144_U179 ; R2144_U181
g7145 nand U2355 R2144_U72 ; R2144_U182
g7146 nand U2766 R2144_U12 ; R2144_U183
g7147 nand R2144_U183 R2144_U182 ; R2144_U184
g7148 nand U2355 R2144_U73 ; R2144_U185
g7149 nand U2767 R2144_U12 ; R2144_U186
g7150 not R2144_U28 ; R2144_U187
g7151 nand U2355 R2144_U74 ; R2144_U188
g7152 nand U2768 R2144_U12 ; R2144_U189
g7153 nand U2355 R2144_U74 ; R2144_U190
g7154 nand U2768 R2144_U12 ; R2144_U191
g7155 nand R2144_U191 R2144_U190 ; R2144_U192
g7156 nand U2355 R2144_U72 ; R2144_U193
g7157 nand U2766 R2144_U12 ; R2144_U194
g7158 nand U2355 R2144_U75 ; R2144_U195
g7159 nand U2765 R2144_U12 ; R2144_U196
g7160 nand U2355 R2144_U75 ; R2144_U197
g7161 nand U2765 R2144_U12 ; R2144_U198
g7162 nand R2144_U198 R2144_U197 ; R2144_U199
g7163 nand U2355 R2144_U71 ; R2144_U200
g7164 nand U2764 R2144_U12 ; R2144_U201
g7165 nand U2355 R2144_U76 ; R2144_U202
g7166 nand U2760 R2144_U12 ; R2144_U203
g7167 not R2144_U29 ; R2144_U204
g7168 nand U2355 R2144_U77 ; R2144_U205
g7169 nand U2759 R2144_U12 ; R2144_U206
g7170 not R2144_U27 ; R2144_U207
g7171 nand R2144_U122 R2144_U207 ; R2144_U208
g7172 nand R2144_U27 R2144_U78 ; R2144_U209
g7173 nand R2144_U121 R2144_U204 ; R2144_U210
g7174 nand R2144_U29 R2144_U79 ; R2144_U211
g7175 nand R2144_U57 R2144_U124 R2144_U23 ; R2144_U212
g7176 nand R2144_U5 R2144_U108 ; R2144_U213
g7177 nand R2144_U102 R2144_U156 ; R2144_U214
g7178 nand R2144_U59 R2144_U160 R2144_U81 ; R2144_U215
g7179 nand R2144_U149 R2144_U83 ; R2144_U216
g7180 nand R2144_U44 R2144_U123 ; R2144_U217
g7181 nand R2144_U150 R2144_U84 ; R2144_U218
g7182 nand R2144_U46 R2144_U119 ; R2144_U219
g7183 nand U2355 R2144_U85 ; R2144_U220
g7184 nand U2754 R2144_U12 ; R2144_U221
g7185 not R2144_U32 ; R2144_U222
g7186 nand U2355 R2144_U86 ; R2144_U223
g7187 nand U2753 R2144_U12 ; R2144_U224
g7188 not R2144_U31 ; R2144_U225
g7189 nand U2355 R2144_U87 ; R2144_U226
g7190 nand U2755 R2144_U12 ; R2144_U227
g7191 not R2144_U33 ; R2144_U228
g7192 nand U2355 R2144_U88 ; R2144_U229
g7193 nand U2756 R2144_U12 ; R2144_U230
g7194 not R2144_U34 ; R2144_U231
g7195 nand U2355 R2144_U89 ; R2144_U232
g7196 nand U2757 R2144_U12 ; R2144_U233
g7197 not R2144_U35 ; R2144_U234
g7198 nand U2355 R2144_U90 ; R2144_U235
g7199 nand U2758 R2144_U12 ; R2144_U236
g7200 not R2144_U36 ; R2144_U237
g7201 nand R2144_U163 R2144_U91 ; R2144_U238
g7202 nand R2144_U48 R2144_U133 ; R2144_U239
g7203 nand R2144_U187 U2751 ; R2144_U240
g7204 nand R2144_U28 R2144_U14 ; R2144_U241
g7205 nand R2144_U187 U2751 ; R2144_U242
g7206 nand R2144_U28 R2144_U14 ; R2144_U243
g7207 nand R2144_U243 R2144_U242 ; R2144_U244
g7208 nand R2144_U92 R2144_U93 ; R2144_U245
g7209 nand R2144_U130 R2144_U244 ; R2144_U246
g7210 nand R2144_U147 R2144_U225 ; R2144_U247
g7211 nand R2144_U31 R2144_U94 ; R2144_U248
g7212 nand R2144_U222 R2144_U143 ; R2144_U249
g7213 nand R2144_U32 R2144_U26 ; R2144_U250
g7214 nand R2144_U142 R2144_U228 ; R2144_U251
g7215 nand R2144_U33 R2144_U95 ; R2144_U252
g7216 nand R2144_U231 R2144_U141 ; R2144_U253
g7217 nand R2144_U34 R2144_U25 ; R2144_U254
g7218 nand R2144_U140 R2144_U234 ; R2144_U255
g7219 nand R2144_U35 R2144_U96 ; R2144_U256
g7220 nand R2144_U139 R2144_U237 ; R2144_U257
g7221 nand R2144_U36 R2144_U97 ; R2144_U258
g7222 nand U2355 R2144_U98 ; R2144_U259
g7223 nand R2144_U148 R2144_U12 ; R2144_U260
g7224 or LT_589_U8 U2673 ; LT_589_U6
g7225 and R584_U7 R584_U6 ; LT_589_U7
g7226 nor LT_589_U7 R584_U9 R584_U8 ; LT_589_U8
g7227 not U2676 ; R584_U6
g7228 not U2677 ; R584_U7
g7229 not U2674 ; R584_U8
g7230 not U2675 ; R584_U9
g7231 not U4178 ; R2099_U4
g7232 not U4177 ; R2099_U5
g7233 not U2678 ; R2099_U6
g7234 nand R2099_U88 R2099_U137 ; R2099_U7
g7235 nand R2099_U89 R2099_U155 ; R2099_U8
g7236 nand R2099_U90 R2099_U157 ; R2099_U9
g7237 nand R2099_U91 R2099_U159 ; R2099_U10
g7238 nand R2099_U92 R2099_U161 ; R2099_U11
g7239 nand R2099_U93 R2099_U163 ; R2099_U12
g7240 nand R2099_U94 R2099_U165 ; R2099_U13
g7241 nand R2099_U95 R2099_U167 ; R2099_U14
g7242 nand R2099_U169 R2099_U55 ; R2099_U15
g7243 nand R2099_U170 R2099_U54 ; R2099_U16
g7244 nand R2099_U171 R2099_U53 ; R2099_U17
g7245 nand R2099_U172 R2099_U52 ; R2099_U18
g7246 nand R2099_U173 R2099_U51 ; R2099_U19
g7247 nand R2099_U174 R2099_U50 ; R2099_U20
g7248 nand R2099_U175 R2099_U49 ; R2099_U21
g7249 nand R2099_U176 R2099_U48 ; R2099_U22
g7250 nand R2099_U177 R2099_U47 ; R2099_U23
g7251 nand R2099_U178 R2099_U46 ; R2099_U24
g7252 nand R2099_U179 R2099_U45 ; R2099_U25
g7253 nand R2099_U210 R2099_U209 ; R2099_U26
g7254 nand R2099_U183 R2099_U182 ; R2099_U27
g7255 nand R2099_U204 R2099_U203 ; R2099_U28
g7256 nand R2099_U207 R2099_U206 ; R2099_U29
g7257 nand R2099_U198 R2099_U197 ; R2099_U30
g7258 nand R2099_U201 R2099_U200 ; R2099_U31
g7259 nand R2099_U186 R2099_U185 ; R2099_U32
g7260 nand R2099_U189 R2099_U188 ; R2099_U33
g7261 nand R2099_U195 R2099_U194 ; R2099_U34
g7262 nand R2099_U192 R2099_U191 ; R2099_U35
g7263 nand R2099_U213 R2099_U212 ; R2099_U36
g7264 nand R2099_U215 R2099_U214 ; R2099_U37
g7265 nand R2099_U217 R2099_U216 ; R2099_U38
g7266 nand R2099_U219 R2099_U218 ; R2099_U39
g7267 nand R2099_U221 R2099_U220 ; R2099_U40
g7268 nand R2099_U223 R2099_U222 ; R2099_U41
g7269 nand R2099_U225 R2099_U224 ; R2099_U42
g7270 nand R2099_U284 R2099_U283 ; R2099_U43
g7271 nand R2099_U287 R2099_U286 ; R2099_U44
g7272 nand R2099_U227 R2099_U226 ; R2099_U45
g7273 nand R2099_U230 R2099_U229 ; R2099_U46
g7274 nand R2099_U233 R2099_U232 ; R2099_U47
g7275 nand R2099_U236 R2099_U235 ; R2099_U48
g7276 nand R2099_U239 R2099_U238 ; R2099_U49
g7277 nand R2099_U242 R2099_U241 ; R2099_U50
g7278 nand R2099_U245 R2099_U244 ; R2099_U51
g7279 nand R2099_U248 R2099_U247 ; R2099_U52
g7280 nand R2099_U251 R2099_U250 ; R2099_U53
g7281 nand R2099_U254 R2099_U253 ; R2099_U54
g7282 nand R2099_U257 R2099_U256 ; R2099_U55
g7283 nand R2099_U278 R2099_U277 ; R2099_U56
g7284 nand R2099_U281 R2099_U280 ; R2099_U57
g7285 nand R2099_U272 R2099_U271 ; R2099_U58
g7286 nand R2099_U275 R2099_U274 ; R2099_U59
g7287 nand R2099_U266 R2099_U265 ; R2099_U60
g7288 nand R2099_U269 R2099_U268 ; R2099_U61
g7289 nand R2099_U260 R2099_U259 ; R2099_U62
g7290 nand R2099_U263 R2099_U262 ; R2099_U63
g7291 nand R2099_U293 R2099_U292 ; R2099_U64
g7292 nand R2099_U295 R2099_U294 ; R2099_U65
g7293 nand R2099_U299 R2099_U298 ; R2099_U66
g7294 nand R2099_U301 R2099_U300 ; R2099_U67
g7295 nand R2099_U303 R2099_U302 ; R2099_U68
g7296 nand R2099_U305 R2099_U304 ; R2099_U69
g7297 nand R2099_U307 R2099_U306 ; R2099_U70
g7298 nand R2099_U309 R2099_U308 ; R2099_U71
g7299 nand R2099_U311 R2099_U310 ; R2099_U72
g7300 nand R2099_U313 R2099_U312 ; R2099_U73
g7301 nand R2099_U315 R2099_U314 ; R2099_U74
g7302 nand R2099_U317 R2099_U316 ; R2099_U75
g7303 nand R2099_U326 R2099_U325 ; R2099_U76
g7304 nand R2099_U328 R2099_U327 ; R2099_U77
g7305 nand R2099_U330 R2099_U329 ; R2099_U78
g7306 nand R2099_U332 R2099_U331 ; R2099_U79
g7307 nand R2099_U334 R2099_U333 ; R2099_U80
g7308 nand R2099_U336 R2099_U335 ; R2099_U81
g7309 nand R2099_U338 R2099_U337 ; R2099_U82
g7310 nand R2099_U340 R2099_U339 ; R2099_U83
g7311 nand R2099_U342 R2099_U341 ; R2099_U84
g7312 nand R2099_U344 R2099_U343 ; R2099_U85
g7313 nand R2099_U349 R2099_U348 ; R2099_U86
g7314 nand R2099_U324 R2099_U323 ; R2099_U87
g7315 and R2099_U34 R2099_U35 ; R2099_U88
g7316 and R2099_U31 R2099_U30 ; R2099_U89
g7317 and R2099_U29 R2099_U28 ; R2099_U90
g7318 and R2099_U26 R2099_U27 ; R2099_U91
g7319 and R2099_U63 R2099_U62 ; R2099_U92
g7320 and R2099_U61 R2099_U60 ; R2099_U93
g7321 and R2099_U59 R2099_U58 ; R2099_U94
g7322 and R2099_U57 R2099_U56 ; R2099_U95
g7323 and R2099_U44 R2099_U43 ; R2099_U96
g7324 nand R2099_U290 R2099_U289 ; R2099_U97
g7325 nand R2099_U346 R2099_U345 ; R2099_U98
g7326 not U2702 ; R2099_U99
g7327 not U2710 ; R2099_U100
g7328 not U2709 ; R2099_U101
g7329 not U2708 ; R2099_U102
g7330 not U2707 ; R2099_U103
g7331 not U2706 ; R2099_U104
g7332 not U2705 ; R2099_U105
g7333 not U2704 ; R2099_U106
g7334 not U2703 ; R2099_U107
g7335 not U2701 ; R2099_U108
g7336 nand R2099_U159 R2099_U27 ; R2099_U109
g7337 nand R2099_U157 R2099_U28 ; R2099_U110
g7338 nand R2099_U155 R2099_U30 ; R2099_U111
g7339 nand R2099_U35 R2099_U137 ; R2099_U112
g7340 not U2682 ; R2099_U113
g7341 not U2683 ; R2099_U114
g7342 not U2684 ; R2099_U115
g7343 not U2685 ; R2099_U116
g7344 not U2686 ; R2099_U117
g7345 not U2687 ; R2099_U118
g7346 not U2688 ; R2099_U119
g7347 not U2689 ; R2099_U120
g7348 not U2690 ; R2099_U121
g7349 not U2691 ; R2099_U122
g7350 not U2692 ; R2099_U123
g7351 not U2700 ; R2099_U124
g7352 not U2699 ; R2099_U125
g7353 not U2698 ; R2099_U126
g7354 not U2697 ; R2099_U127
g7355 not U2696 ; R2099_U128
g7356 not U2695 ; R2099_U129
g7357 not U2694 ; R2099_U130
g7358 not U2693 ; R2099_U131
g7359 not U2680 ; R2099_U132
g7360 not U2681 ; R2099_U133
g7361 not U2679 ; R2099_U134
g7362 nand R2099_U96 R2099_U180 ; R2099_U135
g7363 nand R2099_U180 R2099_U44 ; R2099_U136
g7364 nand R2099_U152 R2099_U151 ; R2099_U137
g7365 and R2099_U297 R2099_U296 ; R2099_U138
g7366 and R2099_U319 R2099_U318 ; R2099_U139
g7367 nand R2099_U148 R2099_U147 ; R2099_U140
g7368 nand R2099_U167 R2099_U56 ; R2099_U141
g7369 nand R2099_U165 R2099_U58 ; R2099_U142
g7370 nand R2099_U163 R2099_U60 ; R2099_U143
g7371 nand R2099_U161 R2099_U62 ; R2099_U144
g7372 not R2099_U135 ; R2099_U145
g7373 or U4178 U4177 ; R2099_U146
g7374 nand R2099_U32 R2099_U146 ; R2099_U147
g7375 nand U4177 U4178 ; R2099_U148
g7376 not R2099_U140 ; R2099_U149
g7377 nand R2099_U190 R2099_U6 ; R2099_U150
g7378 nand R2099_U150 R2099_U140 ; R2099_U151
g7379 nand U2678 R2099_U33 ; R2099_U152
g7380 not R2099_U137 ; R2099_U153
g7381 not R2099_U112 ; R2099_U154
g7382 not R2099_U7 ; R2099_U155
g7383 not R2099_U111 ; R2099_U156
g7384 not R2099_U8 ; R2099_U157
g7385 not R2099_U110 ; R2099_U158
g7386 not R2099_U9 ; R2099_U159
g7387 not R2099_U109 ; R2099_U160
g7388 not R2099_U10 ; R2099_U161
g7389 not R2099_U144 ; R2099_U162
g7390 not R2099_U11 ; R2099_U163
g7391 not R2099_U143 ; R2099_U164
g7392 not R2099_U12 ; R2099_U165
g7393 not R2099_U142 ; R2099_U166
g7394 not R2099_U13 ; R2099_U167
g7395 not R2099_U141 ; R2099_U168
g7396 not R2099_U14 ; R2099_U169
g7397 not R2099_U15 ; R2099_U170
g7398 not R2099_U16 ; R2099_U171
g7399 not R2099_U17 ; R2099_U172
g7400 not R2099_U18 ; R2099_U173
g7401 not R2099_U19 ; R2099_U174
g7402 not R2099_U20 ; R2099_U175
g7403 not R2099_U21 ; R2099_U176
g7404 not R2099_U22 ; R2099_U177
g7405 not R2099_U23 ; R2099_U178
g7406 not R2099_U24 ; R2099_U179
g7407 not R2099_U25 ; R2099_U180
g7408 not R2099_U136 ; R2099_U181
g7409 nand U4178 R2099_U99 ; R2099_U182
g7410 nand U2702 R2099_U4 ; R2099_U183
g7411 not R2099_U27 ; R2099_U184
g7412 nand U4178 R2099_U100 ; R2099_U185
g7413 nand U2710 R2099_U4 ; R2099_U186
g7414 not R2099_U32 ; R2099_U187
g7415 nand U4178 R2099_U101 ; R2099_U188
g7416 nand U2709 R2099_U4 ; R2099_U189
g7417 not R2099_U33 ; R2099_U190
g7418 nand U4178 R2099_U102 ; R2099_U191
g7419 nand U2708 R2099_U4 ; R2099_U192
g7420 not R2099_U35 ; R2099_U193
g7421 nand U4178 R2099_U103 ; R2099_U194
g7422 nand U2707 R2099_U4 ; R2099_U195
g7423 not R2099_U34 ; R2099_U196
g7424 nand U4178 R2099_U104 ; R2099_U197
g7425 nand U2706 R2099_U4 ; R2099_U198
g7426 not R2099_U30 ; R2099_U199
g7427 nand U4178 R2099_U105 ; R2099_U200
g7428 nand U2705 R2099_U4 ; R2099_U201
g7429 not R2099_U31 ; R2099_U202
g7430 nand U4178 R2099_U106 ; R2099_U203
g7431 nand U2704 R2099_U4 ; R2099_U204
g7432 not R2099_U28 ; R2099_U205
g7433 nand U4178 R2099_U107 ; R2099_U206
g7434 nand U2703 R2099_U4 ; R2099_U207
g7435 not R2099_U29 ; R2099_U208
g7436 nand U4178 R2099_U108 ; R2099_U209
g7437 nand U2701 R2099_U4 ; R2099_U210
g7438 not R2099_U26 ; R2099_U211
g7439 nand R2099_U160 R2099_U211 ; R2099_U212
g7440 nand R2099_U26 R2099_U109 ; R2099_U213
g7441 nand R2099_U184 R2099_U159 ; R2099_U214
g7442 nand R2099_U27 R2099_U9 ; R2099_U215
g7443 nand R2099_U158 R2099_U208 ; R2099_U216
g7444 nand R2099_U29 R2099_U110 ; R2099_U217
g7445 nand R2099_U205 R2099_U157 ; R2099_U218
g7446 nand R2099_U28 R2099_U8 ; R2099_U219
g7447 nand R2099_U156 R2099_U202 ; R2099_U220
g7448 nand R2099_U31 R2099_U111 ; R2099_U221
g7449 nand R2099_U199 R2099_U155 ; R2099_U222
g7450 nand R2099_U30 R2099_U7 ; R2099_U223
g7451 nand R2099_U154 R2099_U196 ; R2099_U224
g7452 nand R2099_U34 R2099_U112 ; R2099_U225
g7453 nand U4178 R2099_U113 ; R2099_U226
g7454 nand U2682 R2099_U4 ; R2099_U227
g7455 not R2099_U45 ; R2099_U228
g7456 nand U4178 R2099_U114 ; R2099_U229
g7457 nand U2683 R2099_U4 ; R2099_U230
g7458 not R2099_U46 ; R2099_U231
g7459 nand U4178 R2099_U115 ; R2099_U232
g7460 nand U2684 R2099_U4 ; R2099_U233
g7461 not R2099_U47 ; R2099_U234
g7462 nand U4178 R2099_U116 ; R2099_U235
g7463 nand U2685 R2099_U4 ; R2099_U236
g7464 not R2099_U48 ; R2099_U237
g7465 nand U4178 R2099_U117 ; R2099_U238
g7466 nand U2686 R2099_U4 ; R2099_U239
g7467 not R2099_U49 ; R2099_U240
g7468 nand U4178 R2099_U118 ; R2099_U241
g7469 nand U2687 R2099_U4 ; R2099_U242
g7470 not R2099_U50 ; R2099_U243
g7471 nand U4178 R2099_U119 ; R2099_U244
g7472 nand U2688 R2099_U4 ; R2099_U245
g7473 not R2099_U51 ; R2099_U246
g7474 nand U4178 R2099_U120 ; R2099_U247
g7475 nand U2689 R2099_U4 ; R2099_U248
g7476 not R2099_U52 ; R2099_U249
g7477 nand U4178 R2099_U121 ; R2099_U250
g7478 nand U2690 R2099_U4 ; R2099_U251
g7479 not R2099_U53 ; R2099_U252
g7480 nand U4178 R2099_U122 ; R2099_U253
g7481 nand U2691 R2099_U4 ; R2099_U254
g7482 not R2099_U54 ; R2099_U255
g7483 nand U4178 R2099_U123 ; R2099_U256
g7484 nand U2692 R2099_U4 ; R2099_U257
g7485 not R2099_U55 ; R2099_U258
g7486 nand U4178 R2099_U124 ; R2099_U259
g7487 nand U2700 R2099_U4 ; R2099_U260
g7488 not R2099_U62 ; R2099_U261
g7489 nand U4178 R2099_U125 ; R2099_U262
g7490 nand U2699 R2099_U4 ; R2099_U263
g7491 not R2099_U63 ; R2099_U264
g7492 nand U4178 R2099_U126 ; R2099_U265
g7493 nand U2698 R2099_U4 ; R2099_U266
g7494 not R2099_U60 ; R2099_U267
g7495 nand U4178 R2099_U127 ; R2099_U268
g7496 nand U2697 R2099_U4 ; R2099_U269
g7497 not R2099_U61 ; R2099_U270
g7498 nand U4178 R2099_U128 ; R2099_U271
g7499 nand U2696 R2099_U4 ; R2099_U272
g7500 not R2099_U58 ; R2099_U273
g7501 nand U4178 R2099_U129 ; R2099_U274
g7502 nand U2695 R2099_U4 ; R2099_U275
g7503 not R2099_U59 ; R2099_U276
g7504 nand U4178 R2099_U130 ; R2099_U277
g7505 nand U2694 R2099_U4 ; R2099_U278
g7506 not R2099_U56 ; R2099_U279
g7507 nand U4178 R2099_U131 ; R2099_U280
g7508 nand U2693 R2099_U4 ; R2099_U281
g7509 not R2099_U57 ; R2099_U282
g7510 nand U4178 R2099_U132 ; R2099_U283
g7511 nand U2680 R2099_U4 ; R2099_U284
g7512 not R2099_U43 ; R2099_U285
g7513 nand U4178 R2099_U133 ; R2099_U286
g7514 nand U2681 R2099_U4 ; R2099_U287
g7515 not R2099_U44 ; R2099_U288
g7516 nand U4178 R2099_U134 ; R2099_U289
g7517 nand U2679 R2099_U4 ; R2099_U290
g7518 not R2099_U97 ; R2099_U291
g7519 nand R2099_U145 R2099_U291 ; R2099_U292
g7520 nand R2099_U97 R2099_U135 ; R2099_U293
g7521 nand R2099_U181 R2099_U285 ; R2099_U294
g7522 nand R2099_U43 R2099_U136 ; R2099_U295
g7523 nand R2099_U153 R2099_U193 ; R2099_U296
g7524 nand R2099_U35 R2099_U137 ; R2099_U297
g7525 nand R2099_U288 R2099_U180 ; R2099_U298
g7526 nand R2099_U44 R2099_U25 ; R2099_U299
g7527 nand R2099_U228 R2099_U179 ; R2099_U300
g7528 nand R2099_U45 R2099_U24 ; R2099_U301
g7529 nand R2099_U231 R2099_U178 ; R2099_U302
g7530 nand R2099_U46 R2099_U23 ; R2099_U303
g7531 nand R2099_U234 R2099_U177 ; R2099_U304
g7532 nand R2099_U47 R2099_U22 ; R2099_U305
g7533 nand R2099_U237 R2099_U176 ; R2099_U306
g7534 nand R2099_U48 R2099_U21 ; R2099_U307
g7535 nand R2099_U240 R2099_U175 ; R2099_U308
g7536 nand R2099_U49 R2099_U20 ; R2099_U309
g7537 nand R2099_U243 R2099_U174 ; R2099_U310
g7538 nand R2099_U50 R2099_U19 ; R2099_U311
g7539 nand R2099_U246 R2099_U173 ; R2099_U312
g7540 nand R2099_U51 R2099_U18 ; R2099_U313
g7541 nand R2099_U249 R2099_U172 ; R2099_U314
g7542 nand R2099_U52 R2099_U17 ; R2099_U315
g7543 nand R2099_U252 R2099_U171 ; R2099_U316
g7544 nand R2099_U53 R2099_U16 ; R2099_U317
g7545 nand R2099_U190 U2678 ; R2099_U318
g7546 nand R2099_U33 R2099_U6 ; R2099_U319
g7547 nand R2099_U190 U2678 ; R2099_U320
g7548 nand R2099_U33 R2099_U6 ; R2099_U321
g7549 nand R2099_U321 R2099_U320 ; R2099_U322
g7550 nand R2099_U139 R2099_U140 ; R2099_U323
g7551 nand R2099_U149 R2099_U322 ; R2099_U324
g7552 nand R2099_U255 R2099_U170 ; R2099_U325
g7553 nand R2099_U54 R2099_U15 ; R2099_U326
g7554 nand R2099_U258 R2099_U169 ; R2099_U327
g7555 nand R2099_U55 R2099_U14 ; R2099_U328
g7556 nand R2099_U168 R2099_U282 ; R2099_U329
g7557 nand R2099_U57 R2099_U141 ; R2099_U330
g7558 nand R2099_U279 R2099_U167 ; R2099_U331
g7559 nand R2099_U56 R2099_U13 ; R2099_U332
g7560 nand R2099_U166 R2099_U276 ; R2099_U333
g7561 nand R2099_U59 R2099_U142 ; R2099_U334
g7562 nand R2099_U273 R2099_U165 ; R2099_U335
g7563 nand R2099_U58 R2099_U12 ; R2099_U336
g7564 nand R2099_U164 R2099_U270 ; R2099_U337
g7565 nand R2099_U61 R2099_U143 ; R2099_U338
g7566 nand R2099_U267 R2099_U163 ; R2099_U339
g7567 nand R2099_U60 R2099_U11 ; R2099_U340
g7568 nand R2099_U162 R2099_U264 ; R2099_U341
g7569 nand R2099_U63 R2099_U144 ; R2099_U342
g7570 nand R2099_U261 R2099_U161 ; R2099_U343
g7571 nand R2099_U62 R2099_U10 ; R2099_U344
g7572 nand U4177 R2099_U4 ; R2099_U345
g7573 nand U4178 R2099_U5 ; R2099_U346
g7574 not R2099_U98 ; R2099_U347
g7575 nand R2099_U32 R2099_U347 ; R2099_U348
g7576 nand R2099_U98 R2099_U187 ; R2099_U349
g7577 not U2716 ; R2167_U6
g7578 not U2714 ; R2167_U7
g7579 not U2720 ; R2167_U8
g7580 not U2719 ; R2167_U9
g7581 not U2713 ; R2167_U10
g7582 not U2712 ; R2167_U11
g7583 not U2718 ; R2167_U12
g7584 not U2717 ; R2167_U13
g7585 not U2711 ; R2167_U14
g7586 not U2356 ; R2167_U15
g7587 not STATE2_REG_0__SCAN_IN ; R2167_U16
g7588 nand R2167_U50 R2167_U49 ; R2167_U17
g7589 and R2167_U29 R2167_U30 ; R2167_U18
g7590 and R2167_U32 R2167_U33 ; R2167_U19
g7591 and R2167_U35 R2167_U36 ; R2167_U20
g7592 and R2167_U38 R2167_U39 ; R2167_U21
g7593 not U2721 ; R2167_U22
g7594 not U2722 ; R2167_U23
g7595 nand U2715 R2167_U23 ; R2167_U24
g7596 nand U2715 R2167_U22 ; R2167_U25
g7597 or U2721 U2722 ; R2167_U26
g7598 nand U2714 R2167_U8 ; R2167_U27
g7599 nand R2167_U27 R2167_U26 R2167_U25 R2167_U24 ; R2167_U28
g7600 nand U2720 R2167_U7 ; R2167_U29
g7601 nand U2719 R2167_U10 ; R2167_U30
g7602 nand R2167_U18 R2167_U28 ; R2167_U31
g7603 nand U2713 R2167_U9 ; R2167_U32
g7604 nand U2712 R2167_U12 ; R2167_U33
g7605 nand R2167_U19 R2167_U31 ; R2167_U34
g7606 nand U2718 R2167_U11 ; R2167_U35
g7607 nand U2717 R2167_U14 ; R2167_U36
g7608 nand R2167_U20 R2167_U34 ; R2167_U37
g7609 nand U2711 R2167_U13 ; R2167_U38
g7610 nand U2356 R2167_U6 ; R2167_U39
g7611 nand R2167_U21 R2167_U37 ; R2167_U40
g7612 nand U2716 R2167_U15 ; R2167_U41
g7613 nand R2167_U40 R2167_U41 ; R2167_U42
g7614 nand U2716 R2167_U16 ; R2167_U43
g7615 nand R2167_U42 R2167_U6 ; R2167_U44
g7616 nand R2167_U44 R2167_U43 ; R2167_U45
g7617 nand R2167_U6 STATE2_REG_0__SCAN_IN ; R2167_U46
g7618 nand U2716 R2167_U42 ; R2167_U47
g7619 nand R2167_U47 R2167_U46 ; R2167_U48
g7620 nand R2167_U45 R2167_U15 ; R2167_U49
g7621 nand U2356 R2167_U48 ; R2167_U50
g7622 not U3220 ; SUB_357_U6
g7623 not U3215 ; SUB_357_U7
g7624 not U3221 ; SUB_357_U8
g7625 not U3219 ; SUB_357_U9
g7626 not U3214 ; SUB_357_U10
g7627 not U3217 ; SUB_357_U11
g7628 not U3216 ; SUB_357_U12
g7629 not U3218 ; SUB_357_U13
g7630 and LT_563_1260_U9 LT_563_1260_U8 ; LT_563_1260_U6
g7631 not U2673 ; LT_563_1260_U7
g7632 nand R584_U8 LT_563_1260_U7 ; LT_563_1260_U8
g7633 nand R584_U9 LT_563_1260_U7 ; LT_563_1260_U9
g7634 nand SUB_580_U10 SUB_580_U9 ; SUB_580_U6
g7635 not INSTADDRPOINTER_REG_1__SCAN_IN ; SUB_580_U7
g7636 not INSTADDRPOINTER_REG_0__SCAN_IN ; SUB_580_U8
g7637 nand SUB_580_U8 INSTADDRPOINTER_REG_1__SCAN_IN ; SUB_580_U9
g7638 nand SUB_580_U7 INSTADDRPOINTER_REG_0__SCAN_IN ; SUB_580_U10
g7639 not REIP_REG_1__SCAN_IN ; R2096_U4
g7640 not REIP_REG_2__SCAN_IN ; R2096_U5
g7641 nand REIP_REG_1__SCAN_IN REIP_REG_2__SCAN_IN ; R2096_U6
g7642 not REIP_REG_3__SCAN_IN ; R2096_U7
g7643 nand R2096_U94 REIP_REG_3__SCAN_IN ; R2096_U8
g7644 not REIP_REG_4__SCAN_IN ; R2096_U9
g7645 nand R2096_U95 REIP_REG_4__SCAN_IN ; R2096_U10
g7646 not REIP_REG_5__SCAN_IN ; R2096_U11
g7647 nand R2096_U96 REIP_REG_5__SCAN_IN ; R2096_U12
g7648 not REIP_REG_6__SCAN_IN ; R2096_U13
g7649 nand R2096_U97 REIP_REG_6__SCAN_IN ; R2096_U14
g7650 not REIP_REG_7__SCAN_IN ; R2096_U15
g7651 nand R2096_U98 REIP_REG_7__SCAN_IN ; R2096_U16
g7652 not REIP_REG_8__SCAN_IN ; R2096_U17
g7653 not REIP_REG_9__SCAN_IN ; R2096_U18
g7654 nand R2096_U99 REIP_REG_8__SCAN_IN ; R2096_U19
g7655 nand R2096_U100 REIP_REG_9__SCAN_IN ; R2096_U20
g7656 not REIP_REG_10__SCAN_IN ; R2096_U21
g7657 nand R2096_U101 REIP_REG_10__SCAN_IN ; R2096_U22
g7658 not REIP_REG_11__SCAN_IN ; R2096_U23
g7659 nand R2096_U102 REIP_REG_11__SCAN_IN ; R2096_U24
g7660 not REIP_REG_12__SCAN_IN ; R2096_U25
g7661 nand R2096_U103 REIP_REG_12__SCAN_IN ; R2096_U26
g7662 not REIP_REG_13__SCAN_IN ; R2096_U27
g7663 nand R2096_U104 REIP_REG_13__SCAN_IN ; R2096_U28
g7664 not REIP_REG_14__SCAN_IN ; R2096_U29
g7665 nand R2096_U105 REIP_REG_14__SCAN_IN ; R2096_U30
g7666 not REIP_REG_15__SCAN_IN ; R2096_U31
g7667 nand R2096_U106 REIP_REG_15__SCAN_IN ; R2096_U32
g7668 not REIP_REG_16__SCAN_IN ; R2096_U33
g7669 nand R2096_U107 REIP_REG_16__SCAN_IN ; R2096_U34
g7670 not REIP_REG_17__SCAN_IN ; R2096_U35
g7671 nand R2096_U108 REIP_REG_17__SCAN_IN ; R2096_U36
g7672 not REIP_REG_18__SCAN_IN ; R2096_U37
g7673 nand R2096_U109 REIP_REG_18__SCAN_IN ; R2096_U38
g7674 not REIP_REG_19__SCAN_IN ; R2096_U39
g7675 nand R2096_U110 REIP_REG_19__SCAN_IN ; R2096_U40
g7676 not REIP_REG_20__SCAN_IN ; R2096_U41
g7677 nand R2096_U111 REIP_REG_20__SCAN_IN ; R2096_U42
g7678 not REIP_REG_21__SCAN_IN ; R2096_U43
g7679 nand R2096_U112 REIP_REG_21__SCAN_IN ; R2096_U44
g7680 not REIP_REG_22__SCAN_IN ; R2096_U45
g7681 nand R2096_U113 REIP_REG_22__SCAN_IN ; R2096_U46
g7682 not REIP_REG_23__SCAN_IN ; R2096_U47
g7683 nand R2096_U114 REIP_REG_23__SCAN_IN ; R2096_U48
g7684 not REIP_REG_24__SCAN_IN ; R2096_U49
g7685 nand R2096_U115 REIP_REG_24__SCAN_IN ; R2096_U50
g7686 not REIP_REG_25__SCAN_IN ; R2096_U51
g7687 nand R2096_U116 REIP_REG_25__SCAN_IN ; R2096_U52
g7688 not REIP_REG_26__SCAN_IN ; R2096_U53
g7689 nand R2096_U117 REIP_REG_26__SCAN_IN ; R2096_U54
g7690 not REIP_REG_27__SCAN_IN ; R2096_U55
g7691 nand R2096_U118 REIP_REG_27__SCAN_IN ; R2096_U56
g7692 not REIP_REG_28__SCAN_IN ; R2096_U57
g7693 nand R2096_U119 REIP_REG_28__SCAN_IN ; R2096_U58
g7694 not REIP_REG_29__SCAN_IN ; R2096_U59
g7695 nand R2096_U120 REIP_REG_29__SCAN_IN ; R2096_U60
g7696 not REIP_REG_30__SCAN_IN ; R2096_U61
g7697 nand R2096_U124 R2096_U123 ; R2096_U62
g7698 nand R2096_U126 R2096_U125 ; R2096_U63
g7699 nand R2096_U128 R2096_U127 ; R2096_U64
g7700 nand R2096_U130 R2096_U129 ; R2096_U65
g7701 nand R2096_U132 R2096_U131 ; R2096_U66
g7702 nand R2096_U134 R2096_U133 ; R2096_U67
g7703 nand R2096_U136 R2096_U135 ; R2096_U68
g7704 nand R2096_U138 R2096_U137 ; R2096_U69
g7705 nand R2096_U140 R2096_U139 ; R2096_U70
g7706 nand R2096_U142 R2096_U141 ; R2096_U71
g7707 nand R2096_U144 R2096_U143 ; R2096_U72
g7708 nand R2096_U146 R2096_U145 ; R2096_U73
g7709 nand R2096_U148 R2096_U147 ; R2096_U74
g7710 nand R2096_U150 R2096_U149 ; R2096_U75
g7711 nand R2096_U152 R2096_U151 ; R2096_U76
g7712 nand R2096_U154 R2096_U153 ; R2096_U77
g7713 nand R2096_U156 R2096_U155 ; R2096_U78
g7714 nand R2096_U158 R2096_U157 ; R2096_U79
g7715 nand R2096_U160 R2096_U159 ; R2096_U80
g7716 nand R2096_U162 R2096_U161 ; R2096_U81
g7717 nand R2096_U164 R2096_U163 ; R2096_U82
g7718 nand R2096_U166 R2096_U165 ; R2096_U83
g7719 nand R2096_U168 R2096_U167 ; R2096_U84
g7720 nand R2096_U170 R2096_U169 ; R2096_U85
g7721 nand R2096_U172 R2096_U171 ; R2096_U86
g7722 nand R2096_U174 R2096_U173 ; R2096_U87
g7723 nand R2096_U176 R2096_U175 ; R2096_U88
g7724 nand R2096_U178 R2096_U177 ; R2096_U89
g7725 nand R2096_U180 R2096_U179 ; R2096_U90
g7726 nand R2096_U182 R2096_U181 ; R2096_U91
g7727 not REIP_REG_31__SCAN_IN ; R2096_U92
g7728 nand R2096_U121 REIP_REG_30__SCAN_IN ; R2096_U93
g7729 not R2096_U6 ; R2096_U94
g7730 not R2096_U8 ; R2096_U95
g7731 not R2096_U10 ; R2096_U96
g7732 not R2096_U12 ; R2096_U97
g7733 not R2096_U14 ; R2096_U98
g7734 not R2096_U16 ; R2096_U99
g7735 not R2096_U19 ; R2096_U100
g7736 not R2096_U20 ; R2096_U101
g7737 not R2096_U22 ; R2096_U102
g7738 not R2096_U24 ; R2096_U103
g7739 not R2096_U26 ; R2096_U104
g7740 not R2096_U28 ; R2096_U105
g7741 not R2096_U30 ; R2096_U106
g7742 not R2096_U32 ; R2096_U107
g7743 not R2096_U34 ; R2096_U108
g7744 not R2096_U36 ; R2096_U109
g7745 not R2096_U38 ; R2096_U110
g7746 not R2096_U40 ; R2096_U111
g7747 not R2096_U42 ; R2096_U112
g7748 not R2096_U44 ; R2096_U113
g7749 not R2096_U46 ; R2096_U114
g7750 not R2096_U48 ; R2096_U115
g7751 not R2096_U50 ; R2096_U116
g7752 not R2096_U52 ; R2096_U117
g7753 not R2096_U54 ; R2096_U118
g7754 not R2096_U56 ; R2096_U119
g7755 not R2096_U58 ; R2096_U120
g7756 not R2096_U60 ; R2096_U121
g7757 not R2096_U93 ; R2096_U122
g7758 nand R2096_U19 REIP_REG_9__SCAN_IN ; R2096_U123
g7759 nand R2096_U100 R2096_U18 ; R2096_U124
g7760 nand R2096_U16 REIP_REG_8__SCAN_IN ; R2096_U125
g7761 nand R2096_U99 R2096_U17 ; R2096_U126
g7762 nand R2096_U14 REIP_REG_7__SCAN_IN ; R2096_U127
g7763 nand R2096_U98 R2096_U15 ; R2096_U128
g7764 nand R2096_U12 REIP_REG_6__SCAN_IN ; R2096_U129
g7765 nand R2096_U97 R2096_U13 ; R2096_U130
g7766 nand R2096_U10 REIP_REG_5__SCAN_IN ; R2096_U131
g7767 nand R2096_U96 R2096_U11 ; R2096_U132
g7768 nand R2096_U8 REIP_REG_4__SCAN_IN ; R2096_U133
g7769 nand R2096_U95 R2096_U9 ; R2096_U134
g7770 nand R2096_U6 REIP_REG_3__SCAN_IN ; R2096_U135
g7771 nand R2096_U94 R2096_U7 ; R2096_U136
g7772 nand R2096_U93 REIP_REG_31__SCAN_IN ; R2096_U137
g7773 nand R2096_U122 R2096_U92 ; R2096_U138
g7774 nand R2096_U60 REIP_REG_30__SCAN_IN ; R2096_U139
g7775 nand R2096_U121 R2096_U61 ; R2096_U140
g7776 nand R2096_U4 REIP_REG_2__SCAN_IN ; R2096_U141
g7777 nand R2096_U5 REIP_REG_1__SCAN_IN ; R2096_U142
g7778 nand R2096_U58 REIP_REG_29__SCAN_IN ; R2096_U143
g7779 nand R2096_U120 R2096_U59 ; R2096_U144
g7780 nand R2096_U56 REIP_REG_28__SCAN_IN ; R2096_U145
g7781 nand R2096_U119 R2096_U57 ; R2096_U146
g7782 nand R2096_U54 REIP_REG_27__SCAN_IN ; R2096_U147
g7783 nand R2096_U118 R2096_U55 ; R2096_U148
g7784 nand R2096_U52 REIP_REG_26__SCAN_IN ; R2096_U149
g7785 nand R2096_U117 R2096_U53 ; R2096_U150
g7786 nand R2096_U50 REIP_REG_25__SCAN_IN ; R2096_U151
g7787 nand R2096_U116 R2096_U51 ; R2096_U152
g7788 nand R2096_U48 REIP_REG_24__SCAN_IN ; R2096_U153
g7789 nand R2096_U115 R2096_U49 ; R2096_U154
g7790 nand R2096_U46 REIP_REG_23__SCAN_IN ; R2096_U155
g7791 nand R2096_U114 R2096_U47 ; R2096_U156
g7792 nand R2096_U44 REIP_REG_22__SCAN_IN ; R2096_U157
g7793 nand R2096_U113 R2096_U45 ; R2096_U158
g7794 nand R2096_U42 REIP_REG_21__SCAN_IN ; R2096_U159
g7795 nand R2096_U112 R2096_U43 ; R2096_U160
g7796 nand R2096_U40 REIP_REG_20__SCAN_IN ; R2096_U161
g7797 nand R2096_U111 R2096_U41 ; R2096_U162
g7798 nand R2096_U38 REIP_REG_19__SCAN_IN ; R2096_U163
g7799 nand R2096_U110 R2096_U39 ; R2096_U164
g7800 nand R2096_U36 REIP_REG_18__SCAN_IN ; R2096_U165
g7801 nand R2096_U109 R2096_U37 ; R2096_U166
g7802 nand R2096_U34 REIP_REG_17__SCAN_IN ; R2096_U167
g7803 nand R2096_U108 R2096_U35 ; R2096_U168
g7804 nand R2096_U32 REIP_REG_16__SCAN_IN ; R2096_U169
g7805 nand R2096_U107 R2096_U33 ; R2096_U170
g7806 nand R2096_U30 REIP_REG_15__SCAN_IN ; R2096_U171
g7807 nand R2096_U106 R2096_U31 ; R2096_U172
g7808 nand R2096_U28 REIP_REG_14__SCAN_IN ; R2096_U173
g7809 nand R2096_U105 R2096_U29 ; R2096_U174
g7810 nand R2096_U26 REIP_REG_13__SCAN_IN ; R2096_U175
g7811 nand R2096_U104 R2096_U27 ; R2096_U176
g7812 nand R2096_U24 REIP_REG_12__SCAN_IN ; R2096_U177
g7813 nand R2096_U103 R2096_U25 ; R2096_U178
g7814 nand R2096_U22 REIP_REG_11__SCAN_IN ; R2096_U179
g7815 nand R2096_U102 R2096_U23 ; R2096_U180
g7816 nand R2096_U20 REIP_REG_10__SCAN_IN ; R2096_U181
g7817 nand R2096_U101 R2096_U21 ; R2096_U182
g7818 and LT_563_U27 LT_563_U26 ; LT_563_U6
g7819 not INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; LT_563_U7
g7820 not U3478 ; LT_563_U8
g7821 not U3477 ; LT_563_U9
g7822 not INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; LT_563_U10
g7823 not INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; LT_563_U11
g7824 not U3476 ; LT_563_U12
g7825 and LT_563_U21 LT_563_U22 ; LT_563_U13
g7826 and LT_563_U24 LT_563_U25 ; LT_563_U14
g7827 not U3479 ; LT_563_U15
g7828 not U3480 ; LT_563_U16
g7829 nand LT_563_U16 LT_563_U15 INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; LT_563_U17
g7830 nand LT_563_U15 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; LT_563_U18
g7831 nand LT_563_U8 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; LT_563_U19
g7832 nand LT_563_U28 LT_563_U19 LT_563_U18 LT_563_U17 ; LT_563_U20
g7833 nand U3478 LT_563_U7 ; LT_563_U21
g7834 nand U3477 LT_563_U10 ; LT_563_U22
g7835 nand LT_563_U13 LT_563_U20 ; LT_563_U23
g7836 nand LT_563_U9 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; LT_563_U24
g7837 nand LT_563_U12 INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; LT_563_U25
g7838 nand LT_563_U14 LT_563_U23 ; LT_563_U26
g7839 nand U3476 LT_563_U11 ; LT_563_U27
g7840 nand LT_563_U16 INSTQUEUEWR_ADDR_REG_1__SCAN_IN INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; LT_563_U28
g7841 nand R2238_U45 R2238_U44 ; R2238_U6
g7842 nand R2238_U9 R2238_U46 ; R2238_U7
g7843 not INSTQUEUERD_ADDR_REG_0__SCAN_IN ; R2238_U8
g7844 nand R2238_U18 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; R2238_U9
g7845 not INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; R2238_U10
g7846 not INSTQUEUERD_ADDR_REG_2__SCAN_IN ; R2238_U11
g7847 not INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; R2238_U12
g7848 not INSTQUEUERD_ADDR_REG_3__SCAN_IN ; R2238_U13
g7849 not INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; R2238_U14
g7850 not INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; R2238_U15
g7851 nand R2238_U41 R2238_U40 ; R2238_U16
g7852 not INSTQUEUERD_ADDR_REG_4__SCAN_IN ; R2238_U17
g7853 not INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; R2238_U18
g7854 nand R2238_U51 R2238_U50 ; R2238_U19
g7855 nand R2238_U56 R2238_U55 ; R2238_U20
g7856 nand R2238_U61 R2238_U60 ; R2238_U21
g7857 nand R2238_U66 R2238_U65 ; R2238_U22
g7858 nand R2238_U48 R2238_U47 ; R2238_U23
g7859 nand R2238_U53 R2238_U52 ; R2238_U24
g7860 nand R2238_U58 R2238_U57 ; R2238_U25
g7861 nand R2238_U63 R2238_U62 ; R2238_U26
g7862 nand R2238_U37 R2238_U36 ; R2238_U27
g7863 nand R2238_U33 R2238_U32 ; R2238_U28
g7864 not INSTQUEUERD_ADDR_REG_1__SCAN_IN ; R2238_U29
g7865 not R2238_U9 ; R2238_U30
g7866 nand R2238_U30 R2238_U10 ; R2238_U31
g7867 nand R2238_U31 R2238_U29 ; R2238_U32
g7868 nand R2238_U9 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; R2238_U33
g7869 not R2238_U28 ; R2238_U34
g7870 nand R2238_U12 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; R2238_U35
g7871 nand R2238_U35 R2238_U28 ; R2238_U36
g7872 nand R2238_U11 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; R2238_U37
g7873 not R2238_U27 ; R2238_U38
g7874 nand R2238_U14 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; R2238_U39
g7875 nand R2238_U39 R2238_U27 ; R2238_U40
g7876 nand R2238_U13 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; R2238_U41
g7877 not R2238_U16 ; R2238_U42
g7878 nand R2238_U17 INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; R2238_U43
g7879 nand R2238_U42 R2238_U43 ; R2238_U44
g7880 nand R2238_U15 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; R2238_U45
g7881 nand R2238_U8 INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; R2238_U46
g7882 nand R2238_U15 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; R2238_U47
g7883 nand R2238_U17 INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; R2238_U48
g7884 not R2238_U23 ; R2238_U49
g7885 nand R2238_U49 R2238_U42 ; R2238_U50
g7886 nand R2238_U23 R2238_U16 ; R2238_U51
g7887 nand R2238_U14 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; R2238_U52
g7888 nand R2238_U13 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; R2238_U53
g7889 not R2238_U24 ; R2238_U54
g7890 nand R2238_U38 R2238_U54 ; R2238_U55
g7891 nand R2238_U24 R2238_U27 ; R2238_U56
g7892 nand R2238_U12 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; R2238_U57
g7893 nand R2238_U11 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; R2238_U58
g7894 not R2238_U25 ; R2238_U59
g7895 nand R2238_U34 R2238_U59 ; R2238_U60
g7896 nand R2238_U25 R2238_U28 ; R2238_U61
g7897 nand R2238_U10 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; R2238_U62
g7898 nand R2238_U29 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; R2238_U63
g7899 not R2238_U26 ; R2238_U64
g7900 nand R2238_U64 R2238_U30 ; R2238_U65
g7901 nand R2238_U26 R2238_U9 ; R2238_U66
g7902 nand SUB_450_U45 SUB_450_U44 ; SUB_450_U6
g7903 nand SUB_450_U9 SUB_450_U46 ; SUB_450_U7
g7904 not INSTQUEUERD_ADDR_REG_0__SCAN_IN ; SUB_450_U8
g7905 nand SUB_450_U18 INSTQUEUERD_ADDR_REG_0__SCAN_IN ; SUB_450_U9
g7906 not INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; SUB_450_U10
g7907 not INSTQUEUERD_ADDR_REG_2__SCAN_IN ; SUB_450_U11
g7908 not INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; SUB_450_U12
g7909 not INSTQUEUERD_ADDR_REG_3__SCAN_IN ; SUB_450_U13
g7910 not INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; SUB_450_U14
g7911 not INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; SUB_450_U15
g7912 nand SUB_450_U41 SUB_450_U40 ; SUB_450_U16
g7913 not INSTQUEUERD_ADDR_REG_4__SCAN_IN ; SUB_450_U17
g7914 not INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; SUB_450_U18
g7915 nand SUB_450_U51 SUB_450_U50 ; SUB_450_U19
g7916 nand SUB_450_U56 SUB_450_U55 ; SUB_450_U20
g7917 nand SUB_450_U61 SUB_450_U60 ; SUB_450_U21
g7918 nand SUB_450_U66 SUB_450_U65 ; SUB_450_U22
g7919 nand SUB_450_U48 SUB_450_U47 ; SUB_450_U23
g7920 nand SUB_450_U53 SUB_450_U52 ; SUB_450_U24
g7921 nand SUB_450_U58 SUB_450_U57 ; SUB_450_U25
g7922 nand SUB_450_U63 SUB_450_U62 ; SUB_450_U26
g7923 nand SUB_450_U37 SUB_450_U36 ; SUB_450_U27
g7924 nand SUB_450_U33 SUB_450_U32 ; SUB_450_U28
g7925 not INSTQUEUERD_ADDR_REG_1__SCAN_IN ; SUB_450_U29
g7926 not SUB_450_U9 ; SUB_450_U30
g7927 nand SUB_450_U30 SUB_450_U10 ; SUB_450_U31
g7928 nand SUB_450_U31 SUB_450_U29 ; SUB_450_U32
g7929 nand SUB_450_U9 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; SUB_450_U33
g7930 not SUB_450_U28 ; SUB_450_U34
g7931 nand SUB_450_U12 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; SUB_450_U35
g7932 nand SUB_450_U35 SUB_450_U28 ; SUB_450_U36
g7933 nand SUB_450_U11 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; SUB_450_U37
g7934 not SUB_450_U27 ; SUB_450_U38
g7935 nand SUB_450_U14 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; SUB_450_U39
g7936 nand SUB_450_U39 SUB_450_U27 ; SUB_450_U40
g7937 nand SUB_450_U13 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; SUB_450_U41
g7938 not SUB_450_U16 ; SUB_450_U42
g7939 nand SUB_450_U17 INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; SUB_450_U43
g7940 nand SUB_450_U42 SUB_450_U43 ; SUB_450_U44
g7941 nand SUB_450_U15 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; SUB_450_U45
g7942 nand SUB_450_U8 INSTQUEUEWR_ADDR_REG_0__SCAN_IN ; SUB_450_U46
g7943 nand SUB_450_U15 INSTQUEUERD_ADDR_REG_4__SCAN_IN ; SUB_450_U47
g7944 nand SUB_450_U17 INSTQUEUEWR_ADDR_REG_4__SCAN_IN ; SUB_450_U48
g7945 not SUB_450_U23 ; SUB_450_U49
g7946 nand SUB_450_U49 SUB_450_U42 ; SUB_450_U50
g7947 nand SUB_450_U23 SUB_450_U16 ; SUB_450_U51
g7948 nand SUB_450_U14 INSTQUEUERD_ADDR_REG_3__SCAN_IN ; SUB_450_U52
g7949 nand SUB_450_U13 INSTQUEUEWR_ADDR_REG_3__SCAN_IN ; SUB_450_U53
g7950 not SUB_450_U24 ; SUB_450_U54
g7951 nand SUB_450_U38 SUB_450_U54 ; SUB_450_U55
g7952 nand SUB_450_U24 SUB_450_U27 ; SUB_450_U56
g7953 nand SUB_450_U12 INSTQUEUERD_ADDR_REG_2__SCAN_IN ; SUB_450_U57
g7954 nand SUB_450_U11 INSTQUEUEWR_ADDR_REG_2__SCAN_IN ; SUB_450_U58
g7955 not SUB_450_U25 ; SUB_450_U59
g7956 nand SUB_450_U34 SUB_450_U59 ; SUB_450_U60
g7957 nand SUB_450_U25 SUB_450_U28 ; SUB_450_U61
g7958 nand SUB_450_U10 INSTQUEUERD_ADDR_REG_1__SCAN_IN ; SUB_450_U62
g7959 nand SUB_450_U29 INSTQUEUEWR_ADDR_REG_1__SCAN_IN ; SUB_450_U63
g7960 not SUB_450_U26 ; SUB_450_U64
g7961 nand SUB_450_U64 SUB_450_U30 ; SUB_450_U65
g7962 nand SUB_450_U26 SUB_450_U9 ; SUB_450_U66
g7963 not U3214 ; ADD_371_U4
g7964 nand ADD_371_U24 ADD_371_U32 ; ADD_371_U5
g7965 and ADD_371_U22 ADD_371_U30 ; ADD_371_U6
g7966 not U3215 ; ADD_371_U7
g7967 not U3217 ; ADD_371_U8
g7968 nand U3217 ADD_371_U24 ; ADD_371_U9
g7969 not U3218 ; ADD_371_U10
g7970 nand U3218 ADD_371_U28 ; ADD_371_U11
g7971 not U3219 ; ADD_371_U12
g7972 nand U3219 ADD_371_U29 ; ADD_371_U13
g7973 not U3221 ; ADD_371_U14
g7974 not U3220 ; ADD_371_U15
g7975 not U3216 ; ADD_371_U16
g7976 nand ADD_371_U34 ADD_371_U33 ; ADD_371_U17
g7977 nand ADD_371_U36 ADD_371_U35 ; ADD_371_U18
g7978 nand ADD_371_U38 ADD_371_U37 ; ADD_371_U19
g7979 nand ADD_371_U40 ADD_371_U39 ; ADD_371_U20
g7980 nand ADD_371_U44 ADD_371_U43 ; ADD_371_U21
g7981 and U3221 U3220 ; ADD_371_U22
g7982 nand U3220 ADD_371_U30 ; ADD_371_U23
g7983 nand ADD_371_U16 ADD_371_U26 ; ADD_371_U24
g7984 and ADD_371_U42 ADD_371_U41 ; ADD_371_U25
g7985 nand U3215 U3214 ; ADD_371_U26
g7986 not ADD_371_U24 ; ADD_371_U27
g7987 not ADD_371_U9 ; ADD_371_U28
g7988 not ADD_371_U11 ; ADD_371_U29
g7989 not ADD_371_U13 ; ADD_371_U30
g7990 not ADD_371_U23 ; ADD_371_U31
g7991 nand U3215 U3214 U3216 ; ADD_371_U32
g7992 nand U3221 ADD_371_U23 ; ADD_371_U33
g7993 nand ADD_371_U31 ADD_371_U14 ; ADD_371_U34
g7994 nand U3220 ADD_371_U13 ; ADD_371_U35
g7995 nand ADD_371_U30 ADD_371_U15 ; ADD_371_U36
g7996 nand U3219 ADD_371_U11 ; ADD_371_U37
g7997 nand ADD_371_U29 ADD_371_U12 ; ADD_371_U38
g7998 nand U3218 ADD_371_U9 ; ADD_371_U39
g7999 nand ADD_371_U28 ADD_371_U10 ; ADD_371_U40
g8000 nand U3217 ADD_371_U24 ; ADD_371_U41
g8001 nand ADD_371_U27 ADD_371_U8 ; ADD_371_U42
g8002 nand U3215 ADD_371_U4 ; ADD_371_U43
g8003 nand U3214 ADD_371_U7 ; ADD_371_U44
g8004 not INSTADDRPOINTER_REG_0__SCAN_IN ; ADD_405_U4
g8005 nand ADD_405_U92 ADD_405_U126 ; ADD_405_U5
g8006 not INSTADDRPOINTER_REG_1__SCAN_IN ; ADD_405_U6
g8007 not INSTADDRPOINTER_REG_3__SCAN_IN ; ADD_405_U7
g8008 nand ADD_405_U92 INSTADDRPOINTER_REG_3__SCAN_IN ; ADD_405_U8
g8009 not INSTADDRPOINTER_REG_4__SCAN_IN ; ADD_405_U9
g8010 nand ADD_405_U98 INSTADDRPOINTER_REG_4__SCAN_IN ; ADD_405_U10
g8011 not INSTADDRPOINTER_REG_5__SCAN_IN ; ADD_405_U11
g8012 nand ADD_405_U99 INSTADDRPOINTER_REG_5__SCAN_IN ; ADD_405_U12
g8013 not INSTADDRPOINTER_REG_6__SCAN_IN ; ADD_405_U13
g8014 nand ADD_405_U100 INSTADDRPOINTER_REG_6__SCAN_IN ; ADD_405_U14
g8015 not INSTADDRPOINTER_REG_7__SCAN_IN ; ADD_405_U15
g8016 nand ADD_405_U101 INSTADDRPOINTER_REG_7__SCAN_IN ; ADD_405_U16
g8017 not INSTADDRPOINTER_REG_8__SCAN_IN ; ADD_405_U17
g8018 not INSTADDRPOINTER_REG_9__SCAN_IN ; ADD_405_U18
g8019 nand ADD_405_U102 INSTADDRPOINTER_REG_8__SCAN_IN ; ADD_405_U19
g8020 nand ADD_405_U103 INSTADDRPOINTER_REG_9__SCAN_IN ; ADD_405_U20
g8021 not INSTADDRPOINTER_REG_10__SCAN_IN ; ADD_405_U21
g8022 nand ADD_405_U104 INSTADDRPOINTER_REG_10__SCAN_IN ; ADD_405_U22
g8023 not INSTADDRPOINTER_REG_11__SCAN_IN ; ADD_405_U23
g8024 nand ADD_405_U105 INSTADDRPOINTER_REG_11__SCAN_IN ; ADD_405_U24
g8025 not INSTADDRPOINTER_REG_12__SCAN_IN ; ADD_405_U25
g8026 nand ADD_405_U106 INSTADDRPOINTER_REG_12__SCAN_IN ; ADD_405_U26
g8027 not INSTADDRPOINTER_REG_13__SCAN_IN ; ADD_405_U27
g8028 nand ADD_405_U107 INSTADDRPOINTER_REG_13__SCAN_IN ; ADD_405_U28
g8029 not INSTADDRPOINTER_REG_14__SCAN_IN ; ADD_405_U29
g8030 nand ADD_405_U108 INSTADDRPOINTER_REG_14__SCAN_IN ; ADD_405_U30
g8031 not INSTADDRPOINTER_REG_15__SCAN_IN ; ADD_405_U31
g8032 nand ADD_405_U109 INSTADDRPOINTER_REG_15__SCAN_IN ; ADD_405_U32
g8033 not INSTADDRPOINTER_REG_16__SCAN_IN ; ADD_405_U33
g8034 nand ADD_405_U110 INSTADDRPOINTER_REG_16__SCAN_IN ; ADD_405_U34
g8035 not INSTADDRPOINTER_REG_17__SCAN_IN ; ADD_405_U35
g8036 nand ADD_405_U111 INSTADDRPOINTER_REG_17__SCAN_IN ; ADD_405_U36
g8037 not INSTADDRPOINTER_REG_18__SCAN_IN ; ADD_405_U37
g8038 nand ADD_405_U112 INSTADDRPOINTER_REG_18__SCAN_IN ; ADD_405_U38
g8039 not INSTADDRPOINTER_REG_19__SCAN_IN ; ADD_405_U39
g8040 nand ADD_405_U113 INSTADDRPOINTER_REG_19__SCAN_IN ; ADD_405_U40
g8041 not INSTADDRPOINTER_REG_20__SCAN_IN ; ADD_405_U41
g8042 nand ADD_405_U114 INSTADDRPOINTER_REG_20__SCAN_IN ; ADD_405_U42
g8043 not INSTADDRPOINTER_REG_21__SCAN_IN ; ADD_405_U43
g8044 nand ADD_405_U115 INSTADDRPOINTER_REG_21__SCAN_IN ; ADD_405_U44
g8045 not INSTADDRPOINTER_REG_22__SCAN_IN ; ADD_405_U45
g8046 nand ADD_405_U116 INSTADDRPOINTER_REG_22__SCAN_IN ; ADD_405_U46
g8047 not INSTADDRPOINTER_REG_23__SCAN_IN ; ADD_405_U47
g8048 nand ADD_405_U117 INSTADDRPOINTER_REG_23__SCAN_IN ; ADD_405_U48
g8049 not INSTADDRPOINTER_REG_24__SCAN_IN ; ADD_405_U49
g8050 nand ADD_405_U118 INSTADDRPOINTER_REG_24__SCAN_IN ; ADD_405_U50
g8051 not INSTADDRPOINTER_REG_25__SCAN_IN ; ADD_405_U51
g8052 nand ADD_405_U119 INSTADDRPOINTER_REG_25__SCAN_IN ; ADD_405_U52
g8053 not INSTADDRPOINTER_REG_26__SCAN_IN ; ADD_405_U53
g8054 nand ADD_405_U120 INSTADDRPOINTER_REG_26__SCAN_IN ; ADD_405_U54
g8055 not INSTADDRPOINTER_REG_27__SCAN_IN ; ADD_405_U55
g8056 nand ADD_405_U121 INSTADDRPOINTER_REG_27__SCAN_IN ; ADD_405_U56
g8057 not INSTADDRPOINTER_REG_28__SCAN_IN ; ADD_405_U57
g8058 nand ADD_405_U122 INSTADDRPOINTER_REG_28__SCAN_IN ; ADD_405_U58
g8059 not INSTADDRPOINTER_REG_29__SCAN_IN ; ADD_405_U59
g8060 nand ADD_405_U123 INSTADDRPOINTER_REG_29__SCAN_IN ; ADD_405_U60
g8061 not INSTADDRPOINTER_REG_30__SCAN_IN ; ADD_405_U61
g8062 not INSTADDRPOINTER_REG_2__SCAN_IN ; ADD_405_U62
g8063 nand ADD_405_U128 ADD_405_U127 ; ADD_405_U63
g8064 nand ADD_405_U130 ADD_405_U129 ; ADD_405_U64
g8065 nand ADD_405_U132 ADD_405_U131 ; ADD_405_U65
g8066 nand ADD_405_U134 ADD_405_U133 ; ADD_405_U66
g8067 nand ADD_405_U136 ADD_405_U135 ; ADD_405_U67
g8068 nand ADD_405_U138 ADD_405_U137 ; ADD_405_U68
g8069 nand ADD_405_U142 ADD_405_U141 ; ADD_405_U69
g8070 nand ADD_405_U144 ADD_405_U143 ; ADD_405_U70
g8071 nand ADD_405_U146 ADD_405_U145 ; ADD_405_U71
g8072 nand ADD_405_U148 ADD_405_U147 ; ADD_405_U72
g8073 nand ADD_405_U150 ADD_405_U149 ; ADD_405_U73
g8074 nand ADD_405_U152 ADD_405_U151 ; ADD_405_U74
g8075 nand ADD_405_U154 ADD_405_U153 ; ADD_405_U75
g8076 nand ADD_405_U156 ADD_405_U155 ; ADD_405_U76
g8077 nand ADD_405_U158 ADD_405_U157 ; ADD_405_U77
g8078 nand ADD_405_U160 ADD_405_U159 ; ADD_405_U78
g8079 nand ADD_405_U162 ADD_405_U161 ; ADD_405_U79
g8080 nand ADD_405_U164 ADD_405_U163 ; ADD_405_U80
g8081 nand ADD_405_U166 ADD_405_U165 ; ADD_405_U81
g8082 nand ADD_405_U168 ADD_405_U167 ; ADD_405_U82
g8083 nand ADD_405_U170 ADD_405_U169 ; ADD_405_U83
g8084 nand ADD_405_U172 ADD_405_U171 ; ADD_405_U84
g8085 nand ADD_405_U174 ADD_405_U173 ; ADD_405_U85
g8086 nand ADD_405_U176 ADD_405_U175 ; ADD_405_U86
g8087 nand ADD_405_U178 ADD_405_U177 ; ADD_405_U87
g8088 nand ADD_405_U180 ADD_405_U179 ; ADD_405_U88
g8089 nand ADD_405_U182 ADD_405_U181 ; ADD_405_U89
g8090 nand ADD_405_U184 ADD_405_U183 ; ADD_405_U90
g8091 nand ADD_405_U186 ADD_405_U185 ; ADD_405_U91
g8092 nand ADD_405_U62 ADD_405_U96 ; ADD_405_U92
g8093 and ADD_405_U140 ADD_405_U139 ; ADD_405_U93
g8094 not INSTADDRPOINTER_REG_31__SCAN_IN ; ADD_405_U94
g8095 nand ADD_405_U124 INSTADDRPOINTER_REG_30__SCAN_IN ; ADD_405_U95
g8096 nand INSTADDRPOINTER_REG_0__SCAN_IN INSTADDRPOINTER_REG_1__SCAN_IN ; ADD_405_U96
g8097 not ADD_405_U92 ; ADD_405_U97
g8098 not ADD_405_U8 ; ADD_405_U98
g8099 not ADD_405_U10 ; ADD_405_U99
g8100 not ADD_405_U12 ; ADD_405_U100
g8101 not ADD_405_U14 ; ADD_405_U101
g8102 not ADD_405_U16 ; ADD_405_U102
g8103 not ADD_405_U19 ; ADD_405_U103
g8104 not ADD_405_U20 ; ADD_405_U104
g8105 not ADD_405_U22 ; ADD_405_U105
g8106 not ADD_405_U24 ; ADD_405_U106
g8107 not ADD_405_U26 ; ADD_405_U107
g8108 not ADD_405_U28 ; ADD_405_U108
g8109 not ADD_405_U30 ; ADD_405_U109
g8110 not ADD_405_U32 ; ADD_405_U110
g8111 not ADD_405_U34 ; ADD_405_U111
g8112 not ADD_405_U36 ; ADD_405_U112
g8113 not ADD_405_U38 ; ADD_405_U113
g8114 not ADD_405_U40 ; ADD_405_U114
g8115 not ADD_405_U42 ; ADD_405_U115
g8116 not ADD_405_U44 ; ADD_405_U116
g8117 not ADD_405_U46 ; ADD_405_U117
g8118 not ADD_405_U48 ; ADD_405_U118
g8119 not ADD_405_U50 ; ADD_405_U119
g8120 not ADD_405_U52 ; ADD_405_U120
g8121 not ADD_405_U54 ; ADD_405_U121
g8122 not ADD_405_U56 ; ADD_405_U122
g8123 not ADD_405_U58 ; ADD_405_U123
g8124 not ADD_405_U60 ; ADD_405_U124
g8125 not ADD_405_U95 ; ADD_405_U125
g8126 nand INSTADDRPOINTER_REG_0__SCAN_IN INSTADDRPOINTER_REG_1__SCAN_IN INSTADDRPOINTER_REG_2__SCAN_IN ; ADD_405_U126
g8127 nand ADD_405_U19 INSTADDRPOINTER_REG_9__SCAN_IN ; ADD_405_U127
g8128 nand ADD_405_U103 ADD_405_U18 ; ADD_405_U128
g8129 nand ADD_405_U16 INSTADDRPOINTER_REG_8__SCAN_IN ; ADD_405_U129
g8130 nand ADD_405_U102 ADD_405_U17 ; ADD_405_U130
g8131 nand ADD_405_U14 INSTADDRPOINTER_REG_7__SCAN_IN ; ADD_405_U131
g8132 nand ADD_405_U101 ADD_405_U15 ; ADD_405_U132
g8133 nand ADD_405_U12 INSTADDRPOINTER_REG_6__SCAN_IN ; ADD_405_U133
g8134 nand ADD_405_U100 ADD_405_U13 ; ADD_405_U134
g8135 nand ADD_405_U10 INSTADDRPOINTER_REG_5__SCAN_IN ; ADD_405_U135
g8136 nand ADD_405_U99 ADD_405_U11 ; ADD_405_U136
g8137 nand ADD_405_U8 INSTADDRPOINTER_REG_4__SCAN_IN ; ADD_405_U137
g8138 nand ADD_405_U98 ADD_405_U9 ; ADD_405_U138
g8139 nand ADD_405_U92 INSTADDRPOINTER_REG_3__SCAN_IN ; ADD_405_U139
g8140 nand ADD_405_U97 ADD_405_U7 ; ADD_405_U140
g8141 nand ADD_405_U95 INSTADDRPOINTER_REG_31__SCAN_IN ; ADD_405_U141
g8142 nand ADD_405_U125 ADD_405_U94 ; ADD_405_U142
g8143 nand ADD_405_U60 INSTADDRPOINTER_REG_30__SCAN_IN ; ADD_405_U143
g8144 nand ADD_405_U124 ADD_405_U61 ; ADD_405_U144
g8145 nand ADD_405_U58 INSTADDRPOINTER_REG_29__SCAN_IN ; ADD_405_U145
g8146 nand ADD_405_U123 ADD_405_U59 ; ADD_405_U146
g8147 nand ADD_405_U56 INSTADDRPOINTER_REG_28__SCAN_IN ; ADD_405_U147
g8148 nand ADD_405_U122 ADD_405_U57 ; ADD_405_U148
g8149 nand ADD_405_U54 INSTADDRPOINTER_REG_27__SCAN_IN ; ADD_405_U149
g8150 nand ADD_405_U121 ADD_405_U55 ; ADD_405_U150
g8151 nand ADD_405_U52 INSTADDRPOINTER_REG_26__SCAN_IN ; ADD_405_U151
g8152 nand ADD_405_U120 ADD_405_U53 ; ADD_405_U152
g8153 nand ADD_405_U50 INSTADDRPOINTER_REG_25__SCAN_IN ; ADD_405_U153
g8154 nand ADD_405_U119 ADD_405_U51 ; ADD_405_U154
g8155 nand ADD_405_U48 INSTADDRPOINTER_REG_24__SCAN_IN ; ADD_405_U155
g8156 nand ADD_405_U118 ADD_405_U49 ; ADD_405_U156
g8157 nand ADD_405_U46 INSTADDRPOINTER_REG_23__SCAN_IN ; ADD_405_U157
g8158 nand ADD_405_U117 ADD_405_U47 ; ADD_405_U158
g8159 nand ADD_405_U44 INSTADDRPOINTER_REG_22__SCAN_IN ; ADD_405_U159
g8160 nand ADD_405_U116 ADD_405_U45 ; ADD_405_U160
g8161 nand ADD_405_U42 INSTADDRPOINTER_REG_21__SCAN_IN ; ADD_405_U161
g8162 nand ADD_405_U115 ADD_405_U43 ; ADD_405_U162
g8163 nand ADD_405_U40 INSTADDRPOINTER_REG_20__SCAN_IN ; ADD_405_U163
g8164 nand ADD_405_U114 ADD_405_U41 ; ADD_405_U164
g8165 nand ADD_405_U4 INSTADDRPOINTER_REG_1__SCAN_IN ; ADD_405_U165
g8166 nand ADD_405_U6 INSTADDRPOINTER_REG_0__SCAN_IN ; ADD_405_U166
g8167 nand ADD_405_U38 INSTADDRPOINTER_REG_19__SCAN_IN ; ADD_405_U167
g8168 nand ADD_405_U113 ADD_405_U39 ; ADD_405_U168
g8169 nand ADD_405_U36 INSTADDRPOINTER_REG_18__SCAN_IN ; ADD_405_U169
g8170 nand ADD_405_U112 ADD_405_U37 ; ADD_405_U170
g8171 nand ADD_405_U34 INSTADDRPOINTER_REG_17__SCAN_IN ; ADD_405_U171
g8172 nand ADD_405_U111 ADD_405_U35 ; ADD_405_U172
g8173 nand ADD_405_U32 INSTADDRPOINTER_REG_16__SCAN_IN ; ADD_405_U173
g8174 nand ADD_405_U110 ADD_405_U33 ; ADD_405_U174
g8175 nand ADD_405_U30 INSTADDRPOINTER_REG_15__SCAN_IN ; ADD_405_U175
g8176 nand ADD_405_U109 ADD_405_U31 ; ADD_405_U176
g8177 nand ADD_405_U28 INSTADDRPOINTER_REG_14__SCAN_IN ; ADD_405_U177
g8178 nand ADD_405_U108 ADD_405_U29 ; ADD_405_U178
g8179 nand ADD_405_U26 INSTADDRPOINTER_REG_13__SCAN_IN ; ADD_405_U179
g8180 nand ADD_405_U107 ADD_405_U27 ; ADD_405_U180
g8181 nand ADD_405_U24 INSTADDRPOINTER_REG_12__SCAN_IN ; ADD_405_U181
g8182 nand ADD_405_U106 ADD_405_U25 ; ADD_405_U182
g8183 nand ADD_405_U22 INSTADDRPOINTER_REG_11__SCAN_IN ; ADD_405_U183
g8184 nand ADD_405_U105 ADD_405_U23 ; ADD_405_U184
g8185 nand ADD_405_U20 INSTADDRPOINTER_REG_10__SCAN_IN ; ADD_405_U185
g8186 nand ADD_405_U104 ADD_405_U21 ; ADD_405_U186
g8187 nor R2238_U6 GTE_485_U7 ; GTE_485_U6
g8188 nor R2238_U19 R2238_U20 R2238_U22 R2238_U21 ; GTE_485_U7
g8189 not INSTADDRPOINTER_REG_1__SCAN_IN ; ADD_515_U4
g8190 not INSTADDRPOINTER_REG_2__SCAN_IN ; ADD_515_U5
g8191 nand INSTADDRPOINTER_REG_1__SCAN_IN INSTADDRPOINTER_REG_2__SCAN_IN ; ADD_515_U6
g8192 not INSTADDRPOINTER_REG_3__SCAN_IN ; ADD_515_U7
g8193 nand ADD_515_U94 INSTADDRPOINTER_REG_3__SCAN_IN ; ADD_515_U8
g8194 not INSTADDRPOINTER_REG_4__SCAN_IN ; ADD_515_U9
g8195 nand ADD_515_U95 INSTADDRPOINTER_REG_4__SCAN_IN ; ADD_515_U10
g8196 not INSTADDRPOINTER_REG_5__SCAN_IN ; ADD_515_U11
g8197 nand ADD_515_U96 INSTADDRPOINTER_REG_5__SCAN_IN ; ADD_515_U12
g8198 not INSTADDRPOINTER_REG_6__SCAN_IN ; ADD_515_U13
g8199 nand ADD_515_U97 INSTADDRPOINTER_REG_6__SCAN_IN ; ADD_515_U14
g8200 not INSTADDRPOINTER_REG_7__SCAN_IN ; ADD_515_U15
g8201 nand ADD_515_U98 INSTADDRPOINTER_REG_7__SCAN_IN ; ADD_515_U16
g8202 not INSTADDRPOINTER_REG_8__SCAN_IN ; ADD_515_U17
g8203 not INSTADDRPOINTER_REG_9__SCAN_IN ; ADD_515_U18
g8204 nand ADD_515_U99 INSTADDRPOINTER_REG_8__SCAN_IN ; ADD_515_U19
g8205 nand ADD_515_U100 INSTADDRPOINTER_REG_9__SCAN_IN ; ADD_515_U20
g8206 not INSTADDRPOINTER_REG_10__SCAN_IN ; ADD_515_U21
g8207 nand ADD_515_U101 INSTADDRPOINTER_REG_10__SCAN_IN ; ADD_515_U22
g8208 not INSTADDRPOINTER_REG_11__SCAN_IN ; ADD_515_U23
g8209 nand ADD_515_U102 INSTADDRPOINTER_REG_11__SCAN_IN ; ADD_515_U24
g8210 not INSTADDRPOINTER_REG_12__SCAN_IN ; ADD_515_U25
g8211 nand ADD_515_U103 INSTADDRPOINTER_REG_12__SCAN_IN ; ADD_515_U26
g8212 not INSTADDRPOINTER_REG_13__SCAN_IN ; ADD_515_U27
g8213 nand ADD_515_U104 INSTADDRPOINTER_REG_13__SCAN_IN ; ADD_515_U28
g8214 not INSTADDRPOINTER_REG_14__SCAN_IN ; ADD_515_U29
g8215 nand ADD_515_U105 INSTADDRPOINTER_REG_14__SCAN_IN ; ADD_515_U30
g8216 not INSTADDRPOINTER_REG_15__SCAN_IN ; ADD_515_U31
g8217 nand ADD_515_U106 INSTADDRPOINTER_REG_15__SCAN_IN ; ADD_515_U32
g8218 not INSTADDRPOINTER_REG_16__SCAN_IN ; ADD_515_U33
g8219 nand ADD_515_U107 INSTADDRPOINTER_REG_16__SCAN_IN ; ADD_515_U34
g8220 not INSTADDRPOINTER_REG_17__SCAN_IN ; ADD_515_U35
g8221 nand ADD_515_U108 INSTADDRPOINTER_REG_17__SCAN_IN ; ADD_515_U36
g8222 not INSTADDRPOINTER_REG_18__SCAN_IN ; ADD_515_U37
g8223 nand ADD_515_U109 INSTADDRPOINTER_REG_18__SCAN_IN ; ADD_515_U38
g8224 not INSTADDRPOINTER_REG_19__SCAN_IN ; ADD_515_U39
g8225 nand ADD_515_U110 INSTADDRPOINTER_REG_19__SCAN_IN ; ADD_515_U40
g8226 not INSTADDRPOINTER_REG_20__SCAN_IN ; ADD_515_U41
g8227 nand ADD_515_U111 INSTADDRPOINTER_REG_20__SCAN_IN ; ADD_515_U42
g8228 not INSTADDRPOINTER_REG_21__SCAN_IN ; ADD_515_U43
g8229 nand ADD_515_U112 INSTADDRPOINTER_REG_21__SCAN_IN ; ADD_515_U44
g8230 not INSTADDRPOINTER_REG_22__SCAN_IN ; ADD_515_U45
g8231 nand ADD_515_U113 INSTADDRPOINTER_REG_22__SCAN_IN ; ADD_515_U46
g8232 not INSTADDRPOINTER_REG_23__SCAN_IN ; ADD_515_U47
g8233 nand ADD_515_U114 INSTADDRPOINTER_REG_23__SCAN_IN ; ADD_515_U48
g8234 not INSTADDRPOINTER_REG_24__SCAN_IN ; ADD_515_U49
g8235 nand ADD_515_U115 INSTADDRPOINTER_REG_24__SCAN_IN ; ADD_515_U50
g8236 not INSTADDRPOINTER_REG_25__SCAN_IN ; ADD_515_U51
g8237 nand ADD_515_U116 INSTADDRPOINTER_REG_25__SCAN_IN ; ADD_515_U52
g8238 not INSTADDRPOINTER_REG_26__SCAN_IN ; ADD_515_U53
g8239 nand ADD_515_U117 INSTADDRPOINTER_REG_26__SCAN_IN ; ADD_515_U54
g8240 not INSTADDRPOINTER_REG_27__SCAN_IN ; ADD_515_U55
g8241 nand ADD_515_U118 INSTADDRPOINTER_REG_27__SCAN_IN ; ADD_515_U56
g8242 not INSTADDRPOINTER_REG_28__SCAN_IN ; ADD_515_U57
g8243 nand ADD_515_U119 INSTADDRPOINTER_REG_28__SCAN_IN ; ADD_515_U58
g8244 not INSTADDRPOINTER_REG_29__SCAN_IN ; ADD_515_U59
g8245 nand ADD_515_U120 INSTADDRPOINTER_REG_29__SCAN_IN ; ADD_515_U60
g8246 not INSTADDRPOINTER_REG_30__SCAN_IN ; ADD_515_U61
g8247 nand ADD_515_U124 ADD_515_U123 ; ADD_515_U62
g8248 nand ADD_515_U126 ADD_515_U125 ; ADD_515_U63
g8249 nand ADD_515_U128 ADD_515_U127 ; ADD_515_U64
g8250 nand ADD_515_U130 ADD_515_U129 ; ADD_515_U65
g8251 nand ADD_515_U132 ADD_515_U131 ; ADD_515_U66
g8252 nand ADD_515_U134 ADD_515_U133 ; ADD_515_U67
g8253 nand ADD_515_U136 ADD_515_U135 ; ADD_515_U68
g8254 nand ADD_515_U138 ADD_515_U137 ; ADD_515_U69
g8255 nand ADD_515_U140 ADD_515_U139 ; ADD_515_U70
g8256 nand ADD_515_U142 ADD_515_U141 ; ADD_515_U71
g8257 nand ADD_515_U144 ADD_515_U143 ; ADD_515_U72
g8258 nand ADD_515_U146 ADD_515_U145 ; ADD_515_U73
g8259 nand ADD_515_U148 ADD_515_U147 ; ADD_515_U74
g8260 nand ADD_515_U150 ADD_515_U149 ; ADD_515_U75
g8261 nand ADD_515_U152 ADD_515_U151 ; ADD_515_U76
g8262 nand ADD_515_U154 ADD_515_U153 ; ADD_515_U77
g8263 nand ADD_515_U156 ADD_515_U155 ; ADD_515_U78
g8264 nand ADD_515_U158 ADD_515_U157 ; ADD_515_U79
g8265 nand ADD_515_U160 ADD_515_U159 ; ADD_515_U80
g8266 nand ADD_515_U162 ADD_515_U161 ; ADD_515_U81
g8267 nand ADD_515_U164 ADD_515_U163 ; ADD_515_U82
g8268 nand ADD_515_U166 ADD_515_U165 ; ADD_515_U83
g8269 nand ADD_515_U168 ADD_515_U167 ; ADD_515_U84
g8270 nand ADD_515_U170 ADD_515_U169 ; ADD_515_U85
g8271 nand ADD_515_U172 ADD_515_U171 ; ADD_515_U86
g8272 nand ADD_515_U174 ADD_515_U173 ; ADD_515_U87
g8273 nand ADD_515_U176 ADD_515_U175 ; ADD_515_U88
g8274 nand ADD_515_U178 ADD_515_U177 ; ADD_515_U89
g8275 nand ADD_515_U180 ADD_515_U179 ; ADD_515_U90
g8276 nand ADD_515_U182 ADD_515_U181 ; ADD_515_U91
g8277 not INSTADDRPOINTER_REG_31__SCAN_IN ; ADD_515_U92
g8278 nand ADD_515_U121 INSTADDRPOINTER_REG_30__SCAN_IN ; ADD_515_U93
g8279 not ADD_515_U6 ; ADD_515_U94
g8280 not ADD_515_U8 ; ADD_515_U95
g8281 not ADD_515_U10 ; ADD_515_U96
g8282 not ADD_515_U12 ; ADD_515_U97
g8283 not ADD_515_U14 ; ADD_515_U98
g8284 not ADD_515_U16 ; ADD_515_U99
g8285 not ADD_515_U19 ; ADD_515_U100
g8286 not ADD_515_U20 ; ADD_515_U101
g8287 not ADD_515_U22 ; ADD_515_U102
g8288 not ADD_515_U24 ; ADD_515_U103
g8289 not ADD_515_U26 ; ADD_515_U104
g8290 not ADD_515_U28 ; ADD_515_U105
g8291 not ADD_515_U30 ; ADD_515_U106
g8292 not ADD_515_U32 ; ADD_515_U107
g8293 not ADD_515_U34 ; ADD_515_U108
g8294 not ADD_515_U36 ; ADD_515_U109
g8295 not ADD_515_U38 ; ADD_515_U110
g8296 not ADD_515_U40 ; ADD_515_U111
g8297 not ADD_515_U42 ; ADD_515_U112
g8298 not ADD_515_U44 ; ADD_515_U113
g8299 not ADD_515_U46 ; ADD_515_U114
g8300 not ADD_515_U48 ; ADD_515_U115
g8301 not ADD_515_U50 ; ADD_515_U116
g8302 not ADD_515_U52 ; ADD_515_U117
g8303 not ADD_515_U54 ; ADD_515_U118
g8304 not ADD_515_U56 ; ADD_515_U119
g8305 not ADD_515_U58 ; ADD_515_U120
g8306 not ADD_515_U60 ; ADD_515_U121
g8307 not ADD_515_U93 ; ADD_515_U122
g8308 nand ADD_515_U19 INSTADDRPOINTER_REG_9__SCAN_IN ; ADD_515_U123
g8309 nand ADD_515_U100 ADD_515_U18 ; ADD_515_U124
g8310 nand ADD_515_U16 INSTADDRPOINTER_REG_8__SCAN_IN ; ADD_515_U125
g8311 nand ADD_515_U99 ADD_515_U17 ; ADD_515_U126
g8312 nand ADD_515_U14 INSTADDRPOINTER_REG_7__SCAN_IN ; ADD_515_U127
g8313 nand ADD_515_U98 ADD_515_U15 ; ADD_515_U128
g8314 nand ADD_515_U12 INSTADDRPOINTER_REG_6__SCAN_IN ; ADD_515_U129
g8315 nand ADD_515_U97 ADD_515_U13 ; ADD_515_U130
g8316 nand ADD_515_U10 INSTADDRPOINTER_REG_5__SCAN_IN ; ADD_515_U131
g8317 nand ADD_515_U96 ADD_515_U11 ; ADD_515_U132
g8318 nand ADD_515_U8 INSTADDRPOINTER_REG_4__SCAN_IN ; ADD_515_U133
g8319 nand ADD_515_U95 ADD_515_U9 ; ADD_515_U134
g8320 nand ADD_515_U6 INSTADDRPOINTER_REG_3__SCAN_IN ; ADD_515_U135
g8321 nand ADD_515_U94 ADD_515_U7 ; ADD_515_U136
g8322 nand ADD_515_U93 INSTADDRPOINTER_REG_31__SCAN_IN ; ADD_515_U137
g8323 nand ADD_515_U122 ADD_515_U92 ; ADD_515_U138
g8324 nand ADD_515_U60 INSTADDRPOINTER_REG_30__SCAN_IN ; ADD_515_U139
g8325 nand ADD_515_U121 ADD_515_U61 ; ADD_515_U140
g8326 nand ADD_515_U4 INSTADDRPOINTER_REG_2__SCAN_IN ; ADD_515_U141
g8327 nand ADD_515_U5 INSTADDRPOINTER_REG_1__SCAN_IN ; ADD_515_U142
g8328 nand ADD_515_U58 INSTADDRPOINTER_REG_29__SCAN_IN ; ADD_515_U143
g8329 nand ADD_515_U120 ADD_515_U59 ; ADD_515_U144
g8330 nand ADD_515_U56 INSTADDRPOINTER_REG_28__SCAN_IN ; ADD_515_U145
g8331 nand ADD_515_U119 ADD_515_U57 ; ADD_515_U146
g8332 nand ADD_515_U54 INSTADDRPOINTER_REG_27__SCAN_IN ; ADD_515_U147
g8333 nand ADD_515_U118 ADD_515_U55 ; ADD_515_U148
g8334 nand ADD_515_U52 INSTADDRPOINTER_REG_26__SCAN_IN ; ADD_515_U149
g8335 nand ADD_515_U117 ADD_515_U53 ; ADD_515_U150
g8336 nand ADD_515_U50 INSTADDRPOINTER_REG_25__SCAN_IN ; ADD_515_U151
g8337 nand ADD_515_U116 ADD_515_U51 ; ADD_515_U152
g8338 nand ADD_515_U48 INSTADDRPOINTER_REG_24__SCAN_IN ; ADD_515_U153
g8339 nand ADD_515_U115 ADD_515_U49 ; ADD_515_U154
g8340 nand ADD_515_U46 INSTADDRPOINTER_REG_23__SCAN_IN ; ADD_515_U155
g8341 nand ADD_515_U114 ADD_515_U47 ; ADD_515_U156
g8342 nand ADD_515_U44 INSTADDRPOINTER_REG_22__SCAN_IN ; ADD_515_U157
g8343 nand ADD_515_U113 ADD_515_U45 ; ADD_515_U158
g8344 nand ADD_515_U42 INSTADDRPOINTER_REG_21__SCAN_IN ; ADD_515_U159
g8345 nand ADD_515_U112 ADD_515_U43 ; ADD_515_U160
g8346 nand ADD_515_U40 INSTADDRPOINTER_REG_20__SCAN_IN ; ADD_515_U161
g8347 nand ADD_515_U111 ADD_515_U41 ; ADD_515_U162
g8348 nand ADD_515_U38 INSTADDRPOINTER_REG_19__SCAN_IN ; ADD_515_U163
g8349 nand ADD_515_U110 ADD_515_U39 ; ADD_515_U164
g8350 nand ADD_515_U36 INSTADDRPOINTER_REG_18__SCAN_IN ; ADD_515_U165
g8351 nand ADD_515_U109 ADD_515_U37 ; ADD_515_U166
g8352 nand ADD_515_U34 INSTADDRPOINTER_REG_17__SCAN_IN ; ADD_515_U167
g8353 nand ADD_515_U108 ADD_515_U35 ; ADD_515_U168
g8354 nand ADD_515_U32 INSTADDRPOINTER_REG_16__SCAN_IN ; ADD_515_U169
g8355 nand ADD_515_U107 ADD_515_U33 ; ADD_515_U170
g8356 nand ADD_515_U30 INSTADDRPOINTER_REG_15__SCAN_IN ; ADD_515_U171
g8357 nand ADD_515_U106 ADD_515_U31 ; ADD_515_U172
g8358 nand ADD_515_U28 INSTADDRPOINTER_REG_14__SCAN_IN ; ADD_515_U173
g8359 nand ADD_515_U105 ADD_515_U29 ; ADD_515_U174
g8360 nand ADD_515_U26 INSTADDRPOINTER_REG_13__SCAN_IN ; ADD_515_U175
g8361 nand ADD_515_U104 ADD_515_U27 ; ADD_515_U176
g8362 nand ADD_515_U24 INSTADDRPOINTER_REG_12__SCAN_IN ; ADD_515_U177
g8363 nand ADD_515_U103 ADD_515_U25 ; ADD_515_U178
g8364 nand ADD_515_U22 INSTADDRPOINTER_REG_11__SCAN_IN ; ADD_515_U179
g8365 nand ADD_515_U102 ADD_515_U23 ; ADD_515_U180
g8366 nand ADD_515_U20 INSTADDRPOINTER_REG_10__SCAN_IN ; ADD_515_U181
g8367 nand ADD_515_U101 ADD_515_U21 ; ADD_515_U182
