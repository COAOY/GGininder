name C1908.iscas
i 101(0)
i 104(1)
i 107(2)
i 110(3)
i 113(4)
i 116(5)
i 119(6)
i 122(7)
i 125(8)
i 128(9)
i 131(10)
i 134(11)
i 137(12)
i 140(13)
i 143(14)
i 146(15)
i 210(16)
i 214(17)
i 217(18)
i 221(19)
i 224(20)
i 227(21)
i 234(22)
i 237(23)
i 469(24)
i 472(25)
i 475(26)
i 478(27)
i 898(28)
i 900(29)
i 902(30)
i 952(31)
i 953(32)

o 3(865)
o 6(864)
o 9(863)
o 12(862)
o 30(856)
o 45(851)
o 48(850)
o 15(861)
o 18(860)
o 21(859)
o 24(858)
o 27(857)
o 33(855)
o 36(854)
o 39(853)
o 42(852)
o 75(866)
o 51(899)
o 54(900)
o 60(901)
o 63(902)
o 66(903)
o 69(908)
o 72(909)
o 57(912)

g1 and 953(32) ; 949(33)
g2 and 953(32) ; 947(34)
g3 and 953(32) ; 943(35)
g4 and 953(32) ; 938(36)
g5 and 953(32) ; 934(37)
g6 and 953(32) ; 862(38)
g7 and 953(32) ; 859(39)
g8 and 952(31) ; 932(40)
g9 and 952(31) ; 930(41)
g10 and 952(31) ; 926(42)
g11 and 902(30) ; 922(43)
g12 and 902(30) ; 919(44)
g13 and 902(30) ; 918(45)
g14 and 902(30) ; 911(46)
g15 and 900(29) ; 909(47)
g16 and 898(28) ; 907(48)
g17 and 478(27) ; 553(49)
g18 and 475(26) ; 541(50)
g19 and 472(25) ; 529(51)
g20 and 469(24) ; 517(52)
g21 and 237(23) ; 244(53)
g22 and 237(23) ; 241(54)
g23 and 234(22) ; 248(55)
g24 and 234(22) ; 245(56)
g25 and 900(29) 227(21) ; 233(57)
g26 and 898(28) 224(20) ; 231(58)
g27 and 146(15) ; 206(59)
g28 and 146(15) ; 1626(60)
g29 and 143(14) ; 202(61)
g30 and 143(14) ; 1618(62)
g31 and 140(13) ; 198(63)
g32 and 140(13) ; 1610(64)
g33 and 137(12) ; 194(65)
g34 and 137(12) ; 1602(66)
g35 and 134(11) ; 191(67)
g36 and 134(11) ; 1594(68)
g37 and 131(10) ; 188(69)
g38 and 131(10) ; 1586(70)
g39 and 128(9) ; 184(71)
g40 and 128(9) ; 1578(72)
g41 and 125(8) ; 179(73)
g42 and 125(8) ; 1570(74)
g43 and 122(7) ; 175(75)
g44 and 122(7) ; 1562(76)
g45 and 119(6) ; 171(77)
g46 and 119(6) ; 1554(78)
g47 and 116(5) ; 168(79)
g48 and 116(5) ; 1546(80)
g49 and 113(4) ; 165(81)
g50 and 113(4) ; 1538(82)
g51 and 110(3) ; 160(83)
g52 and 110(3) ; 1530(84)
g53 and 107(2) ; 156(85)
g54 and 107(2) ; 1522(86)
g55 and 104(1) ; 153(87)
g56 and 104(1) ; 1514(88)
g57 and 101(0) ; 149(89)
g58 and 101(0) ; 1506(90)
g59 and 947(34) 930(41) ; 50(91)
g60 and 947(34) 930(41) ; 52(92)
g61 and 947(34) 930(41) ; 56(93)
g62 and 947(34) 930(41) ; 58(94)
g63 and 947(34) 930(41) ; 62(95)
g64 and 947(34) 930(41) ; 64(96)
g65 and 907(48) 943(35) ; 853(97)
g66 and 909(47) 943(35) ; 856(98)
g67 and 934(37) 231(58) ; 1634(99)
g68 and 934(37) 233(57) ; 1644(100)
g69 and 922(43) 248(55) ; 954(101)
g70 and 922(43) 244(53) ; 955(102)
g71 and 553(49) ; 1490(103)
g72 and 553(49) ; 1498(104)
g73 and 541(50) ; 1474(105)
g74 and 541(50) ; 1482(106)
g75 and 529(51) ; 1458(107)
g76 and 529(51) ; 1466(108)
g77 and 517(52) ; 1442(109)
g78 and 517(52) ; 1450(110)
g79 and 237(23) 248(55) ; 893(111)
g80 and 938(36) 227(21) ; 352(112)
g81 and 938(36) 224(20) ; 318(113)
g82 and 938(36) 245(56) 221(19) ; 1335(114)
g83 and 938(36) 245(56) 217(18) ; 1290(115)
g84 and 938(36) 241(54) 214(17) ; 1830(116)
g85 and 938(36) 241(54) 210(16) ; 369(117)
g86 and 206(59) ; 1713(118)
g87 and 206(59) ; 1721(119)
g88 and 206(59) ; 382(120)
g89 and 1626(60) ; 1632(121)
g90 and 202(61) ; 302(122)
g91 and 202(61) ; 1833(123)
g92 and 202(61) ; 1873(124)
g93 and 1618(62) ; 1624(125)
g94 and 198(63) ; 355(126)
g95 and 198(63) ; 1179(127)
g96 and 198(63) ; 385(128)
g97 and 1610(64) ; 1616(129)
g98 and 194(65) ; 1745(130)
g99 and 194(65) ; 1753(131)
g100 and 194(65) ; 1332(132)
g101 and 1602(66) ; 1608(133)
g102 and 191(67) ; 330(134)
g103 and 191(67) ; 1300(135)
g104 and 1594(68) ; 1600(136)
g105 and 188(69) ; 327(137)
g106 and 188(69) ; 1244(138)
g107 and 1586(70) ; 1592(139)
g108 and 184(71) ; 299(140)
g109 and 184(71) ; 1870(141)
g110 and 184(71) ; 1881(142)
g111 and 1578(72) ; 1584(143)
g112 and 179(73) ; 321(144)
g113 and 179(73) ; 1176(145)
g114 and 179(73) ; 1841(146)
g115 and 179(73) ; 1849(147)
g116 and 1570(74) ; 1576(148)
g117 and 175(75) ; 1053(149)
g118 and 175(75) ; 1817(150)
g119 and 175(75) ; 1857(151)
g120 and 1562(76) ; 1568(152)
g121 and 171(77) ; 1697(153)
g122 and 171(77) ; 1705(154)
g123 and 171(77) ; 1878(155)
g124 and 1554(78) ; 1560(156)
g125 and 168(79) ; 291(157)
g126 and 168(79) ; 1854(158)
g127 and 1546(80) ; 1552(159)
g128 and 165(81) ; 288(160)
g129 and 165(81) ; 1814(161)
g130 and 1538(82) ; 1544(162)
g131 and 160(83) ; 1050(163)
g132 and 160(83) ; 1785(164)
g133 and 160(83) ; 1793(165)
g134 and 160(83) ; 1312(166)
g135 and 1530(84) ; 1536(167)
g136 and 156(85) ; 1657(168)
g137 and 156(85) ; 1665(169)
g138 and 156(85) ; 1278(170)
g139 and 1522(86) ; 1528(171)
g140 and 153(87) ; 254(172)
g141 and 153(87) ; 1222(173)
g142 and 1514(88) ; 1520(174)
g143 and 149(89) ; 251(175)
g144 and 149(89) ; 1197(176)
g145 and 149(89) ; 1207(177)
g146 and 1506(90) ; 1512(178)
g147 and 893(111) 949(33) 926(42) ; 979(179)
g148 and 893(111) 949(33) 926(42) ; 978(180)
g149 and 893(111) 943(35) 919(44) 907(48) ; 956(181)
g150 and 893(111) 943(35) 919(44) 909(47) ; 967(182)
g151 and 1634(99) ; 1642(183)
g152 and 1644(100) ; 1652(184)
g153 and 1490(103) ; 1496(185)
g154 and 1498(104) ; 1504(186)
g155 and 1474(105) ; 1480(187)
g156 and 1482(106) ; 1488(188)
g157 and 1458(107) ; 1464(189)
g158 and 1466(108) ; 1472(190)
g159 and 1442(109) ; 1448(191)
g160 and 1450(110) ; 1456(192)
g161 and 352(112) ; 1154(193)
g162 and 352(112) ; 1166(194)
g163 and 318(113) ; 1078(195)
g164 and 318(113) ; 1090(196)
g165 and 954(101) 221(19) ; 487(197)
g166 and 1335(114) ; 1339(198)
g167 and 954(101) 217(18) ; 505(199)
g168 and 954(101) 217(18) ; 459(200)
g169 and 1290(115) ; 1298(201)
g170 and 955(102) 214(17) ; 482(202)
g171 and 1830(116) ; 1836(203)
g172 and 955(102) 210(16) ; 492(204)
g173 and 955(102) 210(16) ; 457(205)
g174 and 369(117) ; 1194(206)
g175 and 369(117) ; 1204(207)
g176 and 1713(118) ; 1717(208)
g177 and 1721(119) ; 1725(209)
g178 and 382(120) ; 1256(210)
g179 and 382(120) ; 1268(211)
g180 and 302(122) ; 1710(212)
g181 and 302(122) ; 1718(213)
g182 and 1833(123) ; 1837(214)
g183 and 1873(124) ; 1877(215)
g184 and 355(126) ; 1782(216)
g185 and 355(126) ; 1790(217)
g186 and 1179(127) ; 1183(218)
g187 and 385(128) ; 1838(219)
g188 and 385(128) ; 1846(220)
g189 and 1745(130) ; 1749(221)
g190 and 1753(131) ; 1757(222)
g191 and 1332(132) ; 1338(223)
g192 and 330(134) ; 1742(224)
g193 and 330(134) ; 1750(225)
g194 and 1300(135) ; 1308(226)
g195 and 327(137) ; 1100(227)
g196 and 327(137) ; 1112(228)
g197 and 1244(138) ; 1252(229)
g198 and 299(140) ; 1058(230)
g199 and 299(140) ; 1068(231)
g200 and 1870(141) ; 1876(232)
g201 and 1881(142) ; 1885(233)
g202 and 321(144) ; 1726(234)
g203 and 321(144) ; 1734(235)
g204 and 1176(145) ; 1182(236)
g205 and 1841(146) ; 1845(237)
g206 and 1849(147) ; 1853(238)
g207 and 1053(149) ; 1057(239)
g208 and 1817(150) ; 1821(240)
g209 and 1857(151) ; 1861(241)
g210 and 1697(153) ; 1701(242)
g211 and 1705(154) ; 1709(243)
g212 and 1878(155) ; 1884(244)
g213 and 291(157) ; 1694(245)
g214 and 291(157) ; 1702(246)
g215 and 1854(158) ; 1860(247)
g216 and 288(160) ; 1030(248)
g217 and 288(160) ; 1040(249)
g218 and 1814(161) ; 1820(250)
g219 and 1050(163) ; 1056(251)
g220 and 1785(164) ; 1789(252)
g221 and 1793(165) ; 1797(253)
g222 and 1312(166) ; 1320(254)
g223 and 1657(168) ; 1661(255)
g224 and 1665(169) ; 1669(256)
g225 and 1278(170) ; 1286(257)
g226 and 254(172) ; 1654(258)
g227 and 254(172) ; 1662(259)
g228 and 1222(173) ; 1230(260)
g229 and 251(175) ; 980(261)
g230 and 251(175) ; 990(262)
g231 and 1197(176) ; 1201(263)
g232 and 1207(177) ; 1211(264)
g233 and 978(180) 956(181) ; 958(265)
g234 and 978(180) 967(182) ; 969(266)
g235 and 1154(193) ; 1162(267)
g236 and 1166(194) ; 1174(268)
g237 and 1078(195) ; 1086(269)
g238 and 1090(196) ; 1098(270)
g239 and 487(197) ; 614(271)
g240 and 487(197) ; 615(272)
g241 and 1338(223) 1335(114) ; 404(273)
g242 and 505(199) ; 1426(274)
g243 and 505(199) ; 1434(275)
g244 and 482(202) ; 565(276)
g245 and 482(202) ; 566(277)
g246 and 1837(214) 1830(116) ; 1248(278)
g247 and 492(204) ; 1410(279)
g248 and 492(204) ; 1418(280)
g249 and 1194(206) ; 1200(281)
g250 and 1201(263) 1194(206) ; 1203(282)
g251 and 1211(264) 1204(207) ; 373(283)
g252 and 1204(207) ; 1210(284)
g253 and 1717(208) 1710(212) ; 1062(285)
g254 and 1725(209) 1718(213) ; 1072(286)
g255 and 1256(210) ; 1264(287)
g256 and 1268(211) ; 1276(288)
g257 and 1710(212) ; 1716(289)
g258 and 1718(213) ; 1724(290)
g259 and 1836(203) 1833(123) ; 1247(291)
g260 and 1876(232) 1873(124) ; 1303(292)
g261 and 1789(252) 1782(216) ; 1158(293)
g262 and 1782(216) ; 1788(294)
g263 and 1797(253) 1790(217) ; 1170(295)
g264 and 1790(217) ; 1796(296)
g265 and 1182(236) 1179(127) ; 361(297)
g266 and 1845(237) 1838(219) ; 1260(298)
g267 and 1838(219) ; 1844(299)
g268 and 1853(238) 1846(220) ; 1272(300)
g269 and 1846(220) ; 1852(301)
g270 and 1749(221) 1742(224) ; 1104(302)
g271 and 1757(222) 1750(225) ; 1116(303)
g272 and 1339(198) 1332(132) ; 405(304)
g273 and 1742(224) ; 1748(305)
g274 and 1750(225) ; 1756(306)
g275 and 1100(227) ; 1108(307)
g276 and 1112(228) ; 1120(308)
g277 and 1058(230) ; 1066(309)
g278 and 1068(231) ; 1076(310)
g279 and 1877(215) 1870(141) ; 1304(311)
g280 and 1884(244) 1881(142) ; 1315(312)
g281 and 1726(234) ; 1732(313)
g282 and 1734(235) ; 1740(314)
g283 and 1183(218) 1176(145) ; 362(315)
g284 and 1056(251) 1053(149) ; 297(316)
g285 and 1820(250) 1817(150) ; 1225(317)
g286 and 1860(247) 1857(151) ; 1281(318)
g287 and 1701(242) 1694(245) ; 1034(319)
g288 and 1709(243) 1702(246) ; 1044(320)
g289 and 1885(233) 1878(155) ; 1316(321)
g290 and 1694(245) ; 1700(322)
g291 and 1702(246) ; 1708(323)
g292 and 1861(241) 1854(158) ; 1282(324)
g293 and 1030(248) ; 1038(325)
g294 and 1040(249) ; 1048(326)
g295 and 1821(240) 1814(161) ; 1226(327)
g296 and 1057(239) 1050(163) ; 298(328)
g297 and 1661(255) 1654(258) ; 984(329)
g298 and 1669(256) 1662(259) ; 994(330)
g299 and 1654(258) ; 1660(331)
g300 and 1662(259) ; 1668(332)
g301 and 980(261) ; 988(333)
g302 and 990(262) ; 998(334)
g303 and 405(304) 404(273) ; 406(335)
g304 and 1426(274) ; 1432(336)
g305 and 1434(275) ; 1440(337)
g306 and 1248(278) 1247(291) ; 1249(338)
g307 and 1410(279) ; 1416(339)
g308 and 1418(280) ; 1424(340)
g309 and 1716(289) 1713(118) ; 1061(341)
g310 and 1724(290) 1721(119) ; 1071(342)
g311 and 1304(311) 1303(292) ; 1305(343)
g312 and 362(315) 361(297) ; 363(344)
g313 and 1748(305) 1745(130) ; 1103(345)
g314 and 1756(306) 1753(131) ; 1115(346)
g315 and 1316(321) 1315(312) ; 1317(347)
g316 and 1844(299) 1841(146) ; 1259(348)
g317 and 1852(301) 1849(147) ; 1271(349)
g318 and 298(328) 297(316) ; 268(350)
g319 and 1226(327) 1225(317) ; 1227(351)
g320 and 1282(324) 1281(318) ; 1283(352)
g321 and 1700(322) 1697(153) ; 1033(353)
g322 and 1708(323) 1705(154) ; 1043(354)
g323 and 1788(294) 1785(164) ; 1157(355)
g324 and 1796(296) 1793(165) ; 1169(356)
g325 and 1660(331) 1657(168) ; 983(357)
g326 and 1668(332) 1665(169) ; 993(358)
g327 and 1200(281) 1197(176) ; 1202(359)
g328 and 1210(284) 1207(177) ; 372(360)
g329 and 406(335) ; 1322(361)
g330 and 1249(338) ; 1253(362)
g331 and 1203(282) 1202(359) ; 1212(363)
g332 and 373(283) 372(360) ; 374(364)
g333 and 1062(285) 1061(341) ; 1063(365)
g334 and 1072(286) 1071(342) ; 1073(366)
g335 and 1305(343) ; 1309(367)
g336 and 1158(293) 1157(355) ; 1159(368)
g337 and 1170(295) 1169(356) ; 1171(369)
g338 and 363(344) ; 1184(370)
g339 and 1260(298) 1259(348) ; 1261(371)
g340 and 1272(300) 1271(349) ; 1273(372)
g341 and 1104(302) 1103(345) ; 1105(373)
g342 and 1116(303) 1115(346) ; 1117(374)
g343 and 1308(226) 1305(343) ; 1310(375)
g344 and 1252(229) 1249(338) ; 1254(376)
g345 and 1317(347) ; 1321(377)
g346 and 268(350) ; 269(378)
g347 and 1227(351) ; 1231(379)
g348 and 1283(352) ; 1287(380)
g349 and 1034(319) 1033(353) ; 1035(381)
g350 and 1044(320) 1043(354) ; 1045(382)
g351 and 1320(254) 1317(347) ; 396(383)
g352 and 984(329) 983(357) ; 985(384)
g353 and 994(330) 993(358) ; 995(385)
g354 and 1286(257) 1283(352) ; 1288(386)
g355 and 1230(260) 1227(351) ; 1232(387)
g356 and 1162(267) 1159(368) ; 1164(388)
g357 and 1174(268) 1171(369) ; 358(389)
g358 and 1322(361) ; 1330(390)
g359 and 1212(363) ; 1220(391)
g360 and 374(364) ; 1381(392)
g361 and 1063(365) ; 1067(393)
g362 and 1073(366) ; 1077(394)
g363 and 1264(287) 1261(371) ; 1266(395)
g364 and 1276(288) 1273(372) ; 388(396)
g365 and 1159(368) ; 1163(397)
g366 and 1171(369) ; 1175(398)
g367 and 1184(370) ; 1192(399)
g368 and 1261(371) ; 1265(400)
g369 and 1273(372) ; 1277(401)
g370 and 1105(373) ; 1109(402)
g371 and 1117(374) ; 1121(403)
g372 and 1309(367) 1300(135) ; 1311(404)
g373 and 1108(307) 1105(373) ; 1110(405)
g374 and 1120(308) 1117(374) ; 333(406)
g375 and 1253(362) 1244(138) ; 1255(407)
g376 and 1066(309) 1063(365) ; 308(408)
g377 and 1076(310) 1073(366) ; 305(409)
g378 and 269(378) ; 1000(410)
g379 and 269(378) ; 1010(411)
g380 and 1035(381) ; 1039(412)
g381 and 1045(382) ; 1049(413)
g382 and 1038(325) 1035(381) ; 272(414)
g383 and 1048(326) 1045(382) ; 294(415)
g384 and 1321(377) 1312(166) ; 397(416)
g385 and 985(384) ; 989(417)
g386 and 995(385) ; 999(418)
g387 and 1287(380) 1278(170) ; 1289(419)
g388 and 1231(379) 1222(173) ; 1233(420)
g389 and 988(333) 985(384) ; 260(421)
g390 and 998(334) 995(385) ; 257(422)
g391 and 1163(397) 1154(193) ; 1165(423)
g392 and 1175(398) 1166(194) ; 359(424)
g393 and 1381(392) ; 1385(425)
g394 and 1265(400) 1256(210) ; 1267(426)
g395 and 1277(401) 1268(211) ; 389(427)
g396 and 1311(404) 1310(375) ; 1862(428)
g397 and 1109(402) 1100(227) ; 1111(429)
g398 and 1121(403) 1112(228) ; 334(430)
g399 and 1255(407) 1254(376) ; 1822(431)
g400 and 1067(393) 1058(230) ; 309(432)
g401 and 1077(394) 1068(231) ; 306(433)
g402 and 1000(410) ; 1008(434)
g403 and 1010(411) ; 1018(435)
g404 and 1039(412) 1030(248) ; 273(436)
g405 and 1049(413) 1040(249) ; 295(437)
g406 and 397(416) 396(383) ; 398(438)
g407 and 1289(419) 1288(386) ; 1865(439)
g408 and 1233(420) 1232(387) ; 1234(440)
g409 and 989(417) 980(261) ; 261(441)
g410 and 999(418) 990(262) ; 258(442)
g411 and 1165(423) 1164(388) ; 1373(443)
g412 and 359(424) 358(389) ; 360(444)
g413 and 1267(426) 1266(395) ; 1825(445)
g414 and 389(427) 388(396) ; 390(446)
g415 and 1862(428) ; 1868(447)
g416 and 1111(429) 1110(405) ; 1798(448)
g417 and 334(430) 333(406) ; 335(449)
g418 and 1822(431) ; 1828(450)
g419 and 309(432) 308(408) ; 310(451)
g420 and 306(433) 305(409) ; 307(452)
g421 and 273(436) 272(414) ; 274(453)
g422 and 295(437) 294(415) ; 296(454)
g423 and 398(438) ; 1886(455)
g424 and 1865(439) ; 1869(456)
g425 and 1234(440) ; 1242(457)
g426 and 261(441) 260(421) ; 262(458)
g427 and 258(442) 257(422) ; 259(459)
g428 and 1373(443) ; 1377(460)
g429 and 360(444) ; 1777(461)
g430 and 1828(450) 1825(445) ; 1237(462)
g431 and 1825(445) ; 1829(463)
g432 and 390(446) ; 1889(464)
g433 and 1869(456) 1862(428) ; 1294(465)
g434 and 1798(448) ; 1804(466)
g435 and 335(449) ; 336(467)
g436 and 310(451) ; 1729(468)
g437 and 310(451) ; 1737(469)
g438 and 310(451) ; 410(470)
g439 and 307(452) ; 314(471)
g440 and 274(453) ; 1670(472)
g441 and 274(453) ; 1678(473)
g442 and 296(454) ; 407(474)
g443 and 1886(455) ; 1892(475)
g444 and 1868(447) 1865(439) ; 1293(476)
g445 and 262(458) ; 1761(477)
g446 and 262(458) ; 1769(478)
g447 and 259(459) ; 265(479)
g448 and 1777(461) ; 1781(480)
g449 and 1892(475) 1889(464) ; 1325(481)
g450 and 1889(464) ; 1893(482)
g451 and 1294(465) 1293(476) ; 1295(483)
g452 and 336(467) ; 340(484)
g453 and 336(467) ; 1897(485)
g454 and 336(467) ; 1905(486)
g455 and 1829(463) 1822(431) ; 1238(487)
g456 and 1729(468) ; 1733(488)
g457 and 1737(469) ; 1741(489)
g458 and 410(470) ; 1894(490)
g459 and 410(470) ; 1902(491)
g460 and 314(471) ; 343(492)
g461 and 314(471) ; 1801(493)
g462 and 1732(313) 1729(468) ; 1081(494)
g463 and 1740(314) 1737(469) ; 1093(495)
g464 and 1670(472) ; 1676(496)
g465 and 1678(473) ; 1684(497)
g466 and 407(474) ; 1340(498)
g467 and 407(474) ; 1352(499)
g468 and 1761(477) ; 1765(500)
g469 and 1769(478) ; 1773(501)
g470 and 265(479) ; 1673(502)
g471 and 265(479) ; 1681(503)
g472 and 1298(201) 1295(483) ; 391(504)
g473 and 1238(487) 1237(462) ; 1239(505)
g474 and 1295(483) ; 1299(506)
g475 and 1804(466) 1801(493) ; 1187(507)
g476 and 340(484) ; 1122(508)
g477 and 340(484) ; 1134(509)
g478 and 1897(485) ; 1901(510)
g479 and 1905(486) ; 1909(511)
g480 and 1894(490) ; 1900(512)
g481 and 1902(491) ; 1908(513)
g482 and 343(492) ; 1758(514)
g483 and 343(492) ; 1766(515)
g484 and 1801(493) ; 1805(516)
g485 and 1733(488) 1726(234) ; 1082(517)
g486 and 1741(489) 1734(235) ; 1094(518)
g487 and 1676(496) 1673(502) ; 1003(519)
g488 and 1684(497) 1681(503) ; 1013(520)
g489 and 1340(498) ; 1348(521)
g490 and 1352(499) ; 1360(522)
g491 and 1893(482) 1886(455) ; 1326(523)
g492 and 1673(502) ; 1677(524)
g493 and 1681(503) ; 1685(525)
g494 and 1299(506) 1290(115) ; 392(526)
g495 and 1239(505) ; 1243(527)
g496 and 1326(523) 1325(481) ; 1327(528)
g497 and 1805(516) 1798(448) ; 1188(529)
g498 and 1122(508) ; 1130(530)
g499 and 1134(509) ; 1142(531)
g500 and 1900(512) 1897(485) ; 1343(532)
g501 and 1908(513) 1905(486) ; 1355(533)
g502 and 1901(510) 1894(490) ; 1344(534)
g503 and 1909(511) 1902(491) ; 1356(535)
g504 and 1758(514) ; 1764(536)
g505 and 1766(515) ; 1772(537)
g506 and 1082(517) 1081(494) ; 1083(538)
g507 and 1094(518) 1093(495) ; 1095(539)
g508 and 1677(524) 1670(472) ; 1004(540)
g509 and 1685(525) 1678(473) ; 1014(541)
g510 and 1242(457) 1239(505) ; 377(542)
g511 and 1765(500) 1758(514) ; 1126(543)
g512 and 1773(501) 1766(515) ; 1138(544)
g513 and 1086(269) 1083(538) ; 1088(545)
g514 and 1098(270) 1095(539) ; 324(546)
g515 and 1330(390) 1327(528) ; 399(547)
g516 and 392(526) 391(504) ; 393(548)
g517 and 1327(528) ; 1331(549)
g518 and 1188(529) 1187(507) ; 1189(550)
g519 and 1344(534) 1343(532) ; 1345(551)
g520 and 1356(535) 1355(533) ; 1357(552)
g521 and 1083(538) ; 1087(553)
g522 and 1095(539) ; 1099(554)
g523 and 1004(540) 1003(519) ; 1005(555)
g524 and 1014(541) 1013(520) ; 1015(556)
g525 and 1243(527) 1234(440) ; 378(557)
g526 and 1764(536) 1761(477) ; 1125(558)
g527 and 1772(537) 1769(478) ; 1137(559)
g528 and 918(45) 393(548) ; 449(560)
g529 and 1087(553) 1078(195) ; 1089(561)
g530 and 1099(554) 1090(196) ; 325(562)
g531 and 1331(549) 1322(361) ; 400(563)
g532 and 393(548) ; 1397(564)
g533 and 1192(399) 1189(550) ; 364(565)
g534 and 1189(550) ; 1193(566)
g535 and 1345(551) ; 1349(567)
g536 and 1357(552) ; 1361(568)
g537 and 1008(434) 1005(555) ; 280(569)
g538 and 1018(435) 1015(556) ; 277(570)
g539 and 1005(555) ; 1009(571)
g540 and 1015(556) ; 1019(572)
g541 and 1348(521) 1345(551) ; 1350(573)
g542 and 1360(522) 1357(552) ; 413(574)
g543 and 378(557) 377(542) ; 379(575)
g544 and 1126(543) 1125(558) ; 1127(576)
g545 and 1138(544) 1137(559) ; 1139(577)
g546 and 918(45) 379(575) ; 445(578)
g547 and 449(560) ; 1493(579)
g548 and 449(560) ; 1501(580)
g549 and 1089(561) 1088(545) ; 1689(581)
g550 and 325(562) 324(546) ; 326(582)
g551 and 400(563) 399(547) ; 401(583)
g552 and 1397(564) ; 1401(584)
g553 and 1193(566) 1184(370) ; 365(585)
g554 and 1130(530) 1127(576) ; 1132(586)
g555 and 1142(531) 1139(577) ; 346(587)
g556 and 1009(571) 1000(410) ; 281(588)
g557 and 1019(572) 1010(411) ; 278(589)
g558 and 1349(567) 1340(498) ; 1351(590)
g559 and 1361(568) 1352(499) ; 414(591)
g560 and 379(575) ; 1389(592)
g561 and 1127(576) ; 1131(593)
g562 and 1139(577) ; 1143(594)
g563 and 445(578) ; 1477(595)
g564 and 445(578) ; 1485(596)
g565 and 1493(579) ; 1497(597)
g566 and 1501(580) ; 1505(598)
g567 and 918(45) 401(583) ; 453(599)
g568 and 1496(185) 1493(579) ; 559(600)
g569 and 1504(186) 1501(580) ; 556(601)
g570 and 1689(581) ; 1693(602)
g571 and 326(582) ; 1365(603)
g572 and 401(583) ; 1405(604)
g573 and 365(585) 364(565) ; 366(605)
g574 and 1131(593) 1122(508) ; 1133(606)
g575 and 1143(594) 1134(509) ; 347(607)
g576 and 281(588) 280(569) ; 282(608)
g577 and 278(589) 277(570) ; 279(609)
g578 and 1351(590) 1350(573) ; 1809(610)
g579 and 414(591) 413(574) ; 415(611)
g580 and 1389(592) ; 1393(612)
g581 and 1477(595) ; 1481(613)
g582 and 1485(596) ; 1489(614)
g583 and 453(599) ; 1429(615)
g584 and 453(599) ; 1437(616)
g585 and 1497(597) 1490(103) ; 560(617)
g586 and 1505(598) 1498(104) ; 557(618)
g587 and 1480(187) 1477(595) ; 547(619)
g588 and 1488(188) 1485(596) ; 544(620)
g589 and 1365(603) ; 1369(621)
g590 and 1405(604) ; 1409(622)
g591 and 366(605) ; 367(623)
g592 and 1133(606) 1132(586) ; 1774(624)
g593 and 347(607) 346(587) ; 348(625)
g594 and 282(608) ; 1686(626)
g595 and 282(608) ; 1362(627)
g596 and 279(609) ; 285(628)
g597 and 1809(610) ; 1813(629)
g598 and 415(611) ; 1378(630)
g599 and 853(97) 285(628) ; 1910(631)
g600 and 367(623) 856(98) ; 1918(632)
g601 and 1429(615) ; 1433(633)
g602 and 1437(616) ; 1441(634)
g603 and 560(617) 559(600) ; 561(635)
g604 and 557(618) 556(601) ; 558(636)
g605 and 1481(613) 1474(105) ; 548(637)
g606 and 1489(614) 1482(106) ; 545(638)
g607 and 1781(480) 1774(624) ; 1148(639)
g608 and 1693(602) 1686(626) ; 1024(640)
g609 and 1369(621) 1362(627) ; 417(641)
g610 and 1432(336) 1429(615) ; 511(642)
g611 and 1440(337) 1437(616) ; 508(643)
g612 and 1385(425) 1378(630) ; 424(644)
g613 and 1774(624) ; 1780(645)
g614 and 348(625) ; 1370(646)
g615 and 1686(626) ; 1692(647)
g616 and 1362(627) ; 1368(648)
g617 and 1378(630) ; 1384(649)
g618 and 1910(631) ; 1916(650)
g619 and 1918(632) ; 1924(651)
g620 and 561(635) ; 719(652)
g621 and 561(635) ; 722(653)
g622 and 558(636) ; 564(654)
g623 and 548(637) 547(619) ; 549(655)
g624 and 545(638) 544(620) ; 546(656)
g625 and 1377(460) 1370(646) ; 421(657)
g626 and 1780(645) 1777(461) ; 1147(658)
g627 and 1692(647) 1689(581) ; 1023(659)
g628 and 1368(648) 1365(603) ; 416(660)
g629 and 1433(633) 1426(274) ; 512(661)
g630 and 1441(634) 1434(275) ; 509(662)
g631 and 1384(649) 1381(392) ; 423(663)
g632 and 1370(646) ; 1376(664)
g633 and 549(655) ; 725(665)
g634 and 549(655) ; 728(666)
g635 and 546(656) ; 552(667)
g636 and 1376(664) 1373(443) ; 420(668)
g637 and 1148(639) 1147(658) ; 1149(669)
g638 and 1024(640) 1023(659) ; 1025(670)
g639 and 417(641) 416(660) ; 418(671)
g640 and 512(661) 511(642) ; 513(672)
g641 and 509(662) 508(643) ; 510(673)
g642 and 424(644) 423(663) ; 425(674)
g643 and 918(45) 425(674) ; 441(675)
g644 and 725(665) 719(652) ; 731(676)
g645 and 728(666) 719(652) ; 756(677)
g646 and 725(665) 722(653) ; 746(678)
g647 and 728(666) 722(653) ; 770(679)
g648 and 421(657) 420(668) ; 422(680)
g649 and 1149(669) ; 1153(681)
g650 and 1025(670) ; 1029(682)
g651 and 418(671) ; 419(683)
g652 and 513(672) ; 663(684)
g653 and 513(672) ; 666(685)
g654 and 510(673) ; 516(686)
g655 and 918(45) 419(683) ; 433(687)
g656 and 918(45) 422(680) ; 437(688)
g657 and 441(675) ; 1461(689)
g658 and 441(675) ; 1469(690)
g659 and 433(687) ; 1413(691)
g660 and 433(687) ; 1421(692)
g661 and 437(688) ; 1445(693)
g662 and 437(688) ; 1453(694)
g663 and 1461(689) ; 1465(695)
g664 and 1469(690) ; 1473(696)
g665 and 1464(189) 1461(689) ; 535(697)
g666 and 1472(190) 1469(690) ; 532(698)
g667 and 1413(691) ; 1417(699)
g668 and 1421(692) ; 1425(700)
g669 and 1445(693) ; 1449(701)
g670 and 1453(694) ; 1457(702)
g671 and 1465(695) 1458(107) ; 536(703)
g672 and 1473(696) 1466(108) ; 533(704)
g673 and 1448(191) 1445(693) ; 523(705)
g674 and 1456(192) 1453(694) ; 520(706)
g675 and 1416(339) 1413(691) ; 498(707)
g676 and 1424(340) 1421(692) ; 495(708)
g677 and 536(703) 535(697) ; 537(709)
g678 and 533(704) 532(698) ; 534(710)
g679 and 1449(701) 1442(109) ; 524(711)
g680 and 1457(702) 1450(110) ; 521(712)
g681 and 1417(699) 1410(279) ; 499(713)
g682 and 1425(700) 1418(280) ; 496(714)
g683 and 537(709) ; 669(715)
g684 and 537(709) ; 672(716)
g685 and 534(710) ; 540(717)
g686 and 524(711) 523(705) ; 525(718)
g687 and 521(712) 520(706) ; 522(719)
g688 and 499(713) 498(707) ; 500(720)
g689 and 496(714) 495(708) ; 497(721)
g690 and 525(718) ; 618(722)
g691 and 522(719) ; 528(723)
g692 and 525(718) 615(272) ; 639(724)
g693 and 669(715) 663(684) ; 675(725)
g694 and 672(716) 663(684) ; 696(726)
g695 and 669(715) 666(685) ; 688(727)
g696 and 672(716) 666(685) ; 710(728)
g697 and 500(720) 566(277) ; 588(729)
g698 and 500(720) ; 569(730)
g699 and 497(721) ; 503(731)
g700 and 618(722) 614(271) ; 621(732)
g701 and 618(722) 615(272) ; 622(733)
g702 and 639(724) ; 639A(734)
g703 and 639(724) ; 639B(735)
g704 and 487(197) 503(731) 528(723) 482(202) 540(717) 552(667) 564(654) 516(686) ; 867(736)
g705 and 569(730) 565(276) ; 572(737)
g706 and 569(730) 566(277) ; 573(738)
g707 and 588(729) ; 588A(739)
g708 and 588(729) ; 588B(740)
g709 and 932(40) 867(736) 949(33) ; 73(741)